C0551559|T185|relax|11488-4|LNC|Consult|Consult note
C0551559|T185|relax|34099-2|LNC|Cardiology Consult|Cardiology Consult note
C0551559|T185|relax|34756-7|LNC|Dentistry Consult|Dentistry Consult note
C0551559|T185|relax|34758-3|LNC|Dermatology Consult|Dermatology Consult note
C0551559|T185|relax|34760-9|LNC|Diabetes Consult|Diabetology Consult note
C0551559|T185|relax|34879-7|LNC|Endocrinology Consult|Endocrinology Consult note
C0551559|T185|relax|34761-7|LNC|Gastroenterology Consult|Gastroenterology Consult note
C0551559|T185|relax|34764-1|LNC|General Medicine Consult|General Medicine Consult note
C0551559|T185|relax|34776-5|LNC|Gerontology Consult|Gerontology Consult note
C0551559|T185|relax|34779-9|LNC|Hematology Medical Oncology Consult|Hematology + Medical Oncology Consult note
C0551559|T185|relax|34781-5|LNC|Infectious Disease Consult|Infectious Disease Consult note
C0551559|T185|relax|72555-6|LNC|Interventional Radiology Consult|Interventional Radiology Consult note
C0551559|T185|relax|34783-1|LNC|Kinesiotherapy Consult|Kinesiotherapy Consult note
C0551559|T185|relax|34785-6|LNC|Mental Health Consult|Mental Health Consult note
C0551559|T185|relax|34795-5|LNC|Nephrology Consult|Nephrology Consult note
C0551559|T185|relax|34798-9|LNC|Neurological Surgery Consult|Neurological Surgery Consult note
C0551559|T185|relax|34797-1|LNC|Neurology Consult|Neurology Consult note
C0551559|T185|relax|34800-3|LNC|Nutrition and Dietetics Consult|Nutrition and Dietetics Consult note
C0551559|T185|relax|34777-3|LNC|Obstetrics and Gynecology Consult|Obstetrics and Gynecology Consult note
C0551559|T185|relax|34803-7|LNC|Occupational Health Consult|Occupational Health Consult note
C0551559|T185|relax|34855-7|LNC|Occupational Therapy Consult|Occupational Therapy Consult note
C0551559|T185|relax|34805-2|LNC|Oncology Consult|Oncology Consult note
C0551559|T185|relax|34807-8|LNC|Ophthalmology Consult|Ophthalmology Consult note
C0551559|T185|relax|34810-2|LNC|Optometry Consult|Optometry Consult note
C0551559|T185|relax|34812-8|LNC|Oromaxillofacial Surgery Consult|Oromaxillofacial Surgery Consult note
C0551559|T185|relax|34814-4|LNC|Orthopedics Consult|Orthopedics Consult note
C0551559|T185|relax|34816-9|LNC|Otorhinolaryngology Consult|Otorhinolaryngology Consult note
C0551559|T185|relax|60570-9|LNC|Pathology Consult|Pathology Consult note
C0551559|T185|relax|34820-1|LNC|Pharmacy Consult|Pharmacy Consult note
C0551559|T185|relax|34822-7|LNC|Physical Medicine and Rehabilitation Consult|Physical Medicine and Rehabilitation Consult note
C0551559|T185|relax|34824-3|LNC|Physical Therapy Consult|Physical Therapy Consult note
C0551559|T185|relax|34826-8|LNC|Plastic Surgery Consult|Plastic Surgery Consult note
C0551559|T185|relax|34828-4|LNC|Podiatry Consult|Podiatry Consult note
C0551559|T185|relax|34788-0|LNC|Psychiatry Consult|Psychiatry Consult note
C0551559|T185|relax|34791-4|LNC|Psychology Consult|Psychology Consult note
C0551559|T185|relax|34103-2|LNC|Pulmonary Consult|Pulmonary Consult note
C0551559|T185|relax|34831-8|LNC|Radiation Oncology Consult|Radiation Oncology Consult note
C0551559|T185|relax|73575-3|LNC|Radiology Consult|Radiology Consult note
C0551559|T185|relax|34833-4|LNC|Recreational Therapy Consult|Recreational Therapy Consult note
C0551559|T185|relax|34835-9|LNC|Rehabilitation Consult|Rehabilitation Consult note
C0551559|T185|relax|34837-5|LNC|Respiratory Therapy Consult|Respiratory Therapy Consult note
C0551559|T185|relax|34839-1|LNC|Rheumatology Consult|Rheumatology Consult note
C0551559|T185|relax|34841-7|LNC|Social Work Consult|Social Work Consult note
C0551559|T185|relax|34845-8|LNC|Speech-language pathology+Audiology Consult|Speech-language pathology+Audiology Consult note
C0551559|T185|relax|34847-4|LNC|Surgery Consult|Surgery Consult note
C0551559|T185|relax|34849-0|LNC|Thoracic surgery Consult|Thoracic surgery Consult note
C0551559|T185|relax|34851-6|LNC|Urology Consult|Urology Consult note
C0551559|T185|relax|34853-2|LNC|Vascular surgery Consult|Vascular surgery Consult note
C0551559|T185|relax|51846-4|LNC|Emergency department Consult|Emergency department Consult note
C0551559|T185|relax|34104-0|LNC|Hospital Consult|Hospital Consult note
C0551559|T185|relax|68619-6|LNC|Adolescent medicine Hospital Consult|Adolescent medicine Hospital Consult note
C0551559|T185|relax|68633-7|LNC|Allergy and immunology Hospital Consult|Allergy and immunology Hospital Consult note
C0551559|T185|relax|68639-4|LNC|Audiology Hospital Consult|Audiology Hospital Consult note
C0551559|T185|relax|68486-0|LNC|Cardiovascular disease.medical student Hospital Consult|Cardiovascular disease.medical student Hospital Consult note
C0551559|T185|relax|68648-5|LNC|Child and adolescent psychiatry Hospital Consult|Child and adolescent psychiatry Hospital Consult note
C0551559|T185|relax|68651-9|LNC|Clinical biochemical genetics Hospital Consult|Clinical biochemical genetics Hospital Consult note
C0551559|T185|relax|68661-8|LNC|Clinical genetics Hospital Consult|Clinical genetics Hospital Consult note
C0551559|T185|relax|64072-2|LNC|Critical care medicine.medical student Hospital Consult|Critical care medicine.medical student Hospital Consult note
C0551559|T185|relax|68551-1|LNC|Dermatology Hospital Consult|Dermatology Hospital Consult note
C0551559|T185|relax|68670-9|LNC|Developmental-behavioral pediatrics Hospital Consult|Developmental-behavioral pediatrics Hospital Consult note
C0551559|T185|relax|64056-5|LNC|General medicine.medical student Hospital Consult|General medicine.medical student Hospital Consult note
C0551559|T185|relax|68681-6|LNC|Multi-specialty program Hospital Consult|Multi-specialty program Hospital Consult note
C0551559|T185|relax|68685-7|LNC|Neonatal perinatal medicine Hospital Consult|Neonatal perinatal medicine Hospital Consult note
C0551559|T185|relax|68694-9|LNC|Neurological surgery Hospital Consult|Neurological surgery Hospital Consult note
C0551559|T185|relax|68705-3|LNC|Neurology with special qualifications in child neurology Hospital Consult|Neurology with special qualifications in child neurology Hospital Consult note
C0551559|T185|relax|68566-9|LNC|Obstetrics and Gynecology Hospital Consult|Obstetrics and Gynecology Hospital Consult note
C0551559|T185|relax|68570-1|LNC|Occupational therapy Hospital Consult|Occupational therapy Hospital Consult note
C0551559|T185|relax|68575-0|LNC|Ophthalmology Hospital Consult|Ophthalmology Hospital Consult note
C0551559|T185|relax|68584-2|LNC|Orthopedic surgery Hospital Consult|Orthopedic surgery Hospital Consult note
C0551559|T185|relax|68716-0|LNC|Pain medicine Hospital Consult|Pain medicine Hospital Consult note
C0551559|T185|relax|68469-6|LNC|Pastoral care Hospital Consult|Pastoral care Hospital Consult note
C0551559|T185|relax|68727-7|LNC|Pediatric cardiology Hospital Consult|Pediatric cardiology Hospital Consult note
C0551559|T185|relax|68892-9|LNC|Pediatric dermatology Hospital Consult|Pediatric dermatology Hospital Consult note
C0551559|T185|relax|68897-8|LNC|Pediatric endocrinology Hospital Consult|Pediatric endocrinology Hospital Consult note
C0551559|T185|relax|68746-7|LNC|Pediatric gastroenterology Hospital Consult|Pediatric gastroenterology Hospital Consult note
C0551559|T185|relax|68757-4|LNC|Pediatric hematology-oncology Hospital Consult|Pediatric hematology-oncology Hospital Consult note
C0551559|T185|relax|68765-7|LNC|Pediatric infectious diseases Hospital Consult|Pediatric infectious diseases Hospital Consult note
C0551559|T185|relax|68869-7|LNC|Pediatric nephrology Hospital Consult|Pediatric nephrology Hospital Consult note
C0551559|T185|relax|68874-7|LNC|Pediatric otolaryngology Hospital Consult|Pediatric otolaryngology Hospital Consult note
C0551559|T185|relax|68787-1|LNC|Pediatric pulmonology Hospital Consult|Pediatric pulmonology Hospital Consult note
C0551559|T185|relax|68879-6|LNC|Pediatric rheumatology Hospital Consult|Pediatric rheumatology Hospital Consult note
C0551559|T185|relax|68802-8|LNC|Pediatric surgery Hospital Consult|Pediatric surgery Hospital Consult note
C0551559|T185|relax|68864-8|LNC|Pediatric transplant hepatology Hospital Consult|Pediatric transplant hepatology Hospital Consult note
C0551559|T185|relax|68812-7|LNC|Pediatric urology Hospital Consult|Pediatric urology Hospital Consult note
C0551559|T185|relax|68821-8|LNC|Pediatrics Hospital Consult|Pediatrics Hospital Consult note
C0551559|T185|relax|68586-7|LNC|Pharmacy Hospital Consult|Pharmacy Hospital Consult note
C0551559|T185|relax|68590-9|LNC|Physical therapy Hospital Consult|Physical therapy Hospital Consult note
C0551559|T185|relax|68597-4|LNC|Plastic surgery Hospital Consult|Plastic surgery Hospital Consult note
C0551559|T185|relax|68837-4|LNC|Primary care Hospital Consult|Primary care Hospital Consult note
C0551559|T185|relax|34102-4|LNC|Psychiatry Hospital Consult|Psychiatry Hospital Consult note
C0551559|T185|relax|64080-5|LNC|Pulmonary disease.medical student Hospital Consult|Pulmonary disease.medical student Hospital Consult note
C0551559|T185|relax|68846-5|LNC|Speech-language pathology Hospital Consult|Speech-language pathology Hospital Consult note
C0551559|T185|relax|64068-0|LNC|Surgery medical student Hospital Consult|Surgery medical student Hospital Consult note
C0551559|T185|relax|64076-3|LNC|Thoracic surgery.medical student Hospital Consult|Thoracic surgery.medical student Hospital Consult note
C0551559|T185|relax|68852-3|LNC|Transplant surgery Hospital Consult|Transplant surgery Hospital Consult note
C0551559|T185|relax|34100-8|LNC|Intensive care unit Consult|Intensive care unit Consult note
C0551559|T185|relax|51854-8|LNC|Long term care facility Consult|Long term care facility Consult note
C0551559|T185|relax|51845-6|LNC|Outpatient Consult|Outpatient Consult note
C0551559|T185|relax|34749-2|LNC|Anesthesiology Outpatient Consult|Anesthesiology Outpatient Consult note
C0551559|T185|relax|34101-6|LNC|General medicine Outpatient Consult|General medicine Outpatient Consult note
C0551559|T185|None|11488-4|LNC|Consult note|None
C0551559|T185|None|34099-2|LNC|Cardiology Consult note|None
C0551559|T185|None|34756-7|LNC|Dentistry Consult note|None
C0551559|T185|None|34758-3|LNC|Dermatology Consult note|None
C0551559|T185|None|34760-9|LNC|Diabetology Consult note|None
C0551559|T185|None|34879-7|LNC|Endocrinology Consult note|None
C0551559|T185|None|34761-7|LNC|Gastroenterology Consult note|None
C0551559|T185|None|34764-1|LNC|General Medicine Consult note|None
C0551559|T185|None|34776-5|LNC|Gerontology Consult note|None
C0551559|T185|None|34779-9|LNC|Hematology + Medical Oncology Consult note|None
C0551559|T185|None|34781-5|LNC|Infectious Disease Consult note|None
C0551559|T185|None|72555-6|LNC|Interventional Radiology Consult note|None
C0551559|T185|None|34783-1|LNC|Kinesiotherapy Consult note|None
C0551559|T185|None|34785-6|LNC|Mental Health Consult note|None
C0551559|T185|None|34795-5|LNC|Nephrology Consult note|None
C0551559|T185|None|34798-9|LNC|Neurological Surgery Consult note|None
C0551559|T185|None|34797-1|LNC|Neurology Consult note|None
C0551559|T185|None|34800-3|LNC|Nutrition and Dietetics Consult note|None
C0551559|T185|None|34777-3|LNC|Obstetrics and Gynecology Consult note|None
C0551559|T185|None|34803-7|LNC|Occupational Health Consult note|None
C0551559|T185|None|34855-7|LNC|Occupational Therapy Consult note|None
C0551559|T185|None|34805-2|LNC|Oncology Consult note|None
C0551559|T185|None|34807-8|LNC|Ophthalmology Consult note|None
C0551559|T185|None|34810-2|LNC|Optometry Consult note|None
C0551559|T185|None|34812-8|LNC|Oromaxillofacial Surgery Consult note|None
C0551559|T185|None|34814-4|LNC|Orthopedics Consult note|None
C0551559|T185|None|34816-9|LNC|Otorhinolaryngology Consult note|None
C0551559|T185|None|60570-9|LNC|Pathology Consult note|None
C0551559|T185|None|34820-1|LNC|Pharmacy Consult note|None
C0551559|T185|None|34822-7|LNC|Physical Medicine and Rehabilitation Consult note|None
C0551559|T185|None|34824-3|LNC|Physical Therapy Consult note|None
C0551559|T185|None|34826-8|LNC|Plastic Surgery Consult note|None
C0551559|T185|None|34828-4|LNC|Podiatry Consult note|None
C0551559|T185|None|34788-0|LNC|Psychiatry Consult note|None
C0551559|T185|None|34791-4|LNC|Psychology Consult note|None
C0551559|T185|None|34103-2|LNC|Pulmonary Consult note|None
C0551559|T185|None|34831-8|LNC|Radiation Oncology Consult note|None
C0551559|T185|None|73575-3|LNC|Radiology Consult note|None
C0551559|T185|None|34833-4|LNC|Recreational Therapy Consult note|None
C0551559|T185|None|34835-9|LNC|Rehabilitation Consult note|None
C0551559|T185|None|34837-5|LNC|Respiratory Therapy Consult note|None
C0551559|T185|None|34839-1|LNC|Rheumatology Consult note|None
C0551559|T185|None|34841-7|LNC|Social Work Consult note|None
C0551559|T185|None|34845-8|LNC|Speech-language pathology+Audiology Consult note|None
C0551559|T185|None|34847-4|LNC|Surgery Consult note|None
C0551559|T185|None|34849-0|LNC|Thoracic surgery Consult note|None
C0551559|T185|None|34851-6|LNC|Urology Consult note|None
C0551559|T185|None|34853-2|LNC|Vascular surgery Consult note|None
C0551559|T185|None|51846-4|LNC|Emergency department Consult note|None
C0551559|T185|None|34104-0|LNC|Hospital Consult note|None
C0551559|T185|None|68619-6|LNC|Adolescent medicine Hospital Consult note|None
C0551559|T185|None|68633-7|LNC|Allergy and immunology Hospital Consult note|None
C0551559|T185|None|68639-4|LNC|Audiology Hospital Consult note|None
C0551559|T185|None|68486-0|LNC|Cardiovascular disease.medical student Hospital Consult note|None
C0551559|T185|None|68648-5|LNC|Child and adolescent psychiatry Hospital Consult note|None
C0551559|T185|None|68651-9|LNC|Clinical biochemical genetics Hospital Consult note|None
C0551559|T185|None|68661-8|LNC|Clinical genetics Hospital Consult note|None
C0551559|T185|None|64072-2|LNC|Critical care medicine.medical student Hospital Consult note|None
C0551559|T185|None|68551-1|LNC|Dermatology Hospital Consult note|None
C0551559|T185|None|68670-9|LNC|Developmental-behavioral pediatrics Hospital Consult note|None
C0551559|T185|None|64056-5|LNC|General medicine.medical student Hospital Consult note|None
C0551559|T185|None|68681-6|LNC|Multi-specialty program Hospital Consult note|None
C0551559|T185|None|68685-7|LNC|Neonatal perinatal medicine Hospital Consult note|None
C0551559|T185|None|68694-9|LNC|Neurological surgery Hospital Consult note|None
C0551559|T185|None|68705-3|LNC|Neurology with special qualifications in child neurology Hospital Consult note|None
C0551559|T185|None|68566-9|LNC|Obstetrics and Gynecology Hospital Consult note|None
C0551559|T185|None|68570-1|LNC|Occupational therapy Hospital Consult note|None
C0551559|T185|None|68575-0|LNC|Ophthalmology Hospital Consult note|None
C0551559|T185|None|68584-2|LNC|Orthopedic surgery Hospital Consult note|None
C0551559|T185|None|68716-0|LNC|Pain medicine Hospital Consult note|None
C0551559|T185|None|68469-6|LNC|Pastoral care Hospital Consult note|None
C0551559|T185|None|68727-7|LNC|Pediatric cardiology Hospital Consult note|None
C0551559|T185|None|68892-9|LNC|Pediatric dermatology Hospital Consult note|None
C0551559|T185|None|68897-8|LNC|Pediatric endocrinology Hospital Consult note|None
C0551559|T185|None|68746-7|LNC|Pediatric gastroenterology Hospital Consult note|None
C0551559|T185|None|68757-4|LNC|Pediatric hematology-oncology Hospital Consult note|None
C0551559|T185|None|68765-7|LNC|Pediatric infectious diseases Hospital Consult note|None
C0551559|T185|None|68869-7|LNC|Pediatric nephrology Hospital Consult note|None
C0551559|T185|None|68874-7|LNC|Pediatric otolaryngology Hospital Consult note|None
C0551559|T185|None|68787-1|LNC|Pediatric pulmonology Hospital Consult note|None
C0551559|T185|None|68879-6|LNC|Pediatric rheumatology Hospital Consult note|None
C0551559|T185|None|68802-8|LNC|Pediatric surgery Hospital Consult note|None
C0551559|T185|None|68864-8|LNC|Pediatric transplant hepatology Hospital Consult note|None
C0551559|T185|None|68812-7|LNC|Pediatric urology Hospital Consult note|None
C0551559|T185|None|68821-8|LNC|Pediatrics Hospital Consult note|None
C0551559|T185|None|68586-7|LNC|Pharmacy Hospital Consult note|None
C0551559|T185|None|68590-9|LNC|Physical therapy Hospital Consult note|None
C0551559|T185|None|68597-4|LNC|Plastic surgery Hospital Consult note|None
C0551559|T185|None|68837-4|LNC|Primary care Hospital Consult note|None
C0551559|T185|None|34102-4|LNC|Psychiatry Hospital Consult note|None
C0551559|T185|None|64080-5|LNC|Pulmonary disease.medical student Hospital Consult note|None
C0551559|T185|None|68846-5|LNC|Speech-language pathology Hospital Consult note|None
C0551559|T185|None|64068-0|LNC|Surgery medical student Hospital Consult note|None
C0551559|T185|None|64076-3|LNC|Thoracic surgery.medical student Hospital Consult note|None
C0551559|T185|None|68852-3|LNC|Transplant surgery Hospital Consult note|None
C0551559|T185|None|34100-8|LNC|Intensive care unit Consult note|None
C0551559|T185|None|51854-8|LNC|Long term care facility Consult note|None
C0551559|T185|None|51845-6|LNC|Outpatient Consult note|None
C0551559|T185|None|34749-2|LNC|Anesthesiology Outpatient Consult note|None
C0551559|T185|None|34101-6|LNC|General medicine Outpatient Consult note|None
C3699344|T077|strict|48765-2|LNC|ALLERGIES, ADVERSE REACTIONS, ALERTS|ALLERGIES, ADVERSE REACTIONS, ALERTS
C3699344|T077|strict|48765-2|LNC|ALLERGIES & ADVERSE REACTIONS|ALLERGIES & ADVERSE REACTIONS
C3699344|T077|strict|48765-2|LNC|ALLERGIES, ADVERSE REACTIONS & ALERTS|ALLERGIES, ADVERSE REACTIONS & ALERTS
C3699344|T077|strict|48765-2|LNC|ALLERGIES AND ADVERSE REACTIONS|ALLERGIES AND ADVERSE REACTIONS
C3699344|T077|strict|48765-2|LNC|ADVERSE DRUG REACTIONS|ADVERSE DRUG REACTIONS
C3699344|T077|strict|48765-2|LNC|ADVERSE REACTIONS|ADVERSE REACTIONS
C3699344|T077|strict|48765-2|LNC|DRUG ALLERGIES|DRUG ALLERGIES
C3699344|T077|strict|48765-2|LNC|POTENTIALLY SERIOUS INTERACTION|POTENTIALLY SERIOUS INTERACTION
C3699344|T077|strict|48765-2|LNC|SERIOUS INTERACTION|SERIOUS INTERACTION
C3699344|T077|strict|48765-2|LNC|ALLERGY LIST|ALLERGY LIST
C3699344|T077|relax|48765-2|LNC|ALERTS|ALERTS
C3699344|T077|relax|48765-2|LNC|ALLERGIES|ALLERGIES
C3699344|T077|relax|48765-2|LNC|ALLERGY|ALLERGY
C3699344|T077|strict|48765-2|LNC|ENVIRONMENTAL ALLERGIES|ENVIRONMENTAL ALLERGIES
C3699344|T077|strict|48765-2|LNC|FOOD ALLERGIES|FOOD ALLERGIES
C3699344|T077|strict|48765-2|LNC|NO KNOWN ALLERGIES|NO KNOWN ALLERGIES
C3699344|T077|strict|48765-2|LNC|NO KNOWN DRUG ALLERGIES|NO KNOWN DRUG ALLERGIES
C3699344|T077|abbr|48765-2|LNC|NKA|NKA
C3699344|T077|abbr|48765-2|LNC|NKDA|NKDA
C3699344|T077|strict|11369-6|LNC|HISTORY OF IMMUNIZATION|HISTORY OF IMMUNIZATION
C3699344|T077|strict|11369-6|LNC|HISTORY OF IMMUNIZATIONS|HISTORY OF IMMUNIZATIONS
C3699344|T077|strict|11369-6|LNC|IMMUNIZATION HISTORY|IMMUNIZATION HISTORY
C3699344|T077|strict|11369-6|LNC|IMMUNIZATIONS AND VACCINES|IMMUNIZATIONS AND VACCINES
C3699344|T077|strict|11369-6|LNC|LIST OF VACCINES|LIST OF VACCINES
C3699344|T077|strict|11369-6|LNC|VACCINES LIST|VACCINES LIST
C3699344|T077|relax|11369-6|LNC|IMMUNIZATIONS LIST|IMMUNIZATIONS LIST
C3699344|T077|relax|11369-6|LNC|IMMUNIZATION|IMMUNIZATION
C3699344|T077|relax|11369-6|LNC|IMMUNIZATIONS|IMMUNIZATIONS
C3699344|T077|relax|11369-6|LNC|VACCINE|VACCINE
C3699344|T077|relax|11369-6|LNC|VACCINES|VACCINES
C3699344|T077|strict|11369-6|LNC|IMMUNIZATIONS RECOMMENDED|IMMUNIZATIONS RECOMMENDED
C3699344|T077|strict|11366-2|LNC|HISTORY OF TOBACCO USE|HISTORY OF TOBACCO USE
C3699344|T077|strict|11366-2|LNC|SMOKING HISTORY|SMOKING HISTORY
C3699344|T077|strict|11366-2|LNC|SMOKING EXPOSURE|SMOKING EXPOSURE
C3699344|T077|strict|11366-2|LNC|SMOKING STATUS|SMOKING STATUS
C3699344|T077|strict|11366-2|LNC|TOBACCO USE|TOBACCO USE
C3699344|T077|strict|11366-2|LNC|TOBACCO USE STATUS|TOBACCO USE STATUS
C3699344|T077|relax|11366-2|LNC|SMOKING|SMOKING
C3699344|T077|relax|11366-2|LNC|TOBACCO|TOBACCO
C3699344|T077|strict|29762-2|LNC|SOCIAL HISTORY|SOCIAL HISTORY
C3699344|T077|strict|29762-2|LNC|SOCIAL HX|SOCIAL HX
C3699344|T077|strict|29762-2|LNC|POVERTY STATUS|POVERTY STATUS
C3699344|T077|relax|29762-2|LNC|DRINKING|DRINKING
C3699344|T077|relax|29762-2|LNC|PHYSICAL EXERCISE|PHYSICAL EXERCISE
C3699344|T077|relax|29762-2|LNC|EXERCISE|EXERCISE
C3699344|T077|relax|29762-2|LNC|SOCIAL|SOCIAL
C3699344|T077|relax|29762-2|LNC|HABITS|HABITS
C3699344|T077|relax|29762-2|LNC|POVERTY|POVERTY
C3699344|T077|relax|29762-2|LNC|HOMELESS|HOMELESS
C3699344|T077|abbr|29762-2|LNC|SHX|SHX
C3699344|T077|abbr|29762-2|LNC|PSH|PSH
C3699344|T077|strict|61144-2|LNC|DIET AND NUTRITION|DIET AND NUTRITION
C3699344|T077|strict|61144-2|LNC|DIET+NUTRITION|DIET+NUTRITION
C3699344|T077|relax|61144-2|LNC|DIET|DIET
C3699344|T077|relax|61144-2|LNC|NUTRITION|NUTRITION
C3699344|T077|strict|42344-2|LNC|DISCHARGE DIET|DISCHARGE DIET
C3699344|T077|strict|42348-3|LNC|ADVANCED DIRECTIVES|ADVANCED DIRECTIVES
C3699344|T077|strict|42348-3|LNC|ADVANCE DIRECTIVES|ADVANCE DIRECTIVES
C3699344|T077|relax|42348-3|LNC|DIRECTIVES|DIRECTIVES
C3699344|T077|strict|45474-4|LNC|ADVANCE DIRECTIVE - DO NOT RESUSCITATE|ADVANCE DIRECTIVE - DO NOT RESUSCITATE
C3699344|T077|strict|45474-4|LNC|DO NOT RESUSCITATE|DO NOT RESUSCITATE
C3699344|T077|abbr|45474-4|LNC|DNR|DNR
C3699344|T077|strict|47420-5|LNC|FUNCTIONAL STATUS ASSESSMENT NOTE|FUNCTIONAL STATUS ASSESSMENT NOTE
C3699344|T077|strict|47420-5|LNC|FUNCTIONAL STATUS ASSESSMENT|FUNCTIONAL STATUS ASSESSMENT
C3699344|T077|strict|47420-5|LNC|FUNCTIONAL STATUS|FUNCTIONAL STATUS
C3699344|T077|strict|47420-5|LNC|CURRENT HEALTH STATUS|CURRENT HEALTH STATUS
C3699344|T077|strict|47420-5|LNC|IMPAIRMENTS|IMPAIRMENTS
C3699344|T077|strict|47420-5|LNC|DISCHARGE CONDITION|DISCHARGE CONDITION
C3699344|T077|strict|47420-5|LNC|DISCHARGED CONDITION ON DISCHARGE|DISCHARGED CONDITION ON DISCHARGE
C3699344|T077|strict|47420-5|LNC|DISCHARGE STATUS|DISCHARGE STATUS
C3699344|T077|strict|47420-5|LNC|CONDITION ON DISCHARGE|CONDITION ON DISCHARGE
C3699344|T077|strict|47420-5|LNC|CONDITION ON TRANSFER|CONDITION ON TRANSFER
C3699344|T077|strict|30954-2|LNC|RELEVANT DIAGNOSTIC TESTS LABORATORY DATA|RELEVANT DIAGNOSTIC TESTS LABORATORY DATA
C3699344|T077|strict|30954-2|LNC|RELEVANT DIAGNOSTIC TESTS OR LABORATORY DATA|RELEVANT DIAGNOSTIC TESTS OR LABORATORY DATA
C3699344|T077|strict|30954-2|LNC|NOTABLE LABS|NOTABLE LABS
C3699344|T077|strict|30954-2|LNC|PERTINENT LAB VALUES|PERTINENT LAB VALUES
C3699344|T077|strict|30954-2|LNC|PERTINENT LABORATORY RESULTS|PERTINENT LABORATORY RESULTS
C3699344|T077|strict|30954-2|LNC|PERTINENT LABORATORY TESTS AND RESULTS|PERTINENT LABORATORY TESTS AND RESULTS
C3699344|T077|strict|30954-2|LNC|PERTINENT LABORATORY TESTS AND STUDIES|PERTINENT LABORATORY TESTS AND STUDIES
C3699344|T077|strict|30954-2|LNC|PERTINENT LABS UPON PRESENTATION|PERTINENT LABS UPON PRESENTATION
C3699344|T077|strict|30954-2|LNC|PERTINENT LABS|PERTINENT LABS
C3699344|T077|strict|30954-2|LNC|RELEVANT LABS|RELEVANT LABS
C3699344|T077|strict|30954-2|LNC|ADMISSION LAB|ADMISSION LAB
C3699344|T077|strict|30954-2|LNC|ADMISSION LABS|ADMISSION LABS
C3699344|T077|strict|30954-2|LNC|ADMISSION LABS AND STUDIES|ADMISSION LABS AND STUDIES
C3699344|T077|strict|30954-2|LNC|ADMISSION LABORATORY|ADMISSION LABORATORY
C3699344|T077|strict|30954-2|LNC|ADMISSION LABORATORIES|ADMISSION LABORATORIES
C3699344|T077|strict|30954-2|LNC|ADMISSION LABORATORY DATA|ADMISSION LABORATORY DATA
C3699344|T077|strict|30954-2|LNC|ADMISSION LABORATORY STUDIES|ADMISSION LABORATORY STUDIES
C3699344|T077|strict|30954-2|LNC|ADMISSION LABORATORY RESULTS|ADMISSION LABORATORY RESULTS
C3699344|T077|strict|30954-2|LNC|ADMISSION LABORATORY VALUES|ADMISSION LABORATORY VALUES
C3699344|T077|strict|30954-2|LNC|ADMISSIONS LABORATORIES|ADMISSIONS LABORATORIES
C3699344|T077|strict|30954-2|LNC|ADMITTING LABORATORY|ADMITTING LABORATORY
C3699344|T077|strict|30954-2|LNC|PREOPERATIVE LAB|PREOPERATIVE LAB
C3699344|T077|strict|30954-2|LNC|ADMIT LABS|ADMIT LABS
C3699344|T077|strict|30954-2|LNC|LAB STUDIES ON ADMISSION|LAB STUDIES ON ADMISSION
C3699344|T077|strict|30954-2|LNC|LABORATORIES ON ADMISSION|LABORATORIES ON ADMISSION
C3699344|T077|strict|30954-2|LNC|LABORATORY DATA AT ADMISSION|LABORATORY DATA AT ADMISSION
C3699344|T077|strict|30954-2|LNC|LABORATORY DATA ON ADMISSION|LABORATORY DATA ON ADMISSION
C3699344|T077|strict|30954-2|LNC|LABORATORY DATA UPON ADMISSION|LABORATORY DATA UPON ADMISSION
C3699344|T077|strict|30954-2|LNC|LABORATORY EXAM ON ADMISSION|LABORATORY EXAM ON ADMISSION
C3699344|T077|strict|30954-2|LNC|LABORATORY EXAMS UPON ADMISSION|LABORATORY EXAMS UPON ADMISSION
C3699344|T077|strict|30954-2|LNC|LABORATORY FINDINGS ON ADMISSION|LABORATORY FINDINGS ON ADMISSION
C3699344|T077|strict|30954-2|LNC|LABORATORY ON ADMISSION|LABORATORY ON ADMISSION
C3699344|T077|strict|30954-2|LNC|LABORATORY STUDIES ON ADMISSION|LABORATORY STUDIES ON ADMISSION
C3699344|T077|strict|30954-2|LNC|LABORATORY STUDIES UPON ADMISSION|LABORATORY STUDIES UPON ADMISSION
C3699344|T077|strict|30954-2|LNC|LABORATORY VALUES ON ADMISSION|LABORATORY VALUES ON ADMISSION
C3699344|T077|strict|30954-2|LNC|LABS AND STUDIES ON ADMISSION|LABS AND STUDIES ON ADMISSION
C3699344|T077|strict|30954-2|LNC|LABS AT ADMISSION|LABS AT ADMISSION
C3699344|T077|strict|30954-2|LNC|LABS ON ADMISSION|LABS ON ADMISSION
C3699344|T077|strict|30954-2|LNC|LABS ON ADMIT|LABS ON ADMIT
C3699344|T077|strict|30954-2|LNC|LABS UPON ADMISSION|LABS UPON ADMISSION
C3699344|T077|strict|30954-2|LNC|NOTABLE LABORATORY VALUES ON ADMISSION|NOTABLE LABORATORY VALUES ON ADMISSION
C3699344|T077|strict|30954-2|LNC|PERTINENT LABORATORY DATA ON ADMISSION|PERTINENT LABORATORY DATA ON ADMISSION
C3699344|T077|strict|30954-2|LNC|PERTINENT LABS ON ADMISSION|PERTINENT LABS ON ADMISSION
C3699344|T077|strict|30954-2|LNC|RELEVANT ADMISSION LABS|RELEVANT ADMISSION LABS
C3699344|T077|strict|30954-2|LNC|SIGNIFICANT LABS ON ADMISSION|SIGNIFICANT LABS ON ADMISSION
C3699344|T077|strict|30954-2|LNC|PREOP LABS|PREOP LABS
C3699344|T077|strict|30954-2|LNC|PREOPERATIVE LABS|PREOPERATIVE LABS
C3699344|T077|strict|30954-2|LNC|PREOPERATIVE LABORATORY DATA|PREOPERATIVE LABORATORY DATA
C3699344|T077|strict|30954-2|LNC|PREOPERATIVE LABORATORY RESULTS|PREOPERATIVE LABORATORY RESULTS
C3699344|T077|strict|30954-2|LNC|PREOPERATIVE LABORATORY VALUES|PREOPERATIVE LABORATORY VALUES
C3699344|T077|strict|30954-2|LNC|LABORATORIES OF NOTE|LABORATORIES OF NOTE
C3699344|T077|multi|30954-2|LNC|RESULTS DIAGNOSTIC FINDINGS|RESULTS DIAGNOSTIC FINDINGS
C3699344|T077|strict|30954-2|LNC|INITIAL LABORATORY DATA|INITIAL LABORATORY DATA
C3699344|T077|strict|30954-2|LNC|INITIAL LABORATORY STUDIES|INITIAL LABORATORY STUDIES
C3699344|T077|strict|30954-2|LNC|LABORATORY DATA|LABORATORY DATA
C3699344|T077|strict|30954-2|LNC|LAB RESULTS|LAB RESULTS
C3699344|T077|strict|30954-2|LNC|LABORATORY EXAM|LABORATORY EXAM
C3699344|T077|strict|30954-2|LNC|LABORATORY EVALUATION|LABORATORY EVALUATION
C3699344|T077|strict|30954-2|LNC|LABORATORY EXAMINATION|LABORATORY EXAMINATION
C3699344|T077|strict|30954-2|LNC|LABORATORY TESTS|LABORATORY TESTS
C3699344|T077|strict|30954-2|LNC|CHEMISTRY STUDIES|CHEMISTRY STUDIES
C3699344|T077|strict|30954-2|LNC|LAB VALUES|LAB VALUES
C3699344|T077|strict|30954-2|LNC|LABORATORY EXAMS|LABORATORY EXAMS
C3699344|T077|strict|30954-2|LNC|LABORATORY INFORMATION|LABORATORY INFORMATION
C3699344|T077|strict|30954-2|LNC|LABORATORY RESULTS|LABORATORY RESULTS
C3699344|T077|strict|30954-2|LNC|LABORATORY STUDIES|LABORATORY STUDIES
C3699344|T077|strict|30954-2|LNC|LABORATORY VALUES|LABORATORY VALUES
C3699344|T077|strict|30954-2|LNC|BENIGN LABS|BENIGN LABS
C3699344|T077|strict|30954-2|LNC|NORMAL LABS|NORMAL LABS
C3699344|T077|multi|30954-2|LNC|LABS AND DIAGNOSTIC STUDIES|LABS AND DIAGNOSTIC STUDIES
C3699344|T077|multi|30954-2|LNC|DIAGNOSTIC STUDIES|DIAGNOSTIC STUDIES
C3699344|T077|multi|30954-2|LNC|DIAGNOSTIC DATA|DIAGNOSTIC DATA
C3699344|T077|multi|30954-2|LNC|SHOWED THE FOLLOWING RESULTS|SHOWED THE FOLLOWING RESULTS
C3699344|T077|multi|30954-2|LNC|RESULTS SUMMARY|RESULTS SUMMARY
C3699344|T077|multi|30954-2|LNC|DIAGNOSTIC TESTS|DIAGNOSTIC TESTS
C3699344|T077|multi|30954-2|LNC|TESTS|TESTS
C3699344|T077|multi|30954-2|LNC|RESULTS|RESULTS
C3699344|T077|multi|30954-2|LNC|OBSERVATIONS|OBSERVATIONS
C3699344|T077|multi|30954-2|LNC|PERTINENT RESULTS|PERTINENT RESULTS
C3699344|T077|multi|30954-2|LNC|RESULTS/INTERPRETATION|RESULTS/INTERPRETATION
C3699344|T077|relax|30954-2|LNC|LAB DATA|LAB DATA
C3699344|T077|relax|30954-2|LNC|LABORATORIES|LABORATORIES
C3699344|T077|relax|30954-2|LNC|LABORATORY|LABORATORY
C3699344|T077|relax|30954-2|LNC|CHEMISTRIES|CHEMISTRIES
C3699344|T077|relax|30954-2|LNC|LABORATORY STUDIES WERE SENT OFF INCLUDING|LABORATORY STUDIES WERE SENT OFF INCLUDING
C3699344|T077|relax|30954-2|LNC|LABS TO FU|LABS TO FU
C3699344|T077|relax|30954-2|LNC|LABS|LABS
C3699344|T077|relax|30954-2|LNC|LAB|LAB
C3699344|T077|relax|30954-2|LNC|LAB NO|LAB NO
C3699344|T077|relax|30954-2|LNC|LAB NO.|LAB NO.
C3699344|T077|strict|664-3|LNC|GRAM STAIN FINAL|GRAM STAIN FINAL
C3699344|T077|strict|664-3|LNC|GRAM STAIN|GRAM STAIN
C3699344|T077|strict|11493-4|LNC|HOSPITAL DISCHARGE STUDIES SUMMARY|HOSPITAL DISCHARGE STUDIES SUMMARY
C3699344|T077|strict|11493-4|LNC|DISCHARGE LAB DATA|DISCHARGE LAB DATA
C3699344|T077|strict|11493-4|LNC|DISCHARGE LABORATORIES|DISCHARGE LABORATORIES
C3699344|T077|strict|11493-4|LNC|DISCHARGE LABORATORY DATA|DISCHARGE LABORATORY DATA
C3699344|T077|strict|11493-4|LNC|DISCHARGE LABORATORY VALUES|DISCHARGE LABORATORY VALUES
C3699344|T077|strict|11493-4|LNC|DISCHARGE LABS|DISCHARGE LABS
C3699344|T077|strict|11493-4|LNC|LAB VALUES ON DAY OF DISCHARGE|LAB VALUES ON DAY OF DISCHARGE
C3699344|T077|strict|11493-4|LNC|LABORATORY DATA AT DISCHARGE|LABORATORY DATA AT DISCHARGE
C3699344|T077|strict|11493-4|LNC|LABORATORY DATA ON DISCHARGE|LABORATORY DATA ON DISCHARGE
C3699344|T077|strict|11493-4|LNC|LABORATORY VALUES ON DISCHARGE|LABORATORY VALUES ON DISCHARGE
C3699344|T077|strict|11493-4|LNC|LABORATORY STUDIES ON DISCHARGE|LABORATORY STUDIES ON DISCHARGE
C3699344|T077|strict|11493-4|LNC|LABORATORY STUDIES UPON DISCHARGE|LABORATORY STUDIES UPON DISCHARGE
C3699344|T077|strict|11493-4|LNC|LABS AT DISCHARGE|LABS AT DISCHARGE
C3699344|T077|strict|11493-4|LNC|LABS AT TIME OF DISCHARGE|LABS AT TIME OF DISCHARGE
C3699344|T077|strict|11493-4|LNC|LABS ON DAY OF DISCHARGE|LABS ON DAY OF DISCHARGE
C3699344|T077|strict|11493-4|LNC|LABS ON TRANSFER|LABS ON TRANSFER
C3699344|T077|strict|11493-4|LNC|LABORATORY PENDING ON DISCHARGE|LABORATORY PENDING ON DISCHARGE
C3699344|T077|multi|61149-1|LNC|OBJECTIVE|OBJECTIVE
C3699344|T077|multi|61149-1|LNC|OBJECTIVE DATA|OBJECTIVE DATA
C3699344|T077|strict|18723-7|LNC|HEMATOLOGY STUDIES|HEMATOLOGY STUDIES
C3699344|T077|relax|18723-7|LNC|HEMATOLOGIC|HEMATOLOGIC
C3699344|T077|relax|18723-7|LNC|HEMATOLOGY|HEMATOLOGY
C3699344|T077|relax|18723-7|LNC|HEME|HEME
C3699344|T077|strict|56846-9|LNC|CARDIAC BIOMARKERS|CARDIAC BIOMARKERS
C3699344|T077|strict|56846-9|LNC|LIPID PANEL|LIPID PANEL
C3699344|T077|strict|56846-9|LNC|METABOLIC PANEL|METABOLIC PANEL
C3699344|T077|relax|56846-9|LNC|CHOLESTEROL|CHOLESTEROL
C3699344|T077|strict|18729-4|LNC|URINALYSIS STUDIES|URINALYSIS STUDIES
C3699344|T077|strict|18729-4|LNC|URINALYSIS|URINALYSIS
C3699344|T077|strict|18729-4|LNC|URINE OUTPUT|URINE OUTPUT
C3699344|T077|strict|18720-3|LNC|COAGULATION STUDIES|COAGULATION STUDIES
C3699344|T077|strict|18728-6|LNC|TOXICOLOGY STUDIES|TOXICOLOGY STUDIES
C3699344|T077|relax|18728-6|LNC|TOXICOLOGY|TOXICOLOGY
C3699344|T077|strict|56874-1|LNC|SEROLOGY AND BLOOD BANK STUDIES|SEROLOGY AND BLOOD BANK STUDIES
C3699344|T077|relax|56874-1|LNC|SEROLOGY|SEROLOGY
C3699344|T077|strict|18725-2|LNC|MICROBIOLOGY STUDIES|MICROBIOLOGY STUDIES
C3699344|T077|relax|18725-2|LNC|MICROBIOLOGY|MICROBIOLOGY
C3699344|T077|relax|56847-7|LNC|CALCULATED AND DERIVED VALUES|CALCULATED AND DERIVED VALUES
C3699344|T077|relax|56847-7|LNC|DERIVED VALUES|DERIVED VALUES
C3699344|T077|strict|10160-0|LNC|HISTORY OF MEDICATION USE|HISTORY OF MEDICATION USE
C3699344|T077|strict|10160-0|LNC|MEDICATION LIST|MEDICATION LIST
C3699344|T077|strict|10160-0|LNC|LIST MEDICATIONS|LIST MEDICATIONS
C3699344|T077|strict|10160-0|LNC|FINAL MEDICATIONS|FINAL MEDICATIONS
C3699344|T077|strict|10160-0|LNC|CONDITION MEDICATIONS|CONDITION MEDICATIONS
C3699344|T077|strict|10160-0|LNC|CURRENT MEDICATIONS|CURRENT MEDICATIONS
C3699344|T077|strict|10160-0|LNC|AS NEEDED MEDICATIONS|AS NEEDED MEDICATIONS
C3699344|T077|strict|10160-0|LNC|THE FOLLOWING MEDICATIONS|THE FOLLOWING MEDICATIONS
C3699344|T077|strict|10160-0|LNC|FOLLOWING MEDICATIONS|FOLLOWING MEDICATIONS
C3699344|T077|strict|10160-0|LNC|DRUG HISTORY|DRUG HISTORY
C3699344|T077|strict|10160-0|LNC|HOME MEDICATIONS|HOME MEDICATIONS
C3699344|T077|strict|10160-0|LNC|MEDICATIONS AT HOME|MEDICATIONS AT HOME
C3699344|T077|strict|10160-0|LNC|INHOSPITAL MEDICATIONS|INHOSPITAL MEDICATIONS
C3699344|T077|strict|10160-0|LNC|MOST RECENT MEDICATIONS|MOST RECENT MEDICATIONS
C3699344|T077|strict|10160-0|LNC|NEW MEDICATIONS|NEW MEDICATIONS
C3699344|T077|strict|10160-0|LNC|MEDICATION CHANGES|MEDICATION CHANGES
C3699344|T077|strict|10160-0|LNC|MEDICATIONS AT REHAB|MEDICATIONS AT REHAB
C3699344|T077|strict|10160-0|LNC|MEDICATIONS AT REHABILITATION|MEDICATIONS AT REHABILITATION
C3699344|T077|strict|10160-0|LNC|MEDICATIONS ON PRESENTATION|MEDICATIONS ON PRESENTATION
C3699344|T077|strict|10160-0|LNC|OUTPATIENT MEDICATIONS|OUTPATIENT MEDICATIONS
C3699344|T077|strict|10160-0|LNC|NUMBER OF DOSES REQUIRED APPROXIMATE|NUMBER OF DOSES REQUIRED APPROXIMATE
C3699344|T077|relax|10160-0|LNC|MEDS AT HOME|MEDS AT HOME
C3699344|T077|relax|10160-0|LNC|MEDS|MEDS
C3699344|T077|relax|10160-0|LNC|PRESCRIPTIONS|PRESCRIPTIONS
C3699344|T077|relax|10160-0|LNC|PRN MEDICATIONS|PRN MEDICATIONS
C3699344|T077|relax|10160-0|LNC|MEDICATIONS|MEDICATIONS
C3699344|T077|relax|10160-0|LNC|MEDICATION|MEDICATION
C3699344|T077|strict|29549-3|LNC|MEDICATIONS ADMINISTERED|MEDICATIONS ADMINISTERED
C3699344|T077|strict|29549-3|LNC|MEDICATION ADMINISTERED|MEDICATION ADMINISTERED
C3699344|T077|strict|29549-3|LNC|FLUIDS RECEIVED|FLUIDS RECEIVED
C3699344|T077|strict|29549-3|LNC|IV FLUIDS|IV FLUIDS
C3699344|T077|relax|29549-3|LNC|FLUIDS|FLUIDS
C3699344|T077|strict|42346-7|LNC|MEDICATIONS ON ADMISSION|MEDICATIONS ON ADMISSION
C3699344|T077|strict|42346-7|LNC|MEDICATIONS AT ADMISSION|MEDICATIONS AT ADMISSION
C3699344|T077|strict|42346-7|LNC|MEDICATIONS AT ADMISSION INCLUDE|MEDICATIONS AT ADMISSION INCLUDE
C3699344|T077|strict|42346-7|LNC|MEDICATIONS UPON ADMISSION|MEDICATIONS UPON ADMISSION
C3699344|T077|strict|42346-7|LNC|MEDICATIONS PRIOR TO ADMISSION|MEDICATIONS PRIOR TO ADMISSION
C3699344|T077|strict|42346-7|LNC|PREADMISSION MEDICATIONS|PREADMISSION MEDICATIONS
C3699344|T077|strict|42346-7|LNC|PREOP MEDICATIONS|PREOP MEDICATIONS
C3699344|T077|strict|42346-7|LNC|PREOPERATIVE MEDICATIONS|PREOPERATIVE MEDICATIONS
C3699344|T077|strict|42346-7|LNC|MEDICATIONS AT THE TIME OF ADMISSION|MEDICATIONS AT THE TIME OF ADMISSION
C3699344|T077|strict|42346-7|LNC|MEDICATIONS AT TIME OF ADMISSION|MEDICATIONS AT TIME OF ADMISSION
C3699344|T077|strict|42346-7|LNC|MEDICATION CHANGES MADE DURING THIS ADMISSION|MEDICATION CHANGES MADE DURING THIS ADMISSION
C3699344|T077|strict|42346-7|LNC|ADMISSION MEDICATIONS|ADMISSION MEDICATIONS
C3699344|T077|strict|42346-7|LNC|HOME MEDICATIONS ON ADMISSION|HOME MEDICATIONS ON ADMISSION
C3699344|T077|strict|42346-7|LNC|BLOCK MEDICATIONS ON ADMISSION|BLOCK MEDICATIONS ON ADMISSION
C3699344|T077|relax|42346-7|LNC|RX ON ADMIT|RX ON ADMIT
C3699344|T077|strict|10183-2|LNC|HOSPITAL DISCHARGE MEDICATIONS|HOSPITAL DISCHARGE MEDICATIONS
C3699344|T077|strict|75311-1|LNC|DISCHARGE MEDICATIONS|DISCHARGE MEDICATIONS
C3699344|T077|strict|75311-1|LNC|DISCHARGE MEDICATIONS INCLUDE|DISCHARGE MEDICATIONS INCLUDE
C3699344|T077|strict|75311-1|LNC|DISCHARGE MEDICATION|DISCHARGE MEDICATION
C3699344|T077|strict|75311-1|LNC|DISCHARGED TO HOME ON THE FOLLOWING MEDICATIONS|DISCHARGED TO HOME ON THE FOLLOWING MEDICATIONS
C3699344|T077|strict|75311-1|LNC|ADDENDUM TO MEDICATIONS ON DISCHARGE|ADDENDUM TO MEDICATIONS ON DISCHARGE
C3699344|T077|strict|75311-1|LNC|REHABILITATION HOSPITAL DISCHARGE MEDICATIONS|REHABILITATION HOSPITAL DISCHARGE MEDICATIONS
C3699344|T077|strict|75311-1|LNC|A REHABILITATION HOSPITAL DISCHARGE MEDICATIONS|A REHABILITATION HOSPITAL DISCHARGE MEDICATIONS
C3699344|T077|strict|75311-1|LNC|MEDICATIONS UPON DISCHARGE|MEDICATIONS UPON DISCHARGE
C3699344|T077|strict|75311-1|LNC|MEDICATION AT THE TIME OF DISCHARGE|MEDICATION AT THE TIME OF DISCHARGE
C3699344|T077|strict|75311-1|LNC|MEDICATION AT TIME OF DISCHARGE|MEDICATION AT TIME OF DISCHARGE
C3699344|T077|strict|75311-1|LNC|MEDICATIONS AT THAT TIME OF DISCHARGE|MEDICATIONS AT THAT TIME OF DISCHARGE
C3699344|T077|strict|75311-1|LNC|MEDICATIONS AT THE TIME OF DISCHARGE|MEDICATIONS AT THE TIME OF DISCHARGE
C3699344|T077|strict|75311-1|LNC|MEDICATIONS AT TIME OF DISCHARGE|MEDICATIONS AT TIME OF DISCHARGE
C3699344|T077|strict|75311-1|LNC|MEDICATIONS ON DISCHARGE|MEDICATIONS ON DISCHARGE
C3699344|T077|strict|75311-1|LNC|MEDICATION ON DISCHARGE|MEDICATION ON DISCHARGE
C3699344|T077|strict|75311-1|LNC|MEDICATIONS AT DISCHARGE|MEDICATIONS AT DISCHARGE
C3699344|T077|strict|75311-1|LNC|MEDICATIONS UPON TRANSFER|MEDICATIONS UPON TRANSFER
C3699344|T077|strict|75311-1|LNC|MEDICATIONS ON TRANSFER|MEDICATIONS ON TRANSFER
C3699344|T077|strict|75311-1|LNC|TRANSFER MEDICATIONS|TRANSFER MEDICATIONS
C3699344|T077|strict|75311-1|LNC|MEDICATIONS AT THE TIME OF TRANSFER|MEDICATIONS AT THE TIME OF TRANSFER
C3699344|T077|strict|75311-1|LNC|MEDICATIONS AT THE TIME OF TRANSFER TO THE CCU|MEDICATIONS AT THE TIME OF TRANSFER TO THE CCU
C3699344|T077|strict|75311-1|LNC|MEDICATIONS AT THE TIME OF TRANSFER TO THE ICU|MEDICATIONS AT THE TIME OF TRANSFER TO THE ICU
C3699344|T077|strict|75311-1|LNC|MEDS ON TRANSFER|MEDS ON TRANSFER
C3699344|T077|strict|10154-3|LNC|CHIEF COMPLAINT|CHIEF COMPLAINT
C3699344|T077|strict|10154-3|LNC|PATIENT STATES COMPLAINT|PATIENT STATES COMPLAINT
C3699344|T077|strict|10154-3|LNC|PATIENT COMPLAINT|PATIENT COMPLAINT
C3699344|T077|multi|10154-3|LNC|COMPLAINTS|COMPLAINTS
C3699344|T077|abbr|10154-3|LNC|CC|CC
C3699344|T077|strict|46239-0|LNC|REASON FOR VISIT AND CHIEF COMPLAINT|REASON FOR VISIT AND CHIEF COMPLAINT
C3699344|T077|strict|46239-0|LNC|REASON FOR VISIT/CHIEF COMPLAINT|REASON FOR VISIT/CHIEF COMPLAINT
C3699344|T077|strict|46239-0|LNC|CHIEF COMPLAINT AND REASON FOR VISIT|CHIEF COMPLAINT AND REASON FOR VISIT
C3699344|T077|strict|46239-0|LNC|CHIEF COMPLAINT REASON FOR VISIT|CHIEF COMPLAINT REASON FOR VISIT
C3699344|T077|strict|29299-5|LNC|REASON FOR VISIT|REASON FOR VISIT
C3699344|T077|strict|29299-5|LNC|REASON FOR CLINIC VISIT|REASON FOR CLINIC VISIT
C3699344|T077|strict|29299-5|LNC|REASON FOR ADMISSION|REASON FOR ADMISSION
C3699344|T077|strict|29299-5|LNC|HISTORY AND REASON FOR HOSPITALIZATION|HISTORY AND REASON FOR HOSPITALIZATION
C3699344|T077|strict|29299-5|LNC|REASON FOR HOSPITALIZATION|REASON FOR HOSPITALIZATION
C3699344|T077|strict|29299-5|LNC|HISTORY AND REASON FOR ADMISSION|HISTORY AND REASON FOR ADMISSION
C3699344|T077|strict|29299-5|LNC|HISTORY REASON FOR HOSPITALIZATION|HISTORY REASON FOR HOSPITALIZATION
C3699344|T077|strict|29299-5|LNC|REASON FOR EXAM|REASON FOR EXAM
C3699344|T077|strict|29299-5|LNC|REASON FOR THIS EXAMINATION|REASON FOR THIS EXAMINATION
C3699344|T077|strict|29299-5|LNC|NEW PROBLEMS|NEW PROBLEMS
C3699344|T077|strict|29299-5|LNC|INDICATIONS|INDICATIONS
C3699344|T077|strict|29299-5|LNC|INDICATION|INDICATION
C3699344|T077|strict|29299-5|LNC|INDICATION FOR SURGERY|INDICATION FOR SURGERY
C3699344|T077|strict|29299-5|LNC|INDICATIONS FOR INDUCTION|INDICATIONS FOR INDUCTION
C3699344|T077|strict|29299-5|LNC|INDICATIONS FOR OPERATION|INDICATIONS FOR OPERATION
C3699344|T077|strict|42349-1|LNC|REASON FOR REFERRAL|REASON FOR REFERRAL
C3699344|T077|strict|42349-1|LNC|REASON FOR CONSULT|REASON FOR CONSULT
C3699344|T077|strict|42349-1|LNC|REASON FOR CONSULTATION|REASON FOR CONSULTATION
C3699344|T077|strict|59768-2|LNC|PROCEDURE INDICATIONS INTERPRETATION|PROCEDURE INDICATIONS INTERPRETATION
C3699344|T077|strict|59768-2|LNC|PROCEDURE INDICATIONS|PROCEDURE INDICATIONS
C3699344|T077|strict|59768-2|LNC|PROCEDURE INDICATION|PROCEDURE INDICATION
C3699344|T077|strict|11450-4|LNC|PROBLEM LIST|PROBLEM LIST
C3699344|T077|strict|11450-4|LNC|ACTIVE PROBLEMS LIST|ACTIVE PROBLEMS LIST
C3699344|T077|strict|11450-4|LNC|ACTIVE PROBLEMS|ACTIVE PROBLEMS
C3699344|T077|strict|11450-4|LNC|PRINCIPAL PROBLEM|PRINCIPAL PROBLEM
C3699344|T077|strict|11450-4|LNC|PRINCIPAL DIAGNOSES|PRINCIPAL DIAGNOSES
C3699344|T077|strict|11450-4|LNC|PROBLEM LIST AND DIAGNOSIS|PROBLEM LIST AND DIAGNOSIS
C3699344|T077|strict|11450-4|LNC|PROBLEMS AND DIAGNOSIS|PROBLEMS AND DIAGNOSIS
C3699344|T077|strict|11450-4|LNC|LIST OF PROBLEM|LIST OF PROBLEM
C3699344|T077|strict|11450-4|LNC|LIST OF PROBLEMS|LIST OF PROBLEMS
C3699344|T077|strict|11450-4|LNC|LIST OF PROBLEMS DURING ADMISSION|LIST OF PROBLEMS DURING ADMISSION
C3699344|T077|strict|11450-4|LNC|LIST OF PROBLEMS DURING HOSPITALIZATION|LIST OF PROBLEMS DURING HOSPITALIZATION
C3699344|T077|strict|11450-4|LNC|BRIEF HOSPITAL COURSE|BRIEF HOSPITAL COURSE
C3699344|T077|strict|11450-4|LNC|EMERGENCY DEPARTMENT COURSE|EMERGENCY DEPARTMENT COURSE
C3699344|T077|strict|11450-4|LNC|HOSPITAL COURSE BY PROBLEM|HOSPITAL COURSE BY PROBLEM
C3699344|T077|strict|11450-4|LNC|HOSPITAL COURSE BY PROBLEMS|HOSPITAL COURSE BY PROBLEMS
C3699344|T077|strict|11450-4|LNC|HOSPITAL COURSE BY SYSTEM AND PROBLEM|HOSPITAL COURSE BY SYSTEM AND PROBLEM
C3699344|T077|strict|11450-4|LNC|SIGNIFICANT PROBLEMS|SIGNIFICANT PROBLEMS
C3699344|T077|strict|11450-4|LNC|SPONTANEOUS CONDITION|SPONTANEOUS CONDITION
C3699344|T077|strict|11450-4|LNC|OTHER SIGNIFICANT PROBLEMS|OTHER SIGNIFICANT PROBLEMS
C3699344|T077|strict|11450-4|LNC|PROBLEM CARDIOVASCULAR|PROBLEM CARDIOVASCULAR
C3699344|T077|multi|11450-4|LNC|SUMMARY OF HOSPITAL COURSE|SUMMARY OF HOSPITAL COURSE
C3699344|T077|strict|11450-4|LNC|COURSE BY PROBLEM|COURSE BY PROBLEM
C3699344|T077|strict|11450-4|LNC|MEDICAL PROBLEMS|MEDICAL PROBLEMS
C3699344|T077|strict|11450-4|LNC|OTHER PROBLEMS|OTHER PROBLEMS
C3699344|T077|strict|11450-4|LNC|OTHER ASSOCIATED PROBLEMS|OTHER ASSOCIATED PROBLEMS
C3699344|T077|strict|11450-4|LNC|PROBLEMS BY SYSTEMS|PROBLEMS BY SYSTEMS
C3699344|T077|strict|11450-4|LNC|UNDERLYING MEDICAL CONDITION|UNDERLYING MEDICAL CONDITION
C3699344|T077|strict|11450-4|LNC|RELATED DIAGNOSES|RELATED DIAGNOSES
C3699344|T077|strict|11450-4|LNC|SYMPTOMS|SYMPTOMS
C3699344|T077|relax|11450-4|LNC|CONDITIONS|CONDITIONS
C3699344|T077|relax|11450-4|LNC|PROBLEMS|PROBLEMS
C3699344|T077|relax|11450-4|LNC|PROBLEM|PROBLEM
C3699344|T077|strict|61133-5|LNC|CLINICAL IMPRESSION|CLINICAL IMPRESSION
C3699344|T077|strict|61133-5|LNC|IMPRESSION|IMPRESSION
C3699344|T077|strict|61133-5|LNC|IMPRESSION ON ADMISSION|IMPRESSION ON ADMISSION
C3699344|T077|strict|61133-5|LNC|PRIMARY PROBLEM INTERPRETATION|PRIMARY PROBLEM INTERPRETATION
C3699344|T077|multi|61133-5|LNC|DIAGNOSTIC IMPRESSION|DIAGNOSTIC IMPRESSION
C3699344|T077|strict|51898-5|LNC|RISK FACTORS|RISK FACTORS
C3699344|T077|strict|51898-5|LNC|CARDIAC RISK FACTORS|CARDIAC RISK FACTORS
C3699344|T077|strict|51898-5|LNC|CORONARY RISK FACTORS|CORONARY RISK FACTORS
C3699344|T077|strict|51898-5|LNC|HYPERTENSIVE URGENCY|HYPERTENSIVE URGENCY
C3699344|T077|strict|51898-5|LNC|HYPERGLYCEMIC SYMPTOMS|HYPERGLYCEMIC SYMPTOMS
C3699344|T077|strict|10157-6|LNC|HISTORY OF FAMILY MEMBER DISEASES|HISTORY OF FAMILY MEMBER DISEASES
C3699344|T077|strict|10157-6|LNC|FAMILY HISTORY|FAMILY HISTORY
C3699344|T077|relax|10157-6|LNC|FATHER|FATHER
C3699344|T077|relax|10157-6|LNC|MOTHER|MOTHER
C3699344|T077|relax|10157-6|LNC|SIBLINGS|SIBLINGS
C3699344|T077|relax|10157-6|LNC|SPOUSE|SPOUSE
C3699344|T077|relax|10157-6|LNC|OFFSPRING|OFFSPRING
C3699344|T077|abbr|10157-6|LNC|FHX|FHX
C3699344|T077|strict|10164-2|LNC|HISTORY OF PRESENT ILLNESS|HISTORY OF PRESENT ILLNESS
C3699344|T077|strict|10164-2|LNC|HISTORY PRESENT ILLNESS|HISTORY PRESENT ILLNESS
C3699344|T077|strict|10164-2|LNC|BRIEF HISTORY OF PHYSICAL ILLNESS|BRIEF HISTORY OF PHYSICAL ILLNESS
C3699344|T077|strict|10164-2|LNC|BRIEF ADMISSION HISTORY OF PRESENT ILLNESS|BRIEF ADMISSION HISTORY OF PRESENT ILLNESS
C3699344|T077|strict|10164-2|LNC|BRIEF HISTORY OF PRESENT ILLNESS|BRIEF HISTORY OF PRESENT ILLNESS
C3699344|T077|strict|10164-2|LNC|HX OF PRES ILLNESS|HX OF PRES ILLNESS
C3699344|T077|strict|10164-2|LNC|HX OF PRESENT ILLNESS|HX OF PRESENT ILLNESS
C3699344|T077|strict|10164-2|LNC|HISTORY OF PRESENT ILLNESS AND HOSPITAL COURSE|HISTORY OF PRESENT ILLNESS AND HOSPITAL COURSE
C3699344|T077|strict|10164-2|LNC|HISTORY OF PRESENT ILLNESS AND REASON FOR HOSPITALIZATION|HISTORY OF PRESENT ILLNESS AND REASON FOR HOSPITALIZATION
C3699344|T077|strict|10164-2|LNC|HISTORY OF PRESENTING ILLNESS|HISTORY OF PRESENTING ILLNESS
C3699344|T077|strict|10164-2|LNC|HISTORY OF THE PRESENT ILLNESS|HISTORY OF THE PRESENT ILLNESS
C3699344|T077|strict|10164-2|LNC|HISTORY AND PHYSICAL HISTORY OF PRESENT ILLNESS|HISTORY AND PHYSICAL HISTORY OF PRESENT ILLNESS
C3699344|T077|multi|10164-2|LNC|HISTORY AND PHYSICAL|HISTORY AND PHYSICAL
C3699344|T077|strict|10164-2|LNC|H&P BY|H&P BY
C3699344|T077|abbr|10164-2|LNC|H&P|H&P
C3699344|T077|relax|10164-2|LNC|PRESENT ILLNESS|PRESENT ILLNESS
C3699344|T077|abbr|10164-2|LNC|HPI|HPI
C3699344|T077|relax|61150-9|LNC|SUBJECTIVE|SUBJECTIVE
C3699344|T077|multi|61150-9|LNC|SUBJECTIVE DATA|SUBJECTIVE DATA
C3699344|T077|strict|10184-0|LNC|HOSPITAL DISCHARGE PHYSICAL FINDINGS|HOSPITAL DISCHARGE PHYSICAL FINDINGS
C3699344|T077|strict|59776-5|LNC|PROCEDURE FINDINGS|PROCEDURE FINDINGS
C3699344|T077|strict|18834-2|LNC|RADIOLOGY COMPARISON STUDY OBSERVATION|RADIOLOGY COMPARISON STUDY OBSERVATION
C3699344|T077|relax|18834-2|LNC|COMPARISON|COMPARISON
C3699344|T077|multi|51848-0|LNC|EVALUATION NOTE|EVALUATION NOTE
C3699344|T077|multi|51848-0|LNC|EVAL NOTE|EVAL NOTE
C3699344|T077|multi|51848-0|LNC|ASSESSMENT/PLAN|ASSESSMENT/PLAN
C3699344|T077|relax|51848-0|LNC|EVALUATION|EVALUATION
C3699344|T077|relax|51848-0|LNC|ASSESSMENT|ASSESSMENT
C3699344|T077|relax|51848-0|LNC|ASSESSMENTS|ASSESSMENTS
C3699344|T077|multi|55108-5|LNC|CLINICAL PRESENTATIONS|CLINICAL PRESENTATIONS
C3699344|T077|multi|55108-5|LNC|CLINICAL PRESENTATION|CLINICAL PRESENTATION
C3699344|T077|strict|55109-3|LNC|COMPLICATIONS DOCUMENT|COMPLICATIONS DOCUMENT
C3699344|T077|relax|55109-3|LNC|COMPLICATIONS|COMPLICATIONS
C3699344|T077|multi|55109-3|LNC|CONCERNS|CONCERNS
C3699344|T077|multi|11329-0|LNC|MEDICAL GENERAL HISTORY|MEDICAL GENERAL HISTORY
C3699344|T077|multi|11329-0|LNC|GENERAL HISTORY|GENERAL HISTORY
C3699344|T077|multi|11329-0|LNC|HISTORY GENERAL|HISTORY GENERAL
C3699344|T077|strict|11329-0|LNC|BRIEF HISTORY|BRIEF HISTORY
C3699344|T077|strict|42347-5|LNC|ADMISSION DIAGNOSIS|ADMISSION DIAGNOSIS
C3699344|T077|strict|42347-5|LNC|ADDITIONAL ADMITTING DIAGNOSIS|ADDITIONAL ADMITTING DIAGNOSIS
C3699344|T077|strict|42347-5|LNC|ADMISSION DIAGNOSES|ADMISSION DIAGNOSES
C3699344|T077|strict|42347-5|LNC|ADMIT DIAGNOSES|ADMIT DIAGNOSES
C3699344|T077|strict|42347-5|LNC|ADMIT DIAGNOSIS|ADMIT DIAGNOSIS
C3699344|T077|strict|42347-5|LNC|ADMITTING DIAGNOSES|ADMITTING DIAGNOSES
C3699344|T077|strict|42347-5|LNC|ADMITTING DIAGNOSIS|ADMITTING DIAGNOSIS
C3699344|T077|strict|42347-5|LNC|LIST OF DIAGNOSIS DURING ADMISSION|LIST OF DIAGNOSIS DURING ADMISSION
C3699344|T077|strict|42347-5|LNC|PRINCIPAL ADMISSION DIAGNOSIS|PRINCIPAL ADMISSION DIAGNOSIS
C3699344|T077|strict|42347-5|LNC|PRINCIPAL DIAGNOSIS FOR ADMISSION|PRINCIPAL DIAGNOSIS FOR ADMISSION
C3699344|T077|strict|42347-5|LNC|PRINCIPAL DIAGNOSIS ON ADMISSION|PRINCIPAL DIAGNOSIS ON ADMISSION
C3699344|T077|strict|42347-5|LNC|PRIMARY ADMISSION DIAGNOSIS|PRIMARY ADMISSION DIAGNOSIS
C3699344|T077|strict|42347-5|LNC|PRIMARY ADMITTING DIAGNOSIS|PRIMARY ADMITTING DIAGNOSIS
C3699344|T077|strict|42347-5|LNC|PRIMARY DIAGNOSIS DURING THIS ADMISSION|PRIMARY DIAGNOSIS DURING THIS ADMISSION
C3699344|T077|strict|42347-5|LNC|PRIMARY DIAGNOSIS ON ADMISSION|PRIMARY DIAGNOSIS ON ADMISSION
C3699344|T077|strict|42347-5|LNC|PRINCIPLE ADMISSION DIAGNOSIS|PRINCIPLE ADMISSION DIAGNOSIS
C3699344|T077|strict|42347-5|LNC|PRINCIPLE DISCHARGE DIAGNOSIS|PRINCIPLE DISCHARGE DIAGNOSIS
C3699344|T077|strict|42347-5|LNC|PRINCIPAL DIAGNOSIS|PRINCIPAL DIAGNOSIS
C3699344|T077|strict|42347-5|LNC|PRINCIPLE DIAGNOSIS|PRINCIPLE DIAGNOSIS
C3699344|T077|strict|42347-5|LNC|PRIMARY DIAGNOSIS|PRIMARY DIAGNOSIS
C3699344|T077|strict|42347-5|LNC|PRIMARY DIAGNOSES|PRIMARY DIAGNOSES
C3699344|T077|relax|42347-5|LNC|CURRENT DIAGNOSIS|CURRENT DIAGNOSIS
C3699344|T077|relax|42347-5|LNC|PRIMARY DX|PRIMARY DX
C3699344|T077|relax|42347-5|LNC|PRIMARY MEDICAL DIAGNOSIS|PRIMARY MEDICAL DIAGNOSIS
C3699344|T077|strict|78375-3|LNC|DISCHARGE DIAGNOSIS|DISCHARGE DIAGNOSIS
C3699344|T077|strict|78375-3|LNC|DISCHARGE DIAGNOSES|DISCHARGE DIAGNOSES
C3699344|T077|strict|78375-3|LNC|DIAGNOSIS AT DISCHARGE|DIAGNOSIS AT DISCHARGE
C3699344|T077|strict|78375-3|LNC|CONDITION AT DISCHARGE|CONDITION AT DISCHARGE
C3699344|T077|strict|78375-3|LNC|ASSOCIATE DISCHARGE DIAGNOSIS|ASSOCIATE DISCHARGE DIAGNOSIS
C3699344|T077|strict|78375-3|LNC|PRINCIPAL DIAGNOSIS ON DISCHARGE|PRINCIPAL DIAGNOSIS ON DISCHARGE
C3699344|T077|strict|78375-3|LNC|PRINCIPAL DIAGNOSIS ON THIS PATIENT|PRINCIPAL DIAGNOSIS ON THIS PATIENT
C3699344|T077|strict|78375-3|LNC|PRIMARY DISCHARGE DIAGNOSIS|PRIMARY DISCHARGE DIAGNOSIS
C3699344|T077|strict|78375-3|LNC|PRINCIPAL DISCHARGE DIAGNOSIS|PRINCIPAL DISCHARGE DIAGNOSIS
C3699344|T077|strict|78375-3|LNC|PRINCIPAL DISCHARGE DIAGNOSES|PRINCIPAL DISCHARGE DIAGNOSES
C3699344|T077|strict|78375-3|LNC|PRELIMINARY DIAGNOSIS|PRELIMINARY DIAGNOSIS
C3699344|T077|strict|78375-3|LNC|PROBLEMS AND DIAGNOSIS|PROBLEMS AND DIAGNOSIS
C3699344|T077|strict|78375-3|LNC|ASSOCIATED DISCHARGE DIAGNOSES|ASSOCIATED DISCHARGE DIAGNOSES
C3699344|T077|strict|78375-3|LNC|OTHER DIAGNOSES ON DISCHARGE|OTHER DIAGNOSES ON DISCHARGE
C3699344|T077|strict|78375-3|LNC|OTHER DIAGNOSIS AT DISCHARGE|OTHER DIAGNOSIS AT DISCHARGE
C3699344|T077|strict|78375-3|LNC|OTHER DISCHARGE DIAGNOSES|OTHER DISCHARGE DIAGNOSES
C3699344|T077|strict|78375-3|LNC|OTHER MEDICAL DIAGNOSIS|OTHER MEDICAL DIAGNOSIS
C3699344|T077|strict|78375-3|LNC|SECONDARY DISCHARGE DIAGNOSES|SECONDARY DISCHARGE DIAGNOSES
C3699344|T077|strict|78375-3|LNC|OTHER DIAGNOSES AND CONDITIONS AFFECTING TREATMENT OR STAY|OTHER DIAGNOSES AND CONDITIONS AFFECTING TREATMENT OR STAY
C3699344|T077|relax|78375-3|LNC|CONDITION|CONDITION
C3699344|T077|relax|78375-3|LNC|DIAGNOSIS|DIAGNOSIS
C3699344|T077|relax|78375-3|LNC|SECONDARY DIAGNOSIS|SECONDARY DIAGNOSIS
C3699344|T077|relax|78375-3|LNC|SECONDARY DIAGNOSES|SECONDARY DIAGNOSES
C3699344|T077|strict|46241-6|LNC|HOSPITAL ADMISSION DIAGNOSIS|HOSPITAL ADMISSION DIAGNOSIS
C3699344|T077|strict|46241-6|LNC|HOSPITAL ADMISSION DX|HOSPITAL ADMISSION DX
C3699344|T077|strict|11535-2|LNC|HOSPITAL DISCHARGE DX|HOSPITAL DISCHARGE DX
C3699344|T077|strict|11535-2|LNC|HOSPITAL DISCHARGE DIAGNOSIS|HOSPITAL DISCHARGE DIAGNOSIS
C3699344|T077|strict|54531-9|LNC|ACTIVE DISEASE DIAGNOSIS|ACTIVE DISEASE DIAGNOSIS
C3699344|T077|strict|54531-9|LNC|ACTIVE DISEASE DIAGNOSES|ACTIVE DISEASE DIAGNOSES
C3699344|T077|strict|54531-9|LNC|ACTIVE DIAGNOSES|ACTIVE DIAGNOSES
C3699344|T077|strict|54531-9|LNC|ACUTE DIAGNOSES|ACUTE DIAGNOSES
C3699344|T077|strict|54531-9|LNC|CHRONIC DIAGNOSES|CHRONIC DIAGNOSES
C3699344|T077|relax|54531-9|LNC|CLINICAL DIAGNOSIS|CLINICAL DIAGNOSIS
C3699344|T077|relax|54531-9|LNC|ACTIVE DIAGNOSIS|ACTIVE DIAGNOSIS
C3699344|T077|strict|54545-9|LNC|DIAGNOSIS LIST|DIAGNOSIS LIST
C3699344|T077|strict|54545-9|LNC|DIAGNOSES LIST|DIAGNOSES LIST
C3699344|T077|strict|54545-9|LNC|LIST OF DIAGNOSES|LIST OF DIAGNOSES
C3699344|T077|strict|54545-9|LNC|LIST OF OTHER DIAGNOSES|LIST OF OTHER DIAGNOSES
C3699344|T077|strict|54545-9|LNC|LIST OF OTHER PROBLEMS AND DIAGNOSES|LIST OF OTHER PROBLEMS AND DIAGNOSES
C3699344|T077|strict|54545-9|LNC|LIST OF PROBLEMS AND DIAGNOSES|LIST OF PROBLEMS AND DIAGNOSES
C3699344|T077|strict|54545-9|LNC|LIST OF PROBLEMS AND OTHER DIAGNOSES|LIST OF PROBLEMS AND OTHER DIAGNOSES
C3699344|T077|strict|54545-9|LNC|LISTS OF PROBLEMS AND DIAGNOSES|LISTS OF PROBLEMS AND DIAGNOSES
C3699344|T077|strict|54545-9|LNC|OTHER SIGNIFICANT DIAGNOSES|OTHER SIGNIFICANT DIAGNOSES
C3699344|T077|relax|54545-9|LNC|OTHER MEDICAL DIAGNOSIS|OTHER MEDICAL DIAGNOSIS
C3699344|T077|relax|54545-9|LNC|OTHER MEDICAL DIAGNOSES|OTHER MEDICAL DIAGNOSES
C3699344|T077|relax|54545-9|LNC|OTHER PROBLEMS AND DIAGNOSES|OTHER PROBLEMS AND DIAGNOSES
C3699344|T077|relax|54545-9|LNC|OTHER PROBLEMS AND DIAGNOSIS|OTHER PROBLEMS AND DIAGNOSIS
C3699344|T077|relax|54545-9|LNC|OTHER DIAGNOSES|OTHER DIAGNOSES
C3699344|T077|relax|54545-9|LNC|OTHER DIAGNOSIS|OTHER DIAGNOSIS
C3699344|T077|relax|54545-9|LNC|ADDITIONAL DIAGNOSES|ADDITIONAL DIAGNOSES
C3699344|T077|relax|54545-9|LNC|ADDITIONAL DIAGNOSIS|ADDITIONAL DIAGNOSIS
C3699344|T077|relax|54545-9|LNC|ASSOCIATED DIAGNOSES|ASSOCIATED DIAGNOSES
C3699344|T077|relax|54545-9|LNC|ASSOCIATED DIAGNOSIS|ASSOCIATED DIAGNOSIS
C3699344|T077|relax|54545-9|LNC|DIAGNOSES|DIAGNOSES
C3699344|T077|relax|54545-9|LNC|DISEASES|DISEASES
C3699344|T077|relax|54545-9|LNC|ADDITIONAL DIAGNOSES INCLUDE|ADDITIONAL DIAGNOSES INCLUDE
C3699344|T077|multi|51847-2|LNC|EVALUATION AND PLAN|EVALUATION AND PLAN
C3699344|T077|multi|51847-2|LNC|ASSESSMENT AND PLAN|ASSESSMENT AND PLAN
C3699344|T077|strict|55110-1|LNC|CONCLUSIONS INTERPRETATION|CONCLUSIONS INTERPRETATION
C3699344|T077|multi|55110-1|LNC|CONCLUSION|CONCLUSION
C3699344|T077|multi|55110-1|LNC|CONCLUSIONS|CONCLUSIONS
C3699344|T077|strict|11348-0|LNC|PAST MEDICAL HISTORY|PAST MEDICAL HISTORY
C3699344|T077|strict|11348-0|LNC|PERSONAL HISTORY|PERSONAL HISTORY
C3699344|T077|strict|11348-0|LNC|HISTORY OF PAST ILLNESS|HISTORY OF PAST ILLNESS
C3699344|T077|strict|11348-0|LNC|PAST GYN HISTORY|PAST GYN HISTORY
C3699344|T077|strict|11348-0|LNC|PAST GYNECOLOGIC HISTORY|PAST GYNECOLOGIC HISTORY
C3699344|T077|strict|11348-0|LNC|PAST PSYCHIATRIC HISTORY|PAST PSYCHIATRIC HISTORY
C3699344|T077|strict|11348-0|LNC|CLINICAL HISTORY|CLINICAL HISTORY
C3699344|T077|multi|11348-0|LNC|PSYCHIATRIC|PSYCHIATRIC
C3699344|T077|abbr|11348-0|LNC|PMH|PMH
C3699344|T077|abbr|11348-0|LNC|PMHX|PMHX
C3699344|T077|strict|10219-4|LNC|SURGICAL OPERATION NOTE PREOPERATIVE DX|SURGICAL OPERATION NOTE PREOPERATIVE DX
C3699344|T077|strict|10219-4|LNC|PREOPERATIVE DX|PREOPERATIVE DX
C3699344|T077|strict|10219-4|LNC|OPERATIVE NOTE PRE-OP DX|OPERATIVE NOTE PRE-OP DX
C3699344|T077|strict|10219-4|LNC|PREOPERATIVE DIAGNOSES|PREOPERATIVE DIAGNOSES
C3699344|T077|relax|10219-4|LNC|PREOPERATIVE DIAGNOSIS|PREOPERATIVE DIAGNOSIS
C3699344|T077|strict|10218-6|LNC|SURGICAL OPERATION NOTE POSTOPERATIVE DIAGNOSIS|SURGICAL OPERATION NOTE POSTOPERATIVE DIAGNOSIS
C3699344|T077|strict|10218-6|LNC|POSTOPERATIVE DIAGNOSES|POSTOPERATIVE DIAGNOSES
C3699344|T077|strict|10218-6|LNC|POSTOPERATIVE DIAGNOSIS|POSTOPERATIVE DIAGNOSIS
C3699344|T077|multi|59769-0|LNC|POSTPROCEDURE DIAGNOSIS|POSTPROCEDURE DIAGNOSIS
C3699344|T077|multi|18785-6|LNC|RADIOLOGY REASON FOR STUDY|RADIOLOGY REASON FOR STUDY
C3699344|T077|multi|19005-8|LNC|RADIOLOGY IMAGING STUDY IMPRESSION|RADIOLOGY IMAGING STUDY IMPRESSION
C3699344|T077|multi|18782-3|LNC|RADIOLOGY STUDY OBSERVATION FINDINGS|RADIOLOGY STUDY OBSERVATION FINDINGS
C3699344|T077|multi|18783-1|LNC|RADIOLOGY STUDY RECOMMENDATION|RADIOLOGY STUDY RECOMMENDATION
C3699344|T077|strict|22029-3|LNC|PHYSICAL EXAM|PHYSICAL EXAM
C3699344|T077|strict|22029-3|LNC|HEAD EYES EARS NOSE THROAT|HEAD EYES EARS NOSE THROAT
C3699344|T077|strict|22029-3|LNC|ADMISSION PHYSICAL EXAMINATION|ADMISSION PHYSICAL EXAMINATION
C3699344|T077|strict|22029-3|LNC|HOSPITAL DISCHARGE PHYSICAL|HOSPITAL DISCHARGE PHYSICAL
C3699344|T077|strict|22029-3|LNC|PHYSICAL EXAM ON ADMISSION|PHYSICAL EXAM ON ADMISSION
C3699344|T077|strict|22029-3|LNC|PHYSICAL EXAMINATION|PHYSICAL EXAMINATION
C3699344|T077|strict|22029-3|LNC|PHYSICAL EXAMINATION ON ADMISSION|PHYSICAL EXAMINATION ON ADMISSION
C3699344|T077|strict|22029-3|LNC|PHYSICAL EXAMINATION ON DISCHARGE|PHYSICAL EXAMINATION ON DISCHARGE
C3699344|T077|strict|22029-3|LNC|PHYSICAL EXAMINATION ON PRESENTATION|PHYSICAL EXAMINATION ON PRESENTATION
C3699344|T077|strict|22029-3|LNC|PHYSICAL EXAMINATION UPON ADMISSION|PHYSICAL EXAMINATION UPON ADMISSION
C3699344|T077|strict|10210-3|LNC|PHYSICAL FINDINGS OF GENERAL STATUS|PHYSICAL FINDINGS OF GENERAL STATUS
C3699344|T077|multi|10210-3|LNC|GENERAL STATUS|GENERAL STATUS
C3699344|T077|strict|8716-3|LNC|VITAL SIGNS|VITAL SIGNS
C3699344|T077|strict|8716-3|LNC|Filed Vitals|Filed Vitals
C3699344|T077|strict|8716-3|LNC|VITALS ON ADMISSION|VITALS ON ADMISSION
C3699344|T077|abbr|8716-3|LNC|VS|VS
C3699344|T077|relax|8716-3|LNC|VITALS|VITALS
C3699344|T077|relax|8716-3|LNC|WEIGHT|WEIGHT
C3699344|T077|relax|8716-3|LNC|BLOOD PRESSURE|BLOOD PRESSURE
C3699344|T077|strict|10187-3|LNC|REVIEW OF SYSTEMS|REVIEW OF SYSTEMS
C3699344|T077|abbr|10187-3|LNC|ROS|ROS
C3699344|T077|strict|10190-7|LNC|MENTAL STATUS|MENTAL STATUS
C3699344|T077|strict|29545-1|LNC|PHYSICAL FINDINGS|PHYSICAL FINDINGS
C3699344|T077|relax|29545-1|LNC|PHYS FIND|PHYS FIND
C3699344|HeaderTUI.T082|body|11384-5|LNC|ABDOMEN|ABDOMEN
C3699344|HeaderTUI.T082|body|11384-5|LNC|ABD|ABD
C3699344|HeaderTUI.T082|body|11384-5|LNC|ADNEXA|ADNEXA
C3699344|HeaderTUI.T082|body|11384-5|LNC|APPEARANCE|APPEARANCE
C3699344|HeaderTUI.T082|body|11384-5|LNC|BACK|BACK
C3699344|HeaderTUI.T082|body|11384-5|LNC|BMI|BMI
C3699344|HeaderTUI.T082|body|11384-5|LNC|BREASTS|BREASTS
C3699344|HeaderTUI.T082|body|11384-5|LNC|CARDIAC|CARDIAC
C3699344|HeaderTUI.T082|body|11384-5|LNC|CARDIAC EXAMINATION|CARDIAC EXAMINATION
C3699344|HeaderTUI.T082|body|11384-5|LNC|CARDIOVASCULAR|CARDIOVASCULAR
C3699344|HeaderTUI.T082|body|11384-5|LNC|CARDIOVASCULAR EXAM|CARDIOVASCULAR EXAM
C3699344|HeaderTUI.T082|body|11384-5|LNC|CARDIOVASCULAR STATUS|CARDIOVASCULAR STATUS
C3699344|HeaderTUI.T082|body|11384-5|LNC|CARDS|CARDS
C3699344|HeaderTUI.T082|body|11384-5|LNC|CAROTIDS|CAROTIDS
C3699344|HeaderTUI.T082|body|11384-5|LNC|CEREBELLAR EXAM|CEREBELLAR EXAM
C3699344|HeaderTUI.T082|body|11384-5|LNC|CHEST|CHEST
C3699344|HeaderTUI.T082|body|11384-5|LNC|COORDINATION|COORDINATION
C3699344|HeaderTUI.T082|body|11384-5|LNC|COR|COR
C3699344|HeaderTUI.T082|body|11384-5|LNC|CRANIAL|CRANIAL
C3699344|HeaderTUI.T082|body|11384-5|LNC|CRANIAL NERVES|CRANIAL NERVES
C3699344|HeaderTUI.T082|body|11384-5|LNC|CVS|CVS
C3699344|HeaderTUI.T082|body|11384-5|LNC|EAR/NOSE/THROAT|EAR/NOSE/THROAT
C3699344|HeaderTUI.T082|body|11384-5|LNC|ENDO|ENDO
C3699344|HeaderTUI.T082|body|11384-5|LNC|ENDOCRINE|ENDOCRINE
C3699344|HeaderTUI.T082|body|11384-5|LNC|EXAM|EXAM
C3699344|HeaderTUI.T082|body|11384-5|LNC|EXAMINATION|EXAMINATION
C3699344|HeaderTUI.T082|body|11384-5|LNC|EXTREMITIES|EXTREMITIES
C3699344|HeaderTUI.T082|body|11384-5|LNC|EXTREMITY EXAM|EXTREMITY EXAM
C3699344|HeaderTUI.T082|body|11384-5|LNC|EYE EXAM|EYE EXAM
C3699344|HeaderTUI.T082|body|11384-5|LNC|EYES|EYES
C3699344|HeaderTUI.T082|body|11384-5|LNC|FOOT EXAM|FOOT EXAM
C3699344|HeaderTUI.T082|body|11384-5|LNC|FUNCTIONAL AND COGNITIVE STATUS|FUNCTIONAL AND COGNITIVE STATUS
C3699344|HeaderTUI.T082|body|11384-5|LNC|GAIT|GAIT
C3699344|HeaderTUI.T082|body|11384-5|LNC|GASTROINTESTINAL|GASTROINTESTINAL
C3699344|HeaderTUI.T082|body|11384-5|LNC|GEN|GEN
C3699344|HeaderTUI.T082|body|11384-5|LNC|GENERAL|GENERAL
C3699344|HeaderTUI.T082|body|11384-5|LNC|GENITOURINARY|GENITOURINARY
C3699344|HeaderTUI.T082|body|11384-5|LNC|GI|GI
C3699344|HeaderTUI.T082|body|11384-5|LNC|GU|GU
C3699344|HeaderTUI.T082|body|11384-5|LNC|HEAD EYES EARS NOSE AND THROAT|HEAD EYES EARS NOSE AND THROAT
C3699344|HeaderTUI.T082|body|11384-5|LNC|HEAD EYES EARS NOSE AND THROAT EXAM|HEAD EYES EARS NOSE AND THROAT EXAM
C3699344|HeaderTUI.T082|body|11384-5|LNC|HEART|HEART
C3699344|HeaderTUI.T082|body|11384-5|LNC|HEENT|HEENT
C3699344|HeaderTUI.T082|body|11384-5|LNC|HEMODYNAMICS|HEMODYNAMICS
C3699344|HeaderTUI.T082|body|11384-5|LNC|INITIAL NEWBORN EXAM|INITIAL NEWBORN EXAM
C3699344|HeaderTUI.T082|body|11384-5|LNC|LUNGS|LUNGS
C3699344|HeaderTUI.T082|body|11384-5|LNC|MENTAL STATUS EXAMINATION|MENTAL STATUS EXAMINATION
C3699344|HeaderTUI.T082|body|11384-5|LNC|MUSCULOSKELETAL|MUSCULOSKELETAL
C3699344|HeaderTUI.T082|body|11384-5|LNC|NECK|NECK
C3699344|HeaderTUI.T082|body|11384-5|LNC|NEURO|NEURO
C3699344|HeaderTUI.T082|body|11384-5|LNC|NEUROLOGIC|NEUROLOGIC
C3699344|HeaderTUI.T082|body|11384-5|LNC|NEUROLOGIC EXAM|NEUROLOGIC EXAM
C3699344|HeaderTUI.T082|body|11384-5|LNC|NEUROLOGICAL|NEUROLOGICAL
C3699344|HeaderTUI.T082|body|11384-5|LNC|NEUROLOGICAL EXAMINATION|NEUROLOGICAL EXAMINATION
C3699344|HeaderTUI.T082|body|11384-5|LNC|NEUROLOGY|NEUROLOGY
C3699344|HeaderTUI.T082|body|11384-5|LNC|NODES|NODES
C3699344|HeaderTUI.T082|body|11384-5|LNC|OPHTHALMOLOGY|OPHTHALMOLOGY
C3699344|HeaderTUI.T082|body|11384-5|LNC|PE|PE
C3699344|HeaderTUI.T082|body|11384-5|LNC|PELVIC|PELVIC
C3699344|HeaderTUI.T082|body|11384-5|LNC|PSYCH|PSYCH
C3699344|HeaderTUI.T082|body|11384-5|LNC|PSYCHOSOCIAL|PSYCHOSOCIAL
C3699344|HeaderTUI.T082|body|11384-5|LNC|PULM|PULM
C3699344|HeaderTUI.T082|body|11384-5|LNC|PULMONARY|PULMONARY
C3699344|HeaderTUI.T082|body|11384-5|LNC|PULSE|PULSE
C3699344|HeaderTUI.T082|body|11384-5|LNC|PULSES|PULSES
C3699344|HeaderTUI.T082|body|11384-5|LNC|PUPILS|PUPILS
C3699344|HeaderTUI.T082|body|11384-5|LNC|RECTAL|RECTAL
C3699344|HeaderTUI.T082|body|11384-5|LNC|REFLEXES|REFLEXES
C3699344|HeaderTUI.T082|body|11384-5|LNC|RENAL|RENAL
C3699344|HeaderTUI.T082|body|11384-5|LNC|RESP|RESP
C3699344|HeaderTUI.T082|body|11384-5|LNC|RESPIRATORY|RESPIRATORY
C3699344|HeaderTUI.T082|body|11384-5|LNC|SENSORY|SENSORY
C3699344|HeaderTUI.T082|body|11384-5|LNC|SENSORY EXAMINATION|SENSORY EXAMINATION
C3699344|HeaderTUI.T082|body|11384-5|LNC|SKIN|SKIN
C3699344|HeaderTUI.T082|body|11384-5|LNC|SPINE|SPINE
C3699344|T077|strict|46062-6|LNC|CURRENT TREATMENT|CURRENT TREATMENT
C3699344|T077|strict|46062-6|LNC|TRANSFUSION SERVICES|TRANSFUSION SERVICES
C3699344|T077|relax|46062-6|LNC|CHEMOTHERAPY|CHEMOTHERAPY
C3699344|T077|relax|46062-6|LNC|DIALYSIS|DIALYSIS
C3699344|T077|relax|46062-6|LNC|IV MEDICATION|IV MEDICATION
C3699344|T077|relax|46062-6|LNC|OSTOMY|OSTOMY
C3699344|T077|relax|46062-6|LNC|OXYGEN THERAPY|OXYGEN THERAPY
C3699344|T077|relax|46062-6|LNC|RADIATION|RADIATION
C3699344|T077|relax|46062-6|LNC|SUCTIONING|SUCTIONING
C3699344|T077|relax|46062-6|LNC|TRACHEOSTOMY|TRACHEOSTOMY
C3699344|T077|relax|46062-6|LNC|TRANSFUSIONS|TRANSFUSIONS
C3699344|T077|relax|46062-6|LNC|VENTILATOR|VENTILATOR
C3699344|T077|relax|46062-6|LNC|RESPIRATOR|RESPIRATOR
C3699344|T077|relax|46062-6|LNC|TREATMENTS|TREATMENTS
C3699344|T077|strict|8648-8|LNC|HOSPITAL COURSE|HOSPITAL COURSE
C3699344|T077|strict|8648-8|LNC|HOSPITAL COURSE BY SYSTEM|HOSPITAL COURSE BY SYSTEM
C3699344|T077|strict|8648-8|LNC|HOSPITAL COURSE BY SYSTEMS|HOSPITAL COURSE BY SYSTEMS
C3699344|T077|strict|8648-8|LNC|HOSPITAL COURSE AND TREATMENT|HOSPITAL COURSE AND TREATMENT
C3699344|T077|strict|8653-8|LNC|HOSPITAL DISCHARGE INSTRUCTIONS|HOSPITAL DISCHARGE INSTRUCTIONS
C3699344|T077|strict|8653-8|LNC|HOSPITAL DISCHARGE INSTRUCTIONS GIVEN BY|HOSPITAL DISCHARGE INSTRUCTIONS GIVEN BY
C3699344|T077|strict|8653-8|LNC|CARE PLAN|CARE PLAN
C3699344|T077|strict|8653-8|LNC|CARE RECOMMENDATIONS|CARE RECOMMENDATIONS
C3699344|T077|strict|8653-8|LNC|CARE AND RECOMMENDATIONS|CARE AND RECOMMENDATIONS
C3699344|T077|strict|8653-8|LNC|CARE AND RECOMMENDATIONS AT THE TIME OF DISCHARGE|CARE AND RECOMMENDATIONS AT THE TIME OF DISCHARGE
C3699344|T077|relax|69730-0|LNC|INSTRUCTIONS|INSTRUCTIONS
C3699344|T077|relax|69730-0|LNC|PLAN|PLAN
C3699344|T077|relax|62387-6|LNC|INTERVENTIONS|INTERVENTIONS
C3699344|T077|strict|62387-6|LNC|INTERVENTIONS PROVIDED|INTERVENTIONS PROVIDED
C3699344|T077|strict|18776-5|LNC|PLAN OF CARE NOTE|PLAN OF CARE NOTE
C3699344|T077|strict|79191-3|LNC|PATIENT DEMOGRAPHICS PANEL|PATIENT DEMOGRAPHICS PANEL
C3699344|T077|strict|79191-3|LNC|PATIENT DEMOGRAPHICS|PATIENT DEMOGRAPHICS
C3699344|T077|strict|79191-3|LNC|DEMOGRAPHICS|DEMOGRAPHICS
C3699344|T077|strict|79191-3|LNC|PATIENT INFORMATION|PATIENT INFORMATION
C3699344|T077|strict|79191-3|LNC|PATIENT INFO|PATIENT INFO
C3699344|T077|relax|79191-3|LNC|PATIENT|PATIENT
C3699344|T077|strict|45392-8|LNC|FIRST NAME|FIRST NAME
C3699344|T077|strict|45392-8|LNC|GIVEN NAME|GIVEN NAME
C3699344|T077|strict|45394-4|LNC|LAST NAME|LAST NAME
C3699344|T077|strict|45394-4|LNC|FAMILY NAME|FAMILY NAME
C3699344|T077|strict|87226-7|LNC|PATIENT NAME|PATIENT NAME
C3699344|T077|strict|87226-7|LNC|LEGAL NAME|LEGAL NAME
C3699344|T077|strict|87226-7|LNC|FULL NAME|FULL NAME
C3699344|T077|relax|87226-7|LNC|NICK NAME|NICK NAME
C3699344|T077|strict|87226-7|LNC|SUBSCRIBER|SUBSCRIBER
C3699344|T077|strict|87226-7|LNC|SUBSCRIBER NAME|SUBSCRIBER NAME
C3699344|T077|strict|87226-7|LNC|INSURANCE SUBSCRIBER NAME|INSURANCE SUBSCRIBER NAME
C3699344|T077|strict|72143-1|LNC|ADMINISTRATIVE GENDER|ADMINISTRATIVE GENDER
C3699344|T077|strict|72143-1|LNC|PATIENT GENDER|PATIENT GENDER
C3699344|T077|strict|72143-1|LNC|GENDER|GENDER
C3699344|T077|strict|72143-1|LNC|PATIENT SEX|PATIENT SEX
C3699344|T077|relax|72143-1|LNC|SEX|SEX
C3699344|T077|strict|21112-8|LNC|BIRTH DATE|BIRTH DATE
C3699344|T077|strict|21112-8|LNC|DATE OF BIRTH|DATE OF BIRTH
C3699344|T077|abbr|21112-8|LNC|DOB|DOB
C3699344|T077|strict|21112-8|LNC|PATIENT DATE OF BIRTH|PATIENT DATE OF BIRTH
C3699344|T077|strict|21112-8|LNC|SUBSCRIBER DATE OF BIRTH|SUBSCRIBER DATE OF BIRTH
C3699344|T077|strict|81954-0|LNC|DATE OF DEATH|DATE OF DEATH
C3699344|T077|relax|81954-0|LNC|DEATH|DEATH
C3699344|T077|strict|21612-7|LNC|PATIENT AGE|PATIENT AGE
C3699344|T077|relax|21612-7|LNC|AGE|AGE
C3699344|T077|strict|80977-2|LNC|PATIENT RACE|PATIENT RACE
C3699344|T077|relax|80977-2|LNC|RACE|RACE
C3699344|T077|strict|80977-2|LNC|TABULATED RACE|TABULATED RACE
C3699344|T077|strict|80977-2|LNC|CDC RACE|CDC RACE
C3699344|T077|strict|80978-0|LNC|PATIENT ETHNICITY|PATIENT ETHNICITY
C3699344|T077|strict|80978-0|LNC|ETHNICITY|ETHNICITY
C3699344|T077|strict|80978-0|LNC|CDC ETHNICITY|CDC ETHNICITY
C3699344|T077|strict|80978-0|LNC|TABULATED ETHNICITY|TABULATED ETHNICITY
C3699344|T077|strict|54899-0|LNC|PREFERRED LANGUAGE|PREFERRED LANGUAGE
C3699344|T077|strict|54899-0|LNC|PREF LANGUAGE|PREF LANGUAGE
C3699344|T077|strict|54899-0|LNC|PATIENT LANGUAGE|PATIENT LANGUAGE
C3699344|T077|strict|54899-0|LNC|LANGUAGE|LANGUAGE
C3699344|T077|strict|42078-6|LNC|FOLLOW-UP CONTACT|FOLLOW-UP CONTACT
C3699344|T077|strict|42078-6|LNC|EMERGENCY CONTACT|EMERGENCY CONTACT
C3699344|T077|relax|42078-6|LNC|CONTACT|CONTACT
C3699344|T077|relax|42078-6|LNC|CONTACT BY|CONTACT BY
C3699344|T077|strict|76458-9|LNC|PATIENT EMAIL ADDRESS|PATIENT EMAIL ADDRESS
C3699344|T077|strict|76458-9|LNC|EMAIL ADDRESS|EMAIL ADDRESS
C3699344|T077|strict|76458-9|LNC|TRUSTED EMAIL|TRUSTED EMAIL
C3699344|T077|multi|76458-9|LNC|EMAIL|EMAIL
C3699344|T077|strict|92634-5|LNC|ADDRESS TYPE|ADDRESS TYPE
C3699344|T077|strict|56799-0|LNC|PATIENT ADDRESS|PATIENT ADDRESS
C3699344|T077|strict|56799-0|LNC|HOME ADDRESS|HOME ADDRESS
C3699344|T077|multi|56799-0|LNC|ADDRESS|ADDRESS
C3699344|T077|strict|56799-0|LNC|WORK ADDRESS|WORK ADDRESS
C3699344|T077|strict|56799-0|LNC|ADDRESS LINE 1|ADDRESS LINE 1
C3699344|T077|strict|56799-0|LNC|ADDRESS LINE 2|ADDRESS LINE 2
C3699344|T077|strict|56799-0|LNC|STREET ADDRESS|STREET ADDRESS
C3699344|T077|multi|56799-0|LNC|STREET|STREET
C3699344|T077|strict|42077-8|LNC|PATIENT PHONE NUMBER|PATIENT PHONE NUMBER
C3699344|T077|strict|42077-8|LNC|CELL PHONE|CELL PHONE
C3699344|T077|strict|42077-8|LNC|HOME PHONE|HOME PHONE
C3699344|T077|multi|42077-8|LNC|PHONE NUMBER|PHONE NUMBER
C3699344|T077|strict|42077-8|LNC|WORK PHONE|WORK PHONE
C3699344|T077|strict|42077-8|LNC|PHONE EXTENSION|PHONE EXTENSION
C3699344|T077|strict|42077-8|LNC|WORK PHONE EXTENSION|WORK PHONE EXTENSION
C3699344|T077|strict|42077-8|LNC|EXTENSION|EXTENSION
C3699344|T077|strict|42077-8|LNC|MOBILE PHONE|MOBILE PHONE
C3699344|T077|relax|42077-8|LNC|MOBILE|MOBILE
C3699344|T077|strict|68997-6|LNC|PATIENT CITY|PATIENT CITY
C3699344|T077|relax|68997-6|LNC|CITY|CITY
C3699344|T077|strict|46499-0|LNC|PATIENT STATE|PATIENT STATE
C3699344|T077|strict|46499-0|LNC|PATIENT HOME STATE|PATIENT HOME STATE
C3699344|T077|strict|46499-0|LNC|STATE OF RESIDENCE|STATE OF RESIDENCE
C3699344|T077|multi|46499-0|LNC|STATE|STATE
C3699344|T077|strict|45401-7|LNC|POSTAL CODE|POSTAL CODE
C3699344|T077|strict|45401-7|LNC|PATIENT ZIP|PATIENT ZIP
C3699344|T077|strict|45401-7|LNC|ZIP CODE|ZIP CODE
C3699344|T077|relax|45401-7|LNC|ZIP|ZIP
C3699344|T077|relax|45401-7|LNC|POSTAL|POSTAL
C3699344|T077|strict|87721-7|LNC|COUNTY OF RESIDENCE|COUNTY OF RESIDENCE
C3699344|T077|multi|87721-7|LNC|COUNTY|COUNTY
C3699344|T077|strict|66477-1|LNC|COUNTRY OF CURRENT RESIDENCE|COUNTRY OF CURRENT RESIDENCE
C3699344|T077|multi|66477-1|LNC|COUNTRY|COUNTRY
C3699344|T077|strict|81365-9|LNC|RELIGIOUS AFFILIATION|RELIGIOUS AFFILIATION
C3699344|T077|strict|81365-9|LNC|PATIENT RELIGION|PATIENT RELIGION
C3699344|T077|relax|81365-9|LNC|RELIGION|RELIGION
C3699344|T077|strict|85658-3|LNC|PROFESSION|PROFESSION
C3699344|T077|strict|85658-3|LNC|OCCUPATION|OCCUPATION
C3699344|T077|strict|85658-3|LNC|OCCUPATION TYPE|OCCUPATION TYPE
C3699344|T077|strict|85658-3|LNC|EMPLOYER NAME|EMPLOYER NAME
C3699344|T077|strict|85658-3|LNC|EMPLOYER ADDRESS|EMPLOYER ADDRESS
C3699344|T077|relax|85658-3|LNC|JOB|JOB
C3699344|T077|strict|46106-1|LNC|MEDICAL RECORD NUMBER|MEDICAL RECORD NUMBER
C3699344|T077|strict|46106-1|LNC|MEDICAL RECORD #|MEDICAL RECORD #
C3699344|T077|abbr|46106-1|LNC|MRN|MRN
C3699344|T077|abbr|45396-9|LNC|SSN|SSN
C3699344|T077|strict|45396-9|LNC|SOCIAL SECURITY NUMBER|SOCIAL SECURITY NUMBER
C3699344|T077|strict|45396-9|LNC|SOCIAL SECURITY NO|SOCIAL SECURITY NO
C3699344|T077|strict|45396-9|LNC|SOCIAL SECURITY NUM|SOCIAL SECURITY NUM
C3699344|T077|strict|45396-9|LNC|SOCIAL SEC NO|SOCIAL SEC NO
C3699344|T077|strict|45396-9|LNC|INSURANCE SUBSCRIBER SSN|INSURANCE SUBSCRIBER SSN
C3699344|T077|strict|45396-9|LNC|SOC SEC NO|SOC SEC NO
C3699344|T077|strict|45396-9|LNC|SOC. SEC. NO|SOC. SEC. NO
C3699344|T077|strict|45396-9|LNC|SOCIAL SECURITY|SOCIAL SECURITY
C3699344|T077|strict|76435-7|LNC|PATIENT ID|PATIENT ID
C3699344|T077|strict|76435-7|LNC|PATIENT IDENTIFIER|PATIENT IDENTIFIER
C3699344|T077|strict|76435-7|LNC|ACC|ACC
C3699344|T077|strict|76435-7|LNC|ACCOUNT|ACCOUNT
C3699344|T077|strict|76435-7|LNC|IDENTIFICATION DATA|IDENTIFICATION DATA
C3699344|T077|strict|76435-7|LNC|IDENTIFYING DATA|IDENTIFYING DATA
C3699344|T077|multi|76435-7|LNC|IDENTIFICATION|IDENTIFICATION
C3699344|T077|strict|76435-7|LNC|INSURANCE ID NUMBER|INSURANCE ID NUMBER
C3699344|T077|strict|76435-7|LNC|EXTERNAL ID|EXTERNAL ID
C3699344|T077|strict|89061-6|LNC|INSURANCE GROUP NUMBER|INSURANCE GROUP NUMBER
C3699344|T077|strict|89061-6|LNC|INSURANCE NUMBER|INSURANCE NUMBER
C3699344|T077|strict|89061-6|LNC|SECONDARY INSURANCE GROUP NUMBER|SECONDARY INSURANCE GROUP NUMBER
C3699344|T077|abbr|89061-6|LNC|INS|INS
C3699344|T077|strict|76437-3|LNC|PRIMARY INSURANCE DATA|PRIMARY INSURANCE DATA
C3699344|T077|strict|76437-3|LNC|PRIMARY INSURANCE|PRIMARY INSURANCE
C3699344|T077|strict|76437-3|LNC|ACTIVE PRIMARY INSURANCE|ACTIVE PRIMARY INSURANCE
C3699344|T077|relax|76437-3|LNC|PAYERS|PAYERS
C3699344|T077|relax|76437-3|LNC|PAYORS|PAYORS
C3699344|T077|relax|76437-3|LNC|INSURANCE|INSURANCE
C3699344|T077|strict|76437-3|LNC|SECONDARY INSURANCE|SECONDARY INSURANCE
C3699344|T077|strict|76437-3|LNC|INSURANCE COMPANY|INSURANCE COMPANY
C3699344|T077|strict|76437-3|LNC|INSURANCE DATA|INSURANCE DATA
C3699344|T077|strict|76437-3|LNC|INSURANCE PROVIDERS|INSURANCE PROVIDERS
C3699344|T077|strict|76437-3|LNC|HEALTH INSURANCE|HEALTH INSURANCE
C3699344|T077|strict|76437-3|LNC|BENEFITS ASSIGNED|BENEFITS ASSIGNED
C3699344|T077|strict|52455-3|LNC|ADMISSION DATE|ADMISSION DATE
C3699344|T077|relax|92707-9|LNC|CARE TEAM|CARE TEAM
C3699344|T077|strict|18770-8|LNC|Dictating practitioner|Dictating practitioner
C3699344|T077|strict|18770-8|LNC|DICTATED BY|DICTATED BY
C3699344|T077|strict|18770-8|LNC|FINAL DIAGNOSIS BY|FINAL DIAGNOSIS BY
C3699344|T077|strict|18770-8|LNC|AUTHOR|AUTHOR
C3699344|T077|strict|18770-8|LNC|COMPLETED BY|COMPLETED BY
C3699344|T077|strict|18770-8|LNC|ENTERED BY|ENTERED BY
C3699344|T077|strict|52525-3|LNC|DISCHARGE DATE|DISCHARGE DATE
C3699344|T077|strict|52525-3|LNC|DISCHARGE TIME|DISCHARGE TIME
C3699344|T077|strict|52525-3|LNC|DISCHARGE DATE TIME|DISCHARGE DATE TIME
C3699344|T077|strict|52525-3|LNC|DISCHARGE DATETIME|DISCHARGE DATETIME
C3699344|T077|strict|52525-3|LNC|DATE OF DISCHARGE|DATE OF DISCHARGE
C3699344|T077|strict|76696-4|LNC|Facility Name|Facility Name
C3699344|T077|strict|76696-4|LNC|Facility|Facility
C3699344|T077|strict|76696-4|LNC|SERVICE|SERVICE
C3699344|T077|strict|76696-4|LNC|BUILDING|BUILDING
C3699344|T077|strict|76696-4|LNC|CAMPUS|CAMPUS
C3699344|T077|strict|76696-4|LNC|DEPARTMENT|DEPARTMENT
C3699344|T077|strict|18841-7|LNC|HOSPITAL CONSULTATIONS|HOSPITAL CONSULTATIONS
C3699344|T077|strict|18841-7|LNC|CONSULT|CONSULT
C3699344|T077|strict|18841-7|LNC|CONSULTATION|CONSULTATION
C3699344|T077|strict|78033-8|LNC|HOSPITAL STAY DURATION|HOSPITAL STAY DURATION
C3699344|T077|strict|78033-8|LNC|LENGTH OF STAY|LENGTH OF STAY
C3699344|T077|abbr|78033-8|LNC|LOS|LOS
C3699344|T077|strict|48768-6|LNC|PAYMENT SOURCES|PAYMENT SOURCES
C3699344|T077|strict|22028-5|LNC|Physician|Physician
C3699344|T077|strict|22028-5|LNC|PROVIDER|PROVIDER
C3699344|T077|strict|22028-5|LNC|DOCTOR|DOCTOR
C3699344|T077|strict|22028-5|LNC|ATTENDING|ATTENDING
C3699344|T077|strict|22028-5|LNC|RESIDENT|RESIDENT
C3699344|T077|strict|22028-5|LNC|PCP|PCP
C3699344|T077|strict|22028-5|LNC|PCP NAME|PCP NAME
C3699344|T077|strict|22028-5|LNC|OBSTETRICIAN|OBSTETRICIAN
C3699344|T077|strict|22028-5|LNC|SUPERVISING|SUPERVISING
C3699344|T077|strict|22028-5|LNC|SEEN BY|SEEN BY
C3699344|T077|strict|75519-9|LNC|ENCOUNTER|ENCOUNTER
C3699344|T077|strict|75519-9|LNC|ENCOUNTER INFO|ENCOUNTER INFO
C3699344|T077|strict|75519-9|LNC|ED VISITS|ED VISITS
C3699344|T077|strict|75519-9|LNC|APPOINTMENT|APPOINTMENT
C3699344|T077|strict|75519-9|LNC|APPOINTMENTS|APPOINTMENTS
C3699344|T077|strict|56816-2|LNC|LOCATION|LOCATION
C3699344|T077|strict|56816-2|LNC|ROOM|ROOM
C3699344|T077|strict|44951-2|LNC|National Provider Identifier|National Provider Identifier
C3699344|T077|abbr|44951-2|LNC|NPI|NPI
C3699344|T077|strict|44951-2|LNC|PROVIDER ID|PROVIDER ID
C3699344|T077|strict|44951-2|LNC|PROVIDER NUMBER|PROVIDER NUMBER
C3699344|T077|strict|11347-2|LNC|History of outpatient visits|History of outpatient visits
C3699344|T077|strict|11347-2|LNC|outpatient visits|outpatient visits
C3699344|T077|strict|11337-3|LNC|HISTORY OF HOSPITALIZATIONS|HISTORY OF HOSPITALIZATIONS
C3699344|T077|strict|11293-8|LNC|Referral source|Referral source
C3699344|T077|strict|11293-8|LNC|REFERRED BY|REFERRED BY
C3699344|T077|strict|85647-6|LNC|SIGNATURE|SIGNATURE
C3699344|T077|strict|85647-6|LNC|SIGNATURE LINE|SIGNATURE LINE
C3699344|T077|strict|85647-6|LNC|ELECTRONICALLY SIGNED|ELECTRONICALLY SIGNED
C3699344|T077|strict|85647-6|LNC|SIGNED|SIGNED
C3699344|T077|strict|85647-6|LNC|SIGNED ELECTRONICALLY BY|SIGNED ELECTRONICALLY BY
C3699344|T077|strict|85647-6|LNC|SIGNATURE ON FILE|SIGNATURE ON FILE
C3699344|T077|strict|19826-7|LNC|INFORMED CONSENT|INFORMED CONSENT
C3699344|T077|relax|19826-7|LNC|CONSENT|CONSENT
C3699344|T077|strict|39289-4|LNC|FOLLOW UP APPOINTMENT|FOLLOW UP APPOINTMENT
C3699344|T077|strict|39289-4|LNC|FOLLOW UP APPOINTMENTS|FOLLOW UP APPOINTMENTS
C3699344|T077|strict|76427-4|LNC|VISIT DATE|VISIT DATE
C3699344|T077|strict|76427-4|LNC|ENCOUNTER DATE|ENCOUNTER DATE
C3699344|T077|strict|76427-4|LNC|DATE TIME|DATE TIME
C3699344|T077|strict|76427-4|LNC|REGISTRATION DATE|REGISTRATION DATE
C3699344|T077|strict|30947-6|LNC|RECORD DATE|RECORD DATE
C3699344|T077|strict|67162-8|LNC|DISPOSITION|DISPOSITION
C3699344|T077|strict|67162-8|LNC|Patient Disposition|Patient Disposition
C3699344|T077|strict|67162-8|LNC|DISPOSITION ON DISCHARGE|DISPOSITION ON DISCHARGE
C3699344|T077|relax|71727-2|LNC|FAX|FAX
C3699344|T077|strict|46240-8|LNC|HISTORY OF HOSPITALIZATIONS+OUTPATIENT VISITS|HISTORY OF HOSPITALIZATIONS+OUTPATIENT VISITS
C3699344|T077|strict|46240-8|LNC|HISTORY OF HOSPITALIZATIONS|HISTORY OF HOSPITALIZATIONS
C3699344|T077|strict|46240-8|LNC|HISTORY OF ENCOUNTERS|HISTORY OF ENCOUNTERS
C3699344|T077|strict|46240-8|LNC|HOSPITALIZATIONS|HOSPITALIZATIONS
C3699344|T077|strict|46240-8|LNC|HOSPITALIZATION|HOSPITALIZATION
C3699344|T077|relax|46240-8|LNC|ENCOUNTERS|ENCOUNTERS
C3699344|T077|strict|55111-9|LNC|CURRENT IMAGING PROCEDURE DESCRIPTIONS|CURRENT IMAGING PROCEDURE DESCRIPTIONS
C3699344|T077|strict|55111-9|LNC|CURRENT IMAGING PROCEDURE|CURRENT IMAGING PROCEDURE
C3699344|T077|strict|47519-4|LNC|HISTORY OF PROCEDURES|HISTORY OF PROCEDURES
C3699344|T077|strict|47519-4|LNC|PROCEDURES HX DOC|PROCEDURES HX DOC
C3699344|T077|strict|47519-4|LNC|PROCEDURES HX|PROCEDURES HX
C3699344|T077|relax|47519-4|LNC|PROCEDURES|PROCEDURES
C3699344|T077|strict|59772-4|LNC|PLANNED PROCEDURE|PLANNED PROCEDURE
C3699344|T077|strict|55114-3|LNC|PRIOR PROCEDURE DESCRIPTIONS|PRIOR PROCEDURE DESCRIPTIONS
C3699344|T077|strict|55114-3|LNC|PRIOR PROCEDURE HISTORY|PRIOR PROCEDURE HISTORY
C3699344|T077|strict|55114-3|LNC|PROCEDURE HISTORY|PROCEDURE HISTORY
C3699344|T077|strict|55114-3|LNC|PROCEDURES HISTORY|PROCEDURES HISTORY
C3699344|T077|strict|29554-3|LNC|PROCEDURE DESCRIPTION|PROCEDURE DESCRIPTION
C3699344|T077|strict|29554-3|LNC|PROCEDURE LIST|PROCEDURE LIST
C3699344|T077|strict|29554-3|LNC|PROCEDURES AND SURGICAL/MEDICAL HISTORY|PROCEDURES AND SURGICAL/MEDICAL HISTORY
C3699344|T077|strict|29554-3|LNC|PRINCIPAL PROCEDURE|PRINCIPAL PROCEDURE
C3699344|T077|relax|29554-3|LNC|PROCEDURE|PROCEDURE
C3699344|T077|strict|59775-7|LNC|PROCEDURE DISPOSITION|PROCEDURE DISPOSITION
C3699344|T077|strict|59773-2|LNC|PROCEDURE SPECIMENS TAKEN|PROCEDURE SPECIMENS TAKEN
C3699344|T077|strict|55115-0|LNC|REQUESTED IMAGING STUDIES INFORMATION|REQUESTED IMAGING STUDIES INFORMATION
C3699344|T077|strict|55115-0|LNC|REQUESTED IMAGING STUDIES|REQUESTED IMAGING STUDIES
C3699344|T077|strict|55115-0|LNC|IMAGING STUDIES|IMAGING STUDIES
C3699344|T077|strict|55115-0|LNC|RADIOGRAPHIC STUDIES|RADIOGRAPHIC STUDIES
C3699344|T077|strict|55115-0|LNC|RADIOLOGIC STUDIES|RADIOLOGIC STUDIES
C3699344|T077|strict|55115-0|LNC|RADIOLOGY IMAGING|RADIOLOGY IMAGING
C3699344|T077|strict|55115-0|LNC|RELEVANT IMAGING|RELEVANT IMAGING
C3699344|T077|relax|55115-0|LNC|RADIOGRAPHIC|RADIOGRAPHIC
C3699344|T077|relax|55115-0|LNC|RADIOLOGY|RADIOLOGY
C3699344|T077|relax|55115-0|LNC|IMAGING|IMAGING
C3699344|T077|abbr|55115-0|LNC|ECG|ECG
C3699344|T077|abbr|55115-0|LNC|EKG|EKG
C3699344|T077|abbr|55115-0|LNC|ECHO|ECHO
C3699344|T077|abbr|55115-0|LNC|EEG|EEG
C3699344|T077|relax|55115-0|LNC|ELECTROCARDIOGRAM|ELECTROCARDIOGRAM
C3699344|T077|relax|55115-0|LNC|CHEST XRAY|CHEST XRAY
C3699344|T077|abbr|55115-0|LNC|CXR|CXR
C3699344|T077|abbr|55115-0|LNC|MRA KIDNEY|MRA KIDNEY
C3699344|T077|abbr|55115-0|LNC|MRI HEAD|MRI HEAD
C3699344|T077|abbr|55115-0|LNC|KUB|KUB
C3699344|T077|strict|59774-0|LNC|PROCEDURE ANESTHESIA|PROCEDURE ANESTHESIA
C3699344|T077|strict|59774-0|LNC|ANESTHESIA SECTION|ANESTHESIA SECTION
C3699344|T077|strict|59774-0|LNC|PRIMARY ANESTHESIA|PRIMARY ANESTHESIA
C3699344|T077|relax|59774-0|LNC|ANESTHESIA|ANESTHESIA
C3699344|T077|strict|8724-7|LNC|DESCRIPTION OF OPERATION|DESCRIPTION OF OPERATION
C3699344|T077|strict|8724-7|LNC|DESCRIPTION OF THE OPERATION|DESCRIPTION OF THE OPERATION
C3699344|T077|strict|8724-7|LNC|TITLE OF OPERATION|TITLE OF OPERATION
C3699344|T077|strict|8724-7|LNC|OPERATION DESCRIPTION|OPERATION DESCRIPTION
C3699344|T077|strict|8724-7|LNC|OPERATION PERFORMED|OPERATION PERFORMED
C3699344|T077|strict|8724-7|LNC|NAME OF OPERATION|NAME OF OPERATION
C3699344|T077|strict|59770-8|LNC|PROCEDURE ESTIMATED BLOOD LOSS|PROCEDURE ESTIMATED BLOOD LOSS
C3699344|T077|multi|59770-8|LNC|BLOOD LOSS|BLOOD LOSS
C3699344|T077|relax|59770-8|LNC|ESTIMATED BLOOD LOSS|ESTIMATED BLOOD LOSS
C3699344|T077|strict|8690-0|LNC|History of Surgical procedures|History of Surgical procedures
C3699344|T077|strict|8690-0|LNC|PAST SURGICAL HISTORY|PAST SURGICAL HISTORY
C3699344|T077|strict|8690-0|LNC|SURGICAL HISTORY|SURGICAL HISTORY
C3699344|T077|relax|8690-0|LNC|OPERATIONS|OPERATIONS
C3699344|T077|relax|8690-0|LNC|OPERATIONS PERFORMED|OPERATIONS PERFORMED
C3699344|T077|relax|8690-0|LNC|OPERATION|OPERATION
C3699344|T077|relax|8690-0|LNC|SURGERIES|SURGERIES
C3699344|T077|strict|11537-8|LNC|SURGICAL DRAINS|SURGICAL DRAINS
C3699344|T077|strict|11537-8|LNC|SURGICAL DRAINS NOTE|SURGICAL DRAINS NOTE
C3699344|T077|strict|59771-6|LNC|PROCEDURE IMPLANTS|PROCEDURE IMPLANTS
C3699344|T077|relax|59771-6|LNC|IMPLANTS|IMPLANTS
C3699344|T077|strict|10216-0|LNC|SURGICAL OPERATION NOTE FLUIDS|SURGICAL OPERATION NOTE FLUIDS
C3699344|T077|strict|10216-0|LNC|OPERATIVE NOTE FLUIDS|OPERATIVE NOTE FLUIDS
C3699344|T077|strict|10223-6|LNC|SURGICAL OPERATION NOTE SURGICAL PROCEDURE|SURGICAL OPERATION NOTE SURGICAL PROCEDURE
C3699344|T077|strict|10223-6|LNC|OPERATIVE NOTE SURGICAL|OPERATIVE NOTE SURGICAL
C3699344|T077|strict|10223-6|LNC|SURGICAL PROCEDURE|SURGICAL PROCEDURE
C3699344|T077|strict|22637-3|LNC|PATHOLOGY REPORT FINAL DIAGNOSIS|PATHOLOGY REPORT FINAL DIAGNOSIS
C3699344|T077|strict|22637-3|LNC|HISTOPATHOLOGICAL DIAGNOSIS|HISTOPATHOLOGICAL DIAGNOSIS
C3699344|T077|strict|22637-3|LNC|PATHOLOGIC DIAGNOSIS|PATHOLOGIC DIAGNOSIS
C3699344|T077|multi|22637-3|LNC|FINAL DIAGNOSES|FINAL DIAGNOSES
C3699344|T077|multi|22637-3|LNC|FINAL DIAGNOSIS|FINAL DIAGNOSIS
C3699344|T077|strict|33746-9|LNC|PATHOLOGIC FINDINGS|PATHOLOGIC FINDINGS
C3699344|T077|strict|33746-9|LNC|ADDITIONAL PATHOLOGIC FINDINGS|ADDITIONAL PATHOLOGIC FINDINGS
C3699344|T077|strict|83321-0|LNC|INTRAOPERATIVE DIAGNOSIS|INTRAOPERATIVE DIAGNOSIS
C3699344|T077|strict|22634-0|LNC|MACROSCOPIC ANATOMIC OBSERVATIONS|MACROSCOPIC ANATOMIC OBSERVATIONS
C3699344|T077|strict|22634-0|LNC|MACROSCOPIC OBSERVATIONS|MACROSCOPIC OBSERVATIONS
C3699344|T077|strict|22634-0|LNC|MACROSCOPIC DESCRIPTION|MACROSCOPIC DESCRIPTION
C3699344|T077|strict|22634-0|LNC|MACROSCOPIC EXAMINATION|MACROSCOPIC EXAMINATION
C3699344|T077|strict|22634-0|LNC|MACROSCOPY|MACROSCOPY
C3699344|T077|strict|22634-0|LNC|SPECIMEN SIZE|SPECIMEN SIZE
C3699344|T077|strict|22634-0|LNC|TUMOR SIZE|TUMOR SIZE
C3699344|T077|strict|22634-0|LNC|TUMOR EXTENT|TUMOR EXTENT
C3699344|T077|strict|22634-0|LNC|PATHOLOGY REPORT GROSS OBSERVATION|PATHOLOGY REPORT GROSS OBSERVATION
C3699344|T077|strict|22634-0|LNC|PATHOLOGY REPORT GROSS DESCRIPTION|PATHOLOGY REPORT GROSS DESCRIPTION
C3699344|T077|strict|22634-0|LNC|GROSS OBSERVATION|GROSS OBSERVATION
C3699344|T077|strict|22634-0|LNC|GROSS DESCRIPTION|GROSS DESCRIPTION
C3699344|T077|strict|22634-0|LNC|GROSS DESCRIPTION TEXT|GROSS DESCRIPTION TEXT
C3699344|T077|strict|22634-0|LNC|GROSS TEXT|GROSS TEXT
C3699344|T077|strict|22634-0|LNC|GROSS FINDINGS|GROSS FINDINGS
C3699344|T077|strict|22634-0|LNC|GROSSLY EVIDENT LESION|GROSSLY EVIDENT LESION
C3699344|T077|strict|22635-7|LNC|MICROSCOPIC OBSERVATION|MICROSCOPIC OBSERVATION
C3699344|T077|strict|22635-7|LNC|MICROSCOPIC DESCRIPTION|MICROSCOPIC DESCRIPTION
C3699344|T077|strict|22635-7|LNC|MICROSCOPIC EXAMINATION|MICROSCOPIC EXAMINATION
C3699344|T077|strict|33732-9|LNC|HISTOLOGIC GRADE|HISTOLOGIC GRADE
C3699344|T077|strict|33732-9|LNC|HISTOLOGIC TYPE|HISTOLOGIC TYPE
C3699344|T077|strict|21859-4|LNC|ANATOMIC SITE|ANATOMIC SITE
C3699344|T077|strict|21859-4|LNC|SITE OF TISSUE|SITE OF TISSUE
C3699344|T077|strict|21859-4|LNC|TISSUE SITE|TISSUE SITE
C3699344|T077|strict|21859-4|LNC|TUMOR LOCATION|TUMOR LOCATION
C3699344|T077|strict|21859-4|LNC|TUMOR SITE|TUMOR SITE
C3699344|T077|strict|21939-4|LNC|SURGICAL MARGINS|SURGICAL MARGINS
C3699344|T077|relax|21939-4|LNC|MARGINS|MARGINS
C3699344|T077|strict|42186-7|LNC|RECEIVED SPECIMEN|RECEIVED SPECIMEN
C3699344|T077|strict|42186-7|LNC|MATERIAL COLLECTED ON|MATERIAL COLLECTED ON
C3699344|T077|strict|42186-7|LNC|MATERIAL RECEIVED ON|MATERIAL RECEIVED ON
C3699344|T077|strict|42186-7|LNC|MATERIAL RECEIVED|MATERIAL RECEIVED
C3699344|T077|strict|66746-9|LNC|SPECIMEN TYPE|SPECIMEN TYPE
C3699344|T077|strict|66746-9|LNC|SPECIMEN|SPECIMEN
C3699344|T077|strict|66746-9|LNC|SPECIMENS|SPECIMENS
C3699344|T077|strict|66746-9|LNC|TISSUE SPECIFICATION|TISSUE SPECIFICATION
C3699344|T077|strict|90041-5|LNC|SPECIMEN COLLECTION|SPECIMEN COLLECTION
C3699344|T077|strict|90041-5|LNC|MATERIAL COLLECTED|MATERIAL COLLECTED
C3699344|T077|strict|90041-5|LNC|SPECIMEN SUBMITTED|SPECIMEN SUBMITTED
C3699344|T077|strict|90041-5|LNC|SPECIMENS SUBMITTED|SPECIMENS SUBMITTED
C3699344|T077|strict|90041-5|LNC|TISSUE SUBMITTED|TISSUE SUBMITTED
C3699344|T077|relax|67203-0|LNC|AJCC CLASSIFICATION|AJCC CLASSIFICATION
C3699344|T077|relax|67203-0|LNC|AJCC STAGING|AJCC STAGING
C3699344|T077|relax|67203-0|LNC|AJCC|AJCC
C3699344|T077|relax|92833-3|LNC|LYMPH NODES|LYMPH NODES
C3699344|T077|strict|75621-3|LNC|TNM PATHOLOGIC STAGING AFTER SURGERY PANEL|TNM PATHOLOGIC STAGING AFTER SURGERY PANEL
C3699344|T077|strict|75621-3|LNC|TNM PATHOLOGIC STAGING|TNM PATHOLOGIC STAGING
C3699344|T077|strict|75621-3|LNC|TNM STAGING|TNM STAGING
C3699344|T077|strict|75621-3|LNC|PATHOLOGIC STAGE|PATHOLOGIC STAGE
C3699344|T077|strict|75621-3|LNC|NOTTINGHAM HISTOLOGIC SCORE|NOTTINGHAM HISTOLOGIC SCORE
C3699344|T077|relax|75621-3|LNC|TNM STAGE|TNM STAGE
C3699344|T077|relax|75621-3|LNC|STAGING|STAGING
C3699344|T077|strict|90947-3|LNC|PATHOLOGY CASE|PATHOLOGY CASE
C3699344|T077|strict|75321-0|LNC|CLINICAL FINDING|CLINICAL FINDING
C3699344|T077|strict|75321-0|LNC|FINDINGS|FINDINGS
C3699344|T077|strict|75321-0|LNC|INTERPRETATION|INTERPRETATION
C3699344|T077|multi|55752-0|LNC|CLINICAL INFORMATION|CLINICAL INFORMATION
C3699344|T077|multi|55752-0|LNC|CLINICAL DATA|CLINICAL DATA
C3699344|T077|strict|55107-7|LNC|ADDENDUM|ADDENDUM
C3699344|T077|strict|55107-7|LNC|AMENDMENTS|AMENDMENTS
C3699344|T077|strict|91582-7|LNC|REPORT STATUS|REPORT STATUS
C3699344|T077|strict|48766-0|LNC|SOURCE|SOURCE
C3699344|T077|multi|55112-7|LNC|DOCUMENT SUMMARY|DOCUMENT SUMMARY
C3699344|T077|relax|55112-7|LNC|SUMMARY|SUMMARY