C0011570|T048|41006004|SNOMEDCT_US|MENTAL DEPRESSION|DEPRESSION (FINDING)
C0011581|T048|192372006|SNOMEDCT_US|DEPRESSIVE DISORDER|[X]DEPRESSIVE DISORDER NOS
C1999266|T048||SNOMEDCT_US|DEPRESSION ADVERSE EVENT
C4049644|T048||SNOMEDCT_US|DEPRESSION SCALE (BASC-2)
C4084909|T048||SNOMEDCT_US|DEPRESSION SUBORDINATE DOMAIN
C4085311|T048||SNOMEDCT_US|DEPRESSION - RECESS
C0743072|T048||SNOMEDCT_US|PSYCHOTIC DEPRESSION
C0743072|T048||SNOMEDCT_US|DEPRESSIVE PSYCHOSIS
C0743072|T048||SNOMEDCT_US|DEPRESSION;PSYCHOTIC
C0743072|T048||SNOMEDCT_US|PSYCHOSIS;DEPRESSIVE
C0743072|T048||SNOMEDCT_US|DEPRESSIVE PSYCHOSES
C0743072|T048||SNOMEDCT_US|DEPRESSION, PSYCHOTIC
C0743072|T048||SNOMEDCT_US|DEPRESSION PSYCHOTIC
C0743072|T048||SNOMEDCT_US|PSYCHOSIS DEPRESSIVE
C0743072|T048||SNOMEDCT_US|DEPRESSION; PSYCHOTIC
C0743072|T048||SNOMEDCT_US|DEPRESSIVE; PSYCHOSIS
C0743072|T048||SNOMEDCT_US|PSYCHOSIS; DEPRESSIVE
C0743072|T048||SNOMEDCT_US|PSYCHOTIC; DEPRESSION
C0541868|T048||SNOMEDCT_US|DEPRESSION FUNCTIONAL
C0541869|T048||SNOMEDCT_US|DEPRESSION WORSENED
C0221074|T048|147016002|SNOMEDCT_US|POSTPARTUM DEPRESSION|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|DEPRESSION, POST-NATAL|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|DEPRESSION, POST-PARTUM|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|DEPRESSION, POSTNATAL|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|DEPRESSION, POSTPARTUM|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|POST NATAL DEPRESSION|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|POST PARTUM DEPRESSION|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|POSTPARTUM DEPRESSION |POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|DEPRESSION, POSTPARTUM [DISEASE/FINDING]|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|POST-NATAL DEPRESSION|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|POST-PARTUM DEPRESSION|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|POSTNATAL DEPRESSION|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|DEPRESSION;POSTNATAL|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|DEPRESSION;PUERPERAL|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|DEPRESSION POSTPARTUM (EXCL PSYCHOSIS)|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|[X]POSTNATAL DEPRESSION NOS|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|[X]POSTPARTUM DEPRESSION NOS|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|DEPRESSION - POSTNATAL|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|POSTNATAL DEPRESSIVE DISORDER |POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|POSTNATAL DEPRESSIVE DISORDER|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|DEPRESSIVE EPISODE WITH POSTPARTUM ONSET|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|MAJOR DEPRESSIVE EPISODE WITH PERIPARTUM ONSET|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|POSTNATAL DEPRESSION (EXCL PSYCHOSIS)|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|DEPRESSION PUERPERAL|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|PUERPERAL DEPRESSION|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|POSTNATAL DEPRESSION (EXCLUDING PSYCHOSIS)|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|POSTPARTUM DEPRESSION |POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|DEPRESSION; POSTNATAL|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|DEPRESSION; POSTPARTUM|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|POSTNATAL; DEPRESSION|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|POSTPARTUM; DEPRESSION|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0221074|T048|147016002|SNOMEDCT_US|DEPRESSION POSTPARTUM (EXCLUDING PSYCHOSIS)|POSTNATAL DEPRESSIVE DISORDER (DISORDER)
C0494397|T048|192367002|SNOMEDCT_US|MILD DEPRESSIVE EPISODE|[X]MILD DEPRESSIVE EPISODE (DISORDER)
C0494397|T048|192367002|SNOMEDCT_US|[X]MILD DEPRESSIVE EPISODE |[X]MILD DEPRESSIVE EPISODE (DISORDER)
C0494397|T048|192367002|SNOMEDCT_US|[X]MILD DEPRESSIVE EPISODE|[X]MILD DEPRESSIVE EPISODE (DISORDER)
C0494397|T048|192367002|SNOMEDCT_US|EPISODE; DEPRESSIVE, MILD|[X]MILD DEPRESSIVE EPISODE (DISORDER)
C0494398|T048|192368007|SNOMEDCT_US|MODERATE DEPRESSIVE EPISODE|[X]MODERATE DEPRESSIVE EPISODE (DISORDER)
C0494398|T048|192368007|SNOMEDCT_US|[X]MODERATE DEPRESSIVE EPISODE |[X]MODERATE DEPRESSIVE EPISODE (DISORDER)
C0494398|T048|192368007|SNOMEDCT_US|[X]MODERATE DEPRESSIVE EPISODE|[X]MODERATE DEPRESSIVE EPISODE (DISORDER)
C0494398|T048|192368007|SNOMEDCT_US|EPISODE; DEPRESSIVE, MODERATE|[X]MODERATE DEPRESSIVE EPISODE (DISORDER)
C0154411|T048|18818009|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, RECURRENT EPISODE, MODERATE DEGREE|MODERATE RECURRENT MAJOR DEPRESSION (DISORDER)
C0154411|T048|18818009|SNOMEDCT_US|RECURRENT DEPRESSIVE DISORDER, CURRENT EPISODE MODERATE|MODERATE RECURRENT MAJOR DEPRESSION (DISORDER)
C0154411|T048|18818009|SNOMEDCT_US|MODERATE RECURRENT MAJOR DEPRESSION |MODERATE RECURRENT MAJOR DEPRESSION (DISORDER)
C0154411|T048|18818009|SNOMEDCT_US|MODERATE RECURRENT MAJOR DEPRESSION|MODERATE RECURRENT MAJOR DEPRESSION (DISORDER)
C0154411|T048|18818009|SNOMEDCT_US|RECURR DEPR PSYCHOS-MOD|MODERATE RECURRENT MAJOR DEPRESSION (DISORDER)
C0154411|T048|18818009|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, RECURRENT, MODERATE|MODERATE RECURRENT MAJOR DEPRESSION (DISORDER)
C0154411|T048|18818009|SNOMEDCT_US|MAJOR DEPRESSIVE AFFECTIVE DISORDER, RECURRENT EPISODE, MODERATE|MODERATE RECURRENT MAJOR DEPRESSION (DISORDER)
C0154411|T048|18818009|SNOMEDCT_US|[X]RECURRENT DEPRESSIVE DISORDER, CURRENT EPISODE MODERATE |MODERATE RECURRENT MAJOR DEPRESSION (DISORDER)
C0154411|T048|18818009|SNOMEDCT_US|[X]RECURRENT DEPRESSIVE DISORDER, CURRENT EPISODE MODERATE|MODERATE RECURRENT MAJOR DEPRESSION (DISORDER)
C0154411|T048|18818009|SNOMEDCT_US|MODERATE RECURRENT MAJOR DEPRESSION |MODERATE RECURRENT MAJOR DEPRESSION (DISORDER)
C0235876|T048||SNOMEDCT_US|DEPRESSION AGGRAVATED
C0236764|T048|33135002|SNOMEDCT_US|RECURRENT MAJOR DEPRESSION IN PARTIAL REMISSION|RECURRENT MAJOR DEPRESSION IN PARTIAL REMISSION (DISORDER)
C0236764|T048|33135002|SNOMEDCT_US|RECURRENT MAJOR DEPRESSION IN PARTIAL REMISSION |RECURRENT MAJOR DEPRESSION IN PARTIAL REMISSION (DISORDER)
C0236764|T048|33135002|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, RECURRENT, IN PARTIAL REMISSION|RECURRENT MAJOR DEPRESSION IN PARTIAL REMISSION (DISORDER)
C0236764|T048|33135002|SNOMEDCT_US|RECURRENT MAJOR DEPRESSION IN PARTIAL REMISSION |RECURRENT MAJOR DEPRESSION IN PARTIAL REMISSION (DISORDER)
C0041696|T048||SNOMEDCT_US|DEPRESSIONS, UNIPOLAR
C0041696|T048||SNOMEDCT_US|UNIPOLAR DEPRESSIONS
C0041696|T048||SNOMEDCT_US|UNIPOLAR DEPRESSION
C0041696|T048||SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER
C0041696|T048||SNOMEDCT_US|MAJOR DEPRESSION
C0041696|T048||SNOMEDCT_US|UNIPOLAR DEPRESSIVE ILLNESS
C0041696|T048||SNOMEDCT_US|DEPRESSION, UNIPOLAR
C0154403|T048|79298009|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE, MILD DEGREE|MILD MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0154403|T048|79298009|SNOMEDCT_US|MILD SINGLE EPISODE MAJOR DEPRESSION |MILD MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0154403|T048|79298009|SNOMEDCT_US|MILD SINGLE EPISODE MAJOR DEPRESSION|MILD MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0154403|T048|79298009|SNOMEDCT_US|DEPRESS PSYCHOSIS-MILD|MILD MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0154403|T048|79298009|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE, MILD|MILD MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0154403|T048|79298009|SNOMEDCT_US|MAJOR DEPRESSIVE AFFECTIVE DISORDER, SINGLE EPISODE, MILD|MILD MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0154403|T048|79298009|SNOMEDCT_US|MILD MAJOR DEPRESSION, SINGLE EPISODE|MILD MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0154403|T048|79298009|SNOMEDCT_US|SINGLE MAJOR DEPRESSIVE EPISODE, MILD|MILD MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0154403|T048|79298009|SNOMEDCT_US|MILD MAJOR DEPRESSION, SINGLE EPISODE |MILD MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0154403|T048|79298009|SNOMEDCT_US|SINGLE MAJOR DEPRESSIVE EPISODE, MILD |MILD MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0154403|T048|79298009|SNOMEDCT_US|DISORDER; DEPRESSIVE, MAJOR, SINGLE EPISODE, MILD|MILD MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0154404|T048|15639000|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE, MODERATE DEGREE|MODERATE MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0154404|T048|15639000|SNOMEDCT_US|MODERATE SINGLE EPISODE MAJOR DEPRESSION |MODERATE MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0154404|T048|15639000|SNOMEDCT_US|MODERATE SINGLE EPISODE MAJOR DEPRESSION|MODERATE MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0154404|T048|15639000|SNOMEDCT_US|DEPRESSIVE PSYCHOSIS-MOD|MODERATE MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0154404|T048|15639000|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE, MODERATE|MODERATE MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0154404|T048|15639000|SNOMEDCT_US|MAJOR DEPRESSIVE AFFECTIVE DISORDER, SINGLE EPISODE, MODERATE|MODERATE MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0154404|T048|15639000|SNOMEDCT_US|MODERATE MAJOR DEPRESSION, SINGLE EPISODE|MODERATE MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0154404|T048|15639000|SNOMEDCT_US|SINGLE MAJOR DEPRESSIVE EPISODE, MODERATE|MODERATE MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0154404|T048|15639000|SNOMEDCT_US|MODERATE MAJOR DEPRESSION, SINGLE EPISODE |MODERATE MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0154404|T048|15639000|SNOMEDCT_US|SINGLE MAJOR DEPRESSIVE EPISODE, MODERATE |MODERATE MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0154404|T048|15639000|SNOMEDCT_US|DISORDER; DEPRESSIVE, MAJOR, SINGLE EPISODE, MODERATE|MODERATE MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C3665435|T048|191610000|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, RECURRENT EPISODE, MILD DEGREE|RECURRENT MAJOR DEPRESSIVE EPISODES, MILD (DISORDER)
C3665435|T048|191610000|SNOMEDCT_US|RECURR DEPR PSYCHOS-MILD|RECURRENT MAJOR DEPRESSIVE EPISODES, MILD (DISORDER)
C3665435|T048|191610000|SNOMEDCT_US|MAJOR DEPRESSIVE AFFECTIVE DISORDER, RECURRENT EPISODE, MILD|RECURRENT MAJOR DEPRESSIVE EPISODES, MILD (DISORDER)
C3665435|T048|191610000|SNOMEDCT_US|MAJOR DEPRESSION, RECURRENT, MILD EPISODE|RECURRENT MAJOR DEPRESSIVE EPISODES, MILD (DISORDER)
C3665435|T048|191610000|SNOMEDCT_US|RECURRENT MAJOR DEPRESSIVE EPISODE, MILD |RECURRENT MAJOR DEPRESSIVE EPISODES, MILD (DISORDER)
C3665435|T048|191610000|SNOMEDCT_US|RECURRENT MAJOR DEPRESSIVE EPISODE, MILD|RECURRENT MAJOR DEPRESSIVE EPISODES, MILD (DISORDER)
C3665435|T048|191610000|SNOMEDCT_US|RECURRENT MAJOR DEPRESSIVE EPISODES, MILD|RECURRENT MAJOR DEPRESSIVE EPISODES, MILD (DISORDER)
C3665435|T048|191610000|SNOMEDCT_US|RECURRENT MAJOR DEPRESSIVE EPISODES, MILD |RECURRENT MAJOR DEPRESSIVE EPISODES, MILD (DISORDER)
C0154412|T048|192377000|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, RECURRENT EPISODE, SEVERE DEGREE, WITHOUT MENTION OF PSYCHOTIC BEHAVIOR|[X]MAJOR DEPRESSION, RECURRENT WITHOUT PSYCHOTIC SYMPTOMS
C0154412|T048|192377000|SNOMEDCT_US|RECURRENT DEPRESSIVE DISORDER, CURRENT EPISODE SEVERE WITHOUT PSYCHOTIC SYMPTOMS|[X]MAJOR DEPRESSION, RECURRENT WITHOUT PSYCHOTIC SYMPTOMS
C0154412|T048|192377000|SNOMEDCT_US|SEVERE RECURRENT MAJOR DEPRESSION WITHOUT PSYCHOTIC FEATURES|[X]MAJOR DEPRESSION, RECURRENT WITHOUT PSYCHOTIC SYMPTOMS
C0154412|T048|192377000|SNOMEDCT_US|SEVERE RECURRENT MAJOR DEPRESSION WITHOUT PSYCHOTIC FEATURES |[X]MAJOR DEPRESSION, RECURRENT WITHOUT PSYCHOTIC SYMPTOMS
C0154412|T048|192377000|SNOMEDCT_US|RECUR DEPR PSYCH-SEVERE|[X]MAJOR DEPRESSION, RECURRENT WITHOUT PSYCHOTIC SYMPTOMS
C0154412|T048|192377000|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, RECURRENT SEVERE WITHOUT PSYCHOTIC FEATURES|[X]MAJOR DEPRESSION, RECURRENT WITHOUT PSYCHOTIC SYMPTOMS
C0154412|T048|192377000|SNOMEDCT_US|MAJOR DEPRESSV DISORDER, RECURRENT SEVERE W/O PSYCH FEATURES|[X]MAJOR DEPRESSION, RECURRENT WITHOUT PSYCHOTIC SYMPTOMS
C0154412|T048|192377000|SNOMEDCT_US|MAJOR DEPRESSIVE AFFECTIVE DISORDER, RECURRENT EPISODE, SEVERE, WITHOUT MENTION OF PSYCHOTIC BEHAVIOR|[X]MAJOR DEPRESSION, RECURRENT WITHOUT PSYCHOTIC SYMPTOMS
C0154412|T048|192377000|SNOMEDCT_US|[X]MAJOR DEPRESSION, RECURRENT WITHOUT PSYCHOTIC SYMPTOMS|[X]MAJOR DEPRESSION, RECURRENT WITHOUT PSYCHOTIC SYMPTOMS
C0154412|T048|192377000|SNOMEDCT_US|[X]RECURRENT DEPRESSIVE DISORDER, CURRENT EPISODE SEVERE WITHOUT PSYCHOTIC SYMPTOMS|[X]MAJOR DEPRESSION, RECURRENT WITHOUT PSYCHOTIC SYMPTOMS
C0154412|T048|192377000|SNOMEDCT_US|[X]RECURRENT DEPRESSIVE DISORDER, CURRENT EPISODE SEVERE WITHOUT PSYCHOTIC SYMPTOMS |[X]MAJOR DEPRESSION, RECURRENT WITHOUT PSYCHOTIC SYMPTOMS
C0154412|T048|192377000|SNOMEDCT_US|SEVERE RECURRENT MAJOR DEPRESSION WITHOUT PSYCHOTIC FEATURES |[X]MAJOR DEPRESSION, RECURRENT WITHOUT PSYCHOTIC SYMPTOMS
C0270455|T048|87512008|SNOMEDCT_US|MILD MAJOR DEPRESSION|MILD MAJOR DEPRESSION (DISORDER)
C0270455|T048|87512008|SNOMEDCT_US|MAJOR DEPRESSION MILD|MILD MAJOR DEPRESSION (DISORDER)
C0270455|T048|87512008|SNOMEDCT_US|MILD MAJOR DEPRESSION |MILD MAJOR DEPRESSION (DISORDER)
C0270455|T048|87512008|SNOMEDCT_US|MILD MAJOR DEPRESSION |MILD MAJOR DEPRESSION (DISORDER)
C0235136|T048|83458005|SNOMEDCT_US|AGITATED DEPRESSION|AGITATED DEPRESSION (DISORDER)
C0235136|T048|83458005|SNOMEDCT_US|AGITATED DEPRESSION |AGITATED DEPRESSION (DISORDER)
C0235136|T048|83458005|SNOMEDCT_US|AGITATED DEPRESSION |AGITATED DEPRESSION (DISORDER)
C0235136|T048|83458005|SNOMEDCT_US|DEPRESSION AGITATED|AGITATED DEPRESSION (DISORDER)
C0235136|T048|83458005|SNOMEDCT_US|DEPRESSION; AGITATED|AGITATED DEPRESSION (DISORDER)
C0235136|T048|83458005|SNOMEDCT_US|AGITATED; DEPRESSION|AGITATED DEPRESSION (DISORDER)
C0011570|T048|41006004|SNOMEDCT_US|DEPRESSION|DEPRESSION (FINDING)
C0011570|T048|41006004|SNOMEDCT_US|MENTAL DEPRESSION|DEPRESSION (FINDING)
C0011570|T048|41006004|SNOMEDCT_US|DEPRESSION PSYCHIC|DEPRESSION (FINDING)
C0011570|T048|41006004|SNOMEDCT_US|MONOPOLAR DEPRESSION NOS|DEPRESSION (FINDING)
C0011570|T048|41006004|SNOMEDCT_US|DEPRESSION NOS|DEPRESSION (FINDING)
C0011570|T048|41006004|SNOMEDCT_US|[X] DEPRESSION NOS|DEPRESSION (FINDING)
C0011570|T048|41006004|SNOMEDCT_US|DEPRESSION NOS |DEPRESSION (FINDING)
C0011570|T048|41006004|SNOMEDCT_US|DEPRESSION |DEPRESSION (FINDING)
C0011570|T048|41006004|SNOMEDCT_US|[X]DEPRESSION NOS|DEPRESSION (FINDING)
C0011570|T048|41006004|SNOMEDCT_US|DEPRESSION, MENTAL|DEPRESSION (FINDING)
C0011570|T048|41006004|SNOMEDCT_US|DEPRESSION MENTAL|DEPRESSION (FINDING)
C0011570|T048|41006004|SNOMEDCT_US|DEPRESSION; MENTAL|DEPRESSION (FINDING)
C0011570|T048|41006004|SNOMEDCT_US|DEPRESSION; MONOPOLAR|DEPRESSION (FINDING)
C0011570|T048|41006004|SNOMEDCT_US|DEPRESSIVE; STATE|DEPRESSION (FINDING)
C0011570|T048|41006004|SNOMEDCT_US|MENTAL; DEPRESSION|DEPRESSION (FINDING)
C0011570|T048|41006004|SNOMEDCT_US|MONOPOLAR; DEPRESSION|DEPRESSION (FINDING)
C0011570|T048|41006004|SNOMEDCT_US|DEPRESSION, NOS|DEPRESSION (FINDING)
C0011570|T048|41006004|SNOMEDCT_US|DEPRESSIVE STATE NOS|DEPRESSION (FINDING)
C0011570|T048|41006004|SNOMEDCT_US|DISORDER;DEPRESSION|DEPRESSION (FINDING)
C1269683|T048|370143000|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER|MAJOR DEPRESSIVE DISORDER (DISORDER)
C1269683|T048|370143000|SNOMEDCT_US|MAJOR DEPRESSION|MAJOR DEPRESSIVE DISORDER (DISORDER)
C1269683|T048|370143000|SNOMEDCT_US|DISORDER, MAJOR DEPRESSIVE|MAJOR DEPRESSIVE DISORDER (DISORDER)
C1269683|T048|370143000|SNOMEDCT_US|DISORDERS, MAJOR DEPRESSIVE|MAJOR DEPRESSIVE DISORDER (DISORDER)
C1269683|T048|370143000|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDERS|MAJOR DEPRESSIVE DISORDER (DISORDER)
C1269683|T048|370143000|SNOMEDCT_US|MDD|MAJOR DEPRESSIVE DISORDER (DISORDER)
C1269683|T048|370143000|SNOMEDCT_US|DEPRESSIVE DIS MAJOR|MAJOR DEPRESSIVE DISORDER (DISORDER)
C1269683|T048|370143000|SNOMEDCT_US|MAJOR DEPRESSIVE DIS|MAJOR DEPRESSIVE DISORDER (DISORDER)
C1269683|T048|370143000|SNOMEDCT_US|MAJOR DEPRESSION NOS|MAJOR DEPRESSIVE DISORDER (DISORDER)
C1269683|T048|370143000|SNOMEDCT_US|DEPRESSIVE DISORDER, MAJOR [DISEASE/FINDING]|MAJOR DEPRESSIVE DISORDER (DISORDER)
C1269683|T048|370143000|SNOMEDCT_US|DEPRESSIVE DISORDER, MAJOR|MAJOR DEPRESSIVE DISORDER (DISORDER)
C1269683|T048|370143000|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER |MAJOR DEPRESSIVE DISORDER (DISORDER)
C1269683|T048|370143000|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER NOS|MAJOR DEPRESSIVE DISORDER (DISORDER)
C1269683|T048|370143000|SNOMEDCT_US|MAJOR DEPRESSIVE ILLNESS|MAJOR DEPRESSIVE DISORDER (DISORDER)
C1269683|T048|370143000|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER |MAJOR DEPRESSIVE DISORDER (DISORDER)
C1269683|T048|370143000|SNOMEDCT_US|MAJOR DEPRESSION, NOS|MAJOR DEPRESSIVE DISORDER (DISORDER)
C1269683|T048|370143000|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, NOS|MAJOR DEPRESSIVE DISORDER (DISORDER)
C1269683|T048|370143000|SNOMEDCT_US|DEPRESSIVE DISORDERS, MAJOR|MAJOR DEPRESSIVE DISORDER (DISORDER)
C0086132|T048|394924000|SNOMEDCT_US|DEPRESSION, EMOTIONAL|SYMPTOMS OF DEPRESSION
C0086132|T048|394924000|SNOMEDCT_US|DEPRESSIONS, EMOTIONAL|SYMPTOMS OF DEPRESSION
C0086132|T048|394924000|SNOMEDCT_US|SYMPTOMS OF DEPRESSION|SYMPTOMS OF DEPRESSION
C0086132|T048|394924000|SNOMEDCT_US|SYMPTOMS OF DEPRESSION |SYMPTOMS OF DEPRESSION
C0086132|T048|394924000|SNOMEDCT_US|EMOTIONAL DEPRESSION|SYMPTOMS OF DEPRESSION
C2700639|T048|192372006|SNOMEDCT_US|[X] (DEPRESSION: [EPISODE, UNSPECIFIED] OR [NOS (& REACTIVE)] OR [DEPRESSIVE DISORDER NOS] |[X] (DEPRESSION: [EPISODE, UNSPECIFIED] OR [NOS (& REACTIVE)] OR [DEPRESSIVE DISORDER NOS] (DISORDER)
C2700639|T048|192372006|SNOMEDCT_US|[X] (DEPRESSION: [EPISODE, UNSPECIFIED] OR [NOS (& REACTIVE)] OR [DEPRESSIVE DISORDER NOS]|[X] (DEPRESSION: [EPISODE, UNSPECIFIED] OR [NOS (& REACTIVE)] OR [DEPRESSIVE DISORDER NOS] (DISORDER)
C2363919|T048||SNOMEDCT_US|CHILDHOOD DEPRESSION
C0270458|T048|73867007|SNOMEDCT_US|SEVERE MAJOR DEPRESSIVE DISORDER WITH PSYCHOTIC FEATURES|SEVERE MAJOR DEPRESSION WITH PSYCHOTIC FEATURES (DISORDER)
C0270458|T048|73867007|SNOMEDCT_US|MAJOR DEPRESSION SEVERE WITH PSYCHOTIC FEATURES|SEVERE MAJOR DEPRESSION WITH PSYCHOTIC FEATURES (DISORDER)
C0270458|T048|73867007|SNOMEDCT_US|SEVERE MAJOR DEPRESSIVE DISORDER WITH PSYCHOTIC FEATURES |SEVERE MAJOR DEPRESSION WITH PSYCHOTIC FEATURES (DISORDER)
C0270458|T048|73867007|SNOMEDCT_US|SEVERE MAJOR DEPRESSION WITH PSYCHOTIC FEATURES|SEVERE MAJOR DEPRESSION WITH PSYCHOTIC FEATURES (DISORDER)
C0270458|T048|73867007|SNOMEDCT_US|PSYCHOTIC DEPRESSION|SEVERE MAJOR DEPRESSION WITH PSYCHOTIC FEATURES (DISORDER)
C0270458|T048|73867007|SNOMEDCT_US|SEVERE MAJOR DEPRESSION WITH PSYCHOTIC FEATURES |SEVERE MAJOR DEPRESSION WITH PSYCHOTIC FEATURES (DISORDER)
C0270458|T048|73867007|SNOMEDCT_US|SEVERE MAJOR DEPRESSION WITH PSYCHOTIC FEATURES, NOS|SEVERE MAJOR DEPRESSION WITH PSYCHOTIC FEATURES (DISORDER)
C0270458|T048|73867007|SNOMEDCT_US|PSYCHOTIC DEPRESSION, NOS|SEVERE MAJOR DEPRESSION WITH PSYCHOTIC FEATURES (DISORDER)
C0011579|T048|87414006|SNOMEDCT_US|DEPRESSIONS, REACTIVE|REACTIVE DEPRESSION (SITUATIONAL) (DISORDER)
C0011579|T048|87414006|SNOMEDCT_US|REACTIVE DEPRESSIONS|REACTIVE DEPRESSION (SITUATIONAL) (DISORDER)
C0011579|T048|87414006|SNOMEDCT_US|NEUROTIC DEPRESSIVE REACTION|REACTIVE DEPRESSION (SITUATIONAL) (DISORDER)
C0011579|T048|87414006|SNOMEDCT_US|REACTIVE DEPRESSION|REACTIVE DEPRESSION (SITUATIONAL) (DISORDER)
C0011579|T048|87414006|SNOMEDCT_US|REACTIVE DEPRESSION (SITUATIONAL) |REACTIVE DEPRESSION (SITUATIONAL) (DISORDER)
C0011579|T048|87414006|SNOMEDCT_US|REACTIVE DEPRESSION (SITUATIONAL) |REACTIVE DEPRESSION (SITUATIONAL) (DISORDER)
C0011579|T048|87414006|SNOMEDCT_US|DEPRESSION;REACTIVE|REACTIVE DEPRESSION (SITUATIONAL) (DISORDER)
C0011579|T048|87414006|SNOMEDCT_US|REACTIVE DEPRESSION |REACTIVE DEPRESSION (SITUATIONAL) (DISORDER)
C0011579|T048|87414006|SNOMEDCT_US|REACTIVE (NEUROTIC) DEPRESSION|REACTIVE DEPRESSION (SITUATIONAL) (DISORDER)
C0011579|T048|87414006|SNOMEDCT_US|[X] REACTIVE DEPRESSION NOS|REACTIVE DEPRESSION (SITUATIONAL) (DISORDER)
C0011579|T048|87414006|SNOMEDCT_US|[X]PROLONGED SINGLE EPISODE OF REACTIVE DEPRESSION|REACTIVE DEPRESSION (SITUATIONAL) (DISORDER)
C0011579|T048|87414006|SNOMEDCT_US|NEUROTIC DEPRESSION REACTIVE TYPE|REACTIVE DEPRESSION (SITUATIONAL) (DISORDER)
C0011579|T048|87414006|SNOMEDCT_US|DEPRESSIVE REACTION|REACTIVE DEPRESSION (SITUATIONAL) (DISORDER)
C0011579|T048|87414006|SNOMEDCT_US|DEPRESSION REACTIVE|REACTIVE DEPRESSION (SITUATIONAL) (DISORDER)
C0011579|T048|87414006|SNOMEDCT_US|REACTIVE DEPRESSION (SITUATIONAL)|REACTIVE DEPRESSION (SITUATIONAL) (DISORDER)
C0011579|T048|87414006|SNOMEDCT_US|DEPRESSION; REACTIVE|REACTIVE DEPRESSION (SITUATIONAL) (DISORDER)
C0011579|T048|87414006|SNOMEDCT_US|DEPRESSIVE; REACTION|REACTIVE DEPRESSION (SITUATIONAL) (DISORDER)
C0011579|T048|87414006|SNOMEDCT_US|REACTION; DEPRESSIVE|REACTIVE DEPRESSION (SITUATIONAL) (DISORDER)
C0011579|T048|87414006|SNOMEDCT_US|REACTIVE; DEPRESSION|REACTIVE DEPRESSION (SITUATIONAL) (DISORDER)
C0011579|T048|87414006|SNOMEDCT_US|DEPRESSIVE REACTION (NEUROTIC)|REACTIVE DEPRESSION (SITUATIONAL) (DISORDER)
C0011579|T048|87414006|SNOMEDCT_US|DEPRESSION, REACTIVE|REACTIVE DEPRESSION (SITUATIONAL) (DISORDER)
C2362914|T048||SNOMEDCT_US|CLINICAL DEPRESSION
C0013415|T048|78667006|SNOMEDCT_US|DYSTHYMIA|DYSTHYMIA (DISORDER)
C0013415|T048|78667006|SNOMEDCT_US|DYSTHYMIC DISORDER|DYSTHYMIA (DISORDER)
C0013415|T048|78667006|SNOMEDCT_US|DYSTHYMIC DISORDERS|DYSTHYMIA (DISORDER)
C0013415|T048|78667006|SNOMEDCT_US|DISORDER, DYSTHYMIC|DYSTHYMIA (DISORDER)
C0013415|T048|78667006|SNOMEDCT_US|DYSTHYMIC DIS|DYSTHYMIA (DISORDER)
C0013415|T048|78667006|SNOMEDCT_US|DYSTHYMIA |DYSTHYMIA (DISORDER)
C0013415|T048|78667006|SNOMEDCT_US|DYSTHYMIC DISORDER [DISEASE/FINDING]|DYSTHYMIA (DISORDER)
C0013415|T048|78667006|SNOMEDCT_US|DYSTHYMIA |DYSTHYMIA (DISORDER)
C0013415|T048|78667006|SNOMEDCT_US|PERSISTENT DEPRESSIVE DISORDER (DYSTHYMIA) |DYSTHYMIA (DISORDER)
C0013415|T048|78667006|SNOMEDCT_US|PERSISTENT DEPRESSIVE DISORDER (DYSTHYMIA)|DYSTHYMIA (DISORDER)
C0013415|T048|78667006|SNOMEDCT_US|DISORDER; DYSTHYMIC|DYSTHYMIA (DISORDER)
C0013415|T048|78667006|SNOMEDCT_US|DYSTHYMIC; DISORDER|DYSTHYMIA (DISORDER)
C0013415|T048|78667006|SNOMEDCT_US|DYSTHYMIA, NOS|DYSTHYMIA (DISORDER)
C0344315|T048|102895009|SNOMEDCT_US|MOOD DEPRESSION|MOROSE MOOD (FINDING)
C1868594|T048|699184009|SNOMEDCT_US|PERRY SYNDROME|PARKINSONISM WITH ALVEOLAR HYPOVENTILATION AND MENTAL DEPRESSION
C1868594|T048|699184009|SNOMEDCT_US|PARKINSONISM WITH ALVEOLAR HYPOVENTILATION AND MENTAL DEPRESSION|PARKINSONISM WITH ALVEOLAR HYPOVENTILATION AND MENTAL DEPRESSION
C1868594|T048|699184009|SNOMEDCT_US|PERRY SYNDROME |PARKINSONISM WITH ALVEOLAR HYPOVENTILATION AND MENTAL DEPRESSION
C0349217|T048|268706007|SNOMEDCT_US|DEPRESSIVE EPISODE, UNSPECIFIED|[X]DEPRESSIVE EPISODE, UNSPECIFIED (DISORDER)
C0349217|T048|268706007|SNOMEDCT_US|DEPRESSIVE EPISODE|[X]DEPRESSIVE EPISODE, UNSPECIFIED (DISORDER)
C0349217|T048|268706007|SNOMEDCT_US|[X]DEPRESSIVE EPISODE, UNSPECIFIED|[X]DEPRESSIVE EPISODE, UNSPECIFIED (DISORDER)
C0349217|T048|268706007|SNOMEDCT_US|[X]DEPRESSIVE EPISODE, UNSPECIFIED |[X]DEPRESSIVE EPISODE, UNSPECIFIED (DISORDER)
C0349217|T048|268706007|SNOMEDCT_US|DEPRESSIVE; EPISODE|[X]DEPRESSIVE EPISODE, UNSPECIFIED (DISORDER)
C0349217|T048|268706007|SNOMEDCT_US|EPISODE; DEPRESSIVE|[X]DEPRESSIVE EPISODE, UNSPECIFIED (DISORDER)
C0812393|T048||SNOMEDCT_US|DEPRESSION
C0812393|T048||SNOMEDCT_US|SUICIDE
C0812393|T048||SNOMEDCT_US|DEPRESSION AND SUICIDE
C0812393|T048||SNOMEDCT_US|SUICIDE AND DEPRESSION
C0494399|T048|268702009|SNOMEDCT_US|SEVERE DEPRESSIVE EPISODE WITHOUT PSYCHOTIC SYMPTOMS|[X]SEVERE DEPRESSIVE EPISODE WITHOUT PSYCHOTIC SYMPTOMS (DISORDER)
C0494399|T048|268702009|SNOMEDCT_US|[X]SEVERE DEPRESSIVE EPISODE WITHOUT PSYCHOTIC SYMPTOMS|[X]SEVERE DEPRESSIVE EPISODE WITHOUT PSYCHOTIC SYMPTOMS (DISORDER)
C0494399|T048|268702009|SNOMEDCT_US|[X]SEVERE DEPRESSIVE EPISODE WITHOUT PSYCHOTIC SYMPTOMS |[X]SEVERE DEPRESSIVE EPISODE WITHOUT PSYCHOTIC SYMPTOMS (DISORDER)
C0494399|T048|268702009|SNOMEDCT_US|DEPRESSIVE; DISORDER, MAJOR, SINGLE EPISODE, MAJOR (WITHOUT PSYCHOTIC SYMPTOMS)|[X]SEVERE DEPRESSIVE EPISODE WITHOUT PSYCHOTIC SYMPTOMS (DISORDER)
C0494399|T048|268702009|SNOMEDCT_US|DEPRESSIVE; EPISODE, SEVERE (WITHOUT PSYCHOTIC SYMPTOMS)|[X]SEVERE DEPRESSIVE EPISODE WITHOUT PSYCHOTIC SYMPTOMS (DISORDER)
C0494399|T048|268702009|SNOMEDCT_US|DISORDER; DEPRESSIVE, MAJOR, SINGLE EPISODE, MAJOR (WITHOUT PSYCHOTIC SYMPTOMS)|[X]SEVERE DEPRESSIVE EPISODE WITHOUT PSYCHOTIC SYMPTOMS (DISORDER)
C0494399|T048|268702009|SNOMEDCT_US|EPISODE; DEPRESSIVE, SEVERE (WITHOUT PSYCHOTIC SYMPTOMS)|[X]SEVERE DEPRESSIVE EPISODE WITHOUT PSYCHOTIC SYMPTOMS (DISORDER)
C0494400|T048|268704005|SNOMEDCT_US|SEVERE DEPRESSIVE EPISODE WITH PSYCHOTIC SYMPTOMS|[X]SEVERE DEPRESSIVE EPISODE WITH PSYCHOTIC SYMPTOMS (DISORDER)
C0494400|T048|268704005|SNOMEDCT_US|[X]SEVERE DEPRESSIVE EPISODE WITH PSYCHOTIC SYMPTOMS|[X]SEVERE DEPRESSIVE EPISODE WITH PSYCHOTIC SYMPTOMS (DISORDER)
C0494400|T048|268704005|SNOMEDCT_US|[X]SEVERE DEPRESSIVE EPISODE WITH PSYCHOTIC SYMPTOMS |[X]SEVERE DEPRESSIVE EPISODE WITH PSYCHOTIC SYMPTOMS (DISORDER)
C0494400|T048|268704005|SNOMEDCT_US|DEPRESSIVE; DISORDER, MAJOR, SINGLE EPISODE, MAJOR, WITH PSYCHOTIC SYMPTOMS|[X]SEVERE DEPRESSIVE EPISODE WITH PSYCHOTIC SYMPTOMS (DISORDER)
C0494400|T048|268704005|SNOMEDCT_US|DEPRESSIVE; EPISODE, SEVERE, WITH PSYCHOTIC SYMPTOMS|[X]SEVERE DEPRESSIVE EPISODE WITH PSYCHOTIC SYMPTOMS (DISORDER)
C0494400|T048|268704005|SNOMEDCT_US|DISORDER; DEPRESSIVE, MAJOR, SINGLE EPISODE, MAJOR, WITH PSYCHOTIC SYMPTOMS|[X]SEVERE DEPRESSIVE EPISODE WITH PSYCHOTIC SYMPTOMS (DISORDER)
C0494400|T048|268704005|SNOMEDCT_US|EPISODE; DEPRESSIVE, SEVERE, WITH PSYCHOTIC SYMPTOMS|[X]SEVERE DEPRESSIVE EPISODE WITH PSYCHOTIC SYMPTOMS (DISORDER)
C0439020|T048|272022009|SNOMEDCT_US|COMPLAINING OF FEELING DEPRESSED|COMPLAINING OF FEELING DEPRESSED
C0439020|T048|272022009|SNOMEDCT_US|C/O - FEELING DEPRESSED|COMPLAINING OF FEELING DEPRESSED
C0439020|T048|272022009|SNOMEDCT_US|C/O - FEELING DEPRESSED (CONTEXT-DEPENDENT CATEGORY)|COMPLAINING OF FEELING DEPRESSED
C0439020|T048|272022009|SNOMEDCT_US|COMPLAINING OF FEELING DEPRESSED |COMPLAINING OF FEELING DEPRESSED
C0005587|T048|191627008|SNOMEDCT_US|BIPOLAR DEPRESSION|BIPOLAR AFFECTIVE DISORDER, CURRENT EPISODE DEPRESSION (DISORDER)
C0005587|T048|191627008|SNOMEDCT_US|BIPOLAR AFFECTIVE DISORDER, CURRENT EPISODE DEPRESSED |BIPOLAR AFFECTIVE DISORDER, CURRENT EPISODE DEPRESSION (DISORDER)
C0005587|T048|191627008|SNOMEDCT_US|BIPOLAR AFFECTIVE DISORDER, CURRENT EPISODE DEPRESSED|BIPOLAR AFFECTIVE DISORDER, CURRENT EPISODE DEPRESSION (DISORDER)
C0005587|T048|191627008|SNOMEDCT_US|BIPOLAR DISORDER AFFECTIVE, CURRENT EPISODE DEPRESSED|BIPOLAR AFFECTIVE DISORDER, CURRENT EPISODE DEPRESSION (DISORDER)
C0005587|T048|191627008|SNOMEDCT_US|BIPOLAR AFFECTIVE DISORDER, DEPRESSED|BIPOLAR AFFECTIVE DISORDER, CURRENT EPISODE DEPRESSION (DISORDER)
C0005587|T048|191627008|SNOMEDCT_US|BIPOLAR AFFECTIVE DISORDER, CURRENT EPISODE DEPRESSION|BIPOLAR AFFECTIVE DISORDER, CURRENT EPISODE DEPRESSION (DISORDER)
C0005587|T048|191627008|SNOMEDCT_US|MANIC-DEPRESSIVE - NOW DEPRESSED|BIPOLAR AFFECTIVE DISORDER, CURRENT EPISODE DEPRESSION (DISORDER)
C0005587|T048|191627008|SNOMEDCT_US|BIPOLAR AFFECTIVE DISORDER, CURRENT EPISODE DEPRESSION |BIPOLAR AFFECTIVE DISORDER, CURRENT EPISODE DEPRESSION (DISORDER)
C0005587|T048|191627008|SNOMEDCT_US|DEPRESSION, BIPOLAR|BIPOLAR AFFECTIVE DISORDER, CURRENT EPISODE DEPRESSION (DISORDER)
C0025193|T048|35489007|SNOMEDCT_US|MELANCHOLIA|MELANCHOLIA
C0025193|T048|35489007|SNOMEDCT_US|MELANCHOLIAS|MELANCHOLIA
C0025193|T048|35489007|SNOMEDCT_US|MELANCHOLIC DEPRESSION|MELANCHOLIA
C0025193|T048|35489007|SNOMEDCT_US|DEPRESSION WITH MELANCHOLIC FEATURES|MELANCHOLIA
C0025193|T048|35489007|SNOMEDCT_US|MELANCHOLIA, NOS|MELANCHOLIA
C0025193|T048|35489007|SNOMEDCT_US|MELANCHOLIA NOS|MELANCHOLIA
C0282126|T048||SNOMEDCT_US|DEPRESSIONS, NEUROTIC
C0282126|T048||SNOMEDCT_US|NEUROTIC DEPRESSIONS
C0282126|T048||SNOMEDCT_US|NEUROTIC DEPRESSION
C0282126|T048||SNOMEDCT_US|DEPRESSION, NEUROTIC
C0282126|T048||SNOMEDCT_US|DEPRESSION NEUROTIC
C0282126|T048||SNOMEDCT_US|DEPRESSION; NEUROTIC
C0282126|T048||SNOMEDCT_US|DEPRESSIVE; STATE, NEUROTIC
C0282126|T048||SNOMEDCT_US|NEUROTIC; DEPRESSION
C0282126|T048||SNOMEDCT_US|STATE; DEPRESSIVE, NEUROTIC
C0282126|T048||SNOMEDCT_US|NEUROTIC DEPRESSIVE STATE
C0011573|T048|300706003|SNOMEDCT_US|DEPRESSIONS, ENDOGENOUS|ENDOGENOUS DEPRESSION (DISORDER)
C0011573|T048|300706003|SNOMEDCT_US|ENDOGENOUS DEPRESSIONS|ENDOGENOUS DEPRESSION (DISORDER)
C0011573|T048|300706003|SNOMEDCT_US|ENDOGENOUS DEPRESSION|ENDOGENOUS DEPRESSION (DISORDER)
C0011573|T048|300706003|SNOMEDCT_US|DEPRESSION;ENDOGENOUS|ENDOGENOUS DEPRESSION (DISORDER)
C0011573|T048|300706003|SNOMEDCT_US|ENDOGENOUS DEPRESSION |ENDOGENOUS DEPRESSION (DISORDER)
C0011573|T048|300706003|SNOMEDCT_US|DEPRESSION ENDOGENOUS|ENDOGENOUS DEPRESSION (DISORDER)
C0011573|T048|300706003|SNOMEDCT_US|ENDOGENOUS DEPRESSION |ENDOGENOUS DEPRESSION (DISORDER)
C0011573|T048|300706003|SNOMEDCT_US|DEPRESSION; ENDOGENOUS|ENDOGENOUS DEPRESSION (DISORDER)
C0011573|T048|300706003|SNOMEDCT_US|ENDOGENOUS; DEPRESSION|ENDOGENOUS DEPRESSION (DISORDER)
C0011573|T048|300706003|SNOMEDCT_US|ENDOGENOUS DEPRESSION [AMBIGUOUS]|ENDOGENOUS DEPRESSION (DISORDER)
C0011573|T048|300706003|SNOMEDCT_US|DEPRESSION, ENDOGENOUS|ENDOGENOUS DEPRESSION (DISORDER)
C0520669|T048|42925002|SNOMEDCT_US|SINGLE EPISODE MAJOR DEPRESSION WITH ATYPICAL FEATURES |MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE WITH ATYPICAL FEATURES (DISORDER)
C0520669|T048|42925002|SNOMEDCT_US|SINGLE EPISODE MAJOR DEPRESSION WITH ATYPICAL FEATURES|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE WITH ATYPICAL FEATURES (DISORDER)
C0520669|T048|42925002|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE WITH ATYPICAL FEATURES|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE WITH ATYPICAL FEATURES (DISORDER)
C0520669|T048|42925002|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE WITH ATYPICAL FEATURES |MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE WITH ATYPICAL FEATURES (DISORDER)
C0154413|T048|192378005|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, RECURRENT EPISODE, SEVERE DEGREE, SPECIFIED AS WITH PSYCHOTIC BEHAVIOR|[X]RECURRENT SEVERE EPISODES OF PSYCHOGENIC DEPRESSIVE PSYCHOSIS
C0154413|T048|192378005|SNOMEDCT_US|RECURRENT DEPRESSIVE DISORDER, CURRENT EPISODE SEVERE WITH PSYCHOTIC SYMPTOMS|[X]RECURRENT SEVERE EPISODES OF PSYCHOGENIC DEPRESSIVE PSYCHOSIS
C0154413|T048|192378005|SNOMEDCT_US|SEVERE RECURRENT MAJOR DEPRESSION WITH PSYCHOTIC FEATURES |[X]RECURRENT SEVERE EPISODES OF PSYCHOGENIC DEPRESSIVE PSYCHOSIS
C0154413|T048|192378005|SNOMEDCT_US|RECURRENT MAJOR DEPRESSION WITH PSYCHOTIC FEATURES |[X]RECURRENT SEVERE EPISODES OF PSYCHOGENIC DEPRESSIVE PSYCHOSIS
C0154413|T048|192378005|SNOMEDCT_US|RECURRENT MAJOR DEPRESSION WITH PSYCHOTIC FEATURES|[X]RECURRENT SEVERE EPISODES OF PSYCHOGENIC DEPRESSIVE PSYCHOSIS
C0154413|T048|192378005|SNOMEDCT_US|SEVERE RECURRENT MAJOR DEPRESSION WITH PSYCHOTIC FEATURES|[X]RECURRENT SEVERE EPISODES OF PSYCHOGENIC DEPRESSIVE PSYCHOSIS
C0154413|T048|192378005|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, RECURRENT EPISODE, SEVERE DEGREE, SPECIFIED AS WITH PSYCHOTIC BEHAVIOUR|[X]RECURRENT SEVERE EPISODES OF PSYCHOGENIC DEPRESSIVE PSYCHOSIS
C0154413|T048|192378005|SNOMEDCT_US|REC DEPR PSYCH-PSYCHOTIC|[X]RECURRENT SEVERE EPISODES OF PSYCHOGENIC DEPRESSIVE PSYCHOSIS
C0154413|T048|192378005|SNOMEDCT_US|MAJOR DEPRESSIVE AFFECTIVE DISORDER, RECURRENT EPISODE, SEVERE, SPECIFIED AS WITH PSYCHOTIC BEHAVIOR|[X]RECURRENT SEVERE EPISODES OF PSYCHOGENIC DEPRESSIVE PSYCHOSIS
C0154413|T048|192378005|SNOMEDCT_US|[X]RECURRENT SEVERE EPISODES OF PSYCHOTIC DEPRESSION|[X]RECURRENT SEVERE EPISODES OF PSYCHOGENIC DEPRESSIVE PSYCHOSIS
C0154413|T048|192378005|SNOMEDCT_US|[X]RECURRENT DEPRESSIVE DISORDER, CURRENT EPISODE SEVERE WITH PSYCHOTIC SYMPTOMS|[X]RECURRENT SEVERE EPISODES OF PSYCHOGENIC DEPRESSIVE PSYCHOSIS
C0154413|T048|192378005|SNOMEDCT_US|[X]RECURRENT DEPRESSIVE DISORDER, CURRENT EPISODE SEVERE WITH PSYCHOTIC SYMPTOMS |[X]RECURRENT SEVERE EPISODES OF PSYCHOGENIC DEPRESSIVE PSYCHOSIS
C0154413|T048|192378005|SNOMEDCT_US|[X]RECURRENT SEVERE EPISODES OF PSYCHOGENIC DEPRESSIVE PSYCHOSIS|[X]RECURRENT SEVERE EPISODES OF PSYCHOGENIC DEPRESSIVE PSYCHOSIS
C0154413|T048|192378005|SNOMEDCT_US|[X]RECURRENT SEVERE EPISODES OF MAJOR DEPRESSION WITH PSYCHOTIC SYMPTOMS|[X]RECURRENT SEVERE EPISODES OF PSYCHOGENIC DEPRESSIVE PSYCHOSIS
C0154413|T048|192378005|SNOMEDCT_US|SEVERE RECURRENT MAJOR DEPRESSION WITH PSYCHOSIS|[X]RECURRENT SEVERE EPISODES OF PSYCHOGENIC DEPRESSIVE PSYCHOSIS
C0154413|T048|192378005|SNOMEDCT_US|SEVERE RECURRENT MAJOR DEPRESSION WITH PSYCHOSIS |[X]RECURRENT SEVERE EPISODES OF PSYCHOGENIC DEPRESSIVE PSYCHOSIS
C0154413|T048|192378005|SNOMEDCT_US|MAJOR DEPRESSION RECURRENT SEVERE WITH PSYCHOSIS|[X]RECURRENT SEVERE EPISODES OF PSYCHOGENIC DEPRESSIVE PSYCHOSIS
C0154413|T048|192378005|SNOMEDCT_US|SEVERE RECURRENT MAJOR DEPRESSION WITH PSYCHOTIC FEATURES |[X]RECURRENT SEVERE EPISODES OF PSYCHOGENIC DEPRESSIVE PSYCHOSIS
C0024517|T048|36923009|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE, UNSPECIFIED DEGREE|MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0024517|T048|36923009|SNOMEDCT_US|SINGLE EPISODE MAJOR DEPRESSION |MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0024517|T048|36923009|SNOMEDCT_US|SINGLE EPISODE MAJOR DEPRESSION|MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0024517|T048|36923009|SNOMEDCT_US|DEPRESS PSYCHOSIS-UNSPEC|MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0024517|T048|36923009|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE, UNSPECIFIED|MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0024517|T048|36923009|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE|MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0024517|T048|36923009|SNOMEDCT_US|SINGLE EPISODE OF MAJOR DEPRESSION|MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0024517|T048|36923009|SNOMEDCT_US|MAJOR DEPRESSIVE AFFECTIVE DISORDER, SINGLE EPISODE, UNSPECIFIED|MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0024517|T048|36923009|SNOMEDCT_US|SINGLE MAJOR DEPRESSIVE EPISODE|MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0024517|T048|36923009|SNOMEDCT_US|SINGLE MAJOR DEPRESSIVE EPISODE, UNSPECIFIED|MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0024517|T048|36923009|SNOMEDCT_US|SINGLE MAJOR DEPRESSIVE EPISODE NOS |MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0024517|T048|36923009|SNOMEDCT_US|SINGLE MAJOR DEPRESSIVE EPISODE |MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0024517|T048|36923009|SNOMEDCT_US|SINGLE MAJOR DEPRESSIVE EPISODE NOS|MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0024517|T048|36923009|SNOMEDCT_US|SINGLE MAJOR DEPRESSIVE EPISODE, UNSPECIFIED |MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0024517|T048|36923009|SNOMEDCT_US|MAJOR DEPRESSION, SINGLE EPISODE |MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0024517|T048|36923009|SNOMEDCT_US|MAJOR DEPRESSION, SINGLE EPISODE|MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0024517|T048|36923009|SNOMEDCT_US|DEPRESSIVE; EPISODE, MAJOR|MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0024517|T048|36923009|SNOMEDCT_US|MAJOR DEPRESSION, SINGLE EPISODE, NOS|MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0024517|T048|36923009|SNOMEDCT_US|SINGLE EPISODE OF MAJOR DEPRESSIVE DISORDER|MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0024517|T048|36923009|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER; SINGLE EPISODE|MAJOR DEPRESSION, SINGLE EPISODE (DISORDER)
C0302874|T048||SNOMEDCT_US|DEPRESSIVE PERSONALITY DISORDER
C0302874|T048||SNOMEDCT_US|PERSONALITY;DEPRESSIVE
C0302874|T048||SNOMEDCT_US|DEPRESSIVE PERSONALITY
C0302874|T048||SNOMEDCT_US|DEPRESSIVE; PERSONALITY DISORDER
C0302874|T048||SNOMEDCT_US|PERSONALITY DISORDER; DEPRESSIVE
C0154405|T048|76441001|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE, SEVERE DEGREE, WITHOUT MENTION OF PSYCHOTIC BEHAVIOR|SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITHOUT PSYCHOTIC FEATURES (DISORDER)
C0154405|T048|76441001|SNOMEDCT_US|SEVERE SINGLE EPISODE MAJOR DEPRESSION WITHOUT PSYCHOTIC FEATURES |SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITHOUT PSYCHOTIC FEATURES (DISORDER)
C0154405|T048|76441001|SNOMEDCT_US|SEVERE SINGLE EPISODE MAJOR DEPRESSION WITHOUT PSYCHOTIC FEATURES|SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITHOUT PSYCHOTIC FEATURES (DISORDER)
C0154405|T048|76441001|SNOMEDCT_US|DEPRESS PSYCHOSIS-SEVERE|SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITHOUT PSYCHOTIC FEATURES (DISORDER)
C0154405|T048|76441001|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE, SEVERE WITHOUT PSYCHOTIC FEATURES|SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITHOUT PSYCHOTIC FEATURES (DISORDER)
C0154405|T048|76441001|SNOMEDCT_US|MAJOR DEPRESSV DISORD, SINGLE EPSD, SEV W/O PSYCH FEATURES|SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITHOUT PSYCHOTIC FEATURES (DISORDER)
C0154405|T048|76441001|SNOMEDCT_US|MAJOR DEPRESSIVE AFFECTIVE DISORDER, SINGLE EPISODE, SEVERE, WITHOUT MENTION OF PSYCHOTIC BEHAVIOR|SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITHOUT PSYCHOTIC FEATURES (DISORDER)
C0154405|T048|76441001|SNOMEDCT_US|SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITHOUT PSYCHOTIC FEATURES|SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITHOUT PSYCHOTIC FEATURES (DISORDER)
C0154405|T048|76441001|SNOMEDCT_US|SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITHOUT PSYCHOTIC FEATURES |SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITHOUT PSYCHOTIC FEATURES (DISORDER)
C0154406|T048|430852001|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE, SEVERE DEGREE, SPECIFIED AS WITH PSYCHOTIC BEHAVIOR|SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITH PSYCHOTIC FEATURES (DISORDER)
C0154406|T048|430852001|SNOMEDCT_US|SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITH PSYCHOTIC FEATURES |SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITH PSYCHOTIC FEATURES (DISORDER)
C0154406|T048|430852001|SNOMEDCT_US|SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITH PSYCHOTIC FEATURES|SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITH PSYCHOTIC FEATURES (DISORDER)
C0154406|T048|430852001|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE, SEVERE WITH PSYCHOTIC FEATURES|SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITH PSYCHOTIC FEATURES (DISORDER)
C0154406|T048|430852001|SNOMEDCT_US|SEVERE SINGLE EPISODE MAJOR DEPRESSION WITH PSYCHOTIC FEATURES|SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITH PSYCHOTIC FEATURES (DISORDER)
C0154406|T048|430852001|SNOMEDCT_US|SEVERE SINGLE EPISODE MAJOR DEPRESSION WITH PSYCHOTIC FEATURES |SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITH PSYCHOTIC FEATURES (DISORDER)
C0154406|T048|430852001|SNOMEDCT_US|DEPR PSYCHOS-SEV W PSYCH|SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITH PSYCHOTIC FEATURES (DISORDER)
C0154406|T048|430852001|SNOMEDCT_US|MAJOR DEPRESSV DISORD, SINGLE EPSD, SEVERE W PSYCH FEATURES|SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITH PSYCHOTIC FEATURES (DISORDER)
C0154406|T048|430852001|SNOMEDCT_US|MAJOR DEPRESSIVE AFFECTIVE DISORDER, SINGLE EPISODE, SEVERE, SPECIFIED AS WITH PSYCHOTIC BEHAVIOR|SEVERE MAJOR DEPRESSION, SINGLE EPISODE, WITH PSYCHOTIC FEATURES (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, RECURRENT EPISODE, UNSPECIFIED DEGREE|RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|RECURRENT MAJOR DEPRESSION|RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|RECURRENT MAJOR DEPRESSION |RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|RECURR DEPR PSYCHOS-UNSP|RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, RECURRENT, UNSPECIFIED|RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, RECURRENT|RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|RECURRENT EPISODES OF MAJOR DEPRESSION|RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|MAJOR DEPRESSIVE AFFECTIVE DISORDER, RECURRENT EPISODE, UNSPECIFIED|RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|RECURRENT MAJOR DEPRESSIVE EPISODE NOS |RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED |RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED|RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|RECURRENT MAJOR DEPRESSIVE EPISODE|RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|RECURRENT MAJOR DEPRESSIVE EPISODE NOS|RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|RECURRENT MAJOR DEPRESSIVE EPISODES|RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|RECURRENT MAJOR DEPRESSIVE EPISODES |RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|MAJOR DEPRESSION RECURRENT EPISODES|RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, RECURRENT EPISODE|RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|RECURRENT MAJOR DEPRESSION |RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|RECURRENT MAJOR DEPRESSIVE DISORDER|RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|RECURRENT MAJOR DEPRESSIVE EPISODES |RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|RECURRENT MAJOR DEPRESSION, NOS|RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|RECURRENT MAJOR DEPRESSIVE DISORDER, NOS|RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154409|T048|191609005|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER; RECURRENT EPISODE|RECURRENT MAJOR DEPRESSIVE EPISODES, UNSPECIFIED (DISORDER)
C0154437|T048|191659001|SNOMEDCT_US|ATYPICAL DEPRESSIVE DISORDER |ATYPICAL DEPRESSIVE DISORDER (DISORDER)
C0154437|T048|191659001|SNOMEDCT_US|ATYPICAL DEPRESSIVE DISORDER|ATYPICAL DEPRESSIVE DISORDER (DISORDER)
C0154437|T048|191659001|SNOMEDCT_US|ATYPICAL DEPRESSIVE DIS|ATYPICAL DEPRESSIVE DISORDER (DISORDER)
C0154437|T048|191659001|SNOMEDCT_US|ATYPICAL DEPRESSION|ATYPICAL DEPRESSIVE DISORDER (DISORDER)
C0154437|T048|191659001|SNOMEDCT_US|ATYPICAL DEPRESSIVE DISORDER |ATYPICAL DEPRESSIVE DISORDER (DISORDER)
C0154437|T048|191659001|SNOMEDCT_US|[X]ATYPICAL DEPRESSION|ATYPICAL DEPRESSIVE DISORDER (DISORDER)
C0154437|T048|191659001|SNOMEDCT_US|ATYPICAL; DEPRESSION|ATYPICAL DEPRESSIVE DISORDER (DISORDER)
C0154437|T048|191659001|SNOMEDCT_US|DEPRESSION; ATYPICAL|ATYPICAL DEPRESSIVE DISORDER (DISORDER)
C0338893|T048|191614009|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, RECURRENT EPISODE, IN PARTIAL OR UNSPECIFIED REMISSION|RECURRENT MAJOR DEPRESSIVE EPISODES, IN PARTIAL OR UNSPECIFIED REMISSION
C0338893|T048|191614009|SNOMEDCT_US|RECUR DEPR PSYC-PART REM|RECURRENT MAJOR DEPRESSIVE EPISODES, IN PARTIAL OR UNSPECIFIED REMISSION
C0338893|T048|191614009|SNOMEDCT_US|MAJOR DEPRESSIVE AFFECTIVE DISORDER, RECURRENT EPISODE, IN PARTIAL OR UNSPECIFIED REMISSION|RECURRENT MAJOR DEPRESSIVE EPISODES, IN PARTIAL OR UNSPECIFIED REMISSION
C0338893|T048|191614009|SNOMEDCT_US|RECURRENT MAJOR DEPRESSIVE EPISODES, IN PARTIAL OR UNSPECIFIED REMISSION|RECURRENT MAJOR DEPRESSIVE EPISODES, IN PARTIAL OR UNSPECIFIED REMISSION
C0338893|T048|191614009|SNOMEDCT_US|RECURRENT MAJOR DEPRESSIVE EPISODES, IN PARTIAL OR UNSPECIFIED REMISSION |RECURRENT MAJOR DEPRESSIVE EPISODES, IN PARTIAL OR UNSPECIFIED REMISSION
C0085159|T048|192374007|SNOMEDCT_US|AFFECTIVE DISORDER, SEASONAL|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|AFFECTIVE DISORDERS, SEASONAL|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|DISORDER, SEASONAL AFFECTIVE|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|DISORDER, SEASONAL MOOD|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|DISORDERS, SEASONAL AFFECTIVE|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|DISORDERS, SEASONAL MOOD|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|MOOD DISORDER, SEASONAL|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|MOOD DISORDERS, SEASONAL|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|SEASONAL AFFECTIVE DISORDER|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|SEASONAL MOOD DISORDERS|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|SAD|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|SEASONAL AFFECTIVE DIS|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|SEASONAL DEPRESSION|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|DEPRESSION IN A SEASONAL PATTERN|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|SEASONAL DEPRESSION |[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|DEPRESSION SEASONAL PATTERN |[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|DEPRESSION SEASONAL PATTERN|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|SEASONAL PATTERN DEPRESSION|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|SEASONAL AFFECTIVE DISORDERS|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|SEASONAL MOOD DISORDER|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|SEASONAL AFFECTIVE DISORDER [DISEASE/FINDING]|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|[X]SEASONAL DEPRESSIVE DISORDER|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|SEASONAL AFFECTIVE DISORDER |[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|[X] SEASONAL DEPRESSIVE DISORDER|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|[X]SAD - SEASONAL AFFECTIVE DISORDER|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|SEASONAL AFFECTIVE DISORDER |[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|SAD - SEASONAL AFFECTIVE DISORDER|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|DEPRESSION; SEASONAL|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0085159|T048|192374007|SNOMEDCT_US|SEASONAL; DEPRESSION|[X]SAD - SEASONAL AFFECTIVE DISORDER
C0011581|T048|192372006|SNOMEDCT_US|DEPRESSIVE NEUROSIS|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|DEPRESSIVE DISORDERS|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|DEPRESSIVE DISORDER|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|DEPRESSIVE NEUROSES|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|DISORDER, DEPRESSIVE|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|DISORDERS, DEPRESSIVE|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|NEUROSES, DEPRESSIVE|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|DEPRESSIVE DIS|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|DEPRESSION|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|DEPRESSION |[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|DEPRESSIVE DISORDER NOS|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|DEPRESSIVE DISORDER [DISEASE/FINDING]|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|NEUROSIS, DEPRESSIVE|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|MOOD DISORDER OF DEPRESSED TYPE|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|[X]DEPRESSIVE DISORDER NOS|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|MOOD DISORDER OF DEPRESSED TYPE |[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|MOOD DISORDER WITH DEPRESSIVE FEATURE|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|-- DEPRESSION|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|DEPRESSIVE ILLNESS|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|DEPRESSIVE DISORDER |[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|DEPRESSION; BEHAVIORAL DISORDER|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|DEPRESSIVE; DISORDER|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|DEPRESSIVE; NEUROSIS|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|DISORDER; DEPRESSIVE|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|NEUROSIS; DEPRESSIVE|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|DEPRESSIVE DISORDER, NOS|[X]DEPRESSIVE DISORDER NOS
C0011581|T048|192372006|SNOMEDCT_US|DISORDER;DEPRESSIVE|[X]DEPRESSIVE DISORDER NOS
C0362037|T048|82218004|SNOMEDCT_US|DEPRESSION POSTOPERATIVE|POSTOPERATIVE DEPRESSION (DISORDER)
C0362037|T048|82218004|SNOMEDCT_US|[D]POSTOPERATIVE DEPRESSION|POSTOPERATIVE DEPRESSION (DISORDER)
C0362037|T048|82218004|SNOMEDCT_US|POSTOPERATIVE DEPRESSION |POSTOPERATIVE DEPRESSION (DISORDER)
C0362037|T048|82218004|SNOMEDCT_US|POSTOPERATIVE DEPRESSION|POSTOPERATIVE DEPRESSION (DISORDER)
C0362037|T048|82218004|SNOMEDCT_US|POSTOPERATIVE DEPRESSION |POSTOPERATIVE DEPRESSION (DISORDER)
C0362037|T048|82218004|SNOMEDCT_US|POSTOPERATIVE DEPRESSION, NOS|POSTOPERATIVE DEPRESSION (DISORDER)
C0221745|T048||SNOMEDCT_US|DEPRESSION SUICIDAL
C0221745|T048||SNOMEDCT_US|SUICIDAL DEPRESSION
C0520665|T048|84788008|SNOMEDCT_US|MENOPAUSAL DEPRESSION|MENOPAUSAL DEPRESSION (DISORDER)
C0520665|T048|84788008|SNOMEDCT_US|DEPRESSION MENOPAUSAL|MENOPAUSAL DEPRESSION (DISORDER)
C0520665|T048|84788008|SNOMEDCT_US|DEPRESSION MENOPAUSAL |MENOPAUSAL DEPRESSION (DISORDER)
C0520665|T048|84788008|SNOMEDCT_US|POSTMENOPAUSAL DEPRESSION|MENOPAUSAL DEPRESSION (DISORDER)
C0520665|T048|84788008|SNOMEDCT_US|DEPRESSION POSTMENOPAUSAL|MENOPAUSAL DEPRESSION (DISORDER)
C0520665|T048|84788008|SNOMEDCT_US|MENOPAUSAL DEPRESSION |MENOPAUSAL DEPRESSION (DISORDER)
C0520665|T048|84788008|SNOMEDCT_US|DEPRESSION; MENOPAUSAL|MENOPAUSAL DEPRESSION (DISORDER)
C0520665|T048|84788008|SNOMEDCT_US|MENOPAUSAL; DEPRESSION|MENOPAUSAL DEPRESSION (DISORDER)
C0520665|T048|84788008|SNOMEDCT_US|MENOPAUSAL DEPRESSION, NOS|MENOPAUSAL DEPRESSION (DISORDER)
C0520665|T048|84788008|SNOMEDCT_US|POSTMENOPAUSAL DEPRESSION, NOS|MENOPAUSAL DEPRESSION (DISORDER)
C3665457|T048|442057004|SNOMEDCT_US|CHRONIC DEPRESSIVE PERSONALITY DISORDER |CHRONIC DEPRESSIVE PERSONALITY DISORDER (DISORDER)
C3665457|T048|442057004|SNOMEDCT_US|CHRONIC DEPRESSIVE PERSONALITY DISORDER|CHRONIC DEPRESSIVE PERSONALITY DISORDER (DISORDER)
C3665457|T048|442057004|SNOMEDCT_US|CHRONIC DEPRESSIVE PERSONALITY DISORDER |CHRONIC DEPRESSIVE PERSONALITY DISORDER (DISORDER)
C3665457|T048|442057004|SNOMEDCT_US|CHR DEPRESSIVE PERSON|CHRONIC DEPRESSIVE PERSONALITY DISORDER (DISORDER)
C3665457|T048|442057004|SNOMEDCT_US|CHRONIC DEPRESSIVE DISORDER|CHRONIC DEPRESSIVE PERSONALITY DISORDER (DISORDER)
C0871610|T048||SNOMEDCT_US|WINTER DEPRESSION
C0871610|T048||SNOMEDCT_US|DEPRESSION MORE IN WINTER 
C0871610|T048||SNOMEDCT_US|DEPRESSION MORE IN WINTER
C2165514|T048||SNOMEDCT_US|SUMMER DEPRESSION
C2165514|T048||SNOMEDCT_US|DEPRESSION MORE IN SUMMER 
C2165514|T048||SNOMEDCT_US|DEPRESSION MORE IN SUMMER
C2165515|T048||SNOMEDCT_US|DEPRESSION PRECEDED BY HIGH ACTIVITY LEVEL
C2165515|T048||SNOMEDCT_US|DEPRESSION PRECEDED BY HIGH ACTIVITY LEVEL 
C2165509|T048||SNOMEDCT_US|DEPRESSION ACCOMPANIED BY EATING MORE
C2165509|T048||SNOMEDCT_US|DEPRESSION ACCOMPANIED BY EATING MORE 
C2165508|T048||SNOMEDCT_US|DEPRESSION ACCOMPANIED BY EATING LESS
C2165508|T048||SNOMEDCT_US|DEPRESSION ACCOMPANIED BY EATING LESS 
C2165511|T048||SNOMEDCT_US|DEPRESSION ACCOMPANIED BY SLEEPING MORE 
C2165511|T048||SNOMEDCT_US|DEPRESSION ACCOMPANIED BY SLEEPING MORE
C2165510|T048||SNOMEDCT_US|DEPRESSION ACCOMPANIED BY SLEEPING LESS 
C2165510|T048||SNOMEDCT_US|DEPRESSION ACCOMPANIED BY SLEEPING LESS
C2165507|T048||SNOMEDCT_US|DEPRESSION ACCOMPANIED BY PERSISTENT WORRY 
C2165507|T048||SNOMEDCT_US|DEPRESSION ACCOMPANIED BY PERSISTENT WORRY
C2165518|T048||SNOMEDCT_US|DEPRESSION RELIEVED BY GOOD NEWS
C2165518|T048||SNOMEDCT_US|DEPRESSION RELIEVED BY GOOD NEWS 
C2165519|T048||SNOMEDCT_US|DEPRESSION RELIEVED BY MEDICATION 
C2165519|T048||SNOMEDCT_US|DEPRESSION RELIEVED BY MEDICATION
C2165517|T048||SNOMEDCT_US|DEPRESSION RELIEVED BY COUNSELING 
C2165517|T048||SNOMEDCT_US|DEPRESSION RELIEVED BY COUNSELING
C2165520|T048||SNOMEDCT_US|DEPRESSION SEASONAL PATTERN WITH FEW NONSEASONAL OCCURRENCES
C2165520|T048||SNOMEDCT_US|DEPRESSION SEASONAL PATTERN W/ FEW NONSEASONAL OCCURRENCES
C2165520|T048||SNOMEDCT_US|DEPRESSION SEASONAL PATTERN WITH FEW NONSEASONAL OCCURRENCES 
C2165520|T048||SNOMEDCT_US|SEASONAL DEPRESSION WITH FEW NONSEASONAL OCCURRENCES
C0338908|T048|192402009|SNOMEDCT_US|MIXED ANXIETY AND DEPRESSIVE DISORDER|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|DEPRESSION WITH ANXIETY|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|DEPRESSION WITH ANXIETY |[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|ANXIETY/DEPRESSION|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|ANXIETY WITH DEPRESSION|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|MIXED ANXIETY AND DEPRESSIVE DISORDER |[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|ANXIETY DEPRESSION|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|ANXIOUS DEPRESSION|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|MIXED ANXIETY & DEPRESSIVE|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|DEPRESSION; ANXIETY|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|DISORDER; MIXED, ANXIETY AND DEPRESSIVE|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|MIXED; DISORDER, ANXIETY AND DEPRESSIVE|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|ANXIETY; DEPRESSION|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C2063289|T048||SNOMEDCT_US|CHRONIC MAJOR DEPRESSION 
C2063289|T048||SNOMEDCT_US|CHRONIC MAJOR DEPRESSION
C2063866|T048||SNOMEDCT_US|RESISTANT DEPRESSION, TREATMENT
C2063866|T048||SNOMEDCT_US|TREATMENT-RESISTANT DEPRESSIVE DISORDERS
C2063866|T048||SNOMEDCT_US|THERAPY-RESISTANT DEPRESSIONS
C2063866|T048||SNOMEDCT_US|DEPRESSIONS, REFRACTORY
C2063866|T048||SNOMEDCT_US|THERAPY RESISTANT DEPRESSION
C2063866|T048||SNOMEDCT_US|DEPRESSION, REFRACTORY
C2063866|T048||SNOMEDCT_US|DEPRESSIVE DISORDER, TREATMENT-RESISTANT
C2063866|T048||SNOMEDCT_US|DISORDERS, TREATMENT-RESISTANT DEPRESSIVE
C2063866|T048||SNOMEDCT_US|DEPRESSION, TREATMENT RESISTANT
C2063866|T048||SNOMEDCT_US|DEPRESSIONS, TREATMENT RESISTANT
C2063866|T048||SNOMEDCT_US|TREATMENT RESISTANT DEPRESSIONS
C2063866|T048||SNOMEDCT_US|DEPRESSIVE DISORDER, TREATMENT RESISTANT
C2063866|T048||SNOMEDCT_US|DEPRESSIVE DISORDERS, TREATMENT-RESISTANT
C2063866|T048||SNOMEDCT_US|DISORDER, TREATMENT-RESISTANT DEPRESSIVE
C2063866|T048||SNOMEDCT_US|TREATMENT-RESISTANT DEPRESSIVE DISORDER
C2063866|T048||SNOMEDCT_US|DEPRESSION, THERAPY-RESISTANT
C2063866|T048||SNOMEDCT_US|DEPRESSIONS, THERAPY-RESISTANT
C2063866|T048||SNOMEDCT_US|RESISTANT DEPRESSIONS, TREATMENT
C2063866|T048||SNOMEDCT_US|REFRACTORY DEPRESSIONS
C2063866|T048||SNOMEDCT_US|REFRACTORY DEPRESSION
C2063866|T048||SNOMEDCT_US|THERAPY-RESISTANT DEPRESSION
C2063866|T048||SNOMEDCT_US|TREATMENT RESISTANT DEPRESSION
C2063866|T048||SNOMEDCT_US|DEPRESSIVE DISORDER, TREATMENT-RESISTANT [DISEASE/FINDING]
C2063866|T048||SNOMEDCT_US|TREATMENT-REFRACTORY DEPRESSION 
C2063866|T048||SNOMEDCT_US|TREATMENT-REFRACTORY DEPRESSION
C2938940|T048||SNOMEDCT_US|POST STROKE DEPRESSION
C0086133|T048||SNOMEDCT_US|DEPRESSIVE SYNDROMES
C0086133|T048||SNOMEDCT_US|SYNDROME, DEPRESSIVE
C0086133|T048||SNOMEDCT_US|SYNDROMES, DEPRESSIVE
C0086133|T048||SNOMEDCT_US|DEPRESSIVE SYNDROME
C0349712|T048|40568001|SNOMEDCT_US|[X]RECURRENT BRIEF DEPRESSIVE EPISODES|RECURRENT BRIEF DEPRESSIVE DISORDER (DISORDER)
C0349712|T048|40568001|SNOMEDCT_US|[X] RECURRENT BRIEF DEPRESSIVE EPISODES|RECURRENT BRIEF DEPRESSIVE DISORDER (DISORDER)
C0349712|T048|40568001|SNOMEDCT_US|DEPRESSION RECURRENT BRIEF|RECURRENT BRIEF DEPRESSIVE DISORDER (DISORDER)
C0349712|T048|40568001|SNOMEDCT_US|RECURRENT BRIEF DEPRESSIVE DISORDER |RECURRENT BRIEF DEPRESSIVE DISORDER (DISORDER)
C0349712|T048|40568001|SNOMEDCT_US|RECURRENT BRIEF DEPRESSIVE DISORDER|RECURRENT BRIEF DEPRESSIVE DISORDER (DISORDER)
C0349712|T048|40568001|SNOMEDCT_US|RECURRENT BRIEF DEPRESSIVE DISORDER |RECURRENT BRIEF DEPRESSIVE DISORDER (DISORDER)
C0349712|T048|40568001|SNOMEDCT_US|DISORDER; RECURRENT BRIEF DEPRESSIVE|RECURRENT BRIEF DEPRESSIVE DISORDER (DISORDER)
C0349712|T048|40568001|SNOMEDCT_US|RECURRENT BRIEF DEPRESSIVE; DISORDER|RECURRENT BRIEF DEPRESSIVE DISORDER (DISORDER)
C0270461|T048|42810003|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, IN REMISSION (MDD)|MAJOR DEPRESSION IN REMISSION (DISORDER)
C0270461|T048|42810003|SNOMEDCT_US|MDD IN REMISSION|MAJOR DEPRESSION IN REMISSION (DISORDER)
C0270461|T048|42810003|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER REMISSION|MAJOR DEPRESSION IN REMISSION (DISORDER)
C0270461|T048|42810003|SNOMEDCT_US|MAJOR DEPRESSION, IN REMISSION|MAJOR DEPRESSION IN REMISSION (DISORDER)
C0270461|T048|42810003|SNOMEDCT_US|MAJOR DEPRESSION - IN REMISSION|MAJOR DEPRESSION IN REMISSION (DISORDER)
C0270461|T048|42810003|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER - IN REMISSION|MAJOR DEPRESSION IN REMISSION (DISORDER)
C0270461|T048|42810003|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, IN REMISSION |MAJOR DEPRESSION IN REMISSION (DISORDER)
C0270461|T048|42810003|SNOMEDCT_US|MAJOR DEPRESSIVE DISORDER, IN REMISSION|MAJOR DEPRESSION IN REMISSION (DISORDER)
C0270461|T048|42810003|SNOMEDCT_US|MAJOR DEPRESSION IN REMISSION |MAJOR DEPRESSION IN REMISSION (DISORDER)
C0270461|T048|42810003|SNOMEDCT_US|MAJOR DEPRESSION IN REMISSION|MAJOR DEPRESSION IN REMISSION (DISORDER)
C0270461|T048|42810003|SNOMEDCT_US|MAJOR DEPRESSION IN REMISSION, NOS|MAJOR DEPRESSION IN REMISSION (DISORDER)
C0270457|T048|75084000|SNOMEDCT_US|MAJOR DEPRESSION SEVERE WITHOUT PSYCHOTIC FEATURES|SEVERE MAJOR DEPRESSION WITHOUT PSYCHOTIC FEATURES (DISORDER)
C0270457|T048|75084000|SNOMEDCT_US|SEVERE MAJOR DEPRESSIVE DISORDER WITHOUT PSYCHOTIC FEATURES |SEVERE MAJOR DEPRESSION WITHOUT PSYCHOTIC FEATURES (DISORDER)
C0270457|T048|75084000|SNOMEDCT_US|SEVERE MAJOR DEPRESSIVE DISORDER WITHOUT PSYCHOTIC FEATURES|SEVERE MAJOR DEPRESSION WITHOUT PSYCHOTIC FEATURES (DISORDER)
C0270457|T048|75084000|SNOMEDCT_US|SEVERE MAJOR DEPRESSION WITHOUT PSYCHOTIC FEATURES|SEVERE MAJOR DEPRESSION WITHOUT PSYCHOTIC FEATURES (DISORDER)
C0270457|T048|75084000|SNOMEDCT_US|SEVERE MAJOR DEPRESSION WITHOUT PSYCHOTIC FEATURES |SEVERE MAJOR DEPRESSION WITHOUT PSYCHOTIC FEATURES (DISORDER)
C0270456|T048|832007|SNOMEDCT_US|MAJOR DEPRESSION MODERATE|MODERATE MAJOR DEPRESSION (DISORDER)
C0270456|T048|832007|SNOMEDCT_US|MODERATE MAJOR DEPRESSION |MODERATE MAJOR DEPRESSION (DISORDER)
C0270456|T048|832007|SNOMEDCT_US|MODERATE MAJOR DEPRESSION|MODERATE MAJOR DEPRESSION (DISORDER)
C0270456|T048|832007|SNOMEDCT_US|MODERATE MAJOR DEPRESSION |MODERATE MAJOR DEPRESSION (DISORDER)
C1282644|T048|320751009|SNOMEDCT_US|MAJOR DEPRESSION, MELANCHOLIC TYPE |MAJOR DEPRESSION, MELANCHOLIC TYPE (DISORDER)
C1282644|T048|320751009|SNOMEDCT_US|MAJOR DEPRESSION, MELANCHOLIC TYPE|MAJOR DEPRESSION, MELANCHOLIC TYPE (DISORDER)
C1282644|T048|320751009|SNOMEDCT_US|MAJOR DEPRESSION MELANCHOLIC TYPE|MAJOR DEPRESSION, MELANCHOLIC TYPE (DISORDER)
C1282644|T048|320751009|SNOMEDCT_US|MAJOR DEPRESSION, MELANCHOLIC TYPE |MAJOR DEPRESSION, MELANCHOLIC TYPE (DISORDER)
C1282644|T048|320751009|SNOMEDCT_US|MAJOR DEPRESSION, MELANCHOLIC TYPE  [AMBIGUOUS]|MAJOR DEPRESSION, MELANCHOLIC TYPE (DISORDER)
C0349218|T048|268707003|SNOMEDCT_US|RECURRENT DEPRESSIVE DISORDER|[X]RECURRENT DEPRESSIVE DISORDER (FINDING)
C0349218|T048|268707003|SNOMEDCT_US|RECURRENT DEPRESSIVE DISORDER, UNSPECIFIED|[X]RECURRENT DEPRESSIVE DISORDER (FINDING)
C0349218|T048|268707003|SNOMEDCT_US|[X]RECURRENT DEPRESSIVE DISORDER, UNSPECIFIED|[X]RECURRENT DEPRESSIVE DISORDER (FINDING)
C0349218|T048|268707003|SNOMEDCT_US|[X]RECURRENT DEPRESSIVE DISORDER|[X]RECURRENT DEPRESSIVE DISORDER (FINDING)
C0349218|T048|268707003|SNOMEDCT_US|[X] RECURRENT EPISODES OF REACTIVE DEPRESSION|[X]RECURRENT DEPRESSIVE DISORDER (FINDING)
C0349218|T048|268707003|SNOMEDCT_US|[X] RECURRENT EPISODES OF DEPRESSIVE REACTION|[X]RECURRENT DEPRESSIVE DISORDER (FINDING)
C0349218|T048|268707003|SNOMEDCT_US|[X]RECURRENT DEPRESSIVE DISORDER, UNSPECIFIED |[X]RECURRENT DEPRESSIVE DISORDER (FINDING)
C0349218|T048|268707003|SNOMEDCT_US|[X]RECURRENT DEPRESSIVE DISORDER |[X]RECURRENT DEPRESSIVE DISORDER (FINDING)
C0349218|T048|268707003|SNOMEDCT_US|[X]RECURRENT EPISODES OF REACTIVE DEPRESSION|[X]RECURRENT DEPRESSIVE DISORDER (FINDING)
C0349218|T048|268707003|SNOMEDCT_US|[X]RECURRENT EPISODES OF DEPRESSIVE REACTION|[X]RECURRENT DEPRESSIVE DISORDER (FINDING)
C0349218|T048|268707003|SNOMEDCT_US|[X]RECURRENT DEPRESSIVE DISORDER |[X]RECURRENT DEPRESSIVE DISORDER (FINDING)
C0701819|T048|319768000|SNOMEDCT_US|RECURRENT MAJOR DEPRESSION WITH MELANCHOLIA|RECURRENT MAJOR DEPRESSIVE DISORDER WITH MELANCHOLIC FEATURES (DISORDER)
C0701819|T048|319768000|SNOMEDCT_US|RECURRENT MAJOR DEPRESSION WITH MELANCHOLIA |RECURRENT MAJOR DEPRESSIVE DISORDER WITH MELANCHOLIC FEATURES (DISORDER)
C0701819|T048|319768000|SNOMEDCT_US|RECURRENT MAJOR DEPRESSIVE DISORDER WITH MELANCHOLIC FEATURES|RECURRENT MAJOR DEPRESSIVE DISORDER WITH MELANCHOLIC FEATURES (DISORDER)
C0701819|T048|319768000|SNOMEDCT_US|RECURRENT MAJOR DEPRESSIVE DISORDER WITH MELANCHOLIC FEATURES |RECURRENT MAJOR DEPRESSIVE DISORDER WITH MELANCHOLIC FEATURES (DISORDER)
C0012706|T048|192078003|SNOMEDCT_US|DEPRESSIVE DISORDER NEC IN SNOMEDCT|DEPRESSIVE DISORDER NEC (DISORDER)
C0012706|T048|192078003|SNOMEDCT_US|DEPRESSIVE DISORDER NEC|DEPRESSIVE DISORDER NEC (DISORDER)
C0012706|T048|192078003|SNOMEDCT_US|DEPRESSIVE DISORDER NEC |DEPRESSIVE DISORDER NEC (DISORDER)
C0588006|T048|390717003|SNOMEDCT_US|MILD DEPRESSION|MILD DEPRESSION -RETIRED-
C0588006|T048|390717003|SNOMEDCT_US|MILD DEPRESSION |MILD DEPRESSION -RETIRED-
C0588006|T048|390717003|SNOMEDCT_US|DEPRESSION MILD|MILD DEPRESSION -RETIRED-
C0588006|T048|390717003|SNOMEDCT_US|MILD DEPRESSION |MILD DEPRESSION -RETIRED-
C0588006|T048|390717003|SNOMEDCT_US|MILD DEPRESSION -RETIRED-|MILD DEPRESSION -RETIRED-
C0338808|T048|231485007|SNOMEDCT_US|POST-SCHIZOPHRENIC DEPRESSION|POST-SCHIZOPHRENIC DEPRESSION (DISORDER)
C0338808|T048|231485007|SNOMEDCT_US|POST-SCHIZOPHRENIC DEPRESSION |POST-SCHIZOPHRENIC DEPRESSION (DISORDER)
C0338808|T048|231485007|SNOMEDCT_US|POST-SCHIZOPHRENIC DEPRESSION |POST-SCHIZOPHRENIC DEPRESSION (DISORDER)
C0338808|T048|231485007|SNOMEDCT_US|DEPRESSION POST-SCHIZOPHRENIC|POST-SCHIZOPHRENIC DEPRESSION (DISORDER)
C0338808|T048|231485007|SNOMEDCT_US|DEPRESSION; POST-SCHIZOPHRENIC|POST-SCHIZOPHRENIC DEPRESSION (DISORDER)
C0338808|T048|231485007|SNOMEDCT_US|POST-SCHIZOPHRENIC; DEPRESSION|POST-SCHIZOPHRENIC DEPRESSION (DISORDER)
C0338808|T048|231485007|SNOMEDCT_US|POSTPSYCHOTIC DEPRESSION; SCHIZOPHRENIC|POST-SCHIZOPHRENIC DEPRESSION (DISORDER)
C0338808|T048|231485007|SNOMEDCT_US|POSTSCHIZOPHRENIC DEPRESSION|POST-SCHIZOPHRENIC DEPRESSION (DISORDER)
C0338808|T048|231485007|SNOMEDCT_US|SCHIZOPHRENIA; POSTPSYCHOTIC DEPRESSION|POST-SCHIZOPHRENIC DEPRESSION (DISORDER)
C0588007|T048|310496002|SNOMEDCT_US|MODERATE DEPRESSION |MODERATE DEPRESSION (DISORDER)
C0588007|T048|310496002|SNOMEDCT_US|MODERATE DEPRESSION|MODERATE DEPRESSION (DISORDER)
C0588007|T048|310496002|SNOMEDCT_US|MODERATE DEPRESSION |MODERATE DEPRESSION (DISORDER)
C0588007|T048|310496002|SNOMEDCT_US|DEPRESSION MODERATE|MODERATE DEPRESSION (DISORDER)
C0270488|T048|79842004|SNOMEDCT_US|DEPRESSION STUPOROUS|STUPOROUS DEPRESSION (DISORDER)
C0270488|T048|79842004|SNOMEDCT_US|STUPOROUS DEPRESSION|STUPOROUS DEPRESSION (DISORDER)
C0270488|T048|79842004|SNOMEDCT_US|STUPOROUS DEPRESSION |STUPOROUS DEPRESSION (DISORDER)
C0270488|T048|79842004|SNOMEDCT_US|STUPOROUS DEPRESSION |STUPOROUS DEPRESSION (DISORDER)
C0588008|T048|310497006|SNOMEDCT_US|SEVERE DEPRESSION|SEVERE DEPRESSION (DISORDER)
C0588008|T048|310497006|SNOMEDCT_US|SEVERE DEPRESSION |SEVERE DEPRESSION (DISORDER)
C0588008|T048|310497006|SNOMEDCT_US|SEVERE DEPRESSION |SEVERE DEPRESSION (DISORDER)
C0588008|T048|310497006|SNOMEDCT_US|DEPRESSION SEVERE|SEVERE DEPRESSION (DISORDER)
C0588008|T048|310497006|SNOMEDCT_US|DEPRESSION; SEVERE|SEVERE DEPRESSION (DISORDER)
C0588008|T048|310497006|SNOMEDCT_US|SEVERE; DEPRESSION|SEVERE DEPRESSION (DISORDER)
C0581391|T048|192080009|SNOMEDCT_US|DEPRESSION CHRONIC|CHRONIC DEPRESSION (DISORDER)
C0581391|T048|192080009|SNOMEDCT_US|CHRONIC DEPRESSION|CHRONIC DEPRESSION (DISORDER)
C0581391|T048|192080009|SNOMEDCT_US|CHRONIC DEPRESSION |CHRONIC DEPRESSION (DISORDER)
C0581391|T048|192080009|SNOMEDCT_US|CHRONIC DEPRESSION |CHRONIC DEPRESSION (DISORDER)
C0581391|T048|192080009|SNOMEDCT_US|CHRONIC DEPRESSION |CHRONIC DEPRESSION (DISORDER)
C0520675|T048|48589009|SNOMEDCT_US|MINOR DEPRESSIVE DISORDER |MINOR DEPRESSIVE DISORDER (DISORDER)
C0520675|T048|48589009|SNOMEDCT_US|MINOR DEPRESSIVE DISORDER|MINOR DEPRESSIVE DISORDER (DISORDER)
C0520675|T048|48589009|SNOMEDCT_US|DEPRESSION MINOR|MINOR DEPRESSIVE DISORDER (DISORDER)
C0520675|T048|48589009|SNOMEDCT_US|MINOR DEPRESSIVE DISORDER |MINOR DEPRESSIVE DISORDER (DISORDER)
C0338897|T048|231500002|SNOMEDCT_US|MASKED DEPRESSION|MASKED DEPRESSION (DISORDER)
C0338897|T048|231500002|SNOMEDCT_US|MASKED DEPRESSION |MASKED DEPRESSION (DISORDER)
C0338897|T048|231500002|SNOMEDCT_US|DEPRESSION MASKED|MASKED DEPRESSION (DISORDER)
C0338897|T048|231500002|SNOMEDCT_US|MASKED DEPRESSION |MASKED DEPRESSION (DISORDER)
C0338897|T048|231500002|SNOMEDCT_US|DEPRESSION; MASKED|MASKED DEPRESSION (DISORDER)
C0338897|T048|231500002|SNOMEDCT_US|MASKED; DEPRESSION|MASKED DEPRESSION (DISORDER)
C0221480|T048|191616006|SNOMEDCT_US|DEPRESSION RECURRENT|RECURRENT DEPRESSION (DISORDER)
C0221480|T048|191616006|SNOMEDCT_US|RECURRENT DEPRESSION|RECURRENT DEPRESSION (DISORDER)
C0221480|T048|191616006|SNOMEDCT_US|RECURRENT DEPRESSION |RECURRENT DEPRESSION (DISORDER)
C0221480|T048|191616006|SNOMEDCT_US|RECURRENT DEPRESSION |RECURRENT DEPRESSION (DISORDER)
C0221480|T048|191616006|SNOMEDCT_US|RECURRENT DEPRESSION |RECURRENT DEPRESSION (DISORDER)
C3697979|T048|698957003|SNOMEDCT_US|DEPRESSIVE DISORDER IN REMISSION|DEPRESSIVE DISORDER IN REMISSION (DISORDER)
C3697979|T048|698957003|SNOMEDCT_US|DEPRESSIVE DISORDER IN REMISSION |DEPRESSIVE DISORDER IN REMISSION (DISORDER)
C3838728|T048|10835871000119104|SNOMEDCT_US|DEPRESSIVE DISORDER IN MOTHER COMPLICATING CHILDBIRTH |DEPRESSION IN CHILDBIRTH
C3838728|T048|10835871000119104|SNOMEDCT_US|DEPRESSIVE DISORDER IN MOTHER COMPLICATING CHILDBIRTH|DEPRESSION IN CHILDBIRTH
C3838728|T048|10835871000119104|SNOMEDCT_US|DEPRESSION IN CHILDBIRTH|DEPRESSION IN CHILDBIRTH
C0520676|T048|596004|SNOMEDCT_US|PREMENSTRUAL DYSPHORIC DISORDER|PREMENSTRUAL DYSPHORIC DISORDER (DISORDER)
C0520676|T048|596004|SNOMEDCT_US|PMDD|PREMENSTRUAL DYSPHORIC DISORDER (DISORDER)
C0520676|T048|596004|SNOMEDCT_US|PREMENSTRUAL DYSPHORIC DISORDER |PREMENSTRUAL DYSPHORIC DISORDER (DISORDER)
C0520676|T048|596004|SNOMEDCT_US|PREMENSTRUAL DISORDER|PREMENSTRUAL DYSPHORIC DISORDER (DISORDER)
C0520676|T048|596004|SNOMEDCT_US|DYSPHORIC DISORDER, PREMENSTRUAL|PREMENSTRUAL DYSPHORIC DISORDER (DISORDER)
C0520676|T048|596004|SNOMEDCT_US|SYNDROME, PREMENSTRUAL DYSPHORIC|PREMENSTRUAL DYSPHORIC DISORDER (DISORDER)
C0520676|T048|596004|SNOMEDCT_US|DISORDER, PREMENSTRUAL DYSPHORIC|PREMENSTRUAL DYSPHORIC DISORDER (DISORDER)
C0520676|T048|596004|SNOMEDCT_US|PREMENSTRUAL DYSPHORIC DISORDER [DISEASE/FINDING]|PREMENSTRUAL DYSPHORIC DISORDER (DISORDER)
C0520676|T048|596004|SNOMEDCT_US|PREMENSTRUAL DYSPHORIC SYNDROME|PREMENSTRUAL DYSPHORIC DISORDER (DISORDER)
C0520676|T048|596004|SNOMEDCT_US|PREMENSTRUAL DYSPHORIC DISORDER |PREMENSTRUAL DYSPHORIC DISORDER (DISORDER)
C3825465|T048||SNOMEDCT_US|DEPRESSION IN INFANTS
C3825452|T048||SNOMEDCT_US|DEPRESSION IN OLD AGE
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR DISORDERS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC DEPRESSIVE ILLNESS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR AFFECTIVE PSYCHOSIS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR DISORDER|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC DEPRESSIVE PSYCHOSIS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESSIVE PSYCHOSES|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|PSYCHOSES, BIPOLAR AFFECTIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|PSYCHOSES, MANIC DEPRESSIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|PSYCHOSIS, BIPOLAR AFFECTIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|PSYCHOSIS, MANIC DEPRESSIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR AFFECTIVE DISORDER|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|DISORDER, BIPOLAR|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESSIVE PSYCHOSIS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR AFFECTIVE DISORDER, UNSPECIFIED|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR DIS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESSION|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC DEPRESSIVE DISORDER|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BPAD|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|UNSPECIFIED BIPOLAR DISORDER|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|UNSPECIFIED BIPOLAR DISORDER |DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR DISORDER NOT OTHERWISE SPECIFIED|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC DEPRESSIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR DISORDER NOS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESSIVE REACTION|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESSIVE ILLNESS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR DISORDER, UNSPECIFIED|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|AFFECTIVE PSYCHOSIS, BIPOLAR|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR DISORDER [DISEASE/FINDING]|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|PSYCHOSES, MANIC-DEPRESSIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|PSYCHOSIS, MANIC-DEPRESSIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|DISORDER;BIPOLAR|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|DEPRESSION;MANIC|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|PSYCHOSIS;MANIC DEPRESSIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BI-POLAR DISORDER|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR DISORDER |DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|UNSPECIFIED BIPOLAR AFFECTIVE DISORDER|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|DEPRESSIVE-MANIC PSYCH.|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|UNSPECIFIED BIPOLAR AFFECTIVE DISORDER |DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|UNSPECIFIED BIPOLAR AFFECTIVE DISORDER, UNSPECIFIED|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|[X]BIPOLAR AFFECTIVE DISORDER, UNSPECIFIED|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|[X]BIPOLAR AFFECTIVE DISORDER, UNSPECIFIED |DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|UNSPECIFIED BIPOLAR AFFECTIVE DISORDER, UNSPECIFIED |DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|UNSPECIFIED BIPOLAR AFFECTIVE DISORDER, NOS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESS.PSYCHOSES|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|UNSPECIFIED BIPOLAR AFFECTIVE DISORDER, NOS |DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC DEPRESSION|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC DEPRESSIVE REACTION|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|REACTION MANIC-DEPRESSIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|PSYCHOSIS MANIC-DEPRESSIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MDI - MANIC-DEPRESSIVE ILLNESS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR; DISORDER, AFFECTIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR; DISORDER|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|DISORDER; BIPOLAR, AFFECTIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|DISORDER; BIPOLAR|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESSIVE; DISORDER|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESSIVE; PSYCHOSIS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESSIVE; SYNDROME|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|PSYCHOSIS; MANIC-DEPRESSIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|SYNDROME; MANIC-DEPRESSIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR DISORDER, NOS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR MOOD DISORDER|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESSIVE REACTION NOS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESSIVE SYNDROME NOS|DEPRESSIVE-MANIC PSYCH.
C4065471|T048|715924009|SNOMEDCT_US|DISRUPTIVE MOOD DYSREGULATION DISORDER |DISRUPTIVE MOOD DYSREGULATION DISORDER (DISORDER)
C4065471|T048|715924009|SNOMEDCT_US|DEPRESSION DISRUPTIVE MOOD DYSREGULATION DISORDER|DISRUPTIVE MOOD DYSREGULATION DISORDER (DISORDER)
C4065471|T048|715924009|SNOMEDCT_US|DISRUPTIVE MOOD DYSREGULATION DISORDER|DISRUPTIVE MOOD DYSREGULATION DISORDER (DISORDER)
C1386135|T048|712823008|SNOMEDCT_US|ACUTE DEPRESSION|ACUTE DEPRESSION (DISORDER)
C1386135|T048|712823008|SNOMEDCT_US|ACUTE DEPRESSION |ACUTE DEPRESSION (DISORDER)
C1386135|T048|712823008|SNOMEDCT_US|DEPRESSION; ACUTE|ACUTE DEPRESSION (DISORDER)
C1386135|T048|712823008|SNOMEDCT_US|ACUTE; DEPRESSION|ACUTE DEPRESSION (DISORDER)
C4074822|T048|94631000119100|SNOMEDCT_US|DEPRESSIVE DISORDER IN MOTHER COMPLICATING PREGNANCY|DEPRESSIVE DISORDER IN MOTHER COMPLICATING PREGNANCY (DISORDER)
C4074822|T048|94631000119100|SNOMEDCT_US|DEPRESSIVE DISORDER IN MOTHER COMPLICATING PREGNANCY |DEPRESSIVE DISORDER IN MOTHER COMPLICATING PREGNANCY (DISORDER)
C1282921|T048|357705009|SNOMEDCT_US|COTARD'S SYNDROME|COTARD'S SYNDROME (DISORDER)
C1282921|T048|357705009|SNOMEDCT_US|COTARD SYNDROME|COTARD'S SYNDROME (DISORDER)
C1282921|T048|357705009|SNOMEDCT_US|COTARD SYNDROME |COTARD'S SYNDROME (DISORDER)
C1282921|T048|357705009|SNOMEDCT_US|COTARD'S SYNDROME |COTARD'S SYNDROME (DISORDER)
C1282921|T048|357705009|SNOMEDCT_US|COTARD'S SYNDROME |COTARD'S SYNDROME (DISORDER)
C1282921|T048|357705009|SNOMEDCT_US|COTARD|COTARD'S SYNDROME (DISORDER)
C0011580|T048|191676002|SNOMEDCT_US|REACTIVE PSYCHOTIC DEPRESSION|REACTIVE DEPRESSIVE PSYCHOSIS (DISORDER)
C0011580|T048|191676002|SNOMEDCT_US|REACTIVE DEPRESSIVE PSYCHOSIS|REACTIVE DEPRESSIVE PSYCHOSIS (DISORDER)
C0011580|T048|191676002|SNOMEDCT_US|REACTIVE DEPRESSIVE PSYCHOSIS |REACTIVE DEPRESSIVE PSYCHOSIS (DISORDER)
C0011580|T048|191676002|SNOMEDCT_US|DEPRESSIVE TYPE PSYCHOSIS (MDD) REACTIVE|REACTIVE DEPRESSIVE PSYCHOSIS (DISORDER)
C0011580|T048|191676002|SNOMEDCT_US|PSYCHOTIC REACTIVE DEPRESSION|REACTIVE DEPRESSIVE PSYCHOSIS (DISORDER)
C0011580|T048|191676002|SNOMEDCT_US|REACTIVE DEPRESSIVE PSYCHOSIS |REACTIVE DEPRESSIVE PSYCHOSIS (DISORDER)
C0011580|T048|191676002|SNOMEDCT_US|DEPRESSION; REACTIVE, PSYCHOTIC|REACTIVE DEPRESSIVE PSYCHOSIS (DISORDER)
C0011580|T048|191676002|SNOMEDCT_US|DEPRESSIVE; REACTION, PSYCHOTIC|REACTIVE DEPRESSIVE PSYCHOSIS (DISORDER)
C0011580|T048|191676002|SNOMEDCT_US|PSYCHOSIS; DEPRESSIVE, REACTIVE|REACTIVE DEPRESSIVE PSYCHOSIS (DISORDER)
C0011580|T048|191676002|SNOMEDCT_US|PSYCHOSIS; REACTIVE, DEPRESSIVE|REACTIVE DEPRESSIVE PSYCHOSIS (DISORDER)
C0011580|T048|191676002|SNOMEDCT_US|REACTION; DEPRESSIVE, PSYCHOTIC|REACTIVE DEPRESSIVE PSYCHOSIS (DISORDER)
C0011580|T048|191676002|SNOMEDCT_US|REACTIVE; DEPRESSION, PSYCHOTIC|REACTIVE DEPRESSIVE PSYCHOSIS (DISORDER)
C0011580|T048|191676002|SNOMEDCT_US|PSYCHOTIC DEPRESSIVE REACTION|REACTIVE DEPRESSIVE PSYCHOSIS (DISORDER)
C0011580|T048|191676002|SNOMEDCT_US|DEPRESSION, REACTIVE, PSYCHOTIC|REACTIVE DEPRESSIVE PSYCHOSIS (DISORDER)
C0270497|T048|84760002|SNOMEDCT_US|SCHIZOAFFECTIVE DISORDER, DEPRESSIVE TYPE|SCHIZOAFFECTIVE DISORDER, DEPRESSIVE TYPE (DISORDER)
C0270497|T048|84760002|SNOMEDCT_US|SCHIZOAFFECTIVE DISORDER DEPRESSIVE TYPE|SCHIZOAFFECTIVE DISORDER, DEPRESSIVE TYPE (DISORDER)
C0270497|T048|84760002|SNOMEDCT_US|SCHIZOPHRENIFORM PSYCHOSIS, DEPRESSIVE TYPE|SCHIZOAFFECTIVE DISORDER, DEPRESSIVE TYPE (DISORDER)
C0270497|T048|84760002|SNOMEDCT_US|SCHIZOAFFECTIVE DISORDER, DEPRESSIVE TYPE |SCHIZOAFFECTIVE DISORDER, DEPRESSIVE TYPE (DISORDER)
C0270497|T048|84760002|SNOMEDCT_US|DISORDER; SCHIZOAFFECTIVE, DEPRESSIVE TYPE|SCHIZOAFFECTIVE DISORDER, DEPRESSIVE TYPE (DISORDER)
C0270497|T048|84760002|SNOMEDCT_US|PSYCHOSIS; SCHIZOPHRENIFORM, DEPRESSIVE TYPE|SCHIZOAFFECTIVE DISORDER, DEPRESSIVE TYPE (DISORDER)
C0339017|T048|231542000|SNOMEDCT_US|DEPRESSIVE CONDUCT DISORDER|DEPRESSIVE CONDUCT DISORDER (DISORDER)
C0339017|T048|231542000|SNOMEDCT_US|DEPRESSIVE CONDUCT DISORDER |DEPRESSIVE CONDUCT DISORDER (DISORDER)
C0339017|T048|231542000|SNOMEDCT_US|DEPRESSIVE CONDUCT DISORDER |DEPRESSIVE CONDUCT DISORDER (DISORDER)
C0339017|T048|231542000|SNOMEDCT_US|BEHAVIORAL DISORDER; DEPRESSIVE|DEPRESSIVE CONDUCT DISORDER (DISORDER)
C0339017|T048|231542000|SNOMEDCT_US|DEPRESSIVE; BEHAVIORAL DISORDER|DEPRESSIVE CONDUCT DISORDER (DISORDER)
C0349216|T048|268705006|SNOMEDCT_US|OTHER DEPRESSIVE EPISODES|[X]OTHER DEPRESSIVE EPISODES (DISORDER)
C0349216|T048|268705006|SNOMEDCT_US|[X]OTHER DEPRESSIVE EPISODES |[X]OTHER DEPRESSIVE EPISODES (DISORDER)
C0349216|T048|268705006|SNOMEDCT_US|[X]OTHER DEPRESSIVE EPISODES|[X]OTHER DEPRESSIVE EPISODES (DISORDER)
C0556016|T048|310465006|SNOMEDCT_US|[X]SINGLE EPISODE AGITATED DEPRESSION WITHOUT PSYCHOTIC SYMPTOMS|[X] SINGLE EPISODE AGITATED DEPRESSION WITHOUT PSYCHOTIC SYMPTOMS (DISORDER)
C0556016|T048|310465006|SNOMEDCT_US|[X] SINGLE EPISODE AGITATED DEPRESSION WITHOUT PSYCHOTIC SYMPTOMS |[X] SINGLE EPISODE AGITATED DEPRESSION WITHOUT PSYCHOTIC SYMPTOMS (DISORDER)
C0556016|T048|310465006|SNOMEDCT_US|[X] SINGLE EPISODE AGITATED DEPRESSION WITHOUT PSYCHOTIC SYMPTOMS|[X] SINGLE EPISODE AGITATED DEPRESSION WITHOUT PSYCHOTIC SYMPTOMS (DISORDER)
C0556018|T048|310462009|SNOMEDCT_US|[X] MANIC-DEPRESSIVE PSYCHOSIS, DEPRESSED TYPE WITHOUT PSYCHOTIC SYMPTOMS|[X] MANIC-DEPRESSIVE PSYCHOSIS, DEPRESSED TYPE WITHOUT PSYCHOTIC SYMPTOMS (DISORDER)
C0556018|T048|310462009|SNOMEDCT_US|[X]MANIC-DEPRESSIVE PSYCHOSIS, DEPRESSED TYPE WITHOUT PSYCHOTIC SYMPTOMS|[X] MANIC-DEPRESSIVE PSYCHOSIS, DEPRESSED TYPE WITHOUT PSYCHOTIC SYMPTOMS (DISORDER)
C0556018|T048|310462009|SNOMEDCT_US|[X] MANIC-DEPRESSIVE PSYCHOSIS, DEPRESSED TYPE WITHOUT PSYCHOTIC SYMPTOMS |[X] MANIC-DEPRESSIVE PSYCHOSIS, DEPRESSED TYPE WITHOUT PSYCHOTIC SYMPTOMS (DISORDER)
C0556018|T048|310462009|SNOMEDCT_US|PSYCHOSIS; MANIC-DEPRESSIVE, DEPRESSED TYPE (WITHOUT PSYCHOTIC SYMPTOMS)|[X] MANIC-DEPRESSIVE PSYCHOSIS, DEPRESSED TYPE WITHOUT PSYCHOTIC SYMPTOMS (DISORDER)
C0556017|T048|192369004|SNOMEDCT_US|[X]SINGLE EPISODE VITAL DEPRESSION WITHOUT PSYCHOTIC SYMPTOMS|[X]SINGLE EPISODE VITAL DEPRESSION WITHOUT PSYCHOTIC SYMPTOMS
C0556017|T048|192369004|SNOMEDCT_US|[X] SINGLE EPISODE MAJOR DEPRESSION WITHOUT PSYCHOTIC SYMPTOMS|[X]SINGLE EPISODE VITAL DEPRESSION WITHOUT PSYCHOTIC SYMPTOMS
C0556017|T048|192369004|SNOMEDCT_US|[X]SINGLE EPISODE MAJOR DEPRESSION WITHOUT PSYCHOTIC SYMPTOMS|[X]SINGLE EPISODE VITAL DEPRESSION WITHOUT PSYCHOTIC SYMPTOMS
C0556017|T048|192369004|SNOMEDCT_US|[X] SINGLE EPISODE MAJOR DEPRESSION WITHOUT PSYCHOTIC SYMPTOMS |[X]SINGLE EPISODE VITAL DEPRESSION WITHOUT PSYCHOTIC SYMPTOMS
C1579931|T048|139480000|SNOMEDCT_US|DEPRESSION|DEPRESSED - SYMPTOM
C3874774|T048|704678007|SNOMEDCT_US|DEPRESSED MOOD WITH POSTPARTUM ONSET |DEPRESSED MOOD IN POSTPARTUM PERIOD
C3874774|T048|704678007|SNOMEDCT_US|DEPRESSED MOOD WITH POSTPARTUM ONSET|DEPRESSED MOOD IN POSTPARTUM PERIOD
C3874774|T048|704678007|SNOMEDCT_US|DEPRESSED MOOD IN POSTPARTUM PERIOD|DEPRESSED MOOD IN POSTPARTUM PERIOD
C3874774|T048|704678007|SNOMEDCT_US|DEPRESSED MOOD DURING POST PARTUM PERIOD|DEPRESSED MOOD IN POSTPARTUM PERIOD
C3698286|T048|142001000119106|SNOMEDCT_US|DEPRESSED MOOD IN ALZHEIMER DISEASE|ALZHEIMERS DEMENTIA WITH DEPRESSED MOOD
C3698286|T048|142001000119106|SNOMEDCT_US|DEPRESSED MOOD IN ALZHEIMER'S DISEASE |ALZHEIMERS DEMENTIA WITH DEPRESSED MOOD
C3698286|T048|142001000119106|SNOMEDCT_US|ALZHEIMERS DEMENTIA WITH DEPRESSED MOOD|ALZHEIMERS DEMENTIA WITH DEPRESSED MOOD
C3698286|T048|142001000119106|SNOMEDCT_US|DEPRESSED MOOD IN ALZHEIMER'S DISEASE|ALZHEIMERS DEMENTIA WITH DEPRESSED MOOD
C2165504|T048||SNOMEDCT_US|DEPRESSED, BUT UNLIKE PREVIOUS GRIEVING FOR A DEATH OR LOSS
C2165504|T048||SNOMEDCT_US|DEPRESSED, BUT UNLIKE PREVIOUS GRIEVING FOR A DEATH OR LOSS (PHYSICAL FINDING)
C3836786|T048||SNOMEDCT_US|MOOD DEPRESSED POSTPARTUM (PHYSICAL FINDING)
C3836786|T048||SNOMEDCT_US|MOOD DEPRESSED POSTPARTUM
C0150041|T048|389335004|SNOMEDCT_US|WILL INCLUDE THIS AS IT'S A BIT MORE CLOSELY CORRELATED WITH DEPRESSION|LOSS OF HOPE FOR THE FUTURE (FINDING)
C0150041|T048|389335004|SNOMEDCT_US|FEELINGS OF HOPELESSNESS|LOSS OF HOPE FOR THE FUTURE (FINDING)
C0150041|T048|389335004|SNOMEDCT_US|FEELING OF HOPELESSNESS|LOSS OF HOPE FOR THE FUTURE (FINDING)
C0150041|T048|389335004|SNOMEDCT_US|HOPELESS|LOSS OF HOPE FOR THE FUTURE (FINDING)
C0150041|T048|389335004|SNOMEDCT_US|RNDX HOPELESSNESS |LOSS OF HOPE FOR THE FUTURE (FINDING)
C0150041|T048|389335004|SNOMEDCT_US|RNDX HOPELESSNESS|LOSS OF HOPE FOR THE FUTURE (FINDING)
C0150041|T048|389335004|SNOMEDCT_US|FEELING;HOPELESS|LOSS OF HOPE FOR THE FUTURE (FINDING)
C0150041|T048|389335004|SNOMEDCT_US|LOSS OF HOPE FOR THE FUTURE|LOSS OF HOPE FOR THE FUTURE (FINDING)
C0150041|T048|389335004|SNOMEDCT_US|FEELING OF HOPELESSNESS |LOSS OF HOPE FOR THE FUTURE (FINDING)
C0150041|T048|389335004|SNOMEDCT_US|LOSS OF HOPE FOR THE FUTURE |LOSS OF HOPE FOR THE FUTURE (FINDING)
C0150041|T048|389335004|SNOMEDCT_US|FEELS THERE IS NO FUTURE|LOSS OF HOPE FOR THE FUTURE (FINDING)
C0150041|T048|389335004|SNOMEDCT_US|NO HOPE FOR THE FUTURE|LOSS OF HOPE FOR THE FUTURE (FINDING)
C0150041|T048|389335004|SNOMEDCT_US|CANNOT SEE A FUTURE|LOSS OF HOPE FOR THE FUTURE (FINDING)
C0150041|T048|389335004|SNOMEDCT_US|FEELING HOPELESS|LOSS OF HOPE FOR THE FUTURE (FINDING)
C0150041|T048|389335004|SNOMEDCT_US|FEELING HOPELESS |LOSS OF HOPE FOR THE FUTURE (FINDING)
C2219873|T048||SNOMEDCT_US|FEELS PESSIMISTIC ABOUT FUTURE OR BROODING ABOUT PAST
C2219873|T048||SNOMEDCT_US|FEELS PESSIMISTIC ABOUT FUTURE OR BROODING ABOUT PAST 
C2219873|T048||SNOMEDCT_US|FEEL PESSIMISTIC ABOUT FUTURE, OR BROODING ABOUT PAST
C2219873|T048||SNOMEDCT_US|PESSIMISTIC ABOUT THE FUTURE, OR BROODING ABOUT THE PAST
C2165505|T048||SNOMEDCT_US|DEPRESSION 1-3 DAYS PRIOR TO MENSTRUATION
C2165505|T048||SNOMEDCT_US|DEPRESSION 1-3 DAYS PRIOR TO MENSTRUATION 
C2165506|T048||SNOMEDCT_US|DEPRESSION ACCOMPANIED BY 
C2165506|T048||SNOMEDCT_US|DEPRESSION ACCOMPANIED BY
C2165506|T048||SNOMEDCT_US|DEPRESSION ACCOMPANIED
C2165516|T048||SNOMEDCT_US|DEPRESSION IS RELIEVED
C2165516|T048||SNOMEDCT_US|FACTORS RELIEVING DEPRESSION
C2165516|T048||SNOMEDCT_US|FACTORS RELIEVING DEPRESSION 
C2051715|T048||SNOMEDCT_US|DEPRESSION OCCURRING
C2051715|T048||SNOMEDCT_US|PATTERN OF DEPRESSION 
C2051715|T048||SNOMEDCT_US|PATTERN OF DEPRESSION
C2169543|T048||SNOMEDCT_US|DEPRESSION RECENTLY
C2169543|T048||SNOMEDCT_US|RECENT DEPRESSION
C2169543|T048||SNOMEDCT_US|RECENT DEPRESSION 
C1561368|T048||SNOMEDCT_US|CTCAE GRADE 3 DEPRESSION
C1561368|T048||SNOMEDCT_US|GRADE 3 DEPRESSION
C1561366|T048||SNOMEDCT_US|CTCAE GRADE 1 DEPRESSION
C1561366|T048||SNOMEDCT_US|GRADE 1 DEPRESSION
C1561367|T048||SNOMEDCT_US|CTCAE GRADE 2 DEPRESSION
C1561367|T048||SNOMEDCT_US|GRADE 2 DEPRESSION
C1561369|T048||SNOMEDCT_US|CTCAE GRADE 4 DEPRESSION
C1561369|T048||SNOMEDCT_US|GRADE 4 DEPRESSION
C1561370|T048||SNOMEDCT_US|CTCAE GRADE 5 DEPRESSION
C1561370|T048||SNOMEDCT_US|GRADE 5 DEPRESSION
