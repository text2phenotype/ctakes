C0086409|T098||CDC|HISPANICS
C3846650|T098||CDC|SPANISH,NOS; HISPANIC,NOS
C0019576|T098||CDC|HISPANIC AMERICANS
C1533017|T098||CDC|HISPANIC BLACK FINDING
C1533018|T098||CDC|HISPANIC BLACK RACIAL GROUP
C1533020|T098||CDC|HISPANIC WHITE FINDING
C1533021|T098||CDC|HISPANIC WHITE RACIAL GROUP
C1881927|T098||CDC|MULTIPLE HISPANIC
C2741637|T098||CDC|HISPANIC OR LATINO:FINDING:POINT IN TIME:^PATIENT:ORDINA
C3844642|T098||CDC|OTHER HISPANIC
C4036190|T098||CDC|YES, ANOTHER HISPANIC, LATINO-A, OR SPANISH ORIGIN
C0086409|T098||CDC|HISPANIC
C0086409|T098||CDC|CENTRAL AMERICAN
C0086409|T098||CDC|CANAL ZONE
C0086409|T098||CDC|CENTRAL AMERICAN INDIAN
C0086409|T098||CDC|COSTA RICAN
C0086409|T098||CDC|GUATEMALAN
C0086409|T098||CDC|HONDURAN
C0086409|T098||CDC|NICARAGUAN
C0086409|T098||CDC|PANAMANIAN
C0086409|T098||CDC|SALVADORAN
C0086409|T098||CDC|CUBAN
C0086409|T098||CDC|DOMINICAN
C0086409|T098||CDC|LATIN AMERICAN
C0086409|T098||CDC|MEXICAN
C0086409|T098||CDC|CHICANO
C0086409|T098||CDC|LA RAZA
C0086409|T098||CDC|MEXICAN AMERICAN INDIAN
C0086409|T098||CDC|MEXICAN AMERICAN
C0086409|T098||CDC|MEXICANO
C0086409|T098||CDC|PUERTO RICAN
C0086409|T098||CDC|SOUTH AMERICAN
C0086409|T098||CDC|ARGENTINEAN
C0086409|T098||CDC|BOLIVIAN
C0086409|T098||CDC|CHILEAN
C0086409|T098||CDC|COLOMBIAN
C0086409|T098||CDC|CRIOLLO
C0086409|T098||CDC|ECUADORIAN
C0086409|T098||CDC|PARAGUAYAN
C0086409|T098||CDC|PERUVIAN
C0086409|T098||CDC|SOUTH AMERICAN INDIAN
C0086409|T098||CDC|URUGUAYAN
C0086409|T098||CDC|VENEZUELAN
C0086409|T098||CDC|SPANIARD
C0086409|T098||CDC|ANDALUSIAN
C0086409|T098||CDC|ASTURIAN
C0086409|T098||CDC|BELEARIC ISLANDER
C0086409|T098||CDC|CANARIAN
C0086409|T098||CDC|CASTILLIAN
C0086409|T098||CDC|CATALONIAN
C0086409|T098||CDC|GALLEGO
C0086409|T098||CDC|SPANISH BASQUE
C0086409|T098||CDC|VALENCIAN
C0019576|T098||CDC|AMERICAN, HISPANIC
C0019576|T098||CDC|AMERICANS, HISPANIC
C0019576|T098||CDC|AMERICANS, SPANISH
C0019576|T098||CDC|HISPANIC AMERICAN
C0019576|T098||CDC|HISPANIC AMERICANS
C0019576|T098||CDC|SPANISH AMERICAN
C0019576|T098||CDC|SPANISH AMERICANS
C1553379|T098||CDC|CUBAN
C1553379|T098||CDC|-- CUBAN
C3829110|T098||CDC|MEXICAN OR MEXICAN AMERICAN
C3828691|T098||CDC|OTHER HISPANIC OR LATINO(A)
C3161473|T098||CDC|SPANISH
C3161473|T098||CDC|SPANISH PERSON
C0086409|T098||CDC|HISPANIC
C0086409|T098||CDC|HISPANICS
C0086409|T098||CDC|HISPANIC OR LATINO
C0086409|T098||CDC|ETHNICITYHISPANIC
C0086409|T098||CDC|HISPANIC ORIGIN
C0086409|T098||CDC|SPANISH
C0086409|T098||CDC|HISPANIC POPULATIONS
C0086409|T098||CDC|HISPANICS OR LATINOS
C0086409|T098||CDC|LATINO POPULATION
C0086409|T098||CDC|SPANISH ORIGIN
C0086409|T098||CDC|HISPANIC (RACIAL GROUP)
C0025884|T098||CDC|AMERICAN, MEXICAN
C0025884|T098||CDC|AMERICANS, MEXICAN
C0025884|T098||CDC|CHICANO
C0025884|T098||CDC|MEXICAN AMERICAN
C0025884|T098||CDC|MEXICAN AMERICANS
C0025884|T098||CDC|CHICANOS
C0025884|T098||CDC|CHICANAS
C0025884|T098||CDC|CHICANA
C0010436|T098||CDC|AMERICANS, CUBAN
C0010436|T098||CDC|CUBAN AMERICAN
C0010436|T098||CDC|CUBAN AMERICANS
C0086528|T098||CDC|LATINO
C0086528|T098||CDC|LATINOS
C0034043|T098||CDC|PUERTO RICAN
C0034043|T098||CDC|PUERTORICAN
C0034043|T098||CDC|-- PUERTO RICAN
C0034043|T098||CDC|PUERTO RICANS
C0935556|T098||CDC|LATINOS/LATINAS
C1533018|T098||CDC|HISPANIC, BLACK (RACIAL GROUP)
C1533018|T098||CDC|HISPANIC, BLACK
C1533018|T098||CDC|HISPANIC BLACK RACIAL GROUP
C1533019|T098||CDC|HISPANIC, COLOR UNKNOWN (RACIAL GROUP)
C1533019|T098||CDC|HISPANIC, COLOR UNKNOWN
C1533019|T098||CDC|HISPANIC, COLOUR UNKNOWN
C1533021|T098||CDC|HISPANIC, WHITE (RACIAL GROUP)
C1533021|T098||CDC|HISPANIC, WHITE
C1533021|T098||CDC|HISPANIC WHITE RACIAL GROUP
C0425359|T098||CDC|SOUTH AMERICAN
C0425359|T098||CDC|-- SOUTH AMERICAN
C0240339|T098||CDC|MEXICAN
C0240339|T098||CDC|ETHNICITYHISPANICMEXICAN
C0240339|T098||CDC|-- MEXICAN
C0238914|T098||CDC|CENTRAL AMERICAN
C0238914|T098||CDC|ETHNICITYHISPANICCENTRALAMERICAN
C0238914|T098||CDC|-- CENTRAL AMERICAN
C1328872|T098||CDC|DOMINICAN
C1328872|T098||CDC|DOMINICAN - ETHNICITY
C1553378|T098||CDC|LATIN AMERICAN
C0337817|T098||CDC|SPANIARDS
C0337817|T098||CDC|SPANIARDS 
C0337817|T098||CDC|SPANIARD
C1881927|T098||CDC|MULTIPLE HISPANIC
C1880193|T098||CDC|CUBAN OR CUBAN AMERICAN
C2135343|T098||CDC|CULTURAL BACKGROUND HISPANIC 
C2135343|T098||CDC|THE CULTURAL BACKGROUND IS HISPANIC
C2135343|T098||CDC|CULTURAL BACKGROUND HISPANIC
C2741637|T098||CDC|HISPANIC OR LATINO:FINDING:POINT IN TIME:^PATIENT:ORDINAL
C2741637|T098||CDC|HISPANIC OR LATINO
C2741637|T098||CDC|HISPANIC OR LATINO:FIND:PT:^PATIENT:ORD
