C0009555|T059|165409003|SNOMEDCT_US|COMPLETE BLOOD COUNT|FULL BLOOD COUNT NOS (PROCEDURE)
C0545131|T059||SNOMEDCT_US|COMPLETE BLOOD COUNT WITH DIFFERENTIAL 
C0545131|T059||SNOMEDCT_US|CBC WITH DIFFERENTIAL
C0545131|T059||SNOMEDCT_US|COMPLETE BLOOD COUNT WITH DIFFERENTIAL
C0545131|T059||SNOMEDCT_US|BLOOD CELL COUNT WITH DIFFERENTIAL
C0545131|T059||SNOMEDCT_US|CBC WITH DIFF
C0009555|T059|165409003|SNOMEDCT_US|COMPLETE BLOOD COUNT|FULL BLOOD COUNT NOS (PROCEDURE)
C0009555|T059|165409003|SNOMEDCT_US|CBC|FULL BLOOD COUNT NOS (PROCEDURE)
C0009555|T059|165409003|SNOMEDCT_US|BLOOD COUNTS, COMPLETE|FULL BLOOD COUNT NOS (PROCEDURE)
C0009555|T059|165409003|SNOMEDCT_US|COMPLETE BLOOD COUNTS|FULL BLOOD COUNT NOS (PROCEDURE)
C0009555|T059|165409003|SNOMEDCT_US|COUNT, COMPLETE BLOOD|FULL BLOOD COUNT NOS (PROCEDURE)
C0009555|T059|165409003|SNOMEDCT_US|COUNTS, COMPLETE BLOOD|FULL BLOOD COUNT NOS (PROCEDURE)
C0009555|T059|165409003|SNOMEDCT_US|FULL BLOOD COUNT|FULL BLOOD COUNT NOS (PROCEDURE)
C0009555|T059|165409003|SNOMEDCT_US|CBC (COMPLETE BLOOD COUNT)|FULL BLOOD COUNT NOS (PROCEDURE)
C0009555|T059|165409003|SNOMEDCT_US|COMPLETE BLOOD COUNT (CBC)|FULL BLOOD COUNT NOS (PROCEDURE)
C0009555|T059|165409003|SNOMEDCT_US|COMPLETE BLOOD COUNT (CBC) |FULL BLOOD COUNT NOS (PROCEDURE)
C0009555|T059|165409003|SNOMEDCT_US|FBC|FULL BLOOD COUNT NOS (PROCEDURE)
C0009555|T059|165409003|SNOMEDCT_US|TEST;FULL BLOOD COUNT|FULL BLOOD COUNT NOS (PROCEDURE)
C0009555|T059|165409003|SNOMEDCT_US|FULL BLOOD COUNT NOS |FULL BLOOD COUNT NOS (PROCEDURE)
C0009555|T059|165409003|SNOMEDCT_US|FULL BLOOD COUNT NOS|FULL BLOOD COUNT NOS (PROCEDURE)
C0009555|T059|165409003|SNOMEDCT_US|FULL BLOOD COUNT |FULL BLOOD COUNT NOS (PROCEDURE)
C0009555|T059|165409003|SNOMEDCT_US|BLOOD CELL COUNT|FULL BLOOD COUNT NOS (PROCEDURE)
C0009555|T059|165409003|SNOMEDCT_US|FBC - FULL BLOOD COUNT|FULL BLOOD COUNT NOS (PROCEDURE)
C0009555|T059|165409003|SNOMEDCT_US|COMPLETE BLOOD COUNT |FULL BLOOD COUNT NOS (PROCEDURE)
C0009555|T059|165409003|SNOMEDCT_US|COMPLETE BLOOD COUNT, NOS|FULL BLOOD COUNT NOS (PROCEDURE)
C0009555|T059|165409003|SNOMEDCT_US|CBC, NOS|FULL BLOOD COUNT NOS (PROCEDURE)
C0009555|T059|165409003|SNOMEDCT_US|BLOOD COUNT, COMPLETE|FULL BLOOD COUNT NOS (PROCEDURE)
C0523113|T059|104102000|SNOMEDCT_US|BLOOD BLAST COUNT|BLAST COUNT, BLOOD (PROCEDURE)
C0523113|T059|104102000|SNOMEDCT_US|BLOOD BLAST COUNT |BLAST COUNT, BLOOD (PROCEDURE)
C0523113|T059|104102000|SNOMEDCT_US|BLAST COUNT|BLAST COUNT, BLOOD (PROCEDURE)
C0523113|T059|104102000|SNOMEDCT_US|BLAST|BLAST COUNT, BLOOD (PROCEDURE)
C0523113|T059|104102000|SNOMEDCT_US|BLASTS|BLAST COUNT, BLOOD (PROCEDURE)
C0523113|T059|104102000|SNOMEDCT_US|BLAST CELLS|BLAST COUNT, BLOOD (PROCEDURE)
C0523113|T059|104102000|SNOMEDCT_US|BLAST CELLS NOS|BLAST COUNT, BLOOD (PROCEDURE)
C0523113|T059|104102000|SNOMEDCT_US|BLAST COUNT, BLOOD|BLAST COUNT, BLOOD (PROCEDURE)
C0523113|T059|104102000|SNOMEDCT_US|BLAST COUNT, BLOOD |BLAST COUNT, BLOOD (PROCEDURE)
C0523113|T059|104102000|SNOMEDCT_US|BLAST COUNT PROCEDURE|BLAST COUNT, BLOOD (PROCEDURE)
C2698870|T059||SNOMEDCT_US|PRECURSOR PLASMA CELL COUNT
C2698870|T059||SNOMEDCT_US|PRECURSOR PLASMA CELLS
C2698870|T059||SNOMEDCT_US|PLSPCE
C2698870|T059||SNOMEDCT_US|PLASMABLAST
C2698029|T059||SNOMEDCT_US|MATURE PLASMA CELL COUNT
C2698029|T059||SNOMEDCT_US|MATURE PLASMA CELLS
C2698029|T059||SNOMEDCT_US|PLASMACYTES
C2698029|T059||SNOMEDCT_US|PLSMCE
C2827509|T059||SNOMEDCT_US|EOSINOPHILIC METAMYELOCYTE COUNT
C2827509|T059||SNOMEDCT_US|EOSINOPHILIC METAMYELOCYTES
C2827509|T059||SNOMEDCT_US|EOSMM
C2827509|T059||SNOMEDCT_US|METAMYELOCYTES.EOSINOPHILIC
C2827510|T059||SNOMEDCT_US|EOSINOPHILIC MYELOCYTE COUNT
C2827510|T059||SNOMEDCT_US|EOSINOPHILIC MYELOCYTES
C2827510|T059||SNOMEDCT_US|EOSMYL
C2827511|T059||SNOMEDCT_US|NEUTROPHILIC METAMYELOCYTE COUNT
C2827511|T059||SNOMEDCT_US|NEUTROPHILIC METAMYELOCYTES
C2827511|T059||SNOMEDCT_US|NEUTMM
C2827512|T059||SNOMEDCT_US|NEUTROPHILIC MYELOCYTE COUNT
C2827512|T059||SNOMEDCT_US|NEUTROPHILIC MYELOCYTES
C2827512|T059||SNOMEDCT_US|NEUTMY
C0014772|T059|142839002|SNOMEDCT_US|COUNT, ERYTHROCYTE|RBC COUNT NOS (PROCEDURE)
C0014772|T059|142839002|SNOMEDCT_US|COUNTS, ERYTHROCYTE|RBC COUNT NOS (PROCEDURE)
C0014772|T059|142839002|SNOMEDCT_US|ERYTHROCYTE COUNT|RBC COUNT NOS (PROCEDURE)
C0014772|T059|142839002|SNOMEDCT_US|ERYTHROCYTE COUNTS|RBC COUNT NOS (PROCEDURE)
C0014772|T059|142839002|SNOMEDCT_US|ERYTHROCYTE NUMBERS|RBC COUNT NOS (PROCEDURE)
C0014772|T059|142839002|SNOMEDCT_US|RED BLOOD CELL COUNT|RBC COUNT NOS (PROCEDURE)
C0014772|T059|142839002|SNOMEDCT_US|RBC COUNT NOS |RBC COUNT NOS (PROCEDURE)
C0014772|T059|142839002|SNOMEDCT_US|ERYTHROCYTE COUNT |RBC COUNT NOS (PROCEDURE)
C0014772|T059|142839002|SNOMEDCT_US|RBC COUNT|RBC COUNT NOS (PROCEDURE)
C0014772|T059|142839002|SNOMEDCT_US|RED CELL COUNT|RBC COUNT NOS (PROCEDURE)
C0014772|T059|142839002|SNOMEDCT_US|RED BLOOD CELL COUNT |RBC COUNT NOS (PROCEDURE)
C0014772|T059|142839002|SNOMEDCT_US|RBC COUNT NOS|RBC COUNT NOS (PROCEDURE)
C0014772|T059|142839002|SNOMEDCT_US|RED BLOOD CELL COUNT NOS |RBC COUNT NOS (PROCEDURE)
C0014772|T059|142839002|SNOMEDCT_US|RED BLOOD CELL COUNT NOS|RBC COUNT NOS (PROCEDURE)
C0014772|T059|142839002|SNOMEDCT_US|ERYTHROCYTES|RBC COUNT NOS (PROCEDURE)
C0014772|T059|142839002|SNOMEDCT_US|RBC|RBC COUNT NOS (PROCEDURE)
C0014772|T059|142839002|SNOMEDCT_US|RED BLOOD CELLS|RBC COUNT NOS (PROCEDURE)
C0014772|T059|142839002|SNOMEDCT_US|ERYTHROCYTE NUMBER|RBC COUNT NOS (PROCEDURE)
C0014772|T059|142839002|SNOMEDCT_US|BLOOD CELL COUNT, RED|RBC COUNT NOS (PROCEDURE)
C0014772|T059|142839002|SNOMEDCT_US|WHOLE BLOOD ERYTHROCYTIC CELL COUNTS|RBC COUNT NOS (PROCEDURE)
C0014772|T059|142839002|SNOMEDCT_US|RBC - RED BLOOD CELL COUNT|RBC COUNT NOS (PROCEDURE)
C0014772|T059|142839002|SNOMEDCT_US|RED BLOOD CELL COUNT MEASUREMENT|RBC COUNT NOS (PROCEDURE)
C0518015|T059|35170002|SNOMEDCT_US|HAEMOGLOBIN|HEMOGLOBIN DETERMINATION (PROCEDURE)
C0518015|T059|35170002|SNOMEDCT_US|HAEM|HEMOGLOBIN DETERMINATION (PROCEDURE)
C0518015|T059|35170002|SNOMEDCT_US|HEMOGLOBIN MEASUREMENT|HEMOGLOBIN DETERMINATION (PROCEDURE)
C0518015|T059|35170002|SNOMEDCT_US|HEMOGLOBIN|HEMOGLOBIN DETERMINATION (PROCEDURE)
C0518015|T059|35170002|SNOMEDCT_US|HEMOGLOBIN MEASUREMENT |HEMOGLOBIN DETERMINATION (PROCEDURE)
C0518015|T059|35170002|SNOMEDCT_US|TEST;HAEMOGLOBIN|HEMOGLOBIN DETERMINATION (PROCEDURE)
C0518015|T059|35170002|SNOMEDCT_US|BLOOD COUNT HEMOGLOBIN|HEMOGLOBIN DETERMINATION (PROCEDURE)
C0518015|T059|35170002|SNOMEDCT_US|HEMOGLOBIN LEVEL|HEMOGLOBIN DETERMINATION (PROCEDURE)
C0518015|T059|35170002|SNOMEDCT_US|MEASUREMENT OF HEMOGLOBIN (HGB)|HEMOGLOBIN DETERMINATION (PROCEDURE)
C0518015|T059|35170002|SNOMEDCT_US|HEMOGLOBIN DETERMINATION |HEMOGLOBIN DETERMINATION (PROCEDURE)
C0518015|T059|35170002|SNOMEDCT_US|HEMOGLOBIN DETERMINATION|HEMOGLOBIN DETERMINATION (PROCEDURE)
C0518015|T059|35170002|SNOMEDCT_US|HAEMOGLOBIN DETERMINATION|HEMOGLOBIN DETERMINATION (PROCEDURE)
C0518015|T059|35170002|SNOMEDCT_US|HGB|HEMOGLOBIN DETERMINATION (PROCEDURE)
C0518015|T059|35170002|SNOMEDCT_US|BLOOD COUNT; HEMOGLOBIN (HGB)|HEMOGLOBIN DETERMINATION (PROCEDURE)
C0518015|T059|35170002|SNOMEDCT_US|FHGB|HEMOGLOBIN DETERMINATION (PROCEDURE)
C0518015|T059|35170002|SNOMEDCT_US|FREE HEMOGLOBIN|HEMOGLOBIN DETERMINATION (PROCEDURE)
C0518015|T059|35170002|SNOMEDCT_US|HEMOGLOBIN DETERMINATION, NOS|HEMOGLOBIN DETERMINATION (PROCEDURE)
C0518015|T059|35170002|SNOMEDCT_US|HAEMOGLOBIN DETERMINATION, NOS|HEMOGLOBIN DETERMINATION (PROCEDURE)
C0518015|T059|35170002|SNOMEDCT_US|TEST;HEMOGLOBIN|HEMOGLOBIN DETERMINATION (PROCEDURE)
C0518015|T059|35170002|SNOMEDCT_US|HAEMOGLOBIN TEST|HEMOGLOBIN DETERMINATION (PROCEDURE)
C0518015|T059|35170002|SNOMEDCT_US|HEMOGLOBIN TEST|HEMOGLOBIN DETERMINATION (PROCEDURE)
C0018935|T059|165418001|SNOMEDCT_US|HCT|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|ERYTHROCYTE VOLUMES, PACKED|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|HEMATOCRIT|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|HEMATOCRITS|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|PACKED ERYTHROCYTE VOLUME|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|PACKED ERYTHROCYTE VOLUMES|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|PACKED RED CELL VOLUME|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|PACKED RED-CELL VOLUMES|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|RED-CELL VOLUME, PACKED|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|RED-CELL VOLUMES, PACKED|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|VOLUME, PACKED ERYTHROCYTE|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|VOLUME, PACKED RED-CELL|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|VOLUMES, PACKED ERYTHROCYTE|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|VOLUMES, PACKED RED-CELL|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|HAEMATOCRIT|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|HEMATOCRIT PROCEDURE|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|HEMATOCRIT |HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|HEMATOCRIT MEASUREMENT|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|BLOOD COUNT HEMATOCRIT|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|MEASUREMENT OF HEMATOCRIT (HCT)|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|PACKED CELL VOLUME (OBSERVABLE ENTITY)|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|HAEMATOCRIT - PCV - NOS|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|PACKED CELL VOLUME|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|HAEMATOCRIT (OBSERVABLE ENTITY)|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|HAEMATOCRIT |HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|HEMATOCRIT - PCV - NOS|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|HAEMATOCRIT - PCV - NOS |HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|HEMATOCRIT - PCV - NOS |HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|HEMATOCRIT PACKED CELL VOLUME |HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|HEMATOCRIT PACKED CELL VOLUME|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|EVF|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|PCV|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|ERYTHROCYTE VOLUME FRACTION|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|BLOOD COUNT; HEMATOCRIT (HCT)|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|PACKED RED-CELL VOLUME|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|ERYTHROCYTE VOLUME, PACKED|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|WHOLE BLOOD HEMATOCRIT TEST|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|HEMATOCRIT DETERMINATION|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|HAEMATOCRIT - PCV|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|HCT - HAEMATOCRIT|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|HCT - HEMATOCRIT|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|HEMATOCRIT - PCV|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|HAEMATOCRIT DETERMINATION|HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|HEMATOCRIT DETERMINATION |HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|PACKED CELL VOLUME MEASUREMENT |HAEMATOCRIT (OBSERVABLE ENTITY)
C0018935|T059|165418001|SNOMEDCT_US|PACKED CELL VOLUME MEASUREMENT|HAEMATOCRIT (OBSERVABLE ENTITY)
C0023508|T059|767002|SNOMEDCT_US|WHITE BLOOD CELL COUNT|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|COUNT, LEUKOCYTE|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|COUNTS, LEUKOCYTE|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|LEUKOCYTE COUNT|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|LEUKOCYTE COUNTS|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|LEUKOCYTE NUMBERS|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|NUMBER, LEUKOCYTE|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|NUMBERS, LEUKOCYTE|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|WHITE BLOOD CELL COUNT PROCEDURE|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|LEUKOCYTE COUNT |WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|WBC COUNT|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|WHITE BLOOD CELL COUNT |WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|LEUKOCYTES|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|WHITE BLOOD CELLS|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|WBC|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|WHITE CELLS|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|LEUKOCYTE COUNT NOS|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|WHITE BLOOD CELL COUNT NOS|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|WHITE BLOOD CELL ANALYSIS|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|LEUCOCYTE COUNT|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|LEUKOCYTE NUMBER|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|BLOOD CELL COUNT, WHITE|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|WHOLE BLOOD LEUKOCYTE COUNTS|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|WBC - WHITE BLOOD CELL COUNT|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|WCC - WHITE BLOOD CELL COUNT|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T059|767002|SNOMEDCT_US|WHITE BLOOD CELL COUNT - OBSERVATION|WHITE BLOOD CELL COUNT - OBSERVATION
C2097083|T059||SNOMEDCT_US|COMPLETE BLOOD COUNT WITH MANUAL DIFFERENTIAL AND INDICES 
C2097083|T059||SNOMEDCT_US|CBC WITH MANUAL DIFFERENTIAL AND INDICES
C2097083|T059||SNOMEDCT_US|MANUAL CBC WITH DIFFERENTIAL AND INDICES
C2097083|T059||SNOMEDCT_US|COMPLETE BLOOD COUNT WITH MANUAL DIFFERENTIAL AND INDICES
C2030595|T059||SNOMEDCT_US|HEMOGRAM INDICES 
C2030595|T059||SNOMEDCT_US|HEMOGRAM INDICES
C2984931|T059||SNOMEDCT_US|MYELOID TO ERYTHROID RATIO MEASUREMENT
C2984931|T059||SNOMEDCT_US|MYPCERPC
C2984931|T059||SNOMEDCT_US|MYELOID/ERYTHROID RATIO
C3272957|T059||SNOMEDCT_US|IMMATURE PLASMA CELL COUNT
C3272957|T059||SNOMEDCT_US|IMMATURE PLASMA CELLS
C3272957|T059||SNOMEDCT_US|PLSIMCE
C0200694|T059|68994006|SNOMEDCT_US|MEASUREMENT OF TOTAL HEMOGLOBIN CONCENTRATION AND HEMATOCRIT |MEASUREMENT OF TOTAL HEMOGLOBIN CONCENTRATION AND HEMATOCRIT (PROCEDURE)
C0200694|T059|68994006|SNOMEDCT_US|HEMOGLOBIN AND HEMATOCRIT DETERMINATION|MEASUREMENT OF TOTAL HEMOGLOBIN CONCENTRATION AND HEMATOCRIT (PROCEDURE)
C0200694|T059|68994006|SNOMEDCT_US|MEASUREMENT OF TOTAL HEMOGLOBIN CONCENTRATION AND HEMATOCRIT|MEASUREMENT OF TOTAL HEMOGLOBIN CONCENTRATION AND HEMATOCRIT (PROCEDURE)
C0200694|T059|68994006|SNOMEDCT_US|MEASUREMENT OF TOTAL HAEMOGLOBIN CONCENTRATION AND HAEMATOCRIT|MEASUREMENT OF TOTAL HEMOGLOBIN CONCENTRATION AND HEMATOCRIT (PROCEDURE)
C0200694|T059|68994006|SNOMEDCT_US|HEMOGLOBIN AND HEMATOCRIT DETERMINATION |MEASUREMENT OF TOTAL HEMOGLOBIN CONCENTRATION AND HEMATOCRIT (PROCEDURE)
C0200694|T059|68994006|SNOMEDCT_US|HAEMOGLOBIN AND HAEMATOCRIT DETERMINATION|MEASUREMENT OF TOTAL HEMOGLOBIN CONCENTRATION AND HEMATOCRIT (PROCEDURE)
C0200694|T059|68994006|SNOMEDCT_US|H & H DETERMINATION|MEASUREMENT OF TOTAL HEMOGLOBIN CONCENTRATION AND HEMATOCRIT (PROCEDURE)
C0200694|T059|68994006|SNOMEDCT_US|TOTAL HEMOGLOBIN CONCENTRATION AND HEMATOCRIT|MEASUREMENT OF TOTAL HEMOGLOBIN CONCENTRATION AND HEMATOCRIT (PROCEDURE)
C0200694|T059|68994006|SNOMEDCT_US|TOTAL HEMOGLOBIN CONCENTRATION AND HEMATOCRIT |MEASUREMENT OF TOTAL HEMOGLOBIN CONCENTRATION AND HEMATOCRIT (PROCEDURE)
C0200694|T059|68994006|SNOMEDCT_US|HAEMOGLOBIN AND HEMATOCRIT DETERMINATION|MEASUREMENT OF TOTAL HEMOGLOBIN CONCENTRATION AND HEMATOCRIT (PROCEDURE)
C2228885|T059||SNOMEDCT_US|MEAN CORPUSCULAR DIAMETER (MCD)
C2228885|T059||SNOMEDCT_US|MEAN CORPUSCULAR DIAMETER (MCD) 
C2228885|T059||SNOMEDCT_US|MEAN CORPUSCULAR DIAMETER
C2228299|T059||SNOMEDCT_US|ERYTHROCYTE VOLUME DISTRIBUTION WIDTH (RDW)
C2228299|T059||SNOMEDCT_US|RBC VOLUME DISTRIBUTION WIDTH (RDW)
C2228299|T059||SNOMEDCT_US|ERYTHROCYTE VOLUME DISTRIBUTION WIDTH (RDW) 
C2228299|T059||SNOMEDCT_US|RBC VOLUME DISTRIBUTION WIDTH
C0883120|T059||SNOMEDCT_US|HEMOGLOBIN & HEMATOCRIT PANEL
C0883120|T059||SNOMEDCT_US|HEMOGLOBIN AND HEMATOCRIT PANEL 
C0883120|T059||SNOMEDCT_US|HEMOGLOBIN AND HEMATOCRIT PANEL
C0369183|T059|142847002|SNOMEDCT_US|MEAN CELL HAEMOGLOBIN|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MCH - NOS |MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|ERYTHROCYTE MEAN CORPUSCULAR HEMOGLOBIN|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|ERYTHROCYTE MEAN CORPUSCULAR HEMOGLOBIN TEST|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MEAN CORPUSCULAR HEMOGLOBIN (MCH)|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MEAN CORPUSCULAR HEMOGLOBIN (MCH) |MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MEAN CORPUSCULAR HAEMOGLOBIN (MCH) - NOS |MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MCH|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MCH - NOS|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MEAN CORPUSCULAR HEMOGLOBIN (MCH) - NOS|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MEAN CELL HAEMOGLOBIN (& LEVEL)|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MEAN CORPUSCULAR HAEMOGLOBIN (MCH) - NOS|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MEAN CELL HAEMOGLOBIN (& LEVEL) |MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MEAN CELL HEMOGLOBIN (& LEVEL)|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MEAN CORPUSCULAR HEMOGLOBIN NOS|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MEAN CELL HEMOGLOBIN|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MEAN CORPUSCULAR HAEMOGLOBIN NOS|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MEAN CORPUSCULAR HEMOGLOBIN NOS |MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|ERY. MEAN CORPUSCULAR HEMOGLOBIN|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MEAN CORPUSCULAR HEMOGLOBIN|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MEAN CORPUSCULAR HAEMOGLOBIN|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MEAN CORPUSCULAR HEMOGLOBIN DETERMINATION|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MCH DETERMINATION|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MCH - MEAN CELL HAEMOGLOBIN|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MCH - MEAN CELL HEMOGLOBIN|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MEAN CORPUSCULAR HAEMOGLOBIN DETERMINATION|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MCH - MEAN CORPUSCULAR HAEMOGLOBIN|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MCH - MEAN CORPUSCULAR HEMOGLOBIN|MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C0369183|T059|142847002|SNOMEDCT_US|MEAN CORPUSCULAR HEMOGLOBIN DETERMINATION |MEAN CELL HAEMOGLOBIN (& LEVEL) (PROCEDURE)
C1948043|T059||SNOMEDCT_US|ERYTHROCYTE MEAN CORPUSCULAR VOLUME
C1948043|T059||SNOMEDCT_US|ERYTHROCYTE MEAN CORPUSCULAR VOLUME MEASUREMENT
C1948043|T059||SNOMEDCT_US|MEAN CORPUSCULAR VOLUME (MCV) 
C1948043|T059||SNOMEDCT_US|MEAN CORPUSCULAR VOLUME (MCV)
C1948043|T059||SNOMEDCT_US|MEAN CORPUSCULAR VOLUME
C1948043|T059||SNOMEDCT_US|ERY. MEAN CORPUSCULAR VOLUME
C1948043|T059||SNOMEDCT_US|RBC MEAN CORPUSCULAR VOLUME
C1948043|T059||SNOMEDCT_US|MCV
C1948043|T059||SNOMEDCT_US|ERYTHROCYTES MEAN CORPUSCULAR VOLUME
C2030597|T059||SNOMEDCT_US|CBC WITH PLATELET COUNT
C2030597|T059||SNOMEDCT_US|CBC WITH PLATELET COUNT 
C4031906|T059||SNOMEDCT_US|CBC AUTOMATED
C4031906|T059||SNOMEDCT_US|AUTOMATED CBC 
C4031906|T059||SNOMEDCT_US|AUTOMATED CBC
C0200665|T059|103214008|SNOMEDCT_US|MEAN PLATELET VOLUME|PLATELET MEAN VOLUME (OBSERVABLE ENTITY)
C0200665|T059|103214008|SNOMEDCT_US|MEAN PLATELET VOLUME (MPV) |PLATELET MEAN VOLUME (OBSERVABLE ENTITY)
C0200665|T059|103214008|SNOMEDCT_US|MEAN PLATELET VOLUME (MPV)|PLATELET MEAN VOLUME (OBSERVABLE ENTITY)
C0200665|T059|103214008|SNOMEDCT_US|MPV|PLATELET MEAN VOLUME (OBSERVABLE ENTITY)
C0200665|T059|103214008|SNOMEDCT_US|MEAN PLATELET VOLUME MEASUREMENT|PLATELET MEAN VOLUME (OBSERVABLE ENTITY)
C0200665|T059|103214008|SNOMEDCT_US|VOLUMES, MEAN PLATELET|PLATELET MEAN VOLUME (OBSERVABLE ENTITY)
C0200665|T059|103214008|SNOMEDCT_US|PLATELET VOLUMES, MEAN|PLATELET MEAN VOLUME (OBSERVABLE ENTITY)
C0200665|T059|103214008|SNOMEDCT_US|PLATELET VOLUME, MEAN|PLATELET MEAN VOLUME (OBSERVABLE ENTITY)
C0200665|T059|103214008|SNOMEDCT_US|VOLUME, MEAN PLATELET|PLATELET MEAN VOLUME (OBSERVABLE ENTITY)
C0200665|T059|103214008|SNOMEDCT_US|MEAN PLATELET VOLUMES|PLATELET MEAN VOLUME (OBSERVABLE ENTITY)
C0200665|T059|103214008|SNOMEDCT_US|MPV - MEAN PLATELET VOLUME|PLATELET MEAN VOLUME (OBSERVABLE ENTITY)
C0200665|T059|103214008|SNOMEDCT_US|PLATELET MEAN VOLUME (OBSERVABLE ENTITY)|PLATELET MEAN VOLUME (OBSERVABLE ENTITY)
C0200665|T059|103214008|SNOMEDCT_US|PLATELET MEAN VOLUME|PLATELET MEAN VOLUME (OBSERVABLE ENTITY)
C0200665|T059|103214008|SNOMEDCT_US|PLATELET MEAN VOLUME DETERMINATION|PLATELET MEAN VOLUME (OBSERVABLE ENTITY)
C0200665|T059|103214008|SNOMEDCT_US|PLATELET MEAN VOLUME DETERMINATION |PLATELET MEAN VOLUME (OBSERVABLE ENTITY)
C4054355|T059||SNOMEDCT_US|NEUTROPHILS BAND FORM/ NEUTROPHILS
C4054355|T059||SNOMEDCT_US|NEUTBNE
C4054355|T059||SNOMEDCT_US|NEUTROPHILS BAND FORM TO NEUTROPHILS RATIO MEASUREMENT
C4054477|T059||SNOMEDCT_US|MONOCYTOID CELLS/LEUKOCYTES
C4054477|T059||SNOMEDCT_US|MONOCYTOID CELLS TO LEUKOCYTES RATIO MEASUREMENT
C4054477|T059||SNOMEDCT_US|MOCYCELE
C4054040|T059||SNOMEDCT_US|NEUTSGNE
C4054040|T059||SNOMEDCT_US|NEUTROPHILS, SEGMENTED/NEUTROPHILS
C4054040|T059||SNOMEDCT_US|SEGMENTED NEUTROPHILS TO NEUTROPHILS RATIO MEASUREMENT
C0200629|T059|35774004|SNOMEDCT_US|COMPLETE BLOOD COUNT WITH MANUAL DIFFERENTIAL|COMPLETE BLOOD COUNT WITH WHITE CELL DIFFERENTIAL, MANUAL (PROCEDURE)
C0200629|T059|35774004|SNOMEDCT_US|COMPLETE BLOOD COUNT WITH MANUAL DIFFERENTIAL |COMPLETE BLOOD COUNT WITH WHITE CELL DIFFERENTIAL, MANUAL (PROCEDURE)
C0200629|T059|35774004|SNOMEDCT_US|CBC WITH MANUAL DIFFERENTIAL|COMPLETE BLOOD COUNT WITH WHITE CELL DIFFERENTIAL, MANUAL (PROCEDURE)
C0200629|T059|35774004|SNOMEDCT_US|COMPLETE BLOOD COUNT WITH WHITE CELL DIFFERENTIAL, MANUAL|COMPLETE BLOOD COUNT WITH WHITE CELL DIFFERENTIAL, MANUAL (PROCEDURE)
C0200629|T059|35774004|SNOMEDCT_US|COMPLETE BLOOD COUNT WITH WHITE CELL DIFFERENTIAL, MANUAL |COMPLETE BLOOD COUNT WITH WHITE CELL DIFFERENTIAL, MANUAL (PROCEDURE)
C0200630|T059|9564003|SNOMEDCT_US|CBC WITH AUTOMATED DIFFERENTIAL|COMPLETE BLOOD COUNT WITH WHITE CELL DIFFERENTIAL, AUTOMATED (PROCEDURE)
C0200630|T059|9564003|SNOMEDCT_US|CBC WITH AUTOMATED DIFFERENTIAL |COMPLETE BLOOD COUNT WITH WHITE CELL DIFFERENTIAL, AUTOMATED (PROCEDURE)
C0200630|T059|9564003|SNOMEDCT_US|COMPLETE BLOOD COUNT WITH WHITE CELL DIFFERENTIAL, AUTOMATED|COMPLETE BLOOD COUNT WITH WHITE CELL DIFFERENTIAL, AUTOMATED (PROCEDURE)
C0200630|T059|9564003|SNOMEDCT_US|COMPLETE BLOOD COUNT WITH WHITE CELL DIFFERENTIAL, AUTOMATED |COMPLETE BLOOD COUNT WITH WHITE CELL DIFFERENTIAL, AUTOMATED (PROCEDURE)
C0200631|T059|43789009|SNOMEDCT_US|HEMOGRAM|COMPLETE BLOOD COUNT WITHOUT DIFFERENTIAL (PROCEDURE)
C0200631|T059|43789009|SNOMEDCT_US|COMPLETE BLOOD COUNT WITHOUT DIFFERENTIAL|COMPLETE BLOOD COUNT WITHOUT DIFFERENTIAL (PROCEDURE)
C0200631|T059|43789009|SNOMEDCT_US|CBC WITHOUT DIFFERENTIAL|COMPLETE BLOOD COUNT WITHOUT DIFFERENTIAL (PROCEDURE)
C0200631|T059|43789009|SNOMEDCT_US|HAEMOGRAM|COMPLETE BLOOD COUNT WITHOUT DIFFERENTIAL (PROCEDURE)
C0200631|T059|43789009|SNOMEDCT_US|COMPLETE BLOOD COUNT WITHOUT DIFFERENTIAL |COMPLETE BLOOD COUNT WITHOUT DIFFERENTIAL (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|BLOOD PLATELET COUNTS|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|BLOOD PLATELET NUMBERS|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|COUNT, BLOOD PLATELET|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|COUNT, PLATELET|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|COUNTS, BLOOD PLATELET|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|COUNTS, PLATELET|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|NUMBER, BLOOD PLATELET|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|NUMBER, PLATELET|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|NUMBERS, BLOOD PLATELET|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|NUMBERS, PLATELET|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|PLATELET COUNT|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|PLATELET COUNT, BLOOD|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|PLATELET COUNTS|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|PLATELET COUNTS, BLOOD|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|PLATELET NUMBER, BLOOD|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|PLATELET NUMBERS|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|PLATELET NUMBERS, BLOOD|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|PLATELETS|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|PLATELET COUNT |PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|PLATELET COUNT NOS |PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|PLATELET COUNT NOS|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|PLATELET COUNT |PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|PLAT|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|ANUCLEATED THROMBOCYTES|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|THROMBOCYTE COUNT|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|PLATELET NUMBER|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|BLOOD PLATELET COUNT|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|BLOOD PLATELET NUMBER|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|WHOLE BLOOD PLATELET COUNTS|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|PLT - PLATELET COUNT|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|PLATELET COUNT - OBSERVATION|PLATELET COUNT (PROCEDURE)
C0032181|T059|61928009|SNOMEDCT_US|PLATELET COUNT MEASUREMENT|PLATELET COUNT (PROCEDURE)
C1879889|T059||SNOMEDCT_US|BLOOD CELL COUNT RATIO MEASUREMENT
