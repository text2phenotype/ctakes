// ID|NAME
0|ABANDA
1|ABBEVILLE
2|ABBOTSFORD
3|ABBOTT
4|ABBOTTSBURG
5|ABBOTTSTOWN
6|ABBYVILLE
7|ABELL
8|ABERCROMBIE
9|ABERDEEN
10|ABERDEEN GARDENS
11|ABERFOIL
12|ABERNANT
13|ABERNATHY
14|ABEYTAS
15|ABIE
16|ABILENE
17|ABINGDON
18|ABINGTON
19|ABIQUIU
20|ABITA SPRINGS
21|ABO
22|ABOITE
23|ABRAHAM
24|ABRAM
25|ABRAMS
26|ABSAROKEE
27|ABSECON
28|ACADEMY
29|ACAMPO
30|ACCOKEEK
31|ACCOMAC
32|ACCORD
33|ACCOVILLE
34|ACEITUNAS
35|ACEITUNAS COMUNIDAD
36|ACEQUIA
37|ACHILLE
38|ACHILLES
39|ACKERLY
40|ACKERMAN
41|ACKERMANVILLE
42|ACKLEY
43|ACKWORTH
44|ACME
45|ACOMA
46|ACOMITA
47|ACOMITA LAKE
48|ACORN
49|ACRA
50|ACREE
51|ACRES GREEN
52|ACTON
53|ACWORTH
54|ACY
55|ADA
56|ADAIR
57|ADAIR VILLAGE
58|ADAIRSVILLE
59|ADAIRVILLE
60|ADAK
61|ADAMS
62|ADAMS CENTER
63|ADAMS CITY
64|ADAMSBURG
65|ADAMSTOWN
66|ADAMSVILLE
67|ADARIO
68|ADDICKS
69|ADDIE
70|ADDIEVILLE
71|ADDINGTON
72|ADDIS
73|ADDISON
74|ADDY
75|ADDYSTON
76|ADEL
77|ADELAIDE
78|ADELANTO
79|ADELINE
80|ADELINO
81|ADELL
82|ADELPHI
83|ADELPHIA
84|ADEN
85|ADENA
86|ADGATEVILLE
87|ADIN
88|ADJUNTAS
89|ADJUNTAS ZONA URBANA
90|ADMIRE
91|ADNA
92|ADOLPHUS
93|ADONA
94|ADRIAN
95|ADVANCE
96|ADWOLF
97|ADY
98|AENEAS
99|AETNA
100|AFFTON
101|AFTON
102|AGAR
103|AGATE
104|AGATE BEACH
105|AGAWAM
106|AGENCY
107|AGENDA
108|AGES
109|AGNES
110|AGNESS
111|AGNEW
112|AGNOS
113|AGOURA
114|AGOURA HILLS
115|AGRA
116|AGRICOLA
117|AGUA DULCE
118|AGUA FRIA
119|AGUA NUEVA
120|AGUADA
121|AGUADA ZONA URBANA
122|AGUADILLA
123|AGUADILLA ZONA URBANA
124|AGUANGA
125|AGUAS BUENAS
126|AGUAS BUENAS ZONA URBANA
127|AGUAS CLARAS
128|AGUAS CLARAS COMUNIDAD
129|AGUDO
130|AGUILA
131|AGUILAR
132|AGUILARES
133|AGUILITA
134|AGUILITA COMUNIDAD
135|AHLOSO
136|AHMEEK
137|AHOSKIE
138|AHTANUM
139|AHWAHNEE
140|AIBONITO
141|AIBONITO ZONA URBANA
142|AIEA
143|AIKEN
144|AILEY
145|AINSWORTH
146|AIRMONT
147|AIRPORT DRIVE
148|AIRPORT ROAD ADDITION
149|AIRWAY HEIGHTS
150|AITKIN
151|AJO
152|AK CHIN
153|AK-CHIN VILLAGE
154|AKASKA
155|AKELEY
156|AKERS
157|AKHIOK
158|AKIACHAK
159|AKIAK
160|AKIN
161|AKINS
162|AKRA
163|AKRON
164|AKUTAN
165|ALABAM
166|ALABASTER
167|ALACHUA
168|ALADDIN
169|ALAFAYA
170|ALAKANUK
171|ALAMANCE
172|ALAMEDA
173|ALAMILLO
174|ALAMO
175|ALAMO ALTO
176|ALAMO HEIGHTS
177|ALAMO OAKS
178|ALAMOGORDO
179|ALAMOSA
180|ALAMOTA
181|ALANREED
182|ALANSON
183|ALAPAHA
184|ALARKA
185|ALATNA
186|ALBA
187|ALBANY
188|ALBEE
189|ALBEMARLE
190|ALBERENE
191|ALBERHILL
192|ALBERS
193|ALBERT
194|ALBERT CITY
195|ALBERT LEA
196|ALBERTA
197|ALBERTON
198|ALBERTSON
199|ALBERTVILLE
200|ALBIA
201|ALBIN
202|ALBION
203|ALBORN
204|ALBRIGHT
205|ALBRIGHTSVILLE
206|ALBUQUERQUE
207|ALBURG
208|ALBURNETT
209|ALBURTIS
210|ALCALDE
211|ALCAN
212|ALCESTER
213|ALCO
214|ALCOA
215|ALCOA CENTER
216|ALCOLU
217|ALCOMA
218|ALCOVA
219|ALDA
220|ALDAN
221|ALDEN
222|ALDEN BRIDGE
223|ALDER
224|ALDER CREEK
225|ALDERDALE
226|ALDERLEY
227|ALDERPOINT
228|ALDERSON
229|ALDERTON
230|ALDERWOOD MANOR
231|ALDINE
232|ALDORA
233|ALDRICH
234|ALEDO
235|ALEKNAGIK
236|ALENEVA
237|ALEX
238|ALEXANDER
239|ALEXANDER CITY
240|ALEXANDER MILLS
241|ALEXANDRIA
242|ALEXANDRIA BAY
243|ALEXIS
244|ALFALFA
245|ALFARATA
246|ALFORD
247|ALFORDSVILLE
248|ALFRED
249|ALGER
250|ALGERITA
251|ALGOA
252|ALGODONES
253|ALGOMA
254|ALGONA
255|ALGONAC
256|ALGONQUIN
257|ALGOOD
258|ALHAMBRA
259|ALI CHUK
260|ALI CHUKSON
261|ALI MOLINA
262|ALIANZA
263|ALIANZA COMUNIDAD
264|ALICE
265|ALICE ACRES
266|ALICEVILLE
267|ALICIA
268|ALINE
269|ALIQUIPPA
270|ALIRE
271|ALISO VIEJO
272|ALIX
273|ALKABO
274|ALLAKAKET
275|ALLAMUCHY
276|ALLANDALE
277|ALLARDT
278|ALLEENE
279|ALLEGAN
280|ALLEGANY
281|ALLEGHANY
282|ALLEGHENYVILLE
283|ALLEGRE
284|ALLEMAN
285|ALLEN
286|ALLEN CITY
287|ALLEN PARK
288|ALLENDALE
289|ALLENFARM
290|ALLENHURST
291|ALLENPORT
292|ALLENSPARK
293|ALLENSVILLE
294|ALLENSWORTH
295|ALLENTON
296|ALLENTOWN
297|ALLENVILLE
298|ALLENWOOD
299|ALLERTON
300|ALLEYTON
301|ALLGOOD
302|ALLIANCE
303|ALLIGATOR
304|ALLISON
305|ALLISON PARK
306|ALLISONIA
307|ALLONS
308|ALLOUEZ
309|ALLOWAY
310|ALLPORT
311|ALLUWE
312|ALLYN
313|ALMA
314|ALMA CENTER
315|ALMANOR
316|ALMEDIA
317|ALMELUND
318|ALMENA
319|ALMERIA
320|ALMIRA
321|ALMO
322|ALMON
323|ALMOND
324|ALMONT
325|ALMONTE
326|ALMOTA
327|ALMY
328|ALMYRA
329|ALNWICK
330|ALOE
331|ALOHA
332|ALONDRA PARK
333|ALORTON
334|ALPAUGH
335|ALPENA
336|ALPHA
337|ALPHARETTA
338|ALPINE
339|ALPINE VILLAGE
340|ALQUINA
341|ALSACE MANOR
342|ALSATIA
343|ALSEA
344|ALSEN
345|ALSEY
346|ALSIP
347|ALSTON
348|ALSTOWN
349|ALSUMA
350|ALTA
351|ALTA LOMA
352|ALTA SIERRA
353|ALTA VISTA
354|ALTADENA
355|ALTAIR
356|ALTAMAHAW
357|ALTAMONT
358|ALTAMONTE SPRINGS
359|ALTAVILLE
360|ALTAVISTA
361|ALTENBURG
362|ALTHA
363|ALTHEIMER
364|ALTMAR
365|ALTO
366|ALTO PASS
367|ALTON
368|ALTONA
369|ALTOONA
370|ALTURA
371|ALTURAS
372|ALTUS
373|ALUM BANK
374|ALUM BRIDGE
375|ALUM CREEK
376|ALUM ROCK
377|ALVA
378|ALVARADO
379|ALVATON
380|ALVIN
381|ALVO
382|ALVORD
383|ALVORDTON
384|ALVWOOD
385|ALZADA
386|AMA
387|AMADO
388|AMADOR CITY
389|AMAGANSETT
390|AMAGON
391|AMALGA
392|AMANA
393|AMANDA
394|AMANDA PARK
395|AMARGOSA COLONIA
396|AMARGOSA VALLEY
397|AMARILLO
398|AMASA
399|AMAWALK
400|AMAYA COLONIA
401|AMAZONIA
402|AMBER
403|AMBERG
404|AMBERLEY
405|AMBIA
406|AMBLER
407|AMBOY
408|AMBRIDGE
409|AMBRIDGE HEIGHTS
410|AMBROSE
411|AMCHITKA
412|AMELIA
413|AMELIA CITY
414|AMELIA COURT HOUSE
415|AMENIA
416|AMERICAN BEACH
417|AMERICAN CANYON
418|AMERICAN FALLS
419|AMERICAN FORK
420|AMERICUS
421|AMERY
422|AMES
423|AMES LAKE
424|AMESTI
425|AMESVILLE
426|AMHERST
427|AMHERST CENTER
428|AMHERST JUNCTION
429|AMHERSTDALE
430|AMIDON
431|AMIRET
432|AMISTAD
433|AMISTAD ACRES
434|AMITE
435|AMITY
436|AMITY GARDENS
437|AMITYVILLE
438|AMMON
439|AMO
440|AMONATE
441|AMORET
442|AMORITA
443|AMORY
444|AMSDEN
445|AMSTERDAM
446|AMY
447|ANACOCO
448|ANACONDA
449|ANACORTES
450|ANADARKO
451|ANAHEIM
452|ANAHOLA
453|ANAHUAC
454|ANAKTUVUK PASS
455|ANAMOOSE
456|ANAMOSA
457|ANANDALE
458|ANATONE
459|ANAWALT
460|ANCENEY
461|ANCHO
462|ANCHOR
463|ANCHOR BAY
464|ANCHOR POINT
465|ANCHORVILLE
466|ANCIENT OAKS
467|ANCOR
468|ANDALE
469|ANDALUSIA
470|ANDERSON
471|ANDERSONVILLE
472|ANDES
473|ANDING
474|ANDOVER
475|ANDREW
476|ANDREWS
477|ANDRIX
478|ANEGAM
479|ANETA
480|ANETH
481|ANGEL FIRE
482|ANGELA
483|ANGELES
484|ANGELICA
485|ANGELS CAMP
486|ANGELUS
487|ANGIE
488|ANGIER
489|ANGIOLA
490|ANGLE INLET
491|ANGLETON
492|ANGOLA
493|ANGOLA ON THE LAKE
494|ANGOON
495|ANGORA
496|ANGUILLA
497|ANGUS
498|ANGWIN
499|ANIAK
500|ANIMAS
501|ANIMAS COMUNIDAD
502|ANITA
503|ANIWA
504|ANKENY
505|ANKENYTOWN
506|ANKONA
507|ANMOORE
508|ANN ARBOR
509|ANNA
510|ANNA MARIA
511|ANNABELLA
512|ANNADA
513|ANNAMORIAH
514|ANNANDALE
515|ANNAPOLIS
516|ANNAWAN
517|ANNETA
518|ANNETTA
519|ANNETTA NORTH
520|ANNETTA SOUTH
521|ANNETTE
522|ANNEX
523|ANNISTON
524|ANNONA
525|ANNSVILLE
526|ANNVILLE
527|ANOKA
528|ANON RAICES COMUNIDAD
529|ANSELMA
530|ANSELMO
531|ANSLEY
532|ANSON
533|ANSONIA
534|ANSONVILLE
535|ANSTED
536|ANSTON
537|ANTARES
538|ANTELOPE
539|ANTELOPE HILLS
540|ANTHEM
541|ANTHON
542|ANTHONY
543|ANTHONYVILLE
544|ANTHOSTON
545|ANTIETAM
546|ANTIGO
547|ANTIMONY
548|ANTIOCH
549|ANTLER
550|ANTLERS
551|ANTOINE
552|ANTON
553|ANTON CHICO
554|ANTONIA
555|ANTONINO
556|ANTONITO
557|ANTREVILLE
558|ANTRIM
559|ANTWERP
560|ANTÓN RUIZ
561|ANTÓN RUÍZ COMUNIDAD
562|ANVIK
563|ANZA
564|APACHE
565|APACHE CREEK
566|APACHE JUNCTION
567|APALACHEE
568|APALACHICOLA
569|APALACHIN
570|APEX
571|APGAR
572|APISON
573|APLIN
574|APLINGTON
575|APOLLO
576|APOLLO BEACH
577|APOPKA
578|APPALACHIA
579|APPLE CANYON LAKE
580|APPLE CREEK
581|APPLE GROVE
582|APPLE MOUNTAIN LAKE
583|APPLE RIVER
584|APPLE SPRINGS
585|APPLE VALLEY
586|APPLEBY
587|APPLEGATE
588|APPLETON
589|APPLETON CITY
590|APPLEWOLD
591|APPLEWOOD
592|APPLING
593|APPOMATTOX
594|APSHAWA
595|APTAKISIC
596|APTOS
597|AQUA PARK
598|AQUADALE
599|AQUASCO
600|AQUEBOGUE
601|AQUIA HARBOUR
602|AQUILLA
603|ARAB
604|ARABI
605|ARABIA
606|ARAGON
607|ARANSAS PASS
608|ARAPAHO
609|ARAPAHOE
610|ARARAT
611|ARBELA
612|ARBOLES
613|ARBON
614|ARBOR HILL
615|ARBOVALE
616|ARBUCKLE
617|ARBURY HILLS
618|ARBUTUS
619|ARBYRD
620|ARCADE
621|ARCADIA
622|ARCADIA LAKES
623|ARCANUM
624|ARCATA
625|ARCH CAPE
626|ARCHBALD
627|ARCHBOLD
628|ARCHDALE
629|ARCHER
630|ARCHER CITY
631|ARCHER LODGE
632|ARCHIBALD
633|ARCHIE
634|ARCHVILLE
635|ARCO
636|ARCOLA
637|ARCTIC VILLAGE
638|ARDARA
639|ARDEN
640|ARDEN HILLS
641|ARDEN ON THE SEVERN
642|ARDEN TOWN
643|ARDENCROFT
644|ARDENTOWN
645|ARDENVOIR
646|ARDMORE
647|ARDOCH
648|ARDSLEY
649|ARECIBO
650|ARECIBO ZONA URBANA
651|AREDALE
652|ARENA
653|ARENAS VALLEY
654|ARENDTSVILLE
655|ARENZVILLE
656|ARGENTA
657|ARGENTINE
658|ARGO
659|ARGONIA
660|ARGONNE
661|ARGOS
662|ARGUSVILLE
663|ARGYLE
664|ARIAL
665|ARIEL
666|ARIMO
667|ARION
668|ARIPEKA
669|ARIPINE
670|ARISPE
671|ARISTA
672|ARISTES
673|ARISTOCRAT RANCHETTES
674|ARITON
675|ARIVACA
676|ARIVACA JUNCTION
677|ARIZONA CITY
678|ARIZONA VILLAGE
679|ARJAY
680|ARKADELPHIA
681|ARKANA
682|ARKANSAS CITY
683|ARKANSAW
684|ARKDALE
685|ARKINDA
686|ARKOE
687|ARKOMA
688|ARKPORT
689|ARLEE
690|ARLETTA
691|ARLEY
692|ARLINGTON
693|ARLINGTON HEIGHTS
694|ARMA
695|ARMADA
696|ARMAGH
697|ARMBRUST
698|ARMIJO
699|ARMINGTON
700|ARMINTO
701|ARMONA
702|ARMONK
703|ARMOR
704|ARMOREL
705|ARMOUR
706|ARMSTRONG
707|ARMSTRONGS MILLS
708|ARNAUDVILLE
709|ARNEGARD
710|ARNETT
711|ARNEY
712|ARNO
713|ARNOLD
714|ARNOLD CITY
715|ARNOLD LINE
716|ARNOLD MILL
717|ARNOLDS PARK
718|ARNOLDSVILLE
719|ARNOT
720|ARNOTT
721|AROCK
722|AROMA PARK
723|AROMAS
724|ARONA
725|AROYA
726|ARP
727|ARPELAR
728|ARPIN
729|ARREDONDO
730|ARREY
731|ARRIBA
732|ARRINGTON
733|ARROW CREEK
734|ARROW POINT
735|ARROW ROCK
736|ARROWBEAR LAKE
737|ARROWHEAD HIGHLANDS
738|ARROWHEAD SPRINGS
739|ARROWSMITH
740|ARROYO
741|ARROYO COLORADO ESTATES COLONIA
742|ARROYO GARDENS
743|ARROYO GRANDE
744|ARROYO HONDO
745|ARROYO SECO
746|ARROYO ZONA URBANA
747|ART
748|ARTAS
749|ARTEMUS
750|ARTESIA
751|ARTESIA WELLS
752|ARTESIAN
753|ARTHUR
754|ARTHUR CITY
755|ARTOIS
756|ARTONDALE
757|ARUNDEL VILLAGE
758|ARVADA
759|ARVANA
760|ARVIN
761|ARVONIA
762|ASBURY
763|ASBURY LAKE
764|ASBURY PARK
765|ASCUTNEY
766|ASH FLAT
767|ASH FORK
768|ASH GROVE
769|ASHAROKEN
770|ASHAWAY
771|ASHBURN
772|ASHBY
773|ASHDOWN
774|ASHEBORO
775|ASHER
776|ASHERTON
777|ASHERVILLE
778|ASHEVILLE
779|ASHFORD
780|ASHIPPUN
781|ASHKUM
782|ASHLAND
783|ASHLAND CITY
784|ASHLAND HEIGHTS
785|ASHLEY
786|ASHLEY HEIGHTS
787|ASHMORE
788|ASHPORT
789|ASHTABULA
790|ASHTOLA
791|ASHTON
792|ASHVILLE
793|ASHWAUBENON
794|ASHWOOD
795|ASKEWVILLE
796|ASKOV
797|ASOTIN
798|ASPEN
799|ASPEN HILL
800|ASPEN PARK
801|ASPEN SPRINGS
802|ASPERMONT
803|ASPERS
804|ASPETUCK
805|ASPINWALL
806|ASSARIA
807|ASSINIPPI
808|ASSUMPTION
809|ASTATULA
810|ASTICO
811|ASTOR
812|ASTOR PARK
813|ASTORIA
814|ATALISSA
815|ATASCADERO
816|ATASCOCITA
817|ATCHISON
818|ATCO
819|ATEN
820|ATGLEN
821|ATHALIA
822|ATHELSTAN
823|ATHENA
824|ATHENS
825|ATHERTON
826|ATHERTONVILLE
827|ATHOL
828|ATHOL SPRINGS
829|ATKA
830|ATKINS
831|ATKINSON
832|ATKINSON MILLS
833|ATLANTA
834|ATLANTIC
835|ATLANTIC BEACH
836|ATLANTIC CITY
837|ATLANTIC HIGHLANDS
838|ATLANTIS
839|ATLAS
840|ATLASBURG
841|ATMAUTLUAK
842|ATMORE
843|ATOKA
844|ATOLIA
845|ATOMIC CITY
846|ATQASUK
847|ATSION
848|ATTALLA
849|ATTAPULGUS
850|ATTICA
851|ATTLEBORO
852|ATTU
853|ATWATER
854|ATWOOD
855|AU GRES
856|AU SABLE
857|AU SABLE FORKS
858|AU TRAIN
859|AUBERRY
860|AUBREY
861|AUBURN
862|AUBURN HILLS
863|AUBURN LAKE TRAILS
864|AUBURNDALE
865|AUBURNTOWN
866|AUCILLA
867|AUDUBON
868|AUDUBON PARK
869|AUGUST
870|AUGUSTA
871|AUGUSTA SPRINGS
872|AUGUSTUS
873|AUKE BAY
874|AULANDER
875|AULLVILLE
876|AULNE
877|AULT
878|AUMSVILLE
879|AURA
880|AURELIA
881|AURORA
882|AURORA CENTER
883|AURORA LODGE
884|AURORAVILLE
885|AUSTELL
886|AUSTIN
887|AUSTINBURG
888|AUSTINTOWN
889|AUSTINVILLE
890|AUSTONIO
891|AUSTWELL
892|AUTAUGAVILLE
893|AUTRYVILLE
894|AUVERGNE
895|AUXIER
896|AUXVASSE
897|AVA
898|AVALON
899|AVALON BEACH
900|AVANT
901|AVARD
902|AVAWAM
903|AVELLA
904|AVENAL
905|AVENEL
906|AVENTURA
907|AVENUE
908|AVERA
909|AVERILL
910|AVERILL PARK
911|AVERY
912|AVERY CREEK
913|AVERY ISLAND
914|AVILA BEACH
915|AVILLA
916|AVINGER
917|AVIS
918|AVISTON
919|AVOCA
920|AVOCADO HEIGHTS
921|AVON
922|AVON HEIGHTS
923|AVON LAKE
924|AVON PARK
925|AVON-BY-THE-SEA
926|AVONDALE
927|AVONDALE ESTATES
928|AVONIA
929|AVONMORE
930|AVRA VALLEY
931|AWENDAW
932|AWOSTING
933|AXIS
934|AXSON
935|AXTELL
936|AXTON
937|AYDEN
938|AYER
939|AYLMER
940|AYNOR
941|AYR
942|AYRSHIRE
943|AZALEA PARK
944|AZALIA
945|AZLE
946|AZTEC
947|AZURE
948|AZUSA
949|AZWELL
950|AÑASCO
951|AÑASCO ZONA URBANA
952|B AND E COLONIA
953|BABB
954|BABBIE
955|BABBITT
956|BABBS
957|BABCOCK
958|BABSON PARK
959|BABYLON
960|BACAVI
961|BACH
962|BACKUS
963|BACKUS BEACH
964|BACLIFF
965|BACONTON
966|BACOVA
967|BACTON
968|BAD AXE
969|BADEN
970|BADGER
971|BADIN
972|BAGDAD
973|BAGGS
974|BAGLEY
975|BAGNELL
976|BAGTOWN
977|BAGWELL
978|BAHAMA
979|BAIDLAND
980|BAIE DE WASAI
981|BAILEY
982|BAILEY LAKE
983|BAILEY PRAIRIE
984|BAILEYS CROSSROADS
985|BAILEYS HARBOR
986|BAILEYTON
987|BAILEYVILLE
988|BAINBRIDGE
989|BAINBRIDGE ISLAND
990|BAINS
991|BAINVILLE
992|BAIRD
993|BAIRDFORD
994|BAIRDSTOWN
995|BAIROA
996|BAIROA LA VEINTICINCO COMUNIDAD
997|BAIROIL
998|BAITING HOLLOW
999|BAJADERO
1000|BAJADERO COMUNIDAD
1001|BAJANDAS
1002|BAJANDAS COMUNIDAD
1003|BAKER
1004|BAKER CITY
1005|BAKER HILL
1006|BAKERS MILL
1007|BAKERSFIELD
1008|BAKERSTOWN
1009|BAKERSTOWN STATION
1010|BAKERSVILLE
1011|BAKERTON
1012|BAL HARBOUR
1013|BALA
1014|BALA-CYNWYD
1015|BALANCE ROCK
1016|BALATON
1017|BALCH SPRINGS
1018|BALCOM
1019|BALCONES HEIGHTS
1020|BALD CREEK
1021|BALD EAGLE
1022|BALD HEAD ISLAND
1023|BALD KNOB
1024|BALDRIDGE
1025|BALDWIN
1026|BALDWIN CITY
1027|BALDWIN HARBOR
1028|BALDWIN PARK
1029|BALDWINSVILLE
1030|BALDWINVILLE
1031|BALDWYN
1032|BALFOUR
1033|BALKO
1034|BALL
1035|BALL CLUB
1036|BALL GROUND
1037|BALLANTINE
1038|BALLARD
1039|BALLARDVALE
1040|BALLENGER CREEK
1041|BALLENTINE
1042|BALLICO
1043|BALLINGER
1044|BALLOU
1045|BALLPLAY
1046|BALLSTON SPA
1047|BALLTOWN
1048|BALLVILLE
1049|BALLWIN
1050|BALLY
1051|BALM
1052|BALMORHEA
1053|BALMVILLE
1054|BALSAM
1055|BALSAM LAKE
1056|BALTA
1057|BALTIC
1058|BALTIMORE
1059|BALTIMORE HIGHLANDS
1060|BAMBERG
1061|BAMMEL
1062|BANCROFT
1063|BANDANA
1064|BANDERA
1065|BANDERA FALLS
1066|BANDON
1067|BANEBERRY
1068|BANGOR
1069|BANGS
1070|BANIDA
1071|BANK LICK
1072|BANKS
1073|BANKS SPRINGS
1074|BANKSTON
1075|BANNACK
1076|BANNER
1077|BANNER ELK
1078|BANNER HILL
1079|BANNERTOWN
1080|BANNING
1081|BANNOCK
1082|BANNOCKBURN
1083|BANQUETE
1084|BANTAM
1085|BANTRY
1086|BAR HARBOR
1087|BAR MILLS
1088|BAR NUNN
1089|BARABOO
1090|BARADA
1091|BARAGA
1092|BARAHONA
1093|BARAHONA COMUNIDAD
1094|BARANOF
1095|BARATARIA
1096|BARBER
1097|BARBERTON
1098|BARBERVILLE
1099|BARBOURMEADE
1100|BARBOURS
1101|BARBOURSVILLE
1102|BARBOURVILLE
1103|BARCELONETA
1104|BARCELONETA ZONA URBANA
1105|BARCLAY
1106|BARCO
1107|BARD
1108|BARDEN
1109|BARDLEY
1110|BARDOLPH
1111|BARDONIA
1112|BARDSTOWN
1113|BARDWELL
1114|BAREVILLE
1115|BARGERSVILLE
1116|BARING
1117|BARK RANCH
1118|BARK RIVER
1119|BARKER
1120|BARKER HEIGHTS
1121|BARKER TEN MILE
1122|BARKEYVILLE
1123|BARKSDALE
1124|BARLING
1125|BARLOW
1126|BARNABUS
1127|BARNARD
1128|BARNEGAT
1129|BARNEGAT LIGHT
1130|BARNES
1131|BARNES CITY
1132|BARNESTON
1133|BARNESVILLE
1134|BARNET
1135|BARNETT
1136|BARNEVELD
1137|BARNEY
1138|BARNHART
1139|BARNHILL
1140|BARNSBORO
1141|BARNSDALL
1142|BARNSTABLE
1143|BARNUM
1144|BARNUM ISLAND
1145|BARNWELL
1146|BARODA
1147|BARON
1148|BARR
1149|BARRACKS
1150|BARRACKVILLE
1151|BARRANQUITAS
1152|BARRANQUITAS ZONA URBANA
1153|BARRE
1154|BARRELVILLE
1155|BARRETTS
1156|BARRINEAU PARK
1157|BARRINGTON
1158|BARRINGTON HILLS
1159|BARRINGTON WOODS
1160|BARRON
1161|BARRONETT
1162|BARROWS
1163|BARRVILLE
1164|BARRY
1165|BARRYTON
1166|BARRYVILLE
1167|BARSTOW
1168|BARTELSO
1169|BARTLES
1170|BARTLESVILLE
1171|BARTLETT
1172|BARTLEY
1173|BARTOLO
1174|BARTOLO COMUNIDAD
1175|BARTON
1176|BARTON CREEK
1177|BARTON HILLS
1178|BARTONSVILLE
1179|BARTONVILLE
1180|BARTOW
1181|BARVIEW
1182|BARWICK
1183|BASALT
1184|BASCO
1185|BASCOM
1186|BASEHOR
1187|BASIC
1188|BASILE
1189|BASIN
1190|BASIN CITY
1191|BASINGER
1192|BASKERVILLE
1193|BASKETT
1194|BASKIN
1195|BASKING RIDGE
1196|BASS HARBOR
1197|BASS LAKE
1198|BASSETT
1199|BASSFIELD
1200|BASSVILLE PARK
1201|BASTIAN
1202|BASTROP
1203|BASYE
1204|BATAVIA
1205|BATCHELOR
1206|BATCHTOWN
1207|BATES
1208|BATES CITY
1209|BATESBURG-LEESVILLE
1210|BATESLAND
1211|BATESVILLE
1212|BATH CORNER
1213|BATHGATE
1214|BATON ROUGE
1215|BATSON
1216|BATTLE CREEK
1217|BATTLE GROUND
1218|BATTLE LAKE
1219|BATTLE MOUNTAIN
1220|BATTLEBORO
1221|BATTLEFIELD
1222|BATTLEMENT MESA
1223|BATTLES
1224|BATTLETOWN
1225|BAUDETTE
1226|BAUERSTOWN
1227|BAUMSTOWN
1228|BAUTISTA
1229|BAUXITE
1230|BAVARIA
1231|BAWCOMVILLE
1232|BAXLEY
1233|BAXTER
1234|BAXTER ESTATES
1235|BAXTER SPRINGS
1236|BAXTERVILLE
1237|BAY
1238|BAY CENTER
1239|BAY CITY
1240|BAY HARBOR ISLANDS
1241|BAY HEAD
1242|BAY HILL
1243|BAY LAKE
1244|BAY MINETTE
1245|BAY PARK
1246|BAY PINES
1247|BAY POINT
1248|BAY PORT
1249|BAY RIDGE
1250|BAY SAINT LOUIS
1251|BAY SHORE
1252|BAY SPRINGS
1253|BAY VIEW
1254|BAY VIEW GARDEN
1255|BAY VILLAGE
1256|BAY WOOD
1257|BAYAMÓN
1258|BAYAMÓN COMUNIDAD
1259|BAYAMÓN ZONA URBANA
1260|BAYARD
1261|BAYBORO
1262|BAYFIELD
1263|BAYLIS
1264|BAYNE
1265|BAYONET POINT
1266|BAYONNE
1267|BAYOU CANE
1268|BAYOU CHICOT
1269|BAYOU CORNE
1270|BAYOU GAUCHE
1271|BAYOU GEORGE
1272|BAYOU GOULA
1273|BAYOU LA BATRE
1274|BAYOU METO
1275|BAYOU SORREL
1276|BAYOU VISTA
1277|BAYPORT
1278|BAYSHORE
1279|BAYSHORE GARDENS
1280|BAYSIDE
1281|BAYSIDE BEACH
1282|BAYSIDE GARDENS
1283|BAYSIDE TERRACE
1284|BAYTOWN
1285|BAYVIEW
1286|BAYVILLE
1287|BAZEMORE
1288|BAZILE MILLS
1289|BAZINE
1290|BEACH CITY
1291|BEACH GLEN
1292|BEACH HAVEN
1293|BEACH HAVEN WEST
1294|BEACH LAKE
1295|BEACH PARK
1296|BEACH RIDGE
1297|BEACHWOOD
1298|BEACON
1299|BEACON HILL
1300|BEACON SQUARE
1301|BEACONSFIELD
1302|BEAGLE
1303|BEAL CITY
1304|BEALETON
1305|BEALLSVILLE
1306|BEAMAN
1307|BEAN STATION
1308|BEAR
1309|BEAR CREEK
1310|BEAR CREEK VILLAGE
1311|BEAR DANCE
1312|BEAR FLAT
1313|BEAR GRASS
1314|BEAR LAKE
1315|BEAR RIVER
1316|BEAR RIVER CITY
1317|BEAR ROCKS
1318|BEAR VALLEY
1319|BEAR VALLEY SPRINGS
1320|BEARCREEK
1321|BEARDEN
1322|BEARDS FORK
1323|BEARDSLEY
1324|BEARDSTOWN
1325|BEARMOUTH
1326|BEASLEY
1327|BEASON
1328|BEATRICE
1329|BEATTIE
1330|BEATTY
1331|BEATTYSTOWN
1332|BEATTYVILLE
1333|BEAUFORT
1334|BEAULIEU
1335|BEAUMONT
1336|BEAUMONT PLACE
1337|BEAUREGARD
1338|BEAUX ARTS VILLAGE
1339|BEAVER
1340|BEAVER BAY
1341|BEAVER CITY
1342|BEAVER CREEK
1343|BEAVER CROSSING
1344|BEAVER DAM
1345|BEAVER DAM LAKE
1346|BEAVER FALLS
1347|BEAVER MEADOWS
1348|BEAVER SPRINGS
1349|BEAVER VALLEY
1350|BEAVERCREEK
1351|BEAVERDALE
1352|BEAVERDAM
1353|BEAVERLICK
1354|BEAVERTON
1355|BEAVERTOWN
1356|BEAVERVILLE
1357|BEBE
1358|BECHTELSVILLE
1359|BECHYN
1360|BECIDA
1361|BECKEMEYER
1362|BECKER
1363|BECKETT
1364|BECKETT RIDGE
1365|BECKLEY
1366|BECKVILLE
1367|BECKWOURTH
1368|BECLABITO
1369|BECTON
1370|BEDA
1371|BEDFORD
1372|BEDFORD CENTER
1373|BEDFORD HEIGHTS
1374|BEDFORD HILLS
1375|BEDFORD PARK
1376|BEDIAS
1377|BEDMINSTER
1378|BEDROCK
1379|BEE BRANCH
1380|BEE CAVE
1381|BEE RIDGE
1382|BEE SPRING
1383|BEEBE
1384|BEECH BLUFF
1385|BEECH BOTTOM
1386|BEECH CREEK
1387|BEECH GROVE
1388|BEECH MOUNTAIN
1389|BEECH MOUNTAIN LAKES
1390|BEECHBURG
1391|BEECHER
1392|BEECHER CITY
1393|BEECHER FALLS
1394|BEECHGROVE
1395|BEECHMONT
1396|BEECHWOOD
1397|BEECHWOOD TRAILS
1398|BEECHWOOD VILLAGE
1399|BEEDEVILLE
1400|BEEKMAN
1401|BEELER
1402|BEEMER
1403|BEEMERVILLE
1404|BEERSHEBA SPRINGS
1405|BEEVILLE
1406|BEGGS
1407|BEIRNE
1408|BEJOU
1409|BEL AIR
1410|BEL ALTON
1411|BEL-NOR
1412|BEL-RIDGE
1413|BELCAMP
1414|BELCHER
1415|BELCHERTOWN
1416|BELCHERVILLE
1417|BELCOURT
1418|BELDEN
1419|BELDING
1420|BELEN
1421|BELFAIR
1422|BELFALLS
1423|BELFAST
1424|BELFIELD
1425|BELFONTE
1426|BELFORD
1427|BELFRY
1428|BELGIQUE
1429|BELGIUM
1430|BELGRADE
1431|BELGREEN
1432|BELHAVEN
1433|BELINDA CITY
1434|BELINGTON
1435|BELK
1436|BELKNAP
1437|BELKOFSKI
1438|BELL ACRES
1439|BELL ARTHUR
1440|BELL BUCKLE
1441|BELL CENTER
1442|BELL CITY
1443|BELL GARDENS
1444|BELL HILL
1445|BELL ISLAND HOT SPRINGS
1446|BELL POINT
1447|BELLA VILLA
1448|BELLA VISTA
1449|BELLAIRE
1450|BELLAMY
1451|BELLBROOK
1452|BELLE
1453|BELLE CENTER
1454|BELLE CHASSE
1455|BELLE FOURCHE
1456|BELLE GLADE
1457|BELLE HAVEN
1458|BELLE ISLE
1459|BELLE MEAD
1460|BELLE MEADE
1461|BELLE PLAINE
1462|BELLE PRAIRIE CITY
1463|BELLE RIVE
1464|BELLE ROSE
1465|BELLE TERRE
1466|BELLE VALLEY
1467|BELLE VERNON
1468|BELLEAIR
1469|BELLEAIR BEACH
1470|BELLEAIR BLUFFS
1471|BELLEAIR SHORES
1472|BELLECHESTER
1473|BELLEFONT
1474|BELLEFONTAINE
1475|BELLEFONTAINE NEIGHBORS
1476|BELLEFONTE
1477|BELLEMEADE
1478|BELLEMONT
1479|BELLEPLAIN
1480|BELLERIVE ACRES
1481|BELLEROSE
1482|BELLEROSE TERRACE
1483|BELLEVIEW
1484|BELLEVILLE
1485|BELLEVUE
1486|BELLEWOOD
1487|BELLFLOWER
1488|BELLFOUNTAIN
1489|BELLINGHAM
1490|BELLMAWR
1491|BELLMEAD
1492|BELLMONT
1493|BELLMORE
1494|BELLOWS FALLS
1495|BELLPORT
1496|BELLTOWN
1497|BELLVALE
1498|BELLVIEW
1499|BELLVILLE
1500|BELLVUE
1501|BELLWOOD
1502|BELMAR
1503|BELMOND
1504|BELMONT
1505|BELMONT ESTATES
1506|BELMORE
1507|BELOIT
1508|BELPRE
1509|BELSPRING
1510|BELTON
1511|BELTRAMI
1512|BELTSVILLE
1513|BELUGA
1514|BELVA
1515|BELVEDERE
1516|BELVEDERE PARK
1517|BELVIDERE
1518|BELVIEW
1519|BELVILLE
1520|BELVOIR
1521|BELVUE
1522|BELWOOD
1523|BELZONI
1524|BEMENT
1525|BEMIDJI
1526|BEMIS
1527|BEMISS
1528|BEMUS POINT
1529|BEN ARNOLD
1530|BEN AVON
1531|BEN AVON HEIGHTS
1532|BEN BOLT
1533|BEN HUR
1534|BEN LOMOND
1535|BEN WHEELER
1536|BENA
1537|BENAVIDES
1538|BENBOW
1539|BENBROOK
1540|BENCHLAND
1541|BENCHLEY
1542|BENDAVIS
1543|BENDENA
1544|BENDERSVILLE
1545|BENDERVILLE
1546|BENDON
1547|BENEDICT
1548|BENEVOLENCE
1549|BENGAL
1550|BENGE
1551|BENHAM
1552|BENICIA
1553|BENITEZ
1554|BENJAMIN
1555|BENKELMAN
1556|BENLD
1557|BENNDALE
1558|BENNET
1559|BENNETT
1560|BENNETT SPRINGS
1561|BENNETTS CORNERS
1562|BENNETTS MILLS
1563|BENNETTSVILLE
1564|BENNINGTON
1565|BENNION
1566|BENNS CHURCH
1567|BENOIT
1568|BENONINE
1569|BENS RUN
1570|BENSALEM
1571|BENSENVILLE
1572|BENSLEY
1573|BENSON
1574|BENT
1575|BENT CREEK
1576|BENTLEY
1577|BENTLEYVILLE
1578|BENTON
1579|BENTON CITY
1580|BENTON HARBOR
1581|BENTON HEIGHTS
1582|BENTON RIDGE
1583|BENTONIA
1584|BENTONVILLE
1585|BENWOOD
1586|BENZONIA
1587|BENÍTEZ COMUNIDAD
1588|BEOWAWE
1589|BERCLAIR
1590|BEREA
1591|BEREAH
1592|BERENDA
1593|BERENICE
1594|BERESFORD
1595|BERGEN
1596|BERGEN PARK
1597|BERGENFIELD
1598|BERGER
1599|BERGHOLTZ
1600|BERGHOLZ
1601|BERGLAND
1602|BERGMAN
1603|BERGOO
1604|BERGTON
1605|BERINO
1606|BERKELEY
1607|BERKELEY LAKE
1608|BERKELEY SPRINGS
1609|BERKEY
1610|BERKLEY
1611|BERLIN
1612|BERLIN HEIGHTS
1613|BERMUDA DUNES
1614|BERMUDA RUN
1615|BERN
1616|BERNALILLO
1617|BERNARD
1618|BERNARDO
1619|BERNARDSVILLE
1620|BERNE
1621|BERNECKER
1622|BERNICE
1623|BERNIE
1624|BERNSTADT
1625|BERNSTEIN
1626|BERNVILLE
1627|BEROUN
1628|BERRIEN SPRINGS
1629|BERRY
1630|BERRY CREEK
1631|BERRY HILL
1632|BERRYDALE
1633|BERRYSBURG
1634|BERRYVILLE
1635|BERTHA
1636|BERTHOLD
1637|BERTHOUD
1638|BERTRAM
1639|BERTRAND
1640|BERTRANDVILLE
1641|BERVILLE
1642|BERWICK
1643|BERWIND
1644|BERWYN
1645|BERWYN HEIGHTS
1646|BERYL
1647|BERYL JUNCTION
1648|BESSEMER
1649|BESSEMER BEND
1650|BESSEMER CITY
1651|BESSIE
1652|BESSMAY
1653|BEST
1654|BETANCES
1655|BETANCES COMUNIDAD
1656|BETE GRISE
1657|BETHALTO
1658|BETHANIA
1659|BETHANY
1660|BETHANY BEACH
1661|BETHAYRES
1662|BETHEDEN
1663|BETHEL
1664|BETHEL ACRES
1665|BETHEL HEIGHTS
1666|BETHEL ISLAND
1667|BETHEL PARK
1668|BETHEL SPRINGS
1669|BETHERA
1670|BETHESDA
1671|BETHLEHEM
1672|BETHPAGE
1673|BETHUNE
1674|BETSY LAYNE
1675|BETTENDORF
1676|BETTERAVIA
1677|BETTERTON
1678|BETTIE
1679|BETTLES
1680|BETTSVILLE
1681|BETWEEN
1682|BEULAH
1683|BEULAH BEACH
1684|BEULAH VALLEY
1685|BEULAVILLE
1686|BEURYS LAKE
1687|BEVERLY
1688|BEVERLY BEACH
1689|BEVERLY HILLS
1690|BEVERLY SHORES
1691|BEVIER
1692|BEVIL OAKS
1693|BEVINGTON
1694|BEVIS
1695|BEWLEYVILLE
1696|BEXAR
1697|BEXLEY
1698|BEYERVILLE
1699|BIBO
1700|BICKLETON
1701|BICKNELL
1702|BIDDEFORD
1703|BIDDLE
1704|BIEBER
1705|BIEHLE
1706|BIENVILLE
1707|BIER
1708|BIG ARM
1709|BIG BAR
1710|BIG BASS LAKE
1711|BIG BAY
1712|BIG BEAR CITY
1713|BIG BEAR LAKE
1714|BIG BEAVER
1715|BIG BEND
1716|BIG BEND CITY
1717|BIG BOW
1718|BIG CABIN
1719|BIG CHIMNEY
1720|BIG CLIFTY
1721|BIG COPPITT KEY
1722|BIG CREEK
1723|BIG DELTA
1724|BIG FALLS
1725|BIG FLAT
1726|BIG FLATS
1727|BIG FORK
1728|BIG HORN
1729|BIG ISLAND
1730|BIG LAGOON
1731|BIG LAKE
1732|BIG MOOSE
1733|BIG OAK FLAT
1734|BIG PINE
1735|BIG PINE KEY
1736|BIG PINEY
1737|BIG PLAIN
1738|BIG POINT
1739|BIG POOL
1740|BIG PRAIRIE
1741|BIG RAPIDS
1742|BIG RIVER
1743|BIG ROCK
1744|BIG RUN
1745|BIG SANDY
1746|BIG SKY
1747|BIG SPRING
1748|BIG SPRINGS
1749|BIG STONE CITY
1750|BIG STONE GAP
1751|BIG SUR
1752|BIG TIMBER
1753|BIG TREE
1754|BIG WATER
1755|BIG WELLS
1756|BIGBEE
1757|BIGBEE VALLEY
1758|BIGELOW
1759|BIGFOOT
1760|BIGFORK
1761|BIGGERS
1762|BIGGERSVILLE
1763|BIGGS
1764|BIGGS JUNCTION
1765|BIGGSVILLE
1766|BIGHORN
1767|BIGLER
1768|BIGLERVILLE
1769|BIJOU HILLS
1770|BILL
1771|BILL MOORES
1772|BILLETT
1773|BILLINGS
1774|BILLINGSLEY
1775|BILLINGTON HEIGHTS
1776|BILOXI
1777|BILTMORE FOREST
1778|BINFORD
1779|BINGEN
1780|BINGER
1781|BINGHAM
1782|BINGHAM FARMS
1783|BINGHAM LAKE
1784|BINGHAMTON
1785|BIOLA
1786|BIORKA
1787|BIPPUS
1788|BIRCH BAY
1789|BIRCH CREEK
1790|BIRCH RIVER
1791|BIRCH RUN
1792|BIRCH TREE
1793|BIRCHWOOD
1794|BIRCHWOOD LAKES
1795|BIRD CITY
1796|BIRD IN HAND
1797|BIRD ISLAND
1798|BIRDS LANDING
1799|BIRDSBORO
1800|BIRDSEYE
1801|BIRDSONG
1802|BIRDSVILLE
1803|BIRMINGHAM
1804|BIRNAMWOOD
1805|BIRNEY
1806|BIRON
1807|BIRTA
1808|BISBEE
1809|BISCAY
1810|BISCAYNE PARK
1811|BISCOE
1812|BISHOP
1813|BISHOP HILL
1814|BISHOP HILLS
1815|BISHOPVILLE
1816|BISMARCK
1817|BISON
1818|BISSELL
1819|BITELY
1820|BITHLO
1821|BITTER CREEK
1822|BITTER SPRINGS
1823|BIVALVE
1824|BIVINS
1825|BIWABIK
1826|BIXBY
1827|BLACK
1828|BLACK BUTTE RANCH
1829|BLACK CANYON CITY
1830|BLACK CREEK
1831|BLACK DIAMOND
1832|BLACK EAGLE
1833|BLACK EARTH
1834|BLACK FOREST
1835|BLACK FORK
1836|BLACK HAWK
1837|BLACK JACK
1838|BLACK LICK
1839|BLACK MOUNTAIN
1840|BLACK OAK
1841|BLACK POINT
1842|BLACK RIVER
1843|BLACK RIVER FALLS
1844|BLACK RIVER VILLAGE
1845|BLACK ROCK
1846|BLACK SPRINGS
1847|BLACK WALNUT
1848|BLACKBERRY
1849|BLACKBURN
1850|BLACKDUCK
1851|BLACKEY
1852|BLACKFOOT
1853|BLACKFORD
1854|BLACKGUM
1855|BLACKHAWK
1856|BLACKHORSE
1857|BLACKLICK ESTATES
1858|BLACKMAN
1859|BLACKSBURG
1860|BLACKSHEAR
1861|BLACKSTOCK
1862|BLACKSTONE
1863|BLACKSVILLE
1864|BLACKTON
1865|BLACKVILLE
1866|BLACKWATER
1867|BLACKWELL
1868|BLACKWELLS
1869|BLACKWELLS MILLS
1870|BLACKWOOD
1871|BLADEN
1872|BLADENBORO
1873|BLADENSBURG
1874|BLADES
1875|BLAIN
1876|BLAINE
1877|BLAINE HILL
1878|BLAIR
1879|BLAIRS
1880|BLAIRS MILLS
1881|BLAIRSBURG
1882|BLAIRSDEN
1883|BLAIRSTOWN
1884|BLAIRSVILLE
1885|BLAIRVILLE
1886|BLAISDELL
1887|BLAKELEY
1888|BLAKELY
1889|BLAKEMAN
1890|BLAKESBURG
1891|BLAKESLEE
1892|BLANCA
1893|BLANCHARD
1894|BLANCHARDVILLE
1895|BLANCHE
1896|BLANCHESTER
1897|BLANCO
1898|BLAND
1899|BLANDBURG
1900|BLANDFORD
1901|BLANDING
1902|BLANDINSVILLE
1903|BLANDON
1904|BLANDVILLE
1905|BLANFORD
1906|BLANKET
1907|BLANTON
1908|BLASDELL
1909|BLAUVELT
1910|BLAWENBURG
1911|BLAWNOX
1912|BLEAKWOOD
1913|BLEDSOE
1914|BLEECKER
1915|BLENCOE
1916|BLENDE
1917|BLENHEIM
1918|BLENNERHASSETT
1919|BLESSING
1920|BLEVINS
1921|BLEWETT
1922|BLISS
1923|BLISS CORNER
1924|BLISSFIELD
1925|BLITCHTON
1926|BLOCHER
1927|BLOCKHOUSE
1928|BLOCKSBURG
1929|BLOCKTON
1930|BLODGETT
1931|BLODGETT LANDING
1932|BLODGETT MILLS
1933|BLOMKEST
1934|BLOOM
1935|BLOOM CITY
1936|BLOOMBURG
1937|BLOOMDALE
1938|BLOOMER
1939|BLOOMFIELD
1940|BLOOMFIELD HILLS
1941|BLOOMING GROVE
1942|BLOOMING PRAIRIE
1943|BLOOMING VALLEY
1944|BLOOMINGBURG
1945|BLOOMINGDALE
1946|BLOOMINGTON
1947|BLOOMSBURG
1948|BLOOMSBURY
1949|BLOOMSDALE
1950|BLOOMVILLE
1951|BLOSSBURG
1952|BLOSSOM
1953|BLOUNTSTOWN
1954|BLOUNTSVILLE
1955|BLOUNTVILLE
1956|BLOWING ROCK
1957|BLOXOM
1958|BLUE ANCHOR
1959|BLUE ASH
1960|BLUE BALL
1961|BLUE BELL
1962|BLUE BERRY HILL
1963|BLUE CANYON
1964|BLUE CREEK
1965|BLUE DIAMOND
1966|BLUE EARTH
1967|BLUE EYE
1968|BLUE GRASS
1969|BLUE HILL
1970|BLUE HILLS
1971|BLUE ISLAND
1972|BLUE JAY
1973|BLUE LAKE
1974|BLUE MOUND
1975|BLUE MOUNDS
1976|BLUE MOUNTAIN
1977|BLUE MOUNTAIN BEACH
1978|BLUE POINT
1979|BLUE RAPIDS
1980|BLUE RIDGE
1981|BLUE RIDGE MANOR
1982|BLUE RIDGE SHORES
1983|BLUE RIDGE SUMMIT
1984|BLUE RIVER
1985|BLUE ROCK
1986|BLUE SPRINGS
1987|BLUEBELL
1988|BLUEBERRY
1989|BLUEFIELD
1990|BLUEJACKET
1991|BLUETOWN
1992|BLUETOWN COLONIA
1993|BLUEWATER
1994|BLUEWELL
1995|BLUFF
1996|BLUFF CITY
1997|BLUFF DALE
1998|BLUFF PARK
1999|BLUFF SPRINGS
2000|BLUFFDALE
2001|BLUFFS
2002|BLUFFSIDE
2003|BLUFFTON
2004|BLUFFVIEW
2005|BLUFORD
2006|BLUM
2007|BLUMENTHAL
2008|BLUNT
2009|BLY
2010|BLYN
2011|BLYTHE
2012|BLYTHEDALE
2013|BLYTHEVILLE
2014|BLYTHEWOOD
2015|BOALSBURG
2016|BOARD CAMP
2017|BOARDMAN
2018|BOATMAN
2019|BOAZ
2020|BOBO
2021|BOBTOWN
2022|BOCA GRANDE
2023|BOCA RATON
2024|BOCK
2025|BODCAW
2026|BODE
2027|BODEGA
2028|BODEGA BAY
2029|BODEN
2030|BODFISH
2031|BOELUS
2032|BOERNE
2033|BOGALUSA
2034|BOGARD
2035|BOGART
2036|BOGATA
2037|BOGER CITY
2038|BOGIA
2039|BOGOTA
2040|BOGUE
2041|BOGUE CHITTO
2042|BOHEMIA
2043|BOHNERS LAKE
2044|BOHON
2045|BOICOURT
2046|BOILING SPRING LAKES
2047|BOILING SPRINGS
2048|BOIS D'ARC
2049|BOISE
2050|BOISE CITY
2051|BOISTFORT
2052|BOKCHITO
2053|BOKEELIA
2054|BOKHOMA
2055|BOKOSHE
2056|BOLAIR
2057|BOLAN
2058|BOLCKOW
2059|BOLD SPRING
2060|BOLES
2061|BOLES ACRES
2062|BOLEY
2063|BOLIGEE
2064|BOLINAS
2065|BOLINDALE
2066|BOLING
2067|BOLINGBROKE
2068|BOLINGBROOK
2069|BOLINGER
2070|BOLIVAR
2071|BOLIVAR PENINSULA
2072|BOLIVIA
2073|BOLLING
2074|BOLT
2075|BOLTON
2076|BOLTON LANDING
2077|BOMA
2078|BOMARTON
2079|BOMBAY BEACH
2080|BON
2081|BON AIR
2082|BON AQUA JUNCTION
2083|BON HOMME COLONY
2084|BON MEADE
2085|BON SECOUR
2086|BON WIER
2087|BONAIRE
2088|BONANZA
2089|BONANZA MOUNTAIN ESTATES
2090|BONAPARTE
2091|BONCARBO
2092|BOND
2093|BONDAD
2094|BONDSVILLE
2095|BONDUEL
2096|BONDURANT
2097|BONDVILLE
2098|BONE GAP
2099|BONEAU
2100|BONESTEEL
2101|BONETRAILL
2102|BONFIELD
2103|BONHAM
2104|BONHOMIE
2105|BONIFAY
2106|BONILLA
2107|BONITA
2108|BONITA SPRINGS
2109|BONLEE
2110|BONNE TERRE
2111|BONNEAU
2112|BONNEAU BEACH
2113|BONNEAUVILLE
2114|BONNER
2115|BONNER SPRINGS
2116|BONNERS FERRY
2117|BONNETSVILLE
2118|BONNEVILLE
2119|BONNEY
2120|BONNEY LAKE
2121|BONNIE
2122|BONNIE DOONE
2123|BONNIEVILLE
2124|BONNOTS MILL
2125|BONNY DOON
2126|BONO
2127|BONSALL
2128|BOODY
2129|BOOKER
2130|BOOMER
2131|BOON
2132|BOONE
2133|BOONES MILL
2134|BOONEVILLE
2135|BOONSBORO
2136|BOONTON
2137|BOONVILLE
2138|BOOTH
2139|BOOTHBAY HARBOR
2140|BOOTHVILLE
2141|BOOTHWYN
2142|BOOTJACK
2143|BOQUERÓN
2144|BOQUERÓN COMUNIDAD
2145|BOQUET
2146|BOQUILLAS CROSSING
2147|BORDEAUX
2148|BORDELONVILLE
2149|BORDEN
2150|BORDEN SPRINGS
2151|BORDENTOWN
2152|BORDER
2153|BORDULAC
2154|BORGER
2155|BORING
2156|BORON
2157|BORONDA
2158|BORREGO SPRINGS
2159|BORTH
2160|BORTON
2161|BORUP
2162|BOSCHERTOWN
2163|BOSCO
2164|BOSCOBEL
2165|BOSLER
2166|BOSQUE
2167|BOSQUE FARMS
2168|BOSS
2169|BOSSIER CITY
2170|BOSTIC
2171|BOSTON
2172|BOSTON HARBOR
2173|BOSTON HEIGHTS
2174|BOSTONIA
2175|BOSTWICK
2176|BOSWELL
2177|BOSWORTH
2178|BOTHELL
2179|BOTHWELL
2180|BOTINES
2181|BOTKINS
2182|BOTNA
2183|BOTTINEAU
2184|BOULDER
2185|BOULDER CITY
2186|BOULDER CREEK
2187|BOULDER FLATS
2188|BOULDER HILL
2189|BOULDER JUNCTION
2190|BOULDER TOWN
2191|BOULEVARD
2192|BOULEVARD GARDENS
2193|BOULEVARD PARK
2194|BOULOGNE
2195|BOUND BROOK
2196|BOUNTIFUL
2197|BOURBON
2198|BOURBONNAIS
2199|BOURG
2200|BOURNE
2201|BOURNEVILLE
2202|BOUSE
2203|BOUTON
2204|BOUTTE
2205|BOVARD
2206|BOVEY
2207|BOVILL
2208|BOVINA
2209|BOW
2210|BOW MAR
2211|BOW VALLEY
2212|BOWBELLS
2213|BOWDEN
2214|BOWDLE
2215|BOWDOIN
2216|BOWDOINHAM
2217|BOWDON
2218|BOWDON JUNCTION
2219|BOWEN
2220|BOWER HILL
2221|BOWERS
2222|BOWERS BEACH
2223|BOWERS MILL
2224|BOWERSTON
2225|BOWERSVILLE
2226|BOWESMONT
2227|BOWIE
2228|BOWLEGS
2229|BOWLER
2230|BOWLES
2231|BOWLEYS QUARTERS
2232|BOWLING GREEN
2233|BOWLUS
2234|BOWMAN
2235|BOWMANS ADDITION
2236|BOWMANSTOWN
2237|BOWMANSVILLE
2238|BOWMONT
2239|BOWMORE
2240|BOWRING
2241|BOX
2242|BOX ELDER
2243|BOXELDER
2244|BOXFORD
2245|BOXHOLM
2246|BOY RIVER
2247|BOYCE
2248|BOYCEVILLE
2249|BOYD
2250|BOYDELL
2251|BOYDEN
2252|BOYDEN ARBOR
2253|BOYDS
2254|BOYDSTON
2255|BOYDSVILLE
2256|BOYDTON
2257|BOYER
2258|BOYERO
2259|BOYERS
2260|BOYERTOWN
2261|BOYES
2262|BOYES HOT SPRINGS
2263|BOYKIN
2264|BOYKINS
2265|BOYLE
2266|BOYNE CITY
2267|BOYNE FALLS
2268|BOYNTON
2269|BOYNTON BEACH
2270|BOYS RANCH
2271|BOYS TOWN
2272|BOYSEN
2273|BOZAR
2274|BOZEMAN
2275|BOZMAN
2276|BRACEVILLE
2277|BRACEY
2278|BRACHFIELD
2279|BRACKEN
2280|BRACKENRIDGE
2281|BRACKETT
2282|BRACKETTVILLE
2283|BRAD
2284|BRADBURY
2285|BRADDOCK
2286|BRADDOCK HEIGHTS
2287|BRADDOCK HILLS
2288|BRADDYVILLE
2289|BRADEN
2290|BRADENTON
2291|BRADENTON BEACH
2292|BRADENVILLE
2293|BRADFORD
2294|BRADFORD HILLS
2295|BRADFORD WOODS
2296|BRADFORDSVILLE
2297|BRADFORDVILLE
2298|BRADGATE
2299|BRADLEY
2300|BRADLEY BEACH
2301|BRADLEY GARDENS
2302|BRADLEY JUNCTION
2303|BRADLEYVILLE
2304|BRADNER
2305|BRADSHAW
2306|BRADY
2307|BRADY LAKE
2308|BRAGG CITY
2309|BRAGGADOCIO
2310|BRAGGS
2311|BRAHAM
2312|BRAIDWOOD
2313|BRAINARD
2314|BRAINARDS
2315|BRAINERD
2316|BRAITHWAITE
2317|BRAMAN
2318|BRAMBLETON
2319|BRAMPTON
2320|BRAMWELL
2321|BRANCH DALE
2322|BRANCH HILL
2323|BRANCHBURG PARK
2324|BRANCHLAND
2325|BRANCHPORT
2326|BRANCHVILLE
2327|BRAND
2328|BRANDENBERG
2329|BRANDENBURG
2330|BRANDERMILL
2331|BRANDON
2332|BRANDONVILLE
2333|BRANDRETH
2334|BRANDSVILLE
2335|BRANDT
2336|BRANDYWINE
2337|BRANDYWINE MANOR
2338|BRANFORD
2339|BRANSFORD
2340|BRANSON
2341|BRANSON WEST
2342|BRANT LAKE
2343|BRANT ROCK
2344|BRANTFORD
2345|BRANTLEY
2346|BRANTLEYVILLE
2347|BRANTON
2348|BRANTWOOD
2349|BRASELTON
2350|BRASFIELD
2351|BRASHEAR
2352|BRASHER FALLS
2353|BRASS CASTLE
2354|BRASSTOWN
2355|BRASWELL
2356|BRATENAHL
2357|BRATT
2358|BRATTLEBORO
2359|BRAVE
2360|BRAWLEY
2361|BRAXTON
2362|BRAY
2363|BRAYMER
2364|BRAYTON
2365|BRAZIL
2366|BRAZILTON
2367|BRAZORIA
2368|BRAZOS
2369|BRAZOS BEND
2370|BRAZOS COUNTRY
2371|BREA
2372|BREATHEDSVILLE
2373|BREAUX BRIDGE
2374|BRECKENRIDGE
2375|BRECKENRIDGE HILLS
2376|BRECKINRIDGE
2377|BRECKINRIDGE CENTER
2378|BRECKSVILLE
2379|BRECON
2380|BREDA
2381|BREEDSVILLE
2382|BREESE
2383|BREESPORT
2384|BREEZY POINT
2385|BREIDABLICK
2386|BREIEN
2387|BREINIGSVILLE
2388|BREMEN
2389|BREMER
2390|BREMERTON
2391|BREMOND
2392|BRENAS
2393|BRENDA
2394|BRENHAM
2395|BRENT
2396|BRENTFORD
2397|BRENTON
2398|BRENTSVILLE
2399|BRENTWOOD
2400|BRENTWOOD LAKE
2401|BRESLAU
2402|BRESSLER
2403|BRETHREN
2404|BREVARD
2405|BREVIG MISSION
2406|BREVORT
2407|BREWER
2408|BREWERTON
2409|BREWSTER
2410|BREWSTER HILL
2411|BREWTON
2412|BREÑAS COMUNIDAD
2413|BRIAN HEAD
2414|BRIAR
2415|BRIAR CREEK
2416|BRIARCLIFF
2417|BRIARCLIFF MANOR
2418|BRIARCLIFFE ACRES
2419|BRIAROAKS
2420|BRIARTOWN
2421|BRIARWOOD
2422|BRICE
2423|BRICE PRAIRIE
2424|BRICELYN
2425|BRICES CREEK
2426|BRICEVILLE
2427|BRICK
2428|BRICKERVILLE
2429|BRICKEYS
2430|BRIDGE
2431|BRIDGE CITY
2432|BRIDGE CREEK
2433|BRIDGEBORO
2434|BRIDGEHAMPTON
2435|BRIDGELAND
2436|BRIDGEPORT
2437|BRIDGER
2438|BRIDGETON
2439|BRIDGETOWN
2440|BRIDGEVIEW
2441|BRIDGEVILLE
2442|BRIDGEWATER
2443|BRIDGMAN
2444|BRIDGTON
2445|BRIELLE
2446|BRIENSBURG
2447|BRIER
2448|BRIER HILL
2449|BRIGANTINE
2450|BRIGGS
2451|BRIGGSDALE
2452|BRIGGSVILLE
2453|BRIGHAM CITY
2454|BRIGHTON
2455|BRIGHTWATERS
2456|BRIGHTWOOD
2457|BRILL
2458|BRILLIANT
2459|BRILLION
2460|BRIMFIELD
2461|BRIMHALL NIZHONI
2462|BRIMLEY
2463|BRIMSON
2464|BRINCKERHOFF
2465|BRINKHAVEN
2466|BRINKLEY
2467|BRINKLOW
2468|BRINKMAN
2469|BRINNON
2470|BRINSMADE
2471|BRINSON
2472|BRINY BREEZES
2473|BRISBANE
2474|BRISBIN
2475|BRISCOE
2476|BRISTOL
2477|BRISTOW
2478|BRITT
2479|BRITTON
2480|BROAD BROOK
2481|BROAD CREEK
2482|BROAD TOP CITY
2483|BROADALBIN
2484|BROADBENT
2485|BROADDUS
2486|BROADFORD
2487|BROADHURST
2488|BROADLAND
2489|BROADLANDS
2490|BROADMOOR
2491|BROADUS
2492|BROADVIEW
2493|BROADVIEW HEIGHTS
2494|BROADVIEW PARK
2495|BROADWATER
2496|BROADWAY
2497|BROADWELL
2498|BROCK
2499|BROCK HALL
2500|BROCKET
2501|BROCKPORT
2502|BROCKTON
2503|BROCKWAY
2504|BROCTON
2505|BRODHEAD
2506|BRODHEADSVILLE
2507|BRODNAX
2508|BROECK POINTE
2509|BROGAN
2510|BROGDEN
2511|BROHARD
2512|BROKAW
2513|BROKEN ARROW
2514|BROKEN BOW
2515|BROKENBURG
2516|BROMIDE
2517|BROMLEY
2518|BRONAUGH
2519|BRONCHO
2520|BRONSON
2521|BRONTE
2522|BRONWOOD
2523|BRONX
2524|BRONXVILLE
2525|BROOK
2526|BROOK HIGHLAND
2527|BROOK PARK
2528|BROOKDALE
2529|BROOKE
2530|BROOKELAND
2531|BROOKER
2532|BROOKESMITH
2533|BROOKEVILLE
2534|BROOKFIELD
2535|BROOKFIELD CENTER
2536|BROOKFORD
2537|BROOKHAVEN
2538|BROOKHURST
2539|BROOKINGS
2540|BROOKLAND
2541|BROOKLAWN
2542|BROOKLET
2543|BROOKLINE
2544|BROOKLYN
2545|BROOKLYN CENTER
2546|BROOKLYN HEIGHTS
2547|BROOKLYN PARK
2548|BROOKMONT
2549|BROOKNEAL
2550|BROOKPORT
2551|BROOKRIDGE
2552|BROOKS
2553|BROOKSBURG
2554|BROOKSHIRE
2555|BROOKSIDE
2556|BROOKSIDE VILLAGE
2557|BROOKSTON
2558|BROOKSVILLE
2559|BROOKTON
2560|BROOKTRAILS
2561|BROOKTREE PARK
2562|BROOKVALE
2563|BROOKVIEW
2564|BROOKVILLE
2565|BROOKWOOD
2566|BROOMALL
2567|BROOMES ISLAND
2568|BROOMFIELD
2569|BROOMTOWN
2570|BROOTEN
2571|BROSELEY
2572|BROSVILLE
2573|BROUGHTON
2574|BROUSSARD
2575|BROWARDALE
2576|BROWERVILLE
2577|BROWN CITY
2578|BROWN DEER
2579|BROWNBRANCH
2580|BROWNDELL
2581|BROWNELL
2582|BROWNFIELD
2583|BROWNING
2584|BROWNINGTON
2585|BROWNLEE
2586|BROWNLEE PARK
2587|BROWNS
2588|BROWNS LAKE
2589|BROWNS MILLS
2590|BROWNS POINT
2591|BROWNS VALLEY
2592|BROWNSBORO
2593|BROWNSBORO FARM
2594|BROWNSBORO VILLAGE
2595|BROWNSBURG
2596|BROWNSDALE
2597|BROWNSFIELD
2598|BROWNSON
2599|BROWNSTOWN
2600|BROWNSVILLE
2601|BROWNTON
2602|BROWNTOWN
2603|BROWNVILLE
2604|BROWNVILLE JUNCTION
2605|BROWNWOOD
2606|BROXTON
2607|BRUCE
2608|BRUCE CROSSING
2609|BRUCETON
2610|BRUCETON MILLS
2611|BRUCETOWN
2612|BRUCEVILLE
2613|BRUCEVILLE-EDDY
2614|BRUIN
2615|BRULE
2616|BRUMLEY
2617|BRUMLEY GAP
2618|BRUNDAGE
2619|BRUNDIDGE
2620|BRUNEAU
2621|BRUNERSBURG
2622|BRUNI
2623|BRUNING
2624|BRUNO
2625|BRUNSON
2626|BRUNSVILLE
2627|BRUNSWICK
2628|BRUNSWICK GARDENS
2629|BRUSETT
2630|BRUSH
2631|BRUSH CREEK
2632|BRUSH FORK
2633|BRUSH PRAIRIE
2634|BRUSHTON
2635|BRUSHVALE
2636|BRUSHY
2637|BRUSHY CREEK
2638|BRUSLY
2639|BRUSLY LANDING
2640|BRUSSELS
2641|BRUTUS
2642|BRYANS ROAD
2643|BRYANT
2644|BRYANT POND
2645|BRYANTOWN
2646|BRYCE
2647|BRYCE CANYON
2648|BRYCE CANYON CITY
2649|BRYCELAND
2650|BRYCEVILLE
2651|BRYDEN
2652|BRYN ATHYN
2653|BRYN MAWR
2654|BRYSON
2655|BRYSON CITY
2656|BUCHANAN
2657|BUCHANAN DAM
2658|BUCHANAN LAKE VILLAGE
2659|BUCHTEL
2660|BUCK CREEK
2661|BUCK GROVE
2662|BUCK MEADOWS
2663|BUCK RUN
2664|BUCKATUNNA
2665|BUCKEYE
2666|BUCKEYE LAKE
2667|BUCKEYSTOWN
2668|BUCKHALL
2669|BUCKHANNON
2670|BUCKHEAD
2671|BUCKHEAD RIDGE
2672|BUCKHOLTS
2673|BUCKHORN
2674|BUCKINGHAM
2675|BUCKLAND
2676|BUCKLEY
2677|BUCKLIN
2678|BUCKMAN
2679|BUCKNER
2680|BUCKS
2681|BUCKS LAKE
2682|BUCKSPORT
2683|BUCKTAIL
2684|BUCKTOWN
2685|BUCODA
2686|BUCYRUS
2687|BUD
2688|BUDA
2689|BUDD LAKE
2690|BUDDTOWN
2691|BUDE
2692|BUELL
2693|BUELLTON
2694|BUENA
2695|BUENA PARK
2696|BUENA VISTA
2697|BUENA VISTA COLONIA
2698|BUENA VISTA COMUNIDAD
2699|BUENAVENTURA LAKES
2700|BUENOS
2701|BUEYEROS
2702|BUFALO
2703|BUFFALO
2704|BUFFALO CENTER
2705|BUFFALO CHIP
2706|BUFFALO CITY
2707|BUFFALO CREEK
2708|BUFFALO GAP
2709|BUFFALO GROVE
2710|BUFFALO LAKE
2711|BUFFALO PRAIRIE
2712|BUFFALO SPRINGS
2713|BUFFALO VALLEY
2714|BUFFINGTON
2715|BUFORD
2716|BUHL
2717|BUHLER
2718|BUIE
2719|BUIES CREEK
2720|BUIST
2721|BULADEAN
2722|BULGER
2723|BULL CREEK
2724|BULL HOLLOW
2725|BULL RUN
2726|BULL RUN MOUNTAIN ESTATES
2727|BULL SHOALS
2728|BULL VALLEY
2729|BULLARD
2730|BULLHEAD
2731|BULLHEAD CITY
2732|BULLITTSVILLE
2733|BULLS GAP
2734|BULPITT
2735|BULVERDE
2736|BUMBLE BEE
2737|BUMPUS MILLS
2738|BUNA
2739|BUNAVISTA
2740|BUNCETON
2741|BUNCOMBE
2742|BUNKER
2743|BUNKER HILL
2744|BUNKER HILL VILLAGE
2745|BUNKERVILLE
2746|BUNKIE
2747|BUNN
2748|BUNNELL
2749|BUNNLEVEL
2750|BURAS
2751|BURBANK
2752|BURCHARD
2753|BURCHINAL
2754|BURDEN
2755|BURDETT
2756|BURDETTE
2757|BURDICK
2758|BURDOCK
2759|BUREAU
2760|BURGAW
2761|BURGDORF
2762|BURGESS
2763|BURGESS JUNCTION
2764|BURGETTSTOWN
2765|BURGIN
2766|BURGOON
2767|BURIEN
2768|BURKBURNETT
2769|BURKE
2770|BURKES GARDEN
2771|BURKESVILLE
2772|BURKET
2773|BURKETT
2774|BURKETTSVILLE
2775|BURKEVILLE
2776|BURKITTSVILLE
2777|BURLEIGH
2778|BURLESON
2779|BURLEY
2780|BURLINGAME
2781|BURLINGTON
2782|BURLINGTON JUNCTION
2783|BURLISON
2784|BURMAH
2785|BURMESTER
2786|BURNA
2787|BURNET
2788|BURNETT
2789|BURNETTOWN
2790|BURNETTSVILLE
2791|BURNEY
2792|BURNEYVILLE
2793|BURNHAM
2794|BURNING SPRINGS
2795|BURNS
2796|BURNS CITY
2797|BURNS FLAT
2798|BURNS HARBOR
2799|BURNSIDE
2800|BURNSTAD
2801|BURNSVILLE
2802|BURNT CORN
2803|BURNT PRAIRIE
2804|BURNT RANCH
2805|BURNT STORE MARINA
2806|BURNTFORK
2807|BURR
2808|BURR FERRY
2809|BURR OAK
2810|BURR RIDGE
2811|BURREL
2812|BURRIS
2813|BURROUGHS
2814|BURROWS
2815|BURRTON
2816|BURRVILLE
2817|BURT
2818|BURTON
2819|BURTONS BRIDGE
2820|BURTONSVILLE
2821|BURTRUM
2822|BURWELL
2823|BUSBY
2824|BUSCH
2825|BUSH
2826|BUSH CITY
2827|BUSHKILL
2828|BUSHLAND
2829|BUSHNELL
2830|BUSHONG
2831|BUSHTON
2832|BUSHYHEAD
2833|BUSSEY
2834|BUSTAMANTE
2835|BUSTI
2836|BUTLER
2837|BUTLER BEACH
2838|BUTLER JUNCTION
2839|BUTLERTOWN
2840|BUTLERVILLE
2841|BUTNER
2842|BUTTE
2843|BUTTE CITY
2844|BUTTE DES MORTS
2845|BUTTE FALLS
2846|BUTTE LA ROSE
2847|BUTTE MEADOWS
2848|BUTTERFIELD
2849|BUTTERNUT
2850|BUTTERS
2851|BUTTEVILLE
2852|BUTTONWILLOW
2853|BUTTZVILLE
2854|BUXTON
2855|BUYCK
2856|BUZZARDS BAY
2857|BYARS
2858|BYER
2859|BYERS
2860|BYERSVILLE
2861|BYESVILLE
2862|BYHALIA
2863|BYLAS
2864|BYNG
2865|BYNUM
2866|BYRAM
2867|BYRDSTOWN
2868|BYRNE
2869|BYRNEDALE
2870|BYRNES MILL
2871|BYROMVILLE
2872|BYRON
2873|BYRON CENTER
2874|BYSTROM
2875|BÚFALO COMUNIDAD
2876|CABALLO
2877|CABAN
2878|CABAZON
2879|CABERY
2880|CABIN JOHN
2881|CABLE
2882|CABO ROJO
2883|CABO ROJO ZONA URBANA
2884|CABOOL
2885|CABORN
2886|CABOT
2887|CABÁN COMUNIDAD
2888|CACAO
2889|CACAO COMUNIDAD
2890|CACHE
2891|CACTUS
2892|CACTUS FLAT
2893|CACTUS FOREST
2894|CADDO
2895|CADDO GAP
2896|CADDO MILLS
2897|CADDO VALLEY
2898|CADDOA
2899|CADE
2900|CADES
2901|CADILLAC
2902|CADIZ
2903|CADLEY
2904|CADOGAN
2905|CADOTT
2906|CADWELL
2907|CADY
2908|CAERNARVON
2909|CAFFEE JUNCTION
2910|CAGUAS
2911|CAGUAS ZONA URBANA
2912|CAHOKIA
2913|CAHONE
2914|CAINEVILLE
2915|CAINSVILLE
2916|CAIRNBROOK
2917|CAIRO
2918|CAJAHS MOUNTAIN
2919|CAJON JUNCTION
2920|CAL-NEV-ARI
2921|CALABASAS
2922|CALABASH
2923|CALAIS
2924|CALAMINE
2925|CALAMUS
2926|CALAVO GARDENS
2927|CALCASIEU
2928|CALCUTTA
2929|CALDWELL
2930|CALE
2931|CALEDONIA
2932|CALERA
2933|CALEXICO
2934|CALHAN
2935|CALHOUN
2936|CALHOUN CITY
2937|CALHOUN FALLS
2938|CALICO ROCK
2939|CALIENTE
2940|CALIFON
2941|CALIFORNIA
2942|CALIFORNIA CITY
2943|CALIFORNIA HOT SPRINGS
2944|CALIFORNIA JUNCTION
2945|CALIFORNIA PINES
2946|CALIMESA
2947|CALIO
2948|CALION
2949|CALIPATRIA
2950|CALISTA
2951|CALISTOGA
2952|CALLAGHAN
2953|CALLAHAN
2954|CALLANDS
2955|CALLAO
2956|CALLAWAY
2957|CALLENDER
2958|CALLENSBURG
2959|CALLERY
2960|CALLICOON
2961|CALLIHAM
2962|CALLIMONT
2963|CALLISBURG
2964|CALMAR
2965|CALN
2966|CALPELLA
2967|CALPINE
2968|CALUMET
2969|CALUMET CITY
2970|CALUMET PARK
2971|CALVA
2972|CALVARY
2973|CALVERT
2974|CALVERT BEACH
2975|CALVERT CITY
2976|CALVERTON
2977|CALVERTON PARK
2978|CALVIN
2979|CALWA
2980|CALYPSO
2981|CALZADA
2982|CALZADA COMUNIDAD
2983|CAMAK
2984|CAMANCHE
2985|CAMANCHE VILLAGE
2986|CAMANO
2987|CAMARGO
2988|CAMARILLO
2989|CAMAS
2990|CAMAS VALLEY
2991|CAMBRIA
2992|CAMBRIA CENTER
2993|CAMBRIAN PARK
2994|CAMBRIDGE
2995|CAMBRIDGE CITY
2996|CAMBRIDGE SPRINGS
2997|CAMDEN
2998|CAMDEN ON GAULEY
2999|CAMDEN POINT
3000|CAMDENTON
3001|CAMEO
3002|CAMERON
3003|CAMERON PARK
3004|CAMERON PARK COLONIA
3005|CAMILLA
3006|CAMILLUS
3007|CAMINO
3008|CAMINO TASSAJARA
3009|CAMMACK VILLAGE
3010|CAMMAL
3011|CAMP
3012|CAMP BIRD
3013|CAMP CREEK
3014|CAMP CROOK
3015|CAMP DENNISON
3016|CAMP DOUGLAS
3017|CAMP HILL
3018|CAMP JO-ANN
3019|CAMP LAKE
3020|CAMP NELSON
3021|CAMP POINT
3022|CAMP SAN SABA
3023|CAMP SHERMAN
3024|CAMP SPRINGS
3025|CAMP SWIFT
3026|CAMP THREE
3027|CAMP VERDE
3028|CAMP WOOD
3029|CAMPAIGN
3030|CAMPANILLA
3031|CAMPANILLA COMUNIDAD
3032|CAMPBELL
3033|CAMPBELL HILL
3034|CAMPBELL STATION
3035|CAMPBELLSBURG
3036|CAMPBELLSPORT
3037|CAMPBELLSTOWN
3038|CAMPBELLSVILLE
3039|CAMPBELLTON
3040|CAMPBELLTOWN
3041|CAMPIA
3042|CAMPO
3043|CAMPO BONITO
3044|CAMPO RICO
3045|CAMPO RICO COMUNIDAD
3046|CAMPOBELLO
3047|CAMPTI
3048|CAMPTON
3049|CAMPTON HILLS
3050|CAMPTONVILLE
3051|CAMPTOWN
3052|CAMPUS
3053|CAMPVILLE
3054|CAMUY
3055|CAMUY ZONA URBANA
3056|CANA
3057|CANAAN
3058|CANADA CREEK RANCH
3059|CANADENSIS
3060|CANADIAN
3061|CANADIAN LAKES
3062|CANADOHTA LAKE
3063|CANADYS
3064|CANAJOHARIE
3065|CANAL FULTON
3066|CANAL LEWISVILLE
3067|CANAL POINT
3068|CANAL WINCHESTER
3069|CANALOU
3070|CANANDAIGUA
3071|CANASERAGA
3072|CANASTOTA
3073|CANBY
3074|CANDELARIA
3075|CANDELARIA ARENAS
3076|CANDELARIA ARENAS COMUNIDAD
3077|CANDELARIA COMUNIDAD
3078|CANDELERO ABAJO COMUNIDAD
3079|CANDELERO ARRIBA
3080|CANDELERO ARRIBA COMUNIDAD
3081|CANDLE
3082|CANDLER
3083|CANDO
3084|CANDOR
3085|CANE BEDS
3086|CANE SAVANNAH
3087|CANE VALLEY
3088|CANEY
3089|CANEY CITY
3090|CANEYVILLE
3091|CANFIELD
3092|CANISTEO
3093|CANISTOTA
3094|CANJILON
3095|CANKTON
3096|CANMER
3097|CANNEL CITY
3098|CANNELBURG
3099|CANNELTON
3100|CANNING
3101|CANNON BALL
3102|CANNON BEACH
3103|CANNON FALLS
3104|CANNON TOWN
3105|CANNONDALE
3106|CANNONSBURG
3107|CANNONVILLE
3108|CANON
3109|CANONSBURG
3110|CANOOCHEE
3111|CANOVA
3112|CANOVANAS
3113|CANTERWOOD
3114|CANTIL
3115|CANTON
3116|CANTON VALLEY
3117|CANTONMENT
3118|CANTRALL
3119|CANTRIL
3120|CANTU ADDITION
3121|CANTUA CREEK
3122|CANTWELL
3123|CANUTE
3124|CANUTILLO
3125|CANYON
3126|CANYON CITY
3127|CANYON COUNTRY
3128|CANYON CREEK
3129|CANYON DAY
3130|CANYON DIABLO
3131|CANYON LAKE
3132|CANYON PARK
3133|CANYON VALLEY
3134|CANYONDAM
3135|CANYONVILLE
3136|CANÓVANAS ZONA URBANA
3137|CAP ROCK
3138|CAPA
3139|CAPAC
3140|CAPE CANAVERAL
3141|CAPE CARTERET
3142|CAPE CHARLES
3143|CAPE CORAL
3144|CAPE FAIR
3145|CAPE GIRARDEAU
3146|CAPE MAY
3147|CAPE MAY COURT HOUSE
3148|CAPE MAY POINT
3149|CAPE MEARES
3150|CAPE NEDDICK
3151|CAPE POLE
3152|CAPE SAINT CLAIRE
3153|CAPE VINCENT
3154|CAPE YAKATAGA
3155|CAPISTRANO BEACH
3156|CAPITAN
3157|CAPITANEJO
3158|CAPITANEJO COMUNIDAD
3159|CAPITOL
3160|CAPITOL HEIGHTS
3161|CAPITOLA
3162|CAPLEVILLE
3163|CAPLINGER MILLS
3164|CAPLIS
3165|CAPON BRIDGE
3166|CAPPS
3167|CAPPS SWITCH
3168|CAPROCK
3169|CAPRON
3170|CAPS
3171|CAPTAIN COOK
3172|CAPTAINS COVE
3173|CAPTINA
3174|CAPTIVA
3175|CAPULIN
3176|CAPUTA
3177|CARAWAY
3178|CARBON
3179|CARBON CLIFF
3180|CARBON HILL
3181|CARBONADO
3182|CARBONDALE
3183|CARBONVILLE
3184|CARBURY
3185|CARDIFF
3186|CARDIFF-BY-THE-SEA
3187|CARDINGTON
3188|CARDWELL
3189|CAREFREE
3190|CARENCRO
3191|CAREY
3192|CAREYWOOD
3193|CARGRAY
3194|CARIBOU
3195|CARL
3196|CARL JUNCTION
3197|CARLE PLACE
3198|CARLETON
3199|CARLILE
3200|CARLIN
3201|CARLINVILLE
3202|CARLISLE
3203|CARLISLE GARDENS
3204|CARLOCK
3205|CARLOS
3206|CARLS CORNER
3207|CARLSBAD
3208|CARLSBORG
3209|CARLSON
3210|CARLSTADT
3211|CARLSVILLE
3212|CARLTON
3213|CARLTON LANDING
3214|CARLYLE
3215|CARLYSS
3216|CARMEL
3217|CARMEL VALLEY
3218|CARMEL VALLEY VILLAGE
3219|CARMEL-BY-THE-SEA
3220|CARMEN
3221|CARMET
3222|CARMI
3223|CARMICHAEL
3224|CARMICHAELS
3225|CARMINE
3226|CARNATION
3227|CARNE
3228|CARNEGIE
3229|CARNEIRO
3230|CARNELIAN BAY
3231|CARNERO
3232|CARNESVILLE
3233|CARNEY
3234|CARNEYS POINT
3235|CARNOT
3236|CARNTOWN
3237|CARNUEL
3238|CARO
3239|CAROGA LAKE
3240|CAROL STREAM
3241|CAROLEEN
3242|CAROLINA
3243|CAROLINA BEACH
3244|CAROLINA SHORES
3245|CAROLINA ZONA URBANA
3246|CAROLINE
3247|CARP
3248|CARP LAKE
3249|CARPENDALE
3250|CARPENTER
3251|CARPENTERSVILLE
3252|CARPENTERVILLE
3253|CARPINTERIA
3254|CARPIO
3255|CARR
3256|CARRABASSETT
3257|CARRABELLE
3258|CARRBORO
3259|CARRICK
3260|CARRIER
3261|CARRIER MILLS
3262|CARRIERE
3263|CARRINGTON
3264|CARRIZALES
3265|CARRIZALES COMUNIDAD
3266|CARRIZO
3267|CARRIZO HILL
3268|CARRIZO SPRINGS
3269|CARRIZOZO
3270|CARROLL
3271|CARROLL VALLEY
3272|CARROLLS
3273|CARROLLTON
3274|CARROLLTON MANOR
3275|CARROLLTOWN
3276|CARROLLWOOD
3277|CARROTHERS
3278|CARRSVILLE
3279|CARSINS
3280|CARSON
3281|CARSON CITY
3282|CARSONVILLE
3283|CARTA VALLEY
3284|CARTAGO
3285|CARTER
3286|CARTER LAKE
3287|CARTERET
3288|CARTERSVILLE
3289|CARTERVILLE
3290|CARTHAGE
3291|CARTWRIGHT
3292|CARUTHERS
3293|CARUTHERSVILLE
3294|CARVER
3295|CARVILLE
3296|CARY
3297|CARYTOWN
3298|CARYVILLE
3299|CASA
3300|CASA BLANCA
3301|CASA COLORADA
3302|CASA CONEJO
3303|CASA DE ORO
3304|CASA GRANDE
3305|CASA PIEDRA
3306|CASAR
3307|CASAS ADOBES
3308|CASCADE
3309|CASCADE LOCKS
3310|CASCADE VALLEY
3311|CASCADIA
3312|CASCO
3313|CASELTON
3314|CASEVILLE
3315|CASEY
3316|CASEYVILLE
3317|CASH
3318|CASHEL
3319|CASHIERS
3320|CASHION
3321|CASHION COMMUNITY
3322|CASHMERE
3323|CASHTON
3324|CASHTOWN
3325|CASITAS SPRINGS
3326|CASKY
3327|CASMALIA
3328|CASNOVIA
3329|CASON
3330|CASPAR
3331|CASPER
3332|CASPER MOUNTAIN
3333|CASPIAN
3334|CASPIANA
3335|CASS
3336|CASS CITY
3337|CASS LAKE
3338|CASSA
3339|CASSADAGA
3340|CASSANDRA
3341|CASSATT
3342|CASSCOE
3343|CASSEL
3344|CASSELBERRY
3345|CASSELMAN
3346|CASSELTON
3347|CASSODAY
3348|CASSOPOLIS
3349|CASSTOWN
3350|CASSVILLE
3351|CASTAIC
3352|CASTALIA
3353|CASTALIAN SPRINGS
3354|CASTANA
3355|CASTANEA
3356|CASTANEDA
3357|CASTELLA
3358|CASTILE
3359|CASTINE
3360|CASTLE
3361|CASTLE DALE
3362|CASTLE DANGER
3363|CASTLE HAYNE
3364|CASTLE HILLS
3365|CASTLE PARK
3366|CASTLE PINES
3367|CASTLE PINES NORTH
3368|CASTLE PINES VILLAGE
3369|CASTLE POINT
3370|CASTLE ROCK
3371|CASTLE SHANNON
3372|CASTLE VALLEY
3373|CASTLEBERRY
3374|CASTLEFORD
3375|CASTLETON
3376|CASTLETON-ON-HUDSON
3377|CASTLEWOOD
3378|CASTOLON
3379|CASTOR
3380|CASTORLAND
3381|CASTRO VALLEY
3382|CASTROVILLE
3383|CASWELL BEACH
3384|CAT CREEK
3385|CAT SPRING
3386|CATAHOULA
3387|CATALINA
3388|CATALINA FOOTHILLS
3389|CATARACT
3390|CATARINA
3391|CATASAUQUA
3392|CATAULA
3393|CATAWBA
3394|CATAWBA ISLAND
3395|CATAWISSA
3396|CATAÑO
3397|CATAÑO ZONA URBANA
3398|CATESBY
3399|CATHARINE
3400|CATHAY
3401|CATHCART
3402|CATHEDRAL
3403|CATHEDRAL CITY
3404|CATHERINE
3405|CATHEYS VALLEY
3406|CATHLAMET
3407|CATLETT
3408|CATLETTSBURG
3409|CATLIN
3410|CATO
3411|CATONSVILLE
3412|CATOOSA
3413|CATRON
3414|CATS BRIDGE
3415|CATSKILL
3416|CATTARAUGUS
3417|CATTLE CREEK
3418|CAULFIELD
3419|CAULKSVILLE
3420|CAUSEY
3421|CAUTHRON
3422|CAVALERO CORNER
3423|CAVALIER
3424|CAVE
3425|CAVE CITY
3426|CAVE CREEK
3427|CAVE JUNCTION
3428|CAVE SPRING
3429|CAVE SPRINGS
3430|CAVE-IN-ROCK
3431|CAVENDISH
3432|CAVETOWN
3433|CAVOUR
3434|CAWKER CITY
3435|CAWOOD
3436|CAYCE
3437|CAYEY
3438|CAYEY ZONA URBANA
3439|CAYLOR
3440|CAYUCO
3441|CAYUCO COMUNIDAD
3442|CAYUCOS
3443|CAYUGA
3444|CAYUGA HEIGHTS
3445|CAYUSE
3446|CAZADERO
3447|CAZENOVIA
3448|CAÑADA DE LOS ALAMOS
3449|CAÑON
3450|CAÑON CITY
3451|CAÑONES
3452|CEARFOSS
3453|CEBOLLA
3454|CECIL
3455|CECILIA
3456|CECILTON
3457|CECILVILLE
3458|CEDAR
3459|CEDAR BLUFF
3460|CEDAR BLUFFS
3461|CEDAR BROOK
3462|CEDAR BUTTE
3463|CEDAR CITY
3464|CEDAR CREEK
3465|CEDAR CREST
3466|CEDAR FALLS
3467|CEDAR FORT
3468|CEDAR GLEN
3469|CEDAR GLEN LAKES
3470|CEDAR GLEN WEST
3471|CEDAR GROVE
3472|CEDAR HIGHLANDS
3473|CEDAR HILL
3474|CEDAR HILL LAKES
3475|CEDAR HILLS
3476|CEDAR KEY
3477|CEDAR KNOLLS
3478|CEDAR LAKE
3479|CEDAR MILL
3480|CEDAR MILLS
3481|CEDAR MOUNTAIN
3482|CEDAR PARK
3483|CEDAR POINT
3484|CEDAR RAPIDS
3485|CEDAR RIDGE
3486|CEDAR RIVER
3487|CEDAR ROCK
3488|CEDAR SLOPE
3489|CEDAR SPRINGS
3490|CEDAR VALE
3491|CEDAR VALLEY
3492|CEDARBURG
3493|CEDAREDGE
3494|CEDARHURST
3495|CEDARPINES PARK
3496|CEDARTOWN
3497|CEDARVILLE
3498|CEDARWOOD
3499|CEDONIA
3500|CEDRO
3501|CEE VEE
3502|CEGO
3503|CEIBA
3504|CEIBA COMUNIDAD
3505|CEIBA ZONA URBANA
3506|CELADA
3507|CELADA COMUNIDAD
3508|CELEBRATION
3509|CELERYVILLE
3510|CELESTE
3511|CELESTINE
3512|CELINA
3513|CELO
3514|CELORON
3515|CEMENT CITY
3516|CEMENTON
3517|CENTENARY
3518|CENTENNIAL
3519|CENTER CITY
3520|CENTER CROSS
3521|CENTER HILL
3522|CENTER JUNCTION
3523|CENTER LINE
3524|CENTER MORICHES
3525|CENTER OSSIPEE
3526|CENTER POINT
3527|CENTER POST
3528|CENTER RIDGE
3529|CENTER SANDWICH
3530|CENTER SQUARE
3531|CENTERBURG
3532|CENTERDALE
3533|CENTEREACH
3534|CENTERFIELD
3535|CENTERPORT
3536|CENTERTON
3537|CENTERTOWN
3538|CENTERVIEW
3539|CENTERVILLE
3540|CENTRAHOMA
3541|CENTRAL AGUIRRE
3542|CENTRAL AGUIRRE COMUNIDAD
3543|CENTRAL BRIDGE
3544|CENTRAL CITY
3545|CENTRAL FALLS
3546|CENTRAL GARAGE
3547|CENTRAL GARDENS
3548|CENTRAL HEIGHTS
3549|CENTRAL HIGH
3550|CENTRAL ISLIP
3551|CENTRAL LAKE
3552|CENTRAL PACOLET
3553|CENTRAL PARK
3554|CENTRAL POINT
3555|CENTRAL SQUARE
3556|CENTRAL VALLEY
3557|CENTRALHATCHEE
3558|CENTRALIA
3559|CENTRE
3560|CENTRE HALL
3561|CENTRE ISLAND
3562|CENTREVILLE
3563|CENTROPOLIS
3564|CENTURIA
3565|CENTURY
3566|CEREDO
3567|CERES
3568|CERESCO
3569|CERRILLOS
3570|CERRILLOS HOYOS COMUNIDAD
3571|CERRITOS
3572|CERRO GORDO
3573|CERULEAN
3574|CESTOS
3575|CETRONIA
3576|CEYLON
3577|CHACKBAY
3578|CHACRA
3579|CHADBOURN
3580|CHADDS FORD
3581|CHADRON
3582|CHADWICK
3583|CHADWICKS
3584|CHAFFEE
3585|CHAGRIN FALLS
3586|CHAIN O' LAKES
3587|CHAIN OF ROCKS
3588|CHAIN-O-LAKES
3589|CHAIRES
3590|CHALCO
3591|CHALFANT
3592|CHALFONT
3593|CHALK MOUNTAIN
3594|CHALKHILL
3595|CHALKYITSIK
3596|CHALLIS
3597|CHALMERS
3598|CHALMETTE
3599|CHALYBEATE SPRINGS
3600|CHAMA
3601|CHAMBERINO
3602|CHAMBERLAIN
3603|CHAMBERLAYNE
3604|CHAMBERLAYNE HEIGHTS
3605|CHAMBERLIN
3606|CHAMBERS
3607|CHAMBERSBURG
3608|CHAMBLEE
3609|CHAMISAL
3610|CHAMITA
3611|CHAMIZAL
3612|CHAMOIS
3613|CHAMP
3614|CHAMPAIGN
3615|CHAMPION
3616|CHAMPLAIN
3617|CHAMPLIN
3618|CHANA
3619|CHANCE
3620|CHANCELLOR
3621|CHANDALAR
3622|CHANDLER
3623|CHANDLER HEIGHTS
3624|CHANDLER SPRINGS
3625|CHANDLERVILLE
3626|CHANEYVILLE
3627|CHANHASSEN
3628|CHANILIUT
3629|CHANNAHON
3630|CHANNEL ISLANDS BEACH
3631|CHANNEL LAKE
3632|CHANNELVIEW
3633|CHANNING
3634|CHANTILLY
3635|CHANUTE
3636|CHAPARRAL
3637|CHAPEL HILL
3638|CHAPIN
3639|CHAPLIN
3640|CHAPMAN
3641|CHAPMAN RANCH
3642|CHAPMANVILLE
3643|CHAPPAQUA
3644|CHAPPELL
3645|CHAPPELL HILL
3646|CHAPPELLS
3647|CHAPTICO
3648|CHARCO
3649|CHARDON
3650|CHARENTON
3651|CHARING
3652|CHARITON
3653|CHARITY
3654|CHARLACK
3655|CHARLEROI
3656|CHARLES
3657|CHARLES CITY
3658|CHARLES TOWN
3659|CHARLESTON
3660|CHARLESTON PARK
3661|CHARLESTOWN
3662|CHARLEVOIX
3663|CHARLO
3664|CHARLOS HEIGHTS
3665|CHARLOTTE
3666|CHARLOTTE AMALIE
3667|CHARLOTTE COURT HOUSE
3668|CHARLOTTE HALL
3669|CHARLOTTE HARBOR
3670|CHARLOTTE PARK
3671|CHARLOTTESVILLE
3672|CHARLTON
3673|CHARLTON HEIGHTS
3674|CHARM
3675|CHARMWOOD
3676|CHARTER OAK
3677|CHARTERS
3678|CHASE
3679|CHASE CITY
3680|CHASE CROSSING
3681|CHASEBURG
3682|CHASELEY
3683|CHASKA
3684|CHASSAHOWITZKA
3685|CHASTANG
3686|CHATAIGNIER
3687|CHATANIKA
3688|CHATAWA
3689|CHATCOLET
3690|CHATEAU WOODS
3691|CHATEAUGAY
3692|CHATFIELD
3693|CHATHAM
3694|CHATMOSS
3695|CHATOM
3696|CHATSWORTH
3697|CHATTAHOOCHEE
3698|CHATTAHOOCHEE HILLS
3699|CHATTANOOGA
3700|CHATTANOOGA VALLEY
3701|CHATTAROY
3702|CHATWOOD
3703|CHAUMONT
3704|CHAUNCEY
3705|CHAUTAUQUA
3706|CHAUVIN
3707|CHAVIES
3708|CHAZY
3709|CHEAT LAKE
3710|CHEBANSE
3711|CHEBOYGAN
3712|CHECOTAH
3713|CHEEKTOWAGA
3714|CHEFORNAK
3715|CHEHALIS
3716|CHELAN
3717|CHELAN FALLS
3718|CHELATCHIE
3719|CHELATNA LODGE
3720|CHELMSFORD
3721|CHELSEA
3722|CHELTENHAM
3723|CHELYAN
3724|CHEMULT
3725|CHEMUNG
3726|CHENA HOT SPRINGS
3727|CHENANGO BRIDGE
3728|CHENEQUA
3729|CHENEY
3730|CHENEYVILLE
3731|CHENOA
3732|CHENOWETH
3733|CHEPACHET
3734|CHERAW
3735|CHERITON
3736|CHERNOFSKI
3737|CHEROKEE
3738|CHEROKEE CITY
3739|CHEROKEE FALLS
3740|CHEROKEE PASS
3741|CHEROKEE STRIP
3742|CHEROKEE VILLAGE
3743|CHERRY
3744|CHERRY CREEK
3745|CHERRY FORK
3746|CHERRY GROVE
3747|CHERRY GROVE BEACH
3748|CHERRY HILL
3749|CHERRY HILL MALL
3750|CHERRY HILLS VILLAGE
3751|CHERRY LOG
3752|CHERRY SPRING
3753|CHERRY TREE
3754|CHERRY VALLEY
3755|CHERRYLAND
3756|CHERRYPLAIN
3757|CHERRYVALE
3758|CHERRYVILLE
3759|CHESANING
3760|CHESAPEAKE
3761|CHESAPEAKE BEACH
3762|CHESAPEAKE CITY
3763|CHESAPEAKE RANCH ESTATES
3764|CHESAW
3765|CHESHIRE
3766|CHESILHURST
3767|CHESNEE
3768|CHEST SPRINGS
3769|CHESTER
3770|CHESTER GAP
3771|CHESTER HEIGHTS
3772|CHESTER HILL
3773|CHESTER SPRINGS
3774|CHESTERBROOK
3775|CHESTERFIELD
3776|CHESTERHILL
3777|CHESTERLAND
3778|CHESTERTON
3779|CHESTERTOWN
3780|CHESTERVILLE
3781|CHESTNUT
3782|CHESTNUT MOUND
3783|CHESTNUT MOUNTAIN
3784|CHESTNUT RIDGE
3785|CHESUNCOOK
3786|CHESWICK
3787|CHESWOLD
3788|CHETEK
3789|CHETOPA
3790|CHEVAK
3791|CHEVAL
3792|CHEVERLY
3793|CHEVIOT
3794|CHEVY CHASE
3795|CHEVY CHASE HEIGHTS
3796|CHEVY CHASE SECTION FIVE
3797|CHEVY CHASE SECTION THREE
3798|CHEVY CHASE VIEW
3799|CHEVY CHASE VILLAGE
3800|CHEWALLA
3801|CHEWELAH
3802|CHEWEY
3803|CHEWSVILLE
3804|CHEWTON
3805|CHEYENNE
3806|CHEYENNE WELLS
3807|CHEYNEY
3808|CHIAWULI TAK
3809|CHICAGO
3810|CHICAGO HEIGHTS
3811|CHICAGO RIDGE
3812|CHICAL
3813|CHICKALAH
3814|CHICKALOON
3815|CHICKAMAUGA
3816|CHICKAMAW BEACH
3817|CHICKASAW
3818|CHICKASHA
3819|CHICKEN
3820|CHICO
3821|CHICO HOT SPRINGS
3822|CHICOPEE
3823|CHICORA
3824|CHICOT
3825|CHIDESTER
3826|CHIEF LAKE
3827|CHIEFLAND
3828|CHIGNIK
3829|CHIGNIK LAGOON
3830|CHIGNIK LAKE
3831|CHILCHINBITO
3832|CHILDERSBURG
3833|CHILDRESS
3834|CHILDS
3835|CHILES
3836|CHILHOWEE
3837|CHILHOWIE
3838|CHILI
3839|CHILILI
3840|CHILLICOTHE
3841|CHILLUM
3842|CHILLY
3843|CHILO
3844|CHILOCCO
3845|CHILOQUIN
3846|CHILSON
3847|CHILTON
3848|CHIMACUM
3849|CHIMAYO
3850|CHIMNEY ROCK
3851|CHINA
3852|CHINA GROVE
3853|CHINA LAKE ACRES
3854|CHINA SPRINGS
3855|CHINCHILLA
3856|CHINCOTEAGUE
3857|CHINESE CAMP
3858|CHINIAK
3859|CHINLE
3860|CHINO
3861|CHINO HILLS
3862|CHINO VALLEY
3863|CHINOOK
3864|CHINQUAPIN
3865|CHIPITA PARK
3866|CHIPLEY
3867|CHIPPEWA FALLS
3868|CHIPPEWA LAKE
3869|CHIPPEWA PARK
3870|CHIRENO
3871|CHISAGO CITY
3872|CHISANA
3873|CHISHOLM
3874|CHISMVILLE
3875|CHISPA
3876|CHISTOCHINA
3877|CHITINA
3878|CHITTENANGO
3879|CHIVINGTON
3880|CHLORIDE
3881|CHOATE
3882|CHOCCOLOCCO
3883|CHOCOWINITY
3884|CHOCTAW
3885|CHOCTAW BLUFF
3886|CHOCTAW LAKE
3887|CHOKIO
3888|CHOKOLOSKEE
3889|CHOLAME
3890|CHOPIN
3891|CHOPTANK
3892|CHOTEAU
3893|CHOUDRANT
3894|CHOUTEAU
3895|CHOWCHILLA
3896|CHRIESMAN
3897|CHRISMAN
3898|CHRISNEY
3899|CHRISTIANA
3900|CHRISTIANSBURG
3901|CHRISTIANSTED
3902|CHRISTIE
3903|CHRISTINA
3904|CHRISTINE
3905|CHRISTMAS
3906|CHRISTOPHER
3907|CHRISTOPHER CREEK
3908|CHRISTOVAL
3909|CHRISTY MANOR
3910|CHROMO
3911|CHRYSLER
3912|CHUALAR
3913|CHUATHBALUK
3914|CHUBBUCK
3915|CHUGCREEK
3916|CHUGIAK
3917|CHUGWATER
3918|CHUICHU
3919|CHULA
3920|CHULA VISTA
3921|CHULA VISTA COLONIA
3922|CHULUOTA
3923|CHUMS CORNER
3924|CHUMUCKLA
3925|CHUNCHULA
3926|CHUNKY
3927|CHUPADERO
3928|CHURCH CREEK
3929|CHURCH HILL
3930|CHURCH POINT
3931|CHURCH ROCK
3932|CHURCHILL
3933|CHURCHS FERRY
3934|CHURCHTON
3935|CHURCHTOWN
3936|CHURCHVILLE
3937|CHURDAN
3938|CHURUBUSCO
3939|CIALES
3940|CIALES ZONA URBANA
3941|CIBECUE
3942|CIBOLA
3943|CIBOLO
3944|CICERO
3945|CIDRA
3946|CIDRA ZONA URBANA
3947|CIENEGA SPRINGS
3948|CIENEGAS TERRACE
3949|CIMA
3950|CIMARRON
3951|CIMARRON CITY
3952|CIMARRON HILLS
3953|CINCINNATI
3954|CINCO BAYOU
3955|CINCO RANCH
3956|CINEBAR
3957|CINNAMINSON
3958|CIRCLE
3959|CIRCLE HOT SPRINGS
3960|CIRCLE PINES
3961|CIRCLEVILLE
3962|CISCO
3963|CISNE
3964|CISSNA PARK
3965|CISTERN
3966|CITRA
3967|CITRONELLE
3968|CITRUS
3969|CITRUS CITY
3970|CITRUS HEIGHTS
3971|CITRUS HILLS
3972|CITRUS PARK
3973|CITRUS SPRINGS
3974|CITY OF MILFORD (BALANCE)
3975|CITY TERRACE
3976|CITY VIEW
3977|CITY VIEW HEIGHTS
3978|CLAFLIN
3979|CLAIBORNE
3980|CLAIRE CITY
3981|CLAIREMONT
3982|CLAIRETTE
3983|CLAIRFIELD
3984|CLAIRTON
3985|CLALLAM BAY
3986|CLAM GULCH
3987|CLAM LAKE
3988|CLANCY
3989|CLANTON
3990|CLARA
3991|CLARA CITY
3992|CLARCONA
3993|CLARE
3994|CLAREMONT
3995|CLAREMORE
3996|CLARENCE
3997|CLARENCE CENTER
3998|CLARENCEVILLE
3999|CLARENDON
4000|CLARENDON HILLS
4001|CLARIDGE
4002|CLARINDA
4003|CLARINGTON
4004|CLARION
4005|CLARISSA
4006|CLARITA
4007|CLARK
4008|CLARK CENTER
4009|CLARK FORK
4010|CLARK MILLS
4011|CLARKDALE
4012|CLARKEDALE
4013|CLARKESVILLE
4014|CLARKFIELD
4015|CLARKLAKE
4016|CLARKRANGE
4017|CLARKRIDGE
4018|CLARKS
4019|CLARKS GREEN
4020|CLARKS GROVE
4021|CLARKS HILL
4022|CLARKS POINT
4023|CLARKS SUMMIT
4024|CLARKSBORO
4025|CLARKSBURG
4026|CLARKSDALE
4027|CLARKSFIELD
4028|CLARKSON
4029|CLARKSON VALLEY
4030|CLARKSTON
4031|CLARKSTON HEIGHTS
4032|CLARKSVILLE
4033|CLARKSVILLE CITY
4034|CLARKTON
4035|CLARKTOWN
4036|CLARYSVILLE
4037|CLARYVILLE
4038|CLATONIA
4039|CLATSKANIE
4040|CLAUDE
4041|CLAUDELL
4042|CLAUENE
4043|CLAUNCH
4044|CLAWSON
4045|CLAXTON
4046|CLAY
4047|CLAY CENTER
4048|CLAY CITY
4049|CLAY SPRINGS
4050|CLAY VILLAGE
4051|CLAYCOMO
4052|CLAYHATCHEE
4053|CLAYMONT
4054|CLAYPOOL
4055|CLAYPOOL HILL
4056|CLAYSBURG
4057|CLAYSVILLE
4058|CLAYTON
4059|CLAYTON LAKE
4060|CLAYVILLE
4061|CLE ELUM
4062|CLEAR CREEK
4063|CLEAR LAKE
4064|CLEAR LAKE CITY
4065|CLEAR LAKE SHORES
4066|CLEAR SPRING
4067|CLEAR SPRINGS
4068|CLEARBROOK
4069|CLEARBROOK PARK
4070|CLEARCO
4071|CLEARFIELD
4072|CLEARLAKE
4073|CLEARLAKE OAKS
4074|CLEARMONT
4075|CLEARVIEW
4076|CLEARVIEW ACRES
4077|CLEARWATER
4078|CLEARWATER LAKE
4079|CLEARY
4080|CLEATON
4081|CLEATOR
4082|CLEBURNE
4083|CLEGHORN
4084|CLEM
4085|CLEMENTON
4086|CLEMENTS
4087|CLEMENTSON
4088|CLEMENTSVILLE
4089|CLEMMONS
4090|CLEMONS
4091|CLEMSON
4092|CLENDENIN
4093|CLEO
4094|CLEO SPRINGS
4095|CLEONA
4096|CLEONE
4097|CLEORA
4098|CLERMONT
4099|CLETA
4100|CLEVELAND
4101|CLEVELAND HEIGHTS
4102|CLEVER
4103|CLEVES
4104|CLEWISTON
4105|CLICQUOT
4106|CLIFF
4107|CLIFF VILLAGE
4108|CLIFFDELL
4109|CLIFFORD
4110|CLIFFSIDE
4111|CLIFFSIDE PARK
4112|CLIFFTOP
4113|CLIFFWOOD
4114|CLIFFWOOD BEACH
4115|CLIFTON
4116|CLIFTON CITY
4117|CLIFTON FORGE
4118|CLIFTON HEIGHTS
4119|CLIFTON HILL
4120|CLIFTON SPRINGS
4121|CLIFTY
4122|CLIMAX
4123|CLIMAX SPRINGS
4124|CLIMBING HILL
4125|CLINCHCO
4126|CLINCHPORT
4127|CLINE
4128|CLINES CORNERS
4129|CLINT
4130|CLINTON
4131|CLINTONDALE
4132|CLINTONVILLE
4133|CLINTWOOD
4134|CLIO
4135|CLIPPER MILLS
4136|CLITHERALL
4137|CLIVE
4138|CLONTARF
4139|CLOPTON
4140|CLOQUET
4141|CLOSPLINT
4142|CLOSTER
4143|CLOUD CREEK
4144|CLOUD LAKE
4145|CLOUDCROFT
4146|CLOVER
4147|CLOVER BANK
4148|CLOVERDALE
4149|CLOVERLEAF
4150|CLOVERLY
4151|CLOVERPORT
4152|CLOVERTON
4153|CLOVIS
4154|CLOW
4155|CLUSTER SPRINGS
4156|CLUTE
4157|CLUTIER
4158|CLYATTVILLE
4159|CLYDE
4160|CLYDE HILL
4161|CLYDE PARK
4162|CLYMAN
4163|CLYMER
4164|CLYO
4165|CO-OPERATIVE
4166|COACHELLA
4167|COADY
4168|COAHOMA
4169|COAL
4170|COAL CENTER
4171|COAL CITY
4172|COAL CREEK
4173|COAL FORK
4174|COAL GROVE
4175|COAL HILL
4176|COAL MOUNTAIN
4177|COAL RUN
4178|COAL RUN VILLAGE
4179|COAL VALLEY
4180|COALDALE
4181|COALFIELD
4182|COALGATE
4183|COALING
4184|COALINGA
4185|COALMONT
4186|COALPORT
4187|COALRIDGE
4188|COALTON
4189|COALVILLE
4190|COALWOOD
4191|COAMO
4192|COAMO ZONA URBANA
4193|COARSEGOLD
4194|COATES
4195|COATESVILLE
4196|COATS
4197|COATSBURG
4198|COBALT
4199|COBALT VILLAGE
4200|COBB
4201|COBB ISLAND
4202|COBBTOWN
4203|COBDEN
4204|COBLE
4205|COBLESKILL
4206|COBRE
4207|COBURG
4208|COBURN
4209|COCHISE
4210|COCHITI
4211|COCHITI LAKE
4212|COCHITUATE
4213|COCHRAN
4214|COCHRANE
4215|COCHRANTON
4216|COCHRANVILLE
4217|COCKEYSVILLE
4218|COCKRELL HILL
4219|COCKRUM
4220|COCO
4221|COCO COMUNIDAD
4222|COCOA
4223|COCOA BEACH
4224|COCODRIE
4225|COCOLALLA
4226|COCONUT
4227|COCONUT CREEK
4228|CODELL
4229|CODMAN
4230|CODY
4231|COE
4232|COEBURN
4233|COELLO
4234|COEUR D'ALENE
4235|COFFEE CITY
4236|COFFEE CREEK
4237|COFFEE SPRINGS
4238|COFFEEN
4239|COFFEEVILLE
4240|COFFEY
4241|COFFEYVILLE
4242|COFFMAN
4243|COFFMAN COVE
4244|COFIELD
4245|COGAR
4246|COGDELL
4247|COGGON
4248|COGSWELL
4249|COHAGEN
4250|COHASSET
4251|COHASSETT BEACH
4252|COHOCTAH
4253|COHOCTON
4254|COHOE
4255|COHOES
4256|COHUTTA
4257|COILA
4258|COIN
4259|COINJOCK
4260|COKATO
4261|COKEBURG
4262|COKEDALE
4263|COKER
4264|COKESBURY
4265|COKETON
4266|COKEVILLE
4267|COLBERT
4268|COLBURN
4269|COLBY
4270|COLCHESTER
4271|COLCORD
4272|COLD BAY
4273|COLD BROOK
4274|COLD SPRING
4275|COLD SPRING HARBOR
4276|COLD SPRINGS
4277|COLDFOOT
4278|COLDIRON
4279|COLDSPRING
4280|COLDSTREAM
4281|COLDWATER
4282|COLE
4283|COLE CAMP
4284|COLEBROOK
4285|COLEHARBOR
4286|COLEMAN
4287|COLEMANS LAKE
4288|COLERAIN
4289|COLERAIN HEIGHTS
4290|COLERAINE
4291|COLERIDGE
4292|COLES
4293|COLESBURG
4294|COLESVILLE
4295|COLETA
4296|COLETOWN
4297|COLEVILLE
4298|COLFAX
4299|COLGATE
4300|COLLBRAN
4301|COLLEGE
4302|COLLEGE CITY
4303|COLLEGE CORNER
4304|COLLEGE GROVE
4305|COLLEGE HEIGHTS
4306|COLLEGE PARK
4307|COLLEGE PLACE
4308|COLLEGE SPRINGS
4309|COLLEGE STATION
4310|COLLEGEDALE
4311|COLLEGEVILLE
4312|COLLETTSVILLE
4313|COLLEYVILLE
4314|COLLIERVILLE
4315|COLLINGDALE
4316|COLLINGS LAKES
4317|COLLINGSWOOD
4318|COLLINGWOOD PARK
4319|COLLINS
4320|COLLINS PARK
4321|COLLINSBURG
4322|COLLINSTON
4323|COLLINSVILLE
4324|COLLINWOOD
4325|COLLIS
4326|COLLISON
4327|COLLYER
4328|COLMA
4329|COLMAN
4330|COLMAR
4331|COLMAR MANOR
4332|COLMESNEIL
4333|COLMOR
4334|COLO
4335|COLOGNE
4336|COLOMA
4337|COLOME
4338|COLONA
4339|COLONIA
4340|COLONIA IGLESIA ANTIGUA
4341|COLONIAL BEACH
4342|COLONIAL HEIGHTS
4343|COLONIAL PARK
4344|COLONIAL PINE HILLS
4345|COLONIAL VILLAGE
4346|COLONIE
4347|COLONY
4348|COLONY PARK
4349|COLORADO
4350|COLORADO CITY
4351|COLORADO SPRINGS
4352|COLP
4353|COLQUITT
4354|COLSON
4355|COLSTRIP
4356|COLT
4357|COLTON
4358|COLTS NECK
4359|COLUMBIA
4360|COLUMBIA CITY
4361|COLUMBIA FALLS
4362|COLUMBIA HEIGHTS
4363|COLUMBIA HILLS CORNERS
4364|COLUMBIA STATION
4365|COLUMBIANA
4366|COLUMBIAVILLE
4367|COLUMBINE
4368|COLUMBINE VALLEY
4369|COLUMBUS
4370|COLUMBUS CITY
4371|COLUMBUS GROVE
4372|COLUMBUS JUNCTION
4373|COLUSA
4374|COLVER
4375|COLVILLE
4376|COLVOS
4377|COLWELL
4378|COLWICH
4379|COLWYN
4380|COMAL
4381|COMANCHE
4382|COMBEE SETTLEMENT
4383|COMBES
4384|COMBINE
4385|COMBINED LOCKS
4386|COMBS
4387|COMER
4388|COMERTOWN
4389|COMERÍO
4390|COMERÍO ZONA URBANA
4391|COMFORT
4392|COMFREY
4393|COMMACK
4394|COMMERCE
4395|COMMERCE CITY
4396|COMMERCIAL POINT
4397|COMMODORE
4398|COMMONWEALTH
4399|COMO
4400|COMOBABI
4401|COMPASS LAKE
4402|COMPETITION
4403|COMPTCHE
4404|COMPTON
4405|COMSTOCK
4406|COMSTOCK PARK
4407|COMUNAS
4408|COMUNAS COMUNIDAD
4409|COMUS
4410|CONASAUGA
4411|CONASHAUGH LAKES
4412|CONATA
4413|CONCAN
4414|CONCEPCION
4415|CONCEPTION
4416|CONCEPTION JUNCTION
4417|CONCESSION
4418|CONCHAS
4419|CONCHO
4420|CONCONULLY
4421|CONCORD
4422|CONCORDIA
4423|CONCORDVILLE
4424|CONCOW
4425|CONCRETE
4426|CONDA
4427|CONDE
4428|CONDIT
4429|CONDON
4430|CONE
4431|CONEHATTA
4432|CONEJO
4433|CONEJOS
4434|CONEMAUGH
4435|CONESTOGA
4436|CONESVILLE
4437|CONETOE
4438|CONEY ISLAND
4439|CONFLUENCE
4440|CONGER
4441|CONGERS
4442|CONGERVILLE
4443|CONGRESS
4444|CONGRUITY
4445|CONIFER
4446|CONKLING PARK
4447|CONLEN
4448|CONLEY
4449|CONNEAUT
4450|CONNEAUT LAKE
4451|CONNEAUTVILLE
4452|CONNELL
4453|CONNELLSVILLE
4454|CONNELLY SPRINGS
4455|CONNER
4456|CONNERSVILLE
4457|CONNERVILLE
4458|CONNOQUENESSING
4459|CONNORSVILLE
4460|CONNORVILLE
4461|CONOVER
4462|CONRAD
4463|CONRATH
4464|CONROE
4465|CONROY
4466|CONSHOHOCKEN
4467|CONSTABLEVILLE
4468|CONSTANTIA
4469|CONSTANTINE
4470|CONTINENTAL
4471|CONTINENTAL DIVIDE
4472|CONTOOCOOK
4473|CONTRA COSTA CENTRE
4474|CONTRERAS
4475|CONVENT
4476|CONVERSE
4477|CONVOY
4478|CONWAY
4479|CONWAY SPRINGS
4480|CONYERS
4481|CONYNGHAM
4482|COOK
4483|COOK STATION
4484|COOKE CITY
4485|COOKEVILLE
4486|COOKIETOWN
4487|COOKS HAMMOCK
4488|COOKSVILLE
4489|COOKVILLE
4490|COOL
4491|COOL SPRINGS
4492|COOL VALLEY
4493|COOLEEMEE
4494|COOLIDGE
4495|COOLIN
4496|COOLVILLE
4497|COON RAPIDS
4498|COON VALLEY
4499|COOPER
4500|COOPER CITY
4501|COOPER HEIGHTS
4502|COOPER LANDING
4503|COOPERDALE
4504|COOPERS PLAINS
4505|COOPERSBURG
4506|COOPERSTOWN
4507|COOPERSVILLE
4508|COOPERTON
4509|COOPERTOWN
4510|COOS BAY
4511|COOSA
4512|COOSADA
4513|COOSAWHATCHIE
4514|COOTER
4515|COPAKE FALLS
4516|COPAKE LAKE
4517|COPALIS BEACH
4518|COPALIS CROSSING
4519|COPAN
4520|COPE
4521|COPELAND
4522|COPEMISH
4523|COPENHAGEN
4524|COPEVILLE
4525|COPIAGUE
4526|COPLAY
4527|COPLEY
4528|COPPELL
4529|COPPER CANYON
4530|COPPER CENTER
4531|COPPER CITY
4532|COPPER HARBOR
4533|COPPER HILL
4534|COPPER MOUNTAIN
4535|COPPERAS COVE
4536|COPPERFIELD
4537|COPPERHILL
4538|COPPEROPOLIS
4539|COPPERTON
4540|COPPOCK
4541|COQUILLE
4542|COQUÍ
4543|COQUÍ COMUNIDAD
4544|CORA
4545|CORAL
4546|CORAL BAY
4547|CORAL GABLES
4548|CORAL HILLS
4549|CORAL SPRINGS
4550|CORAL TERRACE
4551|CORALVILLE
4552|CORAM
4553|CORAOPOLIS
4554|CORAZÓN
4555|CORAZÓN COMUNIDAD
4556|CORBET
4557|CORBETT
4558|CORBIN
4559|CORBIN CITY
4560|CORCORAN
4561|CORCOVADO
4562|CORCOVADO COMUNIDAD
4563|CORDAVILLE
4564|CORDELE
4565|CORDELL
4566|CORDER
4567|CORDES LAKES
4568|CORDOVA
4569|CORDRY SWEETWATER LAKES
4570|CORE
4571|CORFU
4572|CORINNE
4573|CORINTH
4574|CORLEY
4575|CORMORANT
4576|CORN
4577|CORN CREEK
4578|CORNELIA
4579|CORNELIUS
4580|CORNELL
4581|CORNERSTONE
4582|CORNERSVILLE
4583|CORNERVILLE
4584|CORNETTSVILLE
4585|CORNFIELDS
4586|CORNING
4587|CORNISH
4588|CORNLAND
4589|CORNLEA
4590|CORNUCOPIA
4591|CORNUDAS
4592|CORNVILLE
4593|CORNWALL
4594|CORNWALL-ON-HUDSON
4595|CORNWELL
4596|CORNWELLS HEIGHTS
4597|COROLLA
4598|CORONA
4599|CORONA DE TUCSON
4600|CORONACA
4601|CORONADO
4602|COROZAL
4603|COROZAL ZONA URBANA
4604|CORPUS CHRISTI
4605|CORRAL CITY
4606|CORRAL VIEJO
4607|CORRAL VIEJO COMUNIDAD
4608|CORRALES
4609|CORRALITOS
4610|CORRECTIONVILLE
4611|CORRELL
4612|CORREO
4613|CORRIGAN
4614|CORRIGANVILLE
4615|CORRY
4616|CORRYTON
4617|CORSICA
4618|CORSICANA
4619|CORTARO
4620|CORTE MADERA
4621|CORTEZ
4622|CORTLAND
4623|CORUM
4624|CORUNNA
4625|CORVALLIS
4626|CORWIN
4627|CORWIN SPRINGS
4628|CORWITH
4629|CORY
4630|CORYDON
4631|CORYVILLE
4632|COS COB
4633|COSBY
4634|COSGRAVE
4635|COSHOCTON
4636|COSMOPOLIS
4637|COSMOS
4638|COST
4639|COSTA MESA
4640|COSTILLA
4641|COTATI
4642|COTEAU
4643|COTEAU HOLMES
4644|COTESFIELD
4645|COTO DE CAZA
4646|COTO LAUREL
4647|COTO LAUREL COMUNIDAD
4648|COTO NORTE
4649|COTO NORTE COMUNIDAD
4650|COTOPAXI
4651|COTTAGE CITY
4652|COTTAGE GROVE
4653|COTTAGE HILL
4654|COTTAGE HILLS
4655|COTTAGE LAKE
4656|COTTAGEVILLE
4657|COTTER
4658|COTTLEVILLE
4659|COTTON
4660|COTTON CENTER
4661|COTTON CITY
4662|COTTON PLANT
4663|COTTON VALLEY
4664|COTTONDALE
4665|COTTONPORT
4666|COTTONTOWN
4667|COTTONWOOD
4668|COTTONWOOD FALLS
4669|COTTONWOOD HEIGHTS
4670|COTTONWOOD SHORES
4671|COTUIT
4672|COTULLA
4673|COUCHWOOD
4674|COUDERAY
4675|COUDERSPORT
4676|COUGAR
4677|COUGHRAN
4678|COULEE
4679|COULEE CITY
4680|COULEE DAM
4681|COULTER
4682|COULTERVILLE
4683|COUNCE
4684|COUNCIL
4685|COUNCIL BLUFFS
4686|COUNCIL GROVE
4687|COUNCIL HILL
4688|COUNTRY CLUB
4689|COUNTRY CLUB ESTATES
4690|COUNTRY CLUB HEIGHTS
4691|COUNTRY CLUB HILLS
4692|COUNTRY CLUB VILLAGE
4693|COUNTRY HOMES
4694|COUNTRY KNOLLS
4695|COUNTRY LAKE ESTATES
4696|COUNTRY LIFE ACRES
4697|COUNTRY SQUIRE LAKES
4698|COUNTRY WALK
4699|COUNTRYSIDE
4700|COUNTY LINE
4701|COUPEVILLE
4702|COUPLAND
4703|COURTDALE
4704|COURTENAY
4705|COURTLAND
4706|COURTNEY
4707|COUSHATTA
4708|COUSINS ISLAND
4709|COVADA
4710|COVE
4711|COVE CITY
4712|COVE CREEK
4713|COVE NECK
4714|COVEDALE
4715|COVEL
4716|COVELO
4717|COVENANT LIFE
4718|COVENTRY
4719|COVENTRY LAKE
4720|COVERDALE
4721|COVERT
4722|COVESVILLE
4723|COVINA
4724|COVINGTON
4725|COWAN
4726|COWAN HEIGHTS
4727|COWANSBURG
4728|COWARD
4729|COWARTS
4730|COWDEN
4731|COWDREY
4732|COWELL
4733|COWEN
4734|COWETA
4735|COWGILL
4736|COWICHE
4737|COWLES
4738|COWLEY
4739|COWLIC
4740|COWLINGTON
4741|COWPENS
4742|COX
4743|COX CITY
4744|COXS MILLS
4745|COXSACKIE
4746|COXTON
4747|COY
4748|COYANOSA
4749|COYLE
4750|COYNE CENTER
4751|COYOTE
4752|COYOTE ACRES
4753|COYOTE WELLS
4754|COYVILLE
4755|COZAD
4756|CRAB ORCHARD
4757|CRABAPPLE
4758|CRABTREE
4759|CRACKERVILLE
4760|CRAFTON
4761|CRAGFORD
4762|CRAGSMOOR
4763|CRAIG
4764|CRAIG BEACH
4765|CRAIGMONT
4766|CRAIGSVILLE
4767|CRAIGTOWN
4768|CRAIGVILLE
4769|CRAINVILLE
4770|CRAMERTON
4771|CRANBERRY LAKE
4772|CRANBURY
4773|CRANDALL
4774|CRANDON
4775|CRANDON LAKES
4776|CRANE
4777|CRANE LAKE
4778|CRANELL
4779|CRANESVILLE
4780|CRANFILLS GAP
4781|CRANFORD
4782|CRANNELL
4783|CRANSTON
4784|CRARY
4785|CRAWFORD
4786|CRAWFORDSVILLE
4787|CRAWFORDVILLE
4788|CRAYNE
4789|CREAL SPRINGS
4790|CREAM RIDGE
4791|CREEDE
4792|CREEDMOOR
4793|CREEKSIDE
4794|CREELS
4795|CREELSBORO
4796|CREIGHTON
4797|CRELLIN
4798|CRENSHAW
4799|CREOLA
4800|CREOLE
4801|CRESAPTOWN
4802|CRESBARD
4803|CRESCENT
4804|CRESCENT BEACH
4805|CRESCENT CITY
4806|CRESCENT MILLS
4807|CRESCENT PARK
4808|CRESCENT SPRINGS
4809|CRESCENT VALLEY
4810|CRESCO
4811|CRESSEY
4812|CRESSKILL
4813|CRESSON
4814|CRESSONA
4815|CREST
4816|CREST HILL
4817|CRESTED BUTTE
4818|CRESTLINE
4819|CRESTON
4820|CRESTONE
4821|CRESTVIEW
4822|CRESTVIEW HILLS
4823|CRESTWOOD
4824|CRESTWOOD VILLAGE
4825|CRESWELL
4826|CRETA
4827|CRETE
4828|CREVE COEUR
4829|CREWE
4830|CRICKET
4831|CRIDER
4832|CRIDERS CORNERS
4833|CRIDERSVILLE
4834|CRIMORA
4835|CRINER
4836|CRIPPLE CREEK
4837|CRISFIELD
4838|CRISMAN
4839|CRITTENDEN
4840|CRIVITZ
4841|CROCKER
4842|CROCKETT
4843|CROCKETTS BLUFF
4844|CROFT
4845|CROFTON
4846|CROGHAN
4847|CROMBERG
4848|CROMPOND
4849|CROMWELL
4850|CROOK
4851|CROOKED CREEK
4852|CROOKED LAKE PARK
4853|CROOKS
4854|CROOKSTON
4855|CROOKSVILLE
4856|CROOM
4857|CROPPER
4858|CROPSEY
4859|CROSBY
4860|CROSBYTON
4861|CROSS
4862|CROSS ANCHOR
4863|CROSS CITY
4864|CROSS CREEK
4865|CROSS CUT
4866|CROSS HILL
4867|CROSS KEYS
4868|CROSS LAKE
4869|CROSS LANES
4870|CROSS MOUNTAIN
4871|CROSS PLAINS
4872|CROSS ROADS
4873|CROSS TIMBER
4874|CROSS TIMBERS
4875|CROSS VILLAGE
4876|CROSSETT
4877|CROSSGATE
4878|CROSSNORE
4879|CROSSROADS
4880|CROSSTOWN
4881|CROSSVILLE
4882|CROSSWICKS
4883|CROSWELL
4884|CROTHERSVILLE
4885|CROTON
4886|CROTON HEIGHTS
4887|CROTON-ON-HUDSON
4888|CROTONVILLE
4889|CROUCH
4890|CROUSE
4891|CROW AGENCY
4892|CROW RIVER
4893|CROWDER
4894|CROWDERS
4895|CROWELL
4896|CROWHEART
4897|CROWLEY
4898|CROWN
4899|CROWN CITY
4900|CROWN HEIGHTS
4901|CROWN POINT
4902|CROWNPOINT
4903|CROWNSVILLE
4904|CROWS BLUFF
4905|CROWS LANDING
4906|CROWS NEST
4907|CROYDON
4908|CROZET
4909|CROZIER
4910|CRUCERO
4911|CRUCIBLE
4912|CRUGER
4913|CRUGERS
4914|CRUM
4915|CRUMP
4916|CRUMPLER
4917|CRUMSTOWN
4918|CRUSO
4919|CRUTCHFIELD
4920|CRUZ BAY
4921|CRUZVILLE
4922|CRYSTAL
4923|CRYSTAL BAY
4924|CRYSTAL BEACH
4925|CRYSTAL CITY
4926|CRYSTAL FALLS
4927|CRYSTAL HILL
4928|CRYSTAL LAKE
4929|CRYSTAL LAKE PARK
4930|CRYSTAL LAKES
4931|CRYSTAL LAWNS
4932|CRYSTAL RIVER
4933|CRYSTAL ROCK
4934|CRYSTAL SPRINGS
4935|CRYSTOLA
4936|CUBA
4937|CUBA CITY
4938|CUBERO
4939|CUCHARA
4940|CUCUMBER
4941|CUDAHY
4942|CUDJOE KEY
4943|CUERO
4944|CUERVO
4945|CUEVITAS
4946|CULBERSON
4947|CULBERTSON
4948|CULDESAC
4949|CULEBRA
4950|CULEBRA ZONA URBANA
4951|CULLEN
4952|CULLEOKA
4953|CULLISON
4954|CULLMAN
4955|CULLODEN
4956|CULLOM
4957|CULLOMBURG
4958|CULLOWHEE
4959|CULMERVILLE
4960|CULP CREEK
4961|CULPEPER
4962|CULVER
4963|CULVER CITY
4964|CULVERTON
4965|CUMBERLAND
4966|CUMBERLAND CENTER
4967|CUMBERLAND CITY
4968|CUMBERLAND FURNACE
4969|CUMBERLAND GAP
4970|CUMBERLAND HEAD
4971|CUMBERLAND HILL
4972|CUMBOLA
4973|CUMBY
4974|CUMINGS
4975|CUMMING
4976|CUMMINGS
4977|CUMMINSVILLE
4978|CUNDIFF
4979|CUNDIYO
4980|CUNEY
4981|CUNNINGHAM
4982|CUPERTINO
4983|CUPRUM
4984|CURLEW
4985|CURRAN
4986|CURRIE
4987|CURRITUCK
4988|CURRY
4989|CURRYVILLE
4990|CURTICE
4991|CURTIN
4992|CURTIS
4993|CURTISS
4994|CURTISVILLE
4995|CURWENSVILLE
4996|CUSHING
4997|CUSHMAN
4998|CUSICK
4999|CUSSETA
5000|CUSSON
5001|CUSTAR
5002|CUSTER
5003|CUSTER CITY
5004|CUT AND SHOOT
5005|CUT BANK
5006|CUT OFF
5007|CUTCHOGUE
5008|CUTHBERT
5009|CUTLER
5010|CUTLER BAY
5011|CUTLERVILLE
5012|CUTTEN
5013|CUTTER
5014|CUYAHOGA FALLS
5015|CUYAHOGA HEIGHTS
5016|CUYAMA
5017|CUYAMUNGUE
5018|CUYLER
5019|CUYLERVILLE
5020|CUYUNA
5021|CUZCO
5022|CUZZART
5023|CYCLONE
5024|CYGNET
5025|CYLINDER
5026|CYNTHIANA
5027|CYPERT
5028|CYPRESS
5029|CYPRESS GARDENS
5030|CYPRESS INN
5031|CYPRESS LAKE
5032|CYPRESS QUARTERS
5033|CYRIL
5034|CYRUS
5035|CÉSAR CHÁVEZ
5036|D'HANIS
5037|D'IBERVILLE
5038|D'LO
5039|DACOMA
5040|DACONO
5041|DACULA
5042|DADE CITY
5043|DADEVILLE
5044|DAFTER
5045|DAGGETT
5046|DAGMAR
5047|DAGSBORO
5048|DAGUAO
5049|DAGUAO COMUNIDAD
5050|DAHLEN
5051|DAHLGREN
5052|DAHLIA
5053|DAHLONEGA
5054|DAILEY
5055|DAINGERFIELD
5056|DAIRY
5057|DAISETTA
5058|DAISY
5059|DAISYTOWN
5060|DAKOTA
5061|DAKOTA CITY
5062|DAKOTA DUNES
5063|DALARK
5064|DALBO
5065|DALCOUR
5066|DALE
5067|DALE CITY
5068|DALEVILLE
5069|DALEYVILLE
5070|DALHART
5071|DALIES
5072|DALKEITH
5073|DALKENA
5074|DALLARDSVILLE
5075|DALLAS
5076|DALLAS CENTER
5077|DALLAS CITY
5078|DALLASBURG
5079|DALLASTOWN
5080|DALLESPORT
5081|DALMATIA
5082|DALTON
5083|DALTON CITY
5084|DALTON GARDENS
5085|DALWORTHINGTON GARDENS
5086|DALY CITY
5087|DALZELL
5088|DAMAR
5089|DAMARISCOTTA
5090|DAMASCUS
5091|DAMES FERRY
5092|DAMES QUARTER
5093|DAMIANSVILLE
5094|DAMMERON VALLEY
5095|DAMON
5096|DAN
5097|DANA
5098|DANA POINT
5099|DANBURY
5100|DANDRIDGE
5101|DANE
5102|DANEVANG
5103|DANFORTH
5104|DANIA BEACH
5105|DANIEL
5106|DANIELS
5107|DANIELSON
5108|DANIELSVILLE
5109|DANNEBROG
5110|DANNEMORA
5111|DANSVILLE
5112|DANTE
5113|DANUBE
5114|DANVERS
5115|DANVILLE
5116|DAPHNE
5117|DAPHNEDALE PARK
5118|DARBUN
5119|DARBY
5120|DARBYDALE
5121|DARBYVILLE
5122|DARCO
5123|DARDANELLE
5124|DARDEN
5125|DARDENNE PRAIRIE
5126|DARES BEACH
5127|DARFUR
5128|DARGAN
5129|DARIEN
5130|DARLING
5131|DARLINGTON
5132|DARLOVE
5133|DARMSTADT
5134|DARNELL
5135|DARNESTOWN
5136|DARR
5137|DARRAGH
5138|DARRINGTON
5139|DARROUZETT
5140|DARRTOWN
5141|DARWIN
5142|DASH POINT
5143|DASHER
5144|DASSEL
5145|DATELAND
5146|DATIL
5147|DATTO
5148|DAUBERVILLE
5149|DAUFUSKIE LANDING
5150|DAUPHIN
5151|DAUPHIN ISLAND
5152|DAUS
5153|DAVANT
5154|DAVENPORT
5155|DAVENPORT CENTER
5156|DAVEY
5157|DAVID
5158|DAVID CITY
5159|DAVIDSON
5160|DAVIDSON HEIGHTS
5161|DAVIDSONVILLE
5162|DAVIDSVILLE
5163|DAVIE
5164|DAVILLA
5165|DAVIS
5166|DAVIS CITY
5167|DAVIS DAM
5168|DAVIS JUNCTION
5169|DAVISBORO
5170|DAVISON
5171|DAVISTON
5172|DAVISVILLE
5173|DAVY
5174|DAWESVILLE
5175|DAWN
5176|DAWSON
5177|DAWSON SPRINGS
5178|DAWSONVILLE
5179|DAY HEIGHTS
5180|DAY VALLEY
5181|DAYKIN
5182|DAYS CREEK
5183|DAYSVILLE
5184|DAYTON
5185|DAYTON LAKES
5186|DAYTONA BEACH
5187|DAYTONA BEACH SHORES
5188|DAYVILLE
5189|DAZEY
5190|DE ANN
5191|DE BEQUE
5192|DE BERRY
5193|DE BORGIA
5194|DE FOREST
5195|DE FUNIAK SPRINGS
5196|DE GRAFF
5197|DE KALB
5198|DE KALB JUNCTION
5199|DE LAMERE
5200|DE LANCEY
5201|DE LAND
5202|DE LEON
5203|DE LEON SPRINGS
5204|DE LISLE
5205|DE PERE
5206|DE QUEEN
5207|DE ROSSETT
5208|DE SART
5209|DE SMET
5210|DE SOTO
5211|DE SOTO CITY
5212|DE TOUR VILLAGE
5213|DE VALLS BLUFF
5214|DE WITT
5215|DEADHORSE
5216|DEADWOOD
5217|DEAL
5218|DEAL ISLAND
5219|DEALE
5220|DEAN
5221|DEANS
5222|DEANVILLE
5223|DEARBORN
5224|DEARBORN HEIGHTS
5225|DEARING
5226|DEARMANVILLE
5227|DEARY
5228|DEATSVILLE
5229|DEAVER
5230|DEBARY
5231|DECATUR
5232|DECATUR CITY
5233|DECATURVILLE
5234|DECHERD
5235|DECKER
5236|DECKERVILLE
5237|DECLO
5238|DECORAH
5239|DECORDOVA
5240|DECOY
5241|DEDHAM
5242|DEE
5243|DEEMER
5244|DEEMSTON
5245|DEENWOOD
5246|DEEP CREEK
5247|DEEP GAP
5248|DEEP RIVER
5249|DEEP SPRINGS
5250|DEEP WATER
5251|DEEPHAVEN
5252|DEEPSTEP
5253|DEEPWATER
5254|DEER
5255|DEER CREEK
5256|DEER GROVE
5257|DEER ISLAND
5258|DEER LAKE
5259|DEER LODGE
5260|DEER PARK
5261|DEER RANGE
5262|DEER RIVER
5263|DEER TRAIL
5264|DEERBROOK
5265|DEERFIELD
5266|DEERFIELD BEACH
5267|DEERING
5268|DEERSVILLE
5269|DEERTON
5270|DEERWOOD
5271|DEESON
5272|DEETH
5273|DEFERIET
5274|DEFIANCE
5275|DEKALB
5276|DEKLE BEACH
5277|DEL AIRE
5278|DEL CITY
5279|DEL DIOS
5280|DEL MAR
5281|DEL MAR HEIGHTS
5282|DEL MAR WOODS
5283|DEL MONTE FOREST
5284|DEL MUERTO
5285|DEL NORTE
5286|DEL REY
5287|DEL REY OAKS
5288|DEL RIO
5289|DEL ROSA
5290|DEL SOL COLONIA
5291|DEL VALLE
5292|DELAFIELD
5293|DELANCO
5294|DELAND
5295|DELANO
5296|DELANSON
5297|DELAPLAINE
5298|DELAVAN
5299|DELAVAN LAKE
5300|DELAWARE
5301|DELAWARE CITY
5302|DELAWARE WATER GAP
5303|DELBARTON
5304|DELCAMBRE
5305|DELCO
5306|DELEVAN
5307|DELFT
5308|DELFT COLONY
5309|DELHI
5310|DELHI HILLS
5311|DELIA
5312|DELIGHT
5313|DELL
5314|DELL CITY
5315|DELL RAPIDS
5316|DELLEKER
5317|DELLROY
5318|DELLSLOW
5319|DELLVALE
5320|DELLVIEW
5321|DELLWOOD
5322|DELMAR
5323|DELMITA
5324|DELMONT
5325|DELOIT
5326|DELONG
5327|DELPHI
5328|DELPHIA
5329|DELPHOS
5330|DELRAY
5331|DELRAY BEACH
5332|DELTA
5333|DELTA JUNCTION
5334|DELTAVILLE
5335|DELTON
5336|DELTONA
5337|DELWAY
5338|DEMAREST
5339|DEMING
5340|DEMOCRAT
5341|DEMOPOLIS
5342|DEMOREST
5343|DEMOTTE
5344|DEMPSEY
5345|DENAIR
5346|DENALI PARK
5347|DENAUD
5348|DENBIGH
5349|DENBY
5350|DENDRON
5351|DENHAM
5352|DENHAM SPRINGS
5353|DENHOFF
5354|DENIO
5355|DENISON
5356|DENMARK
5357|DENNARD
5358|DENNEHOTSO
5359|DENNING
5360|DENNIS
5361|DENNIS ACRES
5362|DENNIS PORT
5363|DENNISON
5364|DENNISVILLE
5365|DENSMORE
5366|DENT
5367|DENTON
5368|DENTSVILLE
5369|DENVER
5370|DENVER CITY
5371|DENVILLE
5372|DEORA
5373|DEPAUVILLE
5374|DEPAUW
5375|DEPEW
5376|DEPOE BAY
5377|DEPORT
5378|DEPOSIT
5379|DEPUE
5380|DEPUTY
5381|DEQUINCY
5382|DERBY
5383|DERBY ACRES
5384|DERBY CENTER
5385|DERBY LINE
5386|DERIDDER
5387|DERING HARBOR
5388|DERITA
5389|DERMA
5390|DERMOTT
5391|DERRICK CITY
5392|DERRY
5393|DERUYTER
5394|DERWOOD
5395|DES ALLEMANDS
5396|DES ARC
5397|DES LACS
5398|DES MOINES
5399|DES PERES
5400|DES PLAINES
5401|DESCANSO
5402|DESCHUTES RIVER WOODS
5403|DESDEMONA
5404|DESERET
5405|DESERT
5406|DESERT AIRE
5407|DESERT CENTER
5408|DESERT EDGE
5409|DESERT HILLS
5410|DESERT HOT SPRINGS
5411|DESERT SHORES
5412|DESERT VIEW HIGHLANDS
5413|DESHA
5414|DESHLER
5415|DESLOGE
5416|DESOTO
5417|DESOTO LAKES
5418|DESPARD
5419|DESTIN
5420|DESTREHAN
5421|DETMOLD
5422|DETONTI
5423|DETROIT
5424|DETROIT BEACH
5425|DETROIT LAKES
5426|DEVAULT
5427|DEVENS
5428|DEVEREUX
5429|DEVERS
5430|DEVILLE
5431|DEVILS LAKE
5432|DEVILS SLIDE
5433|DEVILS TOWER
5434|DEVINE
5435|DEVOL
5436|DEVOLA
5437|DEVON
5438|DEVORE
5439|DEW
5440|DEWALT
5441|DEWAR
5442|DEWART
5443|DEWEESE
5444|DEWEY
5445|DEWEY BEACH
5446|DEWEY-HUMBOLDT
5447|DEWEYVILLE
5448|DEWITT
5449|DEWY ROSE
5450|DEXTER
5451|DEXTER CITY
5452|DEXTERVILLE
5453|DI GIORGIO
5454|DIABLO
5455|DIABLO GRANDE
5456|DIABLOCK
5457|DIAGONAL
5458|DIALVILLE
5459|DIAMOND
5460|DIAMOND BAR
5461|DIAMOND BEACH
5462|DIAMOND BLUFF
5463|DIAMOND CITY
5464|DIAMOND LAKE
5465|DIAMOND RIDGE
5466|DIAMOND SPRINGS
5467|DIAMONDHEAD
5468|DIAMONDHEAD LAKE
5469|DIAMONDVILLE
5470|DIANA
5471|DIAZ
5472|DIBBLE
5473|DIBOLL
5474|DICKENS
5475|DICKERSON
5476|DICKERSON CITY
5477|DICKEY
5478|DICKEYVILLE
5479|DICKINSON
5480|DICKSON
5481|DICKSON CITY
5482|DICKSONVILLE
5483|DICKWORSHAM
5484|DIEHLSTADT
5485|DIERINGER
5486|DIERKS
5487|DIETERICH
5488|DIETRICH
5489|DIFFICULT
5490|DIGGINS
5491|DIGHTON
5492|DIKE
5493|DILIA
5494|DILKON
5495|DILL CITY
5496|DILLARD
5497|DILLER
5498|DILLEY
5499|DILLINGHAM
5500|DILLON
5501|DILLON BEACH
5502|DILLONVALE
5503|DILLSBORO
5504|DILLSBURG
5505|DILLWYN
5506|DILWORTH
5507|DIME
5508|DIME BOX
5509|DIMMITT
5510|DIMOCK
5511|DIMONDALE
5512|DINERO
5513|DINGMANS FERRY
5514|DINGUS
5515|DINOSAUR
5516|DINUBA
5517|DIOMEDE
5518|DIRGIN
5519|DISAUTEL
5520|DISCOVERY
5521|DISCOVERY BAY
5522|DISCOVERY HARBOUR
5523|DISH
5524|DISHMAN
5525|DISNEY
5526|DISPUTANTA
5527|DISSTON
5528|DISTRICT HEIGHTS
5529|DITTLINGER
5530|DIVERNON
5531|DIVIDE
5532|DIX
5533|DIX HILLS
5534|DIXBORO
5535|DIXFIELD
5536|DIXIE
5537|DIXIE INN
5538|DIXIE UNION
5539|DIXMOOR
5540|DIXON
5541|DIXONS MILLS
5542|DIXONVILLE
5543|DIZNEY
5544|DOBBIN
5545|DOBBINS
5546|DOBBINS HEIGHTS
5547|DOBBS FERRY
5548|DOBSON
5549|DOCK JUNCTION
5550|DOCKTON
5551|DOCTOR PHILLIPS
5552|DOCTORS INLET
5553|DOCTORTOWN
5554|DODD CITY
5555|DODDRIDGE
5556|DODDSVILLE
5557|DODGE
5558|DODGE CENTER
5559|DODGE CITY
5560|DODGE PARK
5561|DODGEVILLE
5562|DODSON
5563|DODSON BRANCH
5564|DODSONVILLE
5565|DOE RUN
5566|DOE VALLEY
5567|DOERING
5568|DOERUN
5569|DOFFING
5570|DOGTOWN
5571|DOLA
5572|DOLAN SPRINGS
5573|DOLAND
5574|DOLES
5575|DOLGEVILLE
5576|DOLLAR BAY
5577|DOLLAR POINT
5578|DOLLIVER
5579|DOLOMITE
5580|DOLORES
5581|DOLTON
5582|DOME
5583|DOMESTIC
5584|DOMINGO
5585|DOMINGUEZ
5586|DOMINION
5587|DOMINO
5588|DONAHUE
5589|DONALD
5590|DONALDS
5591|DONALDSON
5592|DONALDSONVILLE
5593|DONALSONVILLE
5594|DONEGAL
5595|DONGOLA
5596|DONIE
5597|DONIPHAN
5598|DONNA
5599|DONNAN
5600|DONNELLSON
5601|DONNELLY
5602|DONNELSVILLE
5603|DONNER
5604|DONNYBROOK
5605|DONORA
5606|DONOVAN
5607|DOOLE
5608|DOOLING
5609|DOOLITTLE
5610|DOOMS
5611|DOON
5612|DORA
5613|DORADO
5614|DORADO ZONA URBANA
5615|DORAL
5616|DORAN
5617|DORAVILLE
5618|DORCAS
5619|DORCHESTER
5620|DORCHESTER CENTER
5621|DORE
5622|DORENA
5623|DORIS
5624|DORMONT
5625|DORNEYVILLE
5626|DORNSIFE
5627|DOROTHY
5628|DORRANCE
5629|DORRINGTON
5630|DORRIS
5631|DORSET
5632|DORSEY
5633|DORSEYVILLE
5634|DORTCHES
5635|DORTON
5636|DOS CABEZAS
5637|DOS PALOS
5638|DOS PALOS Y
5639|DOS RIOS
5640|DOSSVILLE
5641|DOT LAKE
5642|DOT LAKE VILLAGE
5643|DOTHAN
5644|DOTSERO
5645|DOTY
5646|DOTYVILLE
5647|DOUBLE ADOBE
5648|DOUBLE BAYOU
5649|DOUBLE OAK
5650|DOUBLE SPRINGS
5651|DOUCETTE
5652|DOUDS
5653|DOUGHERTY
5654|DOUGLAS
5655|DOUGLAS CITY
5656|DOUGLASS
5657|DOUGLASS HILLS
5658|DOUGLASSVILLE
5659|DOUGLASVILLE
5660|DOURO
5661|DOUSMAN
5662|DOVE CREEK
5663|DOVE VALLEY
5664|DOVER
5665|DOVER BEACHES NORTH
5666|DOVER BEACHES SOUTH
5667|DOVER HILL
5668|DOVER PLAINS
5669|DOVER-FOXCROFT
5670|DOVRAY
5671|DOW CITY
5672|DOWAGIAC
5673|DOWELL
5674|DOWELLTOWN
5675|DOWLING
5676|DOWLING PARK
5677|DOWNER
5678|DOWNERS GROVE
5679|DOWNEY
5680|DOWNIEVILLE
5681|DOWNING
5682|DOWNINGTOWN
5683|DOWNS
5684|DOWNSVILLE
5685|DOWS
5686|DOYLE
5687|DOYLESTOWN
5688|DOYLEVILLE
5689|DOYLINE
5690|DOZIER
5691|DOÑA ANA
5692|DRACUT
5693|DRAGOON
5694|DRAKE
5695|DRAKES BRANCH
5696|DRAKESBORO
5697|DRAKESVILLE
5698|DRAKETOWN
5699|DRANESVILLE
5700|DRAPER
5701|DRAVOSBURG
5702|DRAYTON
5703|DRESBACH
5704|DRESDEN
5705|DRESSER
5706|DREWRYVILLE
5707|DREXEL
5708|DREXEL HEIGHTS
5709|DREXEL HILL
5710|DRIFTON
5711|DRIFTWOOD
5712|DRIGGS
5713|DRIP ROCK
5714|DRIPPING SPRINGS
5715|DRISCOLL
5716|DRUID HILLS
5717|DRUM POINT
5718|DRUMMOND
5719|DRUMRIGHT
5720|DRY CREEK
5721|DRY FORK
5722|DRY LAKE
5723|DRY PRONG
5724|DRY RIDGE
5725|DRY RUN
5726|DRY TAVERN
5727|DRYDEN
5728|DRYNOB
5729|DRYTOWN
5730|DRYVILLE
5731|DU BOIS
5732|DU PONT
5733|DU QUOIN
5734|DUANE LAKE
5735|DUANESBURG
5736|DUARTE
5737|DUBACH
5738|DUBBERLY
5739|DUBBS
5740|DUBLIN
5741|DUBOIS
5742|DUBOISTOWN
5743|DUBUQUE
5744|DUCHESNE
5745|DUCHESS LANDING
5746|DUCK
5747|DUCK HILL
5748|DUCK KEY
5749|DUCKTOWN
5750|DUCOR
5751|DUDLEY
5752|DUDLEYVILLE
5753|DUE WEST
5754|DUELM
5755|DUENWEG
5756|DUETTE
5757|DUFFIELD
5758|DUFUR
5759|DUGGER
5760|DUGWAY
5761|DUKE
5762|DUKES
5763|DULAC
5764|DULCE
5765|DULLES TOWN CENTER
5766|DULUTH
5767|DUMAS
5768|DUMBARTON
5769|DUMFRIES
5770|DUMONT
5771|DUNBAR
5772|DUNBARTON
5773|DUNCAN
5774|DUNCAN FALLS
5775|DUNCANNON
5776|DUNCANSVILLE
5777|DUNCANVILLE
5778|DUNCOMBE
5779|DUNDALK
5780|DUNDARRACH
5781|DUNDAS
5782|DUNDEE
5783|DUNE ACRES
5784|DUNEAN
5785|DUNEDIN
5786|DUNELLEN
5787|DUNES CITY
5788|DUNFERMLINE
5789|DUNGANNON
5790|DUNGENESS
5791|DUNKEN
5792|DUNKERTON
5793|DUNKINSVILLE
5794|DUNKIRK
5795|DUNLAP
5796|DUNLAP ACRES
5797|DUNLAY
5798|DUNLEVY
5799|DUNLO
5800|DUNLOW
5801|DUNMOR
5802|DUNMORE
5803|DUNN
5804|DUNN CENTER
5805|DUNN LORING
5806|DUNNEGAN
5807|DUNNELL
5808|DUNNELLON
5809|DUNNIGAN
5810|DUNNING
5811|DUNNSTOWN
5812|DUNNVILLE
5813|DUNPHY
5814|DUNREITH
5815|DUNSEITH
5816|DUNSMUIR
5817|DUNTON
5818|DUNWOODY
5819|DUPO
5820|DUPONT
5821|DUPREE
5822|DUPUYER
5823|DUQUE
5824|DUQUE COMUNIDAD
5825|DUQUESNE
5826|DUQUETTE
5827|DUQUOIN
5828|DURAN
5829|DURAND
5830|DURANGO
5831|DURANT
5832|DURBIN
5833|DURHAM
5834|DURHAMVILLE
5835|DURYEA
5836|DUSHORE
5837|DUSON
5838|DUSTER
5839|DUSTIN
5840|DUSTIN ACRES
5841|DUSTY
5842|DUTCH FLAT
5843|DUTCH JOHN
5844|DUTCH MILLS
5845|DUTCHTOWN
5846|DUTTON
5847|DUVALL
5848|DUXBURY
5849|DWALE
5850|DWIGHT
5851|DWIGHT MISSION
5852|DYCKESVILLE
5853|DYCUSBURG
5854|DYER
5855|DYERSBURG
5856|DYERSVILLE
5857|DYESS
5858|DYSART
5859|EADS
5860|EAGAN
5861|EAGAR
5862|EAGERVILLE
5863|EAGLE
5864|EAGLE BEND
5865|EAGLE BUTTE
5866|EAGLE CITY
5867|EAGLE FLAT
5868|EAGLE GROVE
5869|EAGLE HARBOR
5870|EAGLE LAKE
5871|EAGLE MILLS
5872|EAGLE MOUNTAIN
5873|EAGLE NEST
5874|EAGLE PASS
5875|EAGLE POINT
5876|EAGLE RIVER
5877|EAGLE ROCK
5878|EAGLE VALLEY
5879|EAGLE VILLAGE
5880|EAGLEDALE
5881|EAGLEPORT
5882|EAGLES MERE
5883|EAGLETON
5884|EAGLETON VILLAGE
5885|EAGLETOWN
5886|EAGLEVILLE
5887|EAKLY
5888|EARL
5889|EARL PARK
5890|EARLE
5891|EARLHAM
5892|EARLIMART
5893|EARLING
5894|EARLINGTON
5895|EARLSBORO
5896|EARLSTON
5897|EARLTON
5898|EARLVILLE
5899|EARLY BRANCH
5900|EASLEY
5901|EAST ALTON
5902|EAST AMANA
5903|EAST ARCADIA
5904|EAST ATLANTIC BEACH
5905|EAST AURORA
5906|EAST AVON
5907|EAST BANGOR
5908|EAST BANK
5909|EAST BARRE
5910|EAST BEND
5911|EAST BERLIN
5912|EAST BERNARD
5913|EAST BERNSTADT
5914|EAST BERWICK
5915|EAST BETHEL
5916|EAST BRADY
5917|EAST BRANCH
5918|EAST BREWTON
5919|EAST BROOKFIELD
5920|EAST BROOKLYN
5921|EAST BURKE
5922|EAST BUTLER
5923|EAST CAMDEN
5924|EAST CANTON
5925|EAST CAPE GIRARDEAU
5926|EAST CARONDELET
5927|EAST CATHLAMET
5928|EAST CHAIN
5929|EAST CHICAGO
5930|EAST CLARIDON
5931|EAST CLEVELAND
5932|EAST CONEMAUGH
5933|EAST DAILEY
5934|EAST DANVILLE
5935|EAST DENNIS
5936|EAST DOUGLAS
5937|EAST DUBLIN
5938|EAST DUBUQUE
5939|EAST DUNDEE
5940|EAST DUNSEITH
5941|EAST EARL
5942|EAST ELLIJAY
5943|EAST END
5944|EAST ENTERPRISE
5945|EAST FAIRVIEW
5946|EAST FALMOUTH
5947|EAST FARMINGDALE
5948|EAST FARMS
5949|EAST FLAT ROCK
5950|EAST FOOTHILLS
5951|EAST FORK
5952|EAST FREEDOM
5953|EAST FREEHOLD
5954|EAST FULTONHAM
5955|EAST GAFFNEY
5956|EAST GALESBURG
5957|EAST GARDEN CITY
5958|EAST GERMANTOWN
5959|EAST GILLESPIE
5960|EAST GLACIER PARK
5961|EAST GLACIER PARK VILLAGE
5962|EAST GLENVILLE
5963|EAST GRAND FORKS
5964|EAST GRAND RAPIDS
5965|EAST GREENBUSH
5966|EAST GREENVILLE
5967|EAST GRIFFIN
5968|EAST GULL LAKE
5969|EAST HAMPTON
5970|EAST HANOVER
5971|EAST HARTFORD
5972|EAST HARWICH
5973|EAST HAVEN
5974|EAST HAZEL CREST
5975|EAST HELENA
5976|EAST HEMET
5977|EAST HIGHLAND PARK
5978|EAST HIGHLANDS
5979|EAST HILLS
5980|EAST HODGE
5981|EAST HOLDEN
5982|EAST HOPE
5983|EAST ISLIP
5984|EAST ITHACA
5985|EAST JORDAN
5986|EAST JULIETTE
5987|EAST KINGSTON
5988|EAST LA MIRADA
5989|EAST LAKE
5990|EAST LAKE WEIR
5991|EAST LANSDOWNE
5992|EAST LANSING
5993|EAST LAS VEGAS
5994|EAST LAURINBURG
5995|EAST LEAVENWORTH
5996|EAST LEXINGTON
5997|EAST LIBERTY
5998|EAST LIVERPOOL
5999|EAST LOS ANGELES
6000|EAST LYNN
6001|EAST LYNNE
6002|EAST MARION
6003|EAST MASSAPEQUA
6004|EAST MCKEESPORT
6005|EAST MEADOW
6006|EAST MERRIMACK
6007|EAST MIDDLEBURY
6008|EAST MIDDLETOWN
6009|EAST MILLINOCKET
6010|EAST MILLSTONE
6011|EAST MILTON
6012|EAST MISSOULA
6013|EAST MOLINE
6014|EAST MONTPELIER
6015|EAST MORICHES
6016|EAST MOUNTAIN
6017|EAST NAPLES
6018|EAST NASSAU
6019|EAST NEW MARKET
6020|EAST NEWARK
6021|EAST NEWNAN
6022|EAST NICOLAUS
6023|EAST NORTHPORT
6024|EAST NORWICH
6025|EAST OAKDALE
6026|EAST OLYMPIA
6027|EAST ORANGE
6028|EAST OROSI
6029|EAST PALATKA
6030|EAST PALESTINE
6031|EAST PALO ALTO
6032|EAST PASADENA
6033|EAST PATCHOGUE
6034|EAST PECOS
6035|EAST PEORIA
6036|EAST PEPPERELL
6037|EAST PERU
6038|EAST PETERSBURG
6039|EAST PITTSBURGH
6040|EAST POINT
6041|EAST PORT ORCHARD
6042|EAST PORTAL
6043|EAST PORTERVILLE
6044|EAST PRAIRIE
6045|EAST PROSPECT
6046|EAST PROVIDENCE
6047|EAST QUINCY
6048|EAST QUOGUE
6049|EAST RANCHO DOMINGUEZ
6050|EAST RANDOLPH
6051|EAST RENTON HIGHLANDS
6052|EAST RICHMOND HEIGHTS
6053|EAST RIDGE
6054|EAST RINGGOLD
6055|EAST RIVERDALE
6056|EAST ROCHESTER
6057|EAST ROCKAWAY
6058|EAST ROCKINGHAM
6059|EAST ROCKWOOD
6060|EAST RUTHERFORD
6061|EAST SAINT LOUIS
6062|EAST SALEM
6063|EAST SAN GABRIEL
6064|EAST SANDWICH
6065|EAST SETAUKET
6066|EAST SHORE
6067|EAST SHOREHAM
6068|EAST SIDE
6069|EAST SMITHFIELD
6070|EAST SONORA
6071|EAST SPARTA
6072|EAST SPENCER
6073|EAST SPRINGFIELD
6074|EAST STROUDSBURG
6075|EAST SUMTER
6076|EAST SYRACUSE
6077|EAST TAWAKONI
6078|EAST TAWAS
6079|EAST THERMOPOLIS
6080|EAST TRENTON HEIGHTS
6081|EAST TROY
6082|EAST UNIONTOWN
6083|EAST VANDERGRIFT
6084|EAST WALPOLE
6085|EAST WASHINGTON
6086|EAST WATERFORD
6087|EAST WENATCHEE
6088|EAST WHITE PLAINS
6089|EAST WHITTIER
6090|EAST WILLISTON
6091|EAST WILSON
6092|EAST YORK
6093|EASTANOLLEE
6094|EASTBOROUGH
6095|EASTCHESTER
6096|EASTERLY
6097|EASTGATE
6098|EASTHAMPTON
6099|EASTLAKE
6100|EASTLAND
6101|EASTLAWN
6102|EASTLAWN GARDENS
6103|EASTMAN
6104|EASTON
6105|EASTOVER
6106|EASTPOINT
6107|EASTPOINTE
6108|EASTPORT
6109|EASTSOUND
6110|EASTVALE
6111|EASTVIEW
6112|EASTVILLE
6113|EASTWOOD
6114|EASTWOOD MANOR
6115|EATON
6116|EATON ESTATES
6117|EATON PARK
6118|EATON RAPIDS
6119|EATONS NECK
6120|EATONTON
6121|EATONTOWN
6122|EATONVILLE
6123|EAU CLAIRE
6124|EAU GALLIE
6125|EBENEZER
6126|EBENSBURG
6127|EBONY
6128|EBRO
6129|ECCLES
6130|ECHELON
6131|ECHETA
6132|ECKERMAN
6133|ECKHART MINES
6134|ECKLEY
6135|ECKMAN
6136|ECLECTIC
6137|ECONFINA
6138|ECONOMY
6139|ECORSE
6140|ECRU
6141|ECTOR
6142|EDCOUCH
6143|EDDICETON
6144|EDDINGTON
6145|EDDY
6146|EDDYSTONE
6147|EDDYVILLE
6148|EDEN
6149|EDEN ISLE
6150|EDEN PRAIRIE
6151|EDEN ROC
6152|EDEN VALLEY
6153|EDENBORN
6154|EDENBURG
6155|EDENTON
6156|EDENVILLE
6157|EDESVILLE
6158|EDGAR
6159|EDGAR SPRINGS
6160|EDGARD
6161|EDGARTOWN
6162|EDGE
6163|EDGECLIFF VILLAGE
6164|EDGEFIELD
6165|EDGEHILL
6166|EDGELEY
6167|EDGELY
6168|EDGEMERE
6169|EDGEMONT
6170|EDGEMONT PARK
6171|EDGEMOOR
6172|EDGERLY
6173|EDGERTON
6174|EDGEWATER
6175|EDGEWATER ESTATES
6176|EDGEWATER HEIGHTS
6177|EDGEWATER PARK
6178|EDGEWOOD
6179|EDGEWORTH
6180|EDIE
6181|EDINA
6182|EDINBORO
6183|EDINBURG
6184|EDINBURGH
6185|EDISON
6186|EDISTO
6187|EDISTO BEACH
6188|EDISTO ISLAND
6189|EDITH
6190|EDLER
6191|EDMESTON
6192|EDMOND
6193|EDMONDS
6194|EDMONDSON
6195|EDMONSON
6196|EDMONSTON
6197|EDMONTON
6198|EDMORE
6199|EDMUND
6200|EDMUNDSON
6201|EDMUNDSON ACRES
6202|EDNA
6203|EDNA BAY
6204|EDNEYVILLE
6205|EDOM
6206|EDON
6207|EDRAY
6208|EDROY
6209|EDSON
6210|EDWALL
6211|EDWARDS
6212|EDWARDSBURG
6213|EDWARDSPORT
6214|EDWARDSVILLE
6215|EEK
6216|EFFIE
6217|EFFINGHAM
6218|EFFORT
6219|EFLAND
6220|EGAN
6221|EGBERT
6222|EGEGIK
6223|EGELAND
6224|EGG HARBOR
6225|EGG HARBOR CITY
6226|EGGERTSVILLE
6227|EGGLESTON
6228|EGLON
6229|EGNAR
6230|EGYPT
6231|EHRENBERG
6232|EHRENFELD
6233|EHRHARDT
6234|EIDSON ROAD
6235|EIGHTY FOUR
6236|EITZEN
6237|EKALAKA
6238|EKRON
6239|EKWOK
6240|EL CAJON
6241|EL CAMINO ANGOSTO
6242|EL CAMPO
6243|EL CASCO
6244|EL CENIZO
6245|EL CENIZO COLONIA
6246|EL CENTRO
6247|EL CERRITO
6248|EL CERRO
6249|EL COMBATE
6250|EL COMBATE COMUNIDAD
6251|EL DARA
6252|EL DORADO
6253|EL DORADO HILLS
6254|EL DORADO SPRINGS
6255|EL DUENDE
6256|EL GRANADA
6257|EL INDIO
6258|EL JEBEL
6259|EL LAGO
6260|EL MANGÓ
6261|EL MANGÓ COMUNIDAD
6262|EL MIRAGE
6263|EL MONTE
6264|EL MORO
6265|EL NEGRO
6266|EL NEGRO COMUNIDAD
6267|EL NIDO
6268|EL OJO
6269|EL OJO COMUNIDAD
6270|EL PARAISO
6271|EL PARAISO COMUNIDAD
6272|EL PASO
6273|EL PORTAL
6274|EL PORVENIR
6275|EL RANCHO
6276|EL REFUGIO
6277|EL RENO
6278|EL RIO
6279|EL RITO
6280|EL SAUZ
6281|EL SEGUNDO
6282|EL SOBRANTE
6283|EL TORO
6284|EL TUMBAO
6285|EL TUMBAO COMUNIDAD
6286|EL VADO
6287|EL VALLE DE ARROYO SECO
6288|EL VERANO
6289|ELAINE
6290|ELAND
6291|ELBA
6292|ELBE
6293|ELBERFELD
6294|ELBERON
6295|ELBERT
6296|ELBERTA
6297|ELBERTON
6298|ELBING
6299|ELBOW LAKE
6300|ELBRIDGE
6301|ELBURN
6302|ELCHO
6303|ELCO
6304|ELDENA
6305|ELDERON
6306|ELDERSBURG
6307|ELDERTON
6308|ELDERWOOD
6309|ELDON
6310|ELDORA
6311|ELDORADO
6312|ELDORADO AT SANTA FE
6313|ELDORADO SPRINGS
6314|ELDORENDO
6315|ELDRED
6316|ELDRIDGE
6317|ELDRIDGE PARK
6318|ELEANOR
6319|ELECTRA
6320|ELECTRIC CITY
6321|ELECTRIC MILLS
6322|ELEPHANT BUTTE
6323|ELEVA
6324|ELEʻELE
6325|ELFERS
6326|ELFIN COVE
6327|ELFRIDA
6328|ELGIN
6329|ELI
6330|ELIASVILLE
6331|ELIDA
6332|ELIHU
6333|ELIM
6334|ELIMSPORT
6335|ELIZABETH
6336|ELIZABETH CITY
6337|ELIZABETHTON
6338|ELIZABETHTOWN
6339|ELIZABETHVILLE
6340|ELIZAVILLE
6341|ELK
6342|ELK CITY
6343|ELK CREEK
6344|ELK FALLS
6345|ELK GARDEN
6346|ELK GROVE
6347|ELK GROVE VILLAGE
6348|ELK HILL
6349|ELK HORN
6350|ELK MILLS
6351|ELK MOUND
6352|ELK MOUNTAIN
6353|ELK NECK
6354|ELK PARK
6355|ELK PLAIN
6356|ELK POINT
6357|ELK RAPIDS
6358|ELK RIDGE
6359|ELK RIVER
6360|ELK RUN HEIGHTS
6361|ELK SPRINGS
6362|ELK VALLEY
6363|ELKADER
6364|ELKATAWA
6365|ELKHART
6366|ELKHART LAKE
6367|ELKHORN
6368|ELKHORN CITY
6369|ELKIN
6370|ELKINS
6371|ELKINS PARK
6372|ELKLAND
6373|ELKMONT
6374|ELKO
6375|ELKO NEW MARKET
6376|ELKOL
6377|ELKPORT
6378|ELKRIDGE
6379|ELKTON
6380|ELKVIEW
6381|ELKVILLE
6382|ELLA
6383|ELLABELL
6384|ELLAMAR
6385|ELLAMORE
6386|ELLAVILLE
6387|ELLENBORO
6388|ELLENBURG DEPOT
6389|ELLENDALE
6390|ELLENSBURG
6391|ELLENTON
6392|ELLENVILLE
6393|ELLENWOOD
6394|ELLERBE
6395|ELLERSLIE
6396|ELLETTSVILLE
6397|ELLICOTT
6398|ELLICOTT CITY
6399|ELLICOTTVILLE
6400|ELLIJAY
6401|ELLINGER
6402|ELLINGTON
6403|ELLINWOOD
6404|ELLIOTT
6405|ELLIOTTS BLUFF
6406|ELLIS
6407|ELLIS GROVE
6408|ELLISBURG
6409|ELLISFORDE
6410|ELLISON BAY
6411|ELLISPORT
6412|ELLISTON
6413|ELLISVILLE
6414|ELLOREE
6415|ELLPORT
6416|ELLSINORE
6417|ELLSTON
6418|ELLSWORTH
6419|ELLWOOD CITY
6420|ELLZEY
6421|ELM CITY
6422|ELM CREEK
6423|ELM GROVE
6424|ELM MOTT
6425|ELM POINT
6426|ELM SPRINGS
6427|ELMA
6428|ELMA CENTER
6429|ELMDALE
6430|ELMENDORF
6431|ELMER
6432|ELMER CITY
6433|ELMHURST
6434|ELMIRA
6435|ELMIRA HEIGHTS
6436|ELMO
6437|ELMODEL
6438|ELMONT
6439|ELMORE
6440|ELMORE CITY
6441|ELMSFORD
6442|ELMWOOD
6443|ELMWOOD PARK
6444|ELMWOOD PLACE
6445|ELNORA
6446|ELON
6447|ELORA
6448|ELOY
6449|ELRAMA
6450|ELROD
6451|ELROSA
6452|ELROY
6453|ELSA
6454|ELSAH
6455|ELSBERRY
6456|ELSEY
6457|ELSIE
6458|ELSINORE
6459|ELSMERE
6460|ELSMORE
6461|ELTON
6462|ELTOPIA
6463|ELVASTON
6464|ELVERSON
6465|ELVERTA
6466|ELWELL
6467|ELWOOD
6468|ELWYN
6469|ELY
6470|ELYRIA
6471|ELYSBURG
6472|ELYSIAN
6473|EMAJAGUA
6474|EMAJAGUA COMUNIDAD
6475|EMBARRASS
6476|EMBDEN
6477|EMBLEM
6478|EMBREEVILLE
6479|EMBUDO
6480|EMDEN
6481|EMELLE
6482|EMERADO
6483|EMERALD
6484|EMERALD BAY
6485|EMERALD BEACH
6486|EMERALD ISLE
6487|EMERALD LAKE HILLS
6488|EMERALD LAKES
6489|EMERSON
6490|EMERY
6491|EMERYVILLE
6492|EMHOUSE
6493|EMIDA
6494|EMIGRANT
6495|EMIGRANT GAP
6496|EMIGSVILLE
6497|EMILY
6498|EMINENCE
6499|EMINGTON
6500|EMISON
6501|EMLENTON
6502|EMLYN
6503|EMMA
6504|EMMALANE
6505|EMMAUS
6506|EMMET
6507|EMMETSBURG
6508|EMMETT
6509|EMMITSBURG
6510|EMMONAK
6511|EMMONS
6512|EMMORTON
6513|EMORY
6514|EMPIRE
6515|EMPIRE CITY
6516|EMPORIA
6517|EMPORIUM
6518|EMSWORTH
6519|ENAVILLE
6520|ENCAMPMENT
6521|ENCHANTED OAKS
6522|ENCINAL
6523|ENCINITAS
6524|ENCINO
6525|ENDEAVOR
6526|ENDEE
6527|ENDERLIN
6528|ENDERS
6529|ENDICOTT
6530|ENDWELL
6531|ENERGY
6532|ENETAI
6533|ENFIELD
6534|ENGADINE
6535|ENGELHARD
6536|ENGLAND
6537|ENGLE
6538|ENGLEVALE
6539|ENGLEWOOD
6540|ENGLEWOOD CLIFFS
6541|ENGLISH
6542|ENGLISH TURN
6543|ENGLISHTOWN
6544|ENHAUT
6545|ENID
6546|ENIGMA
6547|ENKA
6548|ENLOE
6549|ENLOW
6550|ENNING
6551|ENNIS
6552|ENOCH
6553|ENOCHS
6554|ENOCHVILLE
6555|ENOLA
6556|ENON
6557|ENON VALLEY
6558|ENOREE
6559|ENOS CORNER
6560|ENOSBURG FALLS
6561|ENSENADA
6562|ENSIGN
6563|ENSLEY
6564|ENSOR
6565|ENTERPRISE
6566|ENTIAT
6567|ENUMCLAW
6568|ENVILLE
6569|EOLA
6570|EOLIA
6571|EOLINE
6572|EPES
6573|EPHESUS
6574|EPHRAIM
6575|EPHRATA
6576|EPLEYS
6577|EPPING
6578|EPPS
6579|EPSIE
6580|EPWORTH
6581|EPWORTH HEIGHTS
6582|EQUALITY
6583|ERA
6584|ERATH
6585|ERBACON
6586|ERCILDOUN
6587|ERDA
6588|ERHARD
6589|ERICK
6590|ERICSBURG
6591|ERICSON
6592|ERIDU
6593|ERIE
6594|ERIN
6595|ERIN SPRINGS
6596|ERLANDS POINT
6597|ERLANGER
6598|ERMA
6599|ERNEST
6600|ERNSTVILLE
6601|ERNUL
6602|EROS
6603|EROSE
6604|ERSKINE
6605|ERWIN
6606|ERWINVILLE
6607|ESBON
6608|ESCABOSA
6609|ESCALANTE
6610|ESCALON
6611|ESCANABA
6612|ESCATAWPA
6613|ESCHBACH
6614|ESCOBARES
6615|ESCOBAS
6616|ESCONDIDA
6617|ESCONDIDO
6618|ESKA
6619|ESKO
6620|ESKOTA
6621|ESKRIDGE
6622|ESMOND
6623|ESMONT
6624|ESOFEA
6625|ESOM HILL
6626|ESPANOLA
6627|ESPARTO
6628|ESPAÑOLA
6629|ESPERANCE
6630|ESPERANZA
6631|ESPERANZA COMUNIDAD
6632|ESPINO
6633|ESPINO COMUNIDAD
6634|ESPY
6635|ESSEX
6636|ESSEX FELLS
6637|ESSEX JUNCTION
6638|ESSEXVILLE
6639|ESSINGTON
6640|ESTACADA
6641|ESTANCIA
6642|ESTELL MANOR
6643|ESTELLE
6644|ESTELLINE
6645|ESTER
6646|ESTERBROOK
6647|ESTERO
6648|ESTES
6649|ESTES PARK
6650|ESTHERVILLE
6651|ESTHERWOOD
6652|ESTILL
6653|ESTILL SPRINGS
6654|ESTO
6655|ESTRAL BEACH
6656|ESTRELLA
6657|ETHAN
6658|ETHEL
6659|ETHELSVILLE
6660|ETHETE
6661|ETHRIDGE
6662|ETNA
6663|ETNA GREEN
6664|ETON
6665|ETOWAH
6666|ETRA
6667|ETTA
6668|ETTER
6669|ETTRICK
6670|EUBANK
6671|EUCALYPTUS HILLS
6672|EUCHA
6673|EUCHEEANNA
6674|EUCLID
6675|EUDORA
6676|EUFAULA
6677|EUGENE
6678|EUHARLEE
6679|EULATON
6680|EULESS
6681|EULONIA
6682|EUNICE
6683|EUNOLA
6684|EUPORA
6685|EUREKA
6686|EUREKA MILL
6687|EUREKA ROADHOUSE
6688|EUREKA SPRINGS
6689|EUREN
6690|EUSTACE
6691|EUSTIS
6692|EUTAW
6693|EUTAWVILLE
6694|EVA
6695|EVADALE
6696|EVAN
6697|EVANGELINE
6698|EVANS
6699|EVANS CITY
6700|EVANS MILLS
6701|EVANSBURG
6702|EVANSDALE
6703|EVANSTON
6704|EVANSVILLE
6705|EVANT
6706|EVARO
6707|EVART
6708|EVARTS
6709|EVELETH
6710|EVELYN
6711|EVENDALE
6712|EVENING SHADE
6713|EVENSVILLE
6714|EVEREST
6715|EVERETT
6716|EVERETTS
6717|EVERGLADES CITY
6718|EVERGREEN
6719|EVERGREEN COLONIA
6720|EVERGREEN PARK
6721|EVERLY
6722|EVERMAN
6723|EVERSON
6724|EVERTON
6725|EVESBORO
6726|EVINGTON
6727|EWA BEACH
6728|EWA GENTRY
6729|EWA VILLAGES
6730|EWAN
6731|EWANSVILLE
6732|EWART
6733|EWELL
6734|EWEN
6735|EWING
6736|EXCEL
6737|EXCELLO
6738|EXCELSIOR
6739|EXCELSIOR ESTATES
6740|EXCELSIOR SPRINGS
6741|EXCURSION INLET
6742|EXELAND
6743|EXELL
6744|EXETER
6745|EXETER CORNERS
6746|EXIRA
6747|EXLINE
6748|EXMORE
6749|EXPERIMENT
6750|EXPORT
6751|EXTON
6752|EXUM
6753|EYERS GROVE
6754|EYOTA
6755|EZEL
6756|EZZELL
6757|FABENS
6758|FABIUS
6759|FACEVILLE
6760|FACKLER
6761|FACTORYVILLE
6762|FAGUS
6763|FAIR BLUFF
6764|FAIR GARDEN
6765|FAIR GROVE
6766|FAIR HAVEN
6767|FAIR HILL
6768|FAIR LAWN
6769|FAIR OAKS
6770|FAIR OAKS RANCH
6771|FAIR PLAIN
6772|FAIR PLAY
6773|FAIRACRES
6774|FAIRBANK
6775|FAIRBANKS
6776|FAIRBORN
6777|FAIRBURN
6778|FAIRBURY
6779|FAIRCHANCE
6780|FAIRCHILD
6781|FAIRCHILDS
6782|FAIRDALE
6783|FAIRDEALING
6784|FAIRFAX
6785|FAIRFAX STATION
6786|FAIRFIELD
6787|FAIRFIELD BAY
6788|FAIRFIELD BEACH
6789|FAIRFIELD GLADE
6790|FAIRFIELD HARBOUR
6791|FAIRFORD
6792|FAIRFOREST
6793|FAIRGROVE
6794|FAIRHAVEN
6795|FAIRHOPE
6796|FAIRLAND
6797|FAIRLAWN
6798|FAIRLEA
6799|FAIRLEE
6800|FAIRLESS HILLS
6801|FAIRMEAD
6802|FAIRMONT
6803|FAIRMONT CITY
6804|FAIRMOUNT
6805|FAIRMOUNT HEIGHTS
6806|FAIROAKS
6807|FAIRPLAINS
6808|FAIRPLAY
6809|FAIRPOINT
6810|FAIRPORT
6811|FAIRPORT HARBOR
6812|FAIRTON
6813|FAIRVALLEY
6814|FAIRVIEW
6815|FAIRVIEW BEACH
6816|FAIRVIEW HEIGHTS
6817|FAIRVIEW PARK
6818|FAIRVIEW SHORES
6819|FAIRVILLE
6820|FAIRWATER
6821|FAIRWAY
6822|FAIRWOOD
6823|FAISON
6824|FAITH
6825|FAJARDO
6826|FAJARDO ZONA URBANA
6827|FALCON
6828|FALCON HEIGHTS
6829|FALCON LAKE ESTATES
6830|FALCON MESA
6831|FALCON VILLAGE
6832|FALCONER
6833|FALFURRIAS
6834|FALKIRK
6835|FALKLAND
6836|FALKNER
6837|FALKVILLE
6838|FALL BRANCH
6839|FALL CITY
6840|FALL CREEK
6841|FALL RIVER
6842|FALL RIVER MILLS
6843|FALLBROOK
6844|FALLING SPRING
6845|FALLING WATER
6846|FALLING WATERS
6847|FALLIS
6848|FALLON
6849|FALLS CHURCH
6850|FALLS CITY
6851|FALLS CREEK
6852|FALLS VIEW
6853|FALLS VILLAGE
6854|FALLSBURG
6855|FALLSINGTON
6856|FALLSTON
6857|FALMAN
6858|FALMOUTH
6859|FALMOUTH FORESIDE
6860|FALSE PASS
6861|FALUN
6862|FANCY FARM
6863|FANCY GAP
6864|FANDON
6865|FANNETT
6866|FANNETTSBURG
6867|FANNIN
6868|FANNING
6869|FANNING SPRINGS
6870|FANSHAWE
6871|FANWOOD
6872|FAR HILLS
6873|FAR ROCKAWAY
6874|FARBER
6875|FARGO
6876|FARIBAULT
6877|FARINA
6878|FARLEY
6879|FARLIN
6880|FARLINGTON
6881|FARMER
6882|FARMER CITY
6883|FARMERS
6884|FARMERS BRANCH
6885|FARMERSBURG
6886|FARMERSVILLE
6887|FARMERVILLE
6888|FARMINGDALE
6889|FARMINGTON
6890|FARMINGTON HILLS
6891|FARMINGVILLE
6892|FARMLAND
6893|FARMVILLE
6894|FARNAM
6895|FARNER
6896|FARNHAM
6897|FARNHAMVILLE
6898|FARNSWORTH
6899|FARR WEST
6900|FARRAGUT
6901|FARRANDSVILLE
6902|FARRAR
6903|FARRELL
6904|FARRISTOWN
6905|FARRSVILLE
6906|FARSON
6907|FARTHING
6908|FARWELL
6909|FASHING
6910|FATE
6911|FAUCETT
6912|FAULKNER
6913|FAULKTON
6914|FAUNSDALE
6915|FAUST
6916|FAVORETTA
6917|FAWN GROVE
6918|FAWN LAKE FOREST
6919|FAXON
6920|FAY
6921|FAYETTE
6922|FAYETTE CITY
6923|FAYETTEVILLE
6924|FAYSVILLE
6925|FAYVILLE
6926|FEARISVILLE
6927|FEARRINGTON VILLAGE
6928|FEASTERVILLE
6929|FEATHER SOUND
6930|FEATHERVILLE
6931|FEDERAL
6932|FEDERAL DAM
6933|FEDERAL HEIGHTS
6934|FEDERAL HILL
6935|FEDERAL WAY
6936|FEDERALSBURG
6937|FEDORA
6938|FELCH
6939|FELICITY
6940|FELIDA
6941|FELIXVILLE
6942|FELLOWS
6943|FELLOWSVILLE
6944|FELLSBURG
6945|FELLSMERE
6946|FELSENTHAL
6947|FELTON
6948|FELTS MILLS
6949|FENCE LAKE
6950|FENDERS
6951|FENN
6952|FENNER
6953|FENNIMORE
6954|FENNVILLE
6955|FENTON
6956|FENTRESS
6957|FENWICK
6958|FENWICK ISLAND
6959|FENWOOD
6960|FERDINAND
6961|FERGUS
6962|FERGUS FALLS
6963|FERGUSON
6964|FERN ACRES
6965|FERN CREST VILLAGE
6966|FERN FOREST
6967|FERN PARK
6968|FERN PRAIRIE
6969|FERNALD
6970|FERNAN LAKE VILLAGE
6971|FERNANDINA BEACH
6972|FERNANDO
6973|FERNBROOK
6974|FERNDALE
6975|FERNEY
6976|FERNLEY
6977|FERNVILLE
6978|FERNWAY
6979|FERNWOOD
6980|FERRELLSBURG
6981|FERRELVIEW
6982|FERRIDAY
6983|FERRIS
6984|FERRON
6985|FERRUM
6986|FERRY
6987|FERRY PASS
6988|FERRYSBURG
6989|FERRYVILLE
6990|FERTILE
6991|FESSENDEN
6992|FESTUS
6993|FETTERS HOT SPRINGS
6994|FIDDLETOWN
6995|FIDELIS
6996|FIDELITY
6997|FIELDALE
6998|FIELDBROOK
6999|FIELDING
7000|FIELDON
7001|FIELDS LANDING
7002|FIELDSBORO
7003|FIERRO
7004|FIFE
7005|FIFE HEIGHTS
7006|FIFE LAKE
7007|FIFTH STREET
7008|FIFTH WARD
7009|FIFTY LAKES
7010|FIFTYSIX
7011|FILER
7012|FILER CITY
7013|FILLEY
7014|FILLMORE
7015|FINCASTLE
7016|FINCHFORD
7017|FINCHVILLE
7018|FINDERNE
7019|FINDLAY
7020|FINESVILLE
7021|FINGAL
7022|FINGERVILLE
7023|FINLAND
7024|FINLAY
7025|FINLAYSON
7026|FINLEY
7027|FINLEY POINT
7028|FINLEYSON
7029|FINLEYVILLE
7030|FINNEY
7031|FINNEYTOWN
7032|FINZEL
7033|FIRCREST
7034|FIRE ISLAND
7035|FIREBAUGH
7036|FIREBRICK
7037|FIRECO
7038|FIRESTEEL
7039|FIRESTONE
7040|FIRST COLONY
7041|FIRST MESA
7042|FIRTH
7043|FIRTHCLIFFE
7044|FISCHER
7045|FISH CAMP
7046|FISH CREEK
7047|FISH HAVEN
7048|FISH HAWK
7049|FISH LAKE
7050|FISHER
7051|FISHER ISLAND
7052|FISHERS
7053|FISHERS ISLAND
7054|FISHERS LANDING
7055|FISHERSVILLE
7056|FISHING CREEK
7057|FISHKILL
7058|FISHTAIL
7059|FISK
7060|FISKDALE
7061|FITCHBURG
7062|FITCHVILLE
7063|FITHIAN
7064|FITLER
7065|FITTSTOWN
7066|FITZGERALD
7067|FITZHUGH
7068|FITZPATRICK
7069|FIVE CORNERS
7070|FIVE FORKS
7071|FIVE MILE FORK
7072|FIVE POINTS
7073|FIVEPOINTVILLE
7074|FLAG
7075|FLAGLER
7076|FLAGLER BEACH
7077|FLAGSTAFF
7078|FLAGTOWN
7079|FLAHERTY
7080|FLAMINGO
7081|FLANAGAN
7082|FLANDERS
7083|FLANDREAU
7084|FLANIGAN
7085|FLASHER
7086|FLAT
7087|FLAT LICK
7088|FLAT ROCK
7089|FLAT WOODS
7090|FLATGAP
7091|FLATONIA
7092|FLATS
7093|FLATWILLOW
7094|FLATWOOD
7095|FLATWOODS
7096|FLAXTON
7097|FLAXVILLE
7098|FLEETWOOD
7099|FLEISCHMANNS
7100|FLEMING
7101|FLEMING ISLAND
7102|FLEMING-NEON
7103|FLEMINGSBURG
7104|FLEMINGTON
7105|FLENSBURG
7106|FLETCHER
7107|FLINN SPRINGS
7108|FLINT
7109|FLINT CITY
7110|FLINT CREEK
7111|FLINT HILL
7112|FLINTSTONE
7113|FLINTVILLE
7114|FLIPPEN
7115|FLIPPIN
7116|FLO
7117|FLOM
7118|FLOMATON
7119|FLOMOT
7120|FLOODWOOD
7121|FLORA
7122|FLORA VISTA
7123|FLORADALE
7124|FLORAHOME
7125|FLORAL
7126|FLORAL CITY
7127|FLORAL PARK
7128|FLORALA
7129|FLORAVILLE
7130|FLORDELL HILLS
7131|FLORENCE
7132|FLORENCE HILL
7133|FLORENCE JUNCTION
7134|FLORES
7135|FLORESVILLE
7136|FLOREY
7137|FLORHAM PARK
7138|FLORIDA
7139|FLORIDA CITY
7140|FLORIDA RIDGE
7141|FLORIDA ZONA URBANA
7142|FLORIDATOWN
7143|FLORIEN
7144|FLORIN
7145|FLORIS
7146|FLORISSANT
7147|FLORISTON
7148|FLOSSMOOR
7149|FLOURNOY
7150|FLOURTOWN
7151|FLOVILLA
7152|FLOWELL
7153|FLOWELLA
7154|FLOWER HILL
7155|FLOWER MOUND
7156|FLOWEREE
7157|FLOWERSVILLE
7158|FLOWERY BRANCH
7159|FLOWING SPRINGS
7160|FLOWING WELLS
7161|FLOWOOD
7162|FLOYD
7163|FLOYDADA
7164|FLOYDALE
7165|FLUKER
7166|FLUSHING
7167|FLUTE SPRINGS
7168|FLYING HILLS
7169|FLYNN
7170|FOARD CITY
7171|FOBES HILL
7172|FOGELSVILLE
7173|FOLCROFT
7174|FOLGER
7175|FOLKSTON
7176|FOLLANSBEE
7177|FOLLETT
7178|FOLLETTS
7179|FOLLY BEACH
7180|FOLSOM
7181|FOND DU LAC
7182|FONDA
7183|FONDE
7184|FONTANA
7185|FONTANA VILLAGE
7186|FONTANELLE
7187|FONTANET
7188|FONTENELLE
7189|FOOSLAND
7190|FOOT OF TEN
7191|FOOTHILL FARMS
7192|FOOTS CREEK
7193|FOOTVILLE
7194|FORADA
7195|FORAKER
7196|FORBES
7197|FORBES ROAD
7198|FORBESTOWN
7199|FORBING
7200|FORBUS
7201|FORD
7202|FORD CITY
7203|FORD CLIFF
7204|FORD HEIGHTS
7205|FORDLAND
7206|FORDOCHE
7207|FORDS
7208|FORDS PRAIRIE
7209|FORDSVILLE
7210|FORDVILLE
7211|FORDYCE
7212|FOREMAN
7213|FOREST
7214|FOREST ACRES
7215|FOREST CENTER
7216|FOREST CITY
7217|FOREST GLADE
7218|FOREST GLEN
7219|FOREST GROVE
7220|FOREST HEIGHTS
7221|FOREST HILL
7222|FOREST HILL VILLAGE
7223|FOREST HILLS
7224|FOREST HOME
7225|FOREST JUNCTION
7226|FOREST KNOLLS
7227|FOREST LAKE
7228|FOREST LAKES ESTATES
7229|FOREST MEADOWS
7230|FOREST OAKS
7231|FOREST PARK
7232|FOREST RANCH
7233|FOREST RIVER
7234|FOREST VIEW
7235|FORESTBROOK
7236|FORESTBURG
7237|FORESTDALE
7238|FORESTHILL
7239|FORESTON
7240|FORESTVILLE
7241|FORGAN
7242|FORGE VILLAGE
7243|FORISTELL
7244|FORK
7245|FORK MOUNTAIN
7246|FORK UNION
7247|FORKED ISLAND
7248|FORKED RIVER
7249|FORKLAND
7250|FORKS
7251|FORKSVILLE
7252|FORKVILLE
7253|FORMAN
7254|FORMOSA
7255|FORMOSO
7256|FORNEY
7257|FORREST
7258|FORREST CITY
7259|FORRESTON
7260|FORSAN
7261|FORSYTH
7262|FORT ADAMS
7263|FORT ANN
7264|FORT APACHE
7265|FORT ASHBY
7266|FORT ATKINSON
7267|FORT BARNWELL
7268|FORT BASINGER
7269|FORT BELKNAP AGENCY
7270|FORT BELLEFONTAINE
7271|FORT BENTON
7272|FORT BIDWELL
7273|FORT BLACKMORE
7274|FORT BRAGG
7275|FORT BRANCH
7276|FORT BRIDGER
7277|FORT CALHOUN
7278|FORT CARSON
7279|FORT CHADBOURNE
7280|FORT CHISWELL
7281|FORT CLARK
7282|FORT CLARK SPRINGS
7283|FORT COBB
7284|FORT COFFEE
7285|FORT COLLINS
7286|FORT DAVIS
7287|FORT DEFIANCE
7288|FORT DEPOSIT
7289|FORT DICK
7290|FORT DIX
7291|FORT DODGE
7292|FORT DOUGLAS
7293|FORT DRUM
7294|FORT DUCHESNE
7295|FORT EDWARD
7296|FORT FAIRFIELD
7297|FORT GAINES
7298|FORT GARLAND
7299|FORT GATES
7300|FORT GAY
7301|FORT GIBSON
7302|FORT GREEN
7303|FORT GREEN SPRINGS
7304|FORT GRIFFIN
7305|FORT HALL
7306|FORT HANCOCK
7307|FORT HILL CENSUS DESIGNATED PLACE
7308|FORT HUNT
7309|FORT INDIANTOWN GAP
7310|FORT IRWIN
7311|FORT JENNINGS
7312|FORT JESUP
7313|FORT JOHNSON
7314|FORT JONES
7315|FORT KENT
7316|FORT KLAMATH
7317|FORT LARAMIE
7318|FORT LAUDERDALE
7319|FORT LAWN
7320|FORT LEE
7321|FORT LORAMIE
7322|FORT LOUDON
7323|FORT LUPTON
7324|FORT MADISON
7325|FORT MEADE
7326|FORT MILL
7327|FORT MITCHELL
7328|FORT MONTGOMERY
7329|FORT MORGAN
7330|FORT MOTTE
7331|FORT MYERS
7332|FORT MYERS BEACH
7333|FORT MYERS SHORES
7334|FORT OGDEN
7335|FORT OGLETHORPE
7336|FORT PAYNE
7337|FORT PECK
7338|FORT PIERCE
7339|FORT PIERRE
7340|FORT PLAIN
7341|FORT RANSOM
7342|FORT RECOVERY
7343|FORT RIPLEY
7344|FORT SALONGA
7345|FORT SCOTT
7346|FORT SENECA
7347|FORT SHAW
7348|FORT SHAWNEE
7349|FORT SMITH
7350|FORT STANTON
7351|FORT STOCKTON
7352|FORT SUMNER
7353|FORT SUPPLY
7354|FORT THOMAS
7355|FORT THOMPSON
7356|FORT TOTTEN
7357|FORT TOWSON
7358|FORT VALLEY
7359|FORT WALTON BEACH
7360|FORT WASHAKIE
7361|FORT WASHINGTON
7362|FORT WAYNE
7363|FORT WHITE
7364|FORT WINGATE
7365|FORT WORTH
7366|FORT WRIGHT
7367|FORT YATES
7368|FORT YUKON
7369|FORTESCUE
7370|FORTINE
7371|FORTSON
7372|FORTSONIA
7373|FORTUNA
7374|FORTUNA FOOTHILLS
7375|FORTVILLE
7376|FORTY FORT
7377|FOSCOE
7378|FOSS
7379|FOSSIL
7380|FOSSTON
7381|FOSSUM
7382|FOSTER
7383|FOSTER BROOK
7384|FOSTER CENTER
7385|FOSTER CITY
7386|FOSTERS
7387|FOSTORIA
7388|FOUKE
7389|FOUNDRYVILLE
7390|FOUNTAIN
7391|FOUNTAIN CITY
7392|FOUNTAIN GREEN
7393|FOUNTAIN HILL
7394|FOUNTAIN HILLS
7395|FOUNTAIN INN
7396|FOUNTAIN LAKE
7397|FOUNTAIN N' LAKES
7398|FOUNTAIN RUN
7399|FOUNTAIN SPRINGS
7400|FOUNTAIN VALLEY
7401|FOUNTAINEBLEAU
7402|FOUR BEARS VILLAGE
7403|FOUR BUTTES
7404|FOUR CORNERS
7405|FOUR LAKES
7406|FOUR OAKS
7407|FOUR POINTS COLONIA
7408|FOUR SEASONS
7409|FOUR STATES
7410|FOUR TOWN
7411|FOUR WAY
7412|FOURCHE
7413|FOWLER
7414|FOWLERTON
7415|FOWLERVILLE
7416|FOWLKES
7417|FOWLSTOWN
7418|FOX
7419|FOX CHAPEL
7420|FOX CHASE
7421|FOX CREEK
7422|FOX CROSSING
7423|FOX ISLAND
7424|FOX LAKE
7425|FOX LAKE HILLS
7426|FOX POINT
7427|FOX RIVER
7428|FOX RIVER GROVE
7429|FOX RUN
7430|FOXBORO
7431|FOXBOROUGH
7432|FOXBURG
7433|FOXFIELD
7434|FOXFIRE
7435|FOXHOLM
7436|FOXHOME
7437|FOXPARK
7438|FOXWORTH
7439|FOYIL
7440|FRACKVILLE
7441|FRAGARIA
7442|FRAMINGHAM
7443|FRANCES
7444|FRANCESVILLE
7445|FRANCIS
7446|FRANCIS CREEK
7447|FRANCIS MILLS
7448|FRANCISCO
7449|FRANCISVILLE
7450|FRANCITAS
7451|FRANCONIA
7452|FRANK
7453|FRANKCLAY
7454|FRANKENMUTH
7455|FRANKEWING
7456|FRANKFORD
7457|FRANKFORT
7458|FRANKFORT SPRINGS
7459|FRANKFORT SQUARE
7460|FRANKLIN
7461|FRANKLIN FURNACE
7462|FRANKLIN GROVE
7463|FRANKLIN LAKES
7464|FRANKLIN PARK
7465|FRANKLIN SPRINGS
7466|FRANKLIN SQUARE
7467|FRANKLINTON
7468|FRANKLINTOWN
7469|FRANKLINVILLE
7470|FRANKSTON
7471|FRANKSVILLE
7472|FRANKTON
7473|FRANKTOWN
7474|FRANKVILLE
7475|FRANNIE
7476|FRANQUEZ
7477|FRASER
7478|FRAZEE
7479|FRAZER
7480|FRAZEYSBURG
7481|FRAZIER PARK
7482|FRED
7483|FREDA
7484|FREDERIC
7485|FREDERICA
7486|FREDERICK
7487|FREDERICKSBURG
7488|FREDERICKSON
7489|FREDERICKTOWN
7490|FREDERIKA
7491|FREDERIKSTED
7492|FREDONIA
7493|FREE HOME
7494|FREE SOIL
7495|FREE UNION
7496|FREEBORN
7497|FREEBURG
7498|FREEBURN
7499|FREEDHEM
7500|FREEDOM
7501|FREEDOM ACRES
7502|FREEDOM PLAINS
7503|FREEDOM STATION
7504|FREEHOLD
7505|FREELAND
7506|FREELANDVILLE
7507|FREEMAN
7508|FREEMAN SPUR
7509|FREEMANSBURG
7510|FREEMONT
7511|FREENY
7512|FREEPORT
7513|FREER
7514|FREETOWN
7515|FREEVILLE
7516|FREEWOOD ACRES
7517|FREISTATT
7518|FREMONT
7519|FREMONT HILLS
7520|FRENCH
7521|FRENCH CAMP
7522|FRENCH GULCH
7523|FRENCH ISLAND
7524|FRENCH LICK
7525|FRENCH RIVER
7526|FRENCH SETTLEMENT
7527|FRENCH VILLAGE
7528|FRENCHBURG
7529|FRENCHGLEN
7530|FRENCHMAN
7531|FRENCHTON
7532|FRENCHTOWN
7533|FRENIER
7534|FRESNO
7535|FREWSBURG
7536|FRIANT
7537|FRIARS POINT
7538|FRIDAY
7539|FRIDAY HARBOR
7540|FRIDLEY
7541|FRIEDENS
7542|FRIEDENSBURG
7543|FRIEND
7544|FRIENDLY
7545|FRIENDSHIP
7546|FRIENDSVILLE
7547|FRIENDSWOOD
7548|FRIERSON
7549|FRIES
7550|FRIES MILL
7551|FRIESLAND
7552|FRINK
7553|FRIONA
7554|FRISCO
7555|FRISCO CITY
7556|FRISTOE
7557|FRITCH
7558|FRITZ
7559|FRITZ CREEK
7560|FRIZZLEBURG
7561|FROGMORE
7562|FROHNA
7563|FROID
7564|FROMBERG
7565|FRONT ROYAL
7566|FRONTENAC
7567|FRONTIER
7568|FRONTON
7569|FROST
7570|FROSTBURG
7571|FROSTPROOF
7572|FRUIT COVE
7573|FRUIT HEIGHTS
7574|FRUIT HILL
7575|FRUITA
7576|FRUITDALE
7577|FRUITHURST
7578|FRUITLAND
7579|FRUITLAND PARK
7580|FRUITPORT
7581|FRUITVALE
7582|FRUITVILLE
7583|FRYBURG
7584|FRYEBURG
7585|FRYSTOWN
7586|FRYTOWN
7587|FRÁNQUEZ COMUNIDAD
7588|FT MITCHELL
7589|FUIG
7590|FUIG COMUNIDAD
7591|FULDA
7592|FULFORD
7593|FULKS RUN
7594|FULLER ACRES
7595|FULLER HEIGHTS
7596|FULLERTON
7597|FULLERVILLE
7598|FULSHEAR
7599|FULTON
7600|FULTONDALE
7601|FULTONHAM
7602|FULTONVILLE
7603|FULTS
7604|FUNK
7605|FUNKLEY
7606|FUNKSTOWN
7607|FUNNY RIVER
7608|FUNSTON
7609|FUNTER
7610|FUQUAY-VARINA
7611|FURLEY
7612|FURMAN
7613|FURNACE
7614|FURNACE BRANCH
7615|FURNACE CREEK
7616|FURNACE WOODS
7617|FUSSELS CORNER
7618|FYFFE
7619|G. L. GARCIA
7620|G. L. GARCÍA COMUNIDAD
7621|GAASTRA
7622|GABBETTVILLE
7623|GABBS
7624|GACKLE
7625|GADSDEN
7626|GAFFNEY
7627|GAGE
7628|GAGEBY
7629|GAGEN
7630|GAGES LAKE
7631|GAGETOWN
7632|GAHANNA
7633|GAIL
7634|GAINES
7635|GAINESBORO
7636|GAINESVILLE
7637|GAITHERSBURG
7638|GAKONA
7639|GALATA
7640|GALATEO
7641|GALATEO COMUNIDAD
7642|GALATIA
7643|GALAX
7644|GALBRAITH
7645|GALENA
7646|GALENA PARK
7647|GALES FERRY
7648|GALESBURG
7649|GALESTOWN
7650|GALESVILLE
7651|GALETON
7652|GALEVILLE
7653|GALIEN
7654|GALION
7655|GALISTEO
7656|GALIVANTS FERRY
7657|GALLANT
7658|GALLATIN
7659|GALLATIN GATEWAY
7660|GALLAWAY
7661|GALLIANO
7662|GALLINA
7663|GALLINAS
7664|GALLION
7665|GALLIPOLIS
7666|GALLIPOLIS FERRY
7667|GALLITZIN
7668|GALLMAN
7669|GALLOWAY
7670|GALLUP
7671|GALT
7672|GALVA
7673|GALVESTON
7674|GALWAY
7675|GAMALIEL
7676|GAMBELL
7677|GAMBIER
7678|GAMBRILLS
7679|GAME CREEK
7680|GAMERCO
7681|GAMEWELL
7682|GANADO
7683|GANDEEVILLE
7684|GANDY
7685|GANG MILLS
7686|GANNETT
7687|GANO
7688|GANS
7689|GANSEVOORT
7690|GANTT
7691|GAP MILLS
7692|GAPLAND
7693|GARBER
7694|GARBERVILLE
7695|GARCENO
7696|GARCIA
7697|GARCIASVILLE
7698|GARD
7699|GARDAR
7700|GARDEN
7701|GARDEN ACRES
7702|GARDEN CITY
7703|GARDEN CITY PARK
7704|GARDEN CITY SOUTH
7705|GARDEN FARMS
7706|GARDEN GROVE
7707|GARDEN LAKES
7708|GARDEN PLAIN
7709|GARDEN PRAIRIE
7710|GARDEN RIDGE
7711|GARDEN VALLEY
7712|GARDEN VIEW
7713|GARDENA
7714|GARDENDALE
7715|GARDERE
7716|GARDI
7717|GARDINER
7718|GARDNER
7719|GARDNERS
7720|GARDNERTOWN
7721|GARDNERVILLE
7722|GARDNERVILLE RANCHOS
7723|GAREY
7724|GARFIELD
7725|GARFIELD HEIGHTS
7726|GARGATHA
7727|GARIBALDI
7728|GARLAND
7729|GARLIN
7730|GARLOCK
7731|GARNAVILLO
7732|GARNEILL
7733|GARNER
7734|GARNET
7735|GARNETT
7736|GARO
7737|GARRETSON
7738|GARRETT
7739|GARRETT PARK
7740|GARRETTS MILL
7741|GARRETTSVILLE
7742|GARRISON
7743|GARROCHALES
7744|GARROCHALES COMUNIDAD
7745|GARRYOWEN
7746|GARVIN
7747|GARWIN
7748|GARWOOD
7749|GARY
7750|GARYSBURG
7751|GARYVILLE
7752|GAS CITY
7753|GASBURG
7754|GASCON
7755|GASCONADE
7756|GASCOYNE
7757|GASKIN
7758|GASPER
7759|GASPORT
7760|GASQUE
7761|GASQUET
7762|GASSAWAY
7763|GASSOWAY
7764|GASSVILLE
7765|GASTON
7766|GASTONIA
7767|GASTONVILLE
7768|GATE
7769|GATE CITY
7770|GATES
7771|GATES CENTER
7772|GATES MILLS
7773|GATESVILLE
7774|GATEWAY
7775|GATLIFF
7776|GATLINBURG
7777|GATTMAN
7778|GAULEY BRIDGE
7779|GAUSE
7780|GAUTIER
7781|GAVIOTA
7782|GAY
7783|GAYLE MILL
7784|GAYLESVILLE
7785|GAYLORD
7786|GAYLY
7787|GAYS
7788|GAYS MILLS
7789|GAYVILLE
7790|GAZA
7791|GAZELLE
7792|GEARHART
7793|GEARY
7794|GEDDES
7795|GEEVILLE
7796|GEFF
7797|GEIGER
7798|GEIGERTOWN
7799|GEISMAR
7800|GEISTOWN
7801|GEM
7802|GEM LAKE
7803|GEM VILLAGE
7804|GEMMELL
7805|GENE AUTRY
7806|GENESEE
7807|GENESEE DEPOT
7808|GENESEO
7809|GENEVA
7810|GENEVA-ON-THE-LAKE
7811|GENOA
7812|GENOA CITY
7813|GENOLA
7814|GENTRY
7815|GENTRYVILLE
7816|GEORGE
7817|GEORGE WEST
7818|GEORGES MILLS
7819|GEORGETOWN
7820|GEORGIANA
7821|GEORGIAVILLE
7822|GERALD
7823|GERALDINE
7824|GERBER
7825|GERING
7826|GERLACH
7827|GERMAN VALLEY
7828|GERMANIA
7829|GERMANO
7830|GERMANTON
7831|GERMANTOWN
7832|GERMANTOWN HILLS
7833|GERMFASK
7834|GERONIMO
7835|GERRARD
7836|GERSTER
7837|GERTON
7838|GERTY
7839|GERVAIS
7840|GESSIE
7841|GETTYSBURG
7842|GETZVILLE
7843|GEUDA SPRINGS
7844|GEYSER
7845|GEYSERVILLE
7846|GHEEN
7847|GHENT
7848|GHOLSON
7849|GIBBON
7850|GIBBONSVILLE
7851|GIBBS
7852|GIBBSBORO
7853|GIBBSTOWN
7854|GIBBSVILLE
7855|GIBRALTAR
7856|GIBSLAND
7857|GIBSON
7858|GIBSON CITY
7859|GIBSON FLATS
7860|GIBSON ISLAND
7861|GIBSONBURG
7862|GIBSONIA
7863|GIBSONTON
7864|GIBSONVILLE
7865|GIDDINGS
7866|GIDEON
7867|GIFFORD
7868|GIG HARBOR
7869|GILA
7870|GILA BEND
7871|GILA CROSSING
7872|GILARK
7873|GILBERT
7874|GILBERT CREEK
7875|GILBERTON
7876|GILBERTOWN
7877|GILBERTS
7878|GILBERTSVILLE
7879|GILBERTVILLE
7880|GILBOA
7881|GILBY
7882|GILCHRIST
7883|GILCREST
7884|GILDFORD
7885|GILEAD
7886|GILES
7887|GILFORD PARK
7888|GILL
7889|GILLESPIE
7890|GILLETT
7891|GILLETT GROVE
7892|GILLETTE
7893|GILLHAM
7894|GILLIAM
7895|GILLIATT
7896|GILLIS
7897|GILLS ROCK
7898|GILLSVILLE
7899|GILLULY
7900|GILMAN
7901|GILMAN CITY
7902|GILMANTON
7903|GILMER
7904|GILMORE
7905|GILMORE CITY
7906|GILPIN
7907|GILROY
7908|GILSON
7909|GILT EDGE
7910|GILTNER
7911|GINGER BLUE
7912|GIRARD
7913|GIRARDVILLE
7914|GIRDLETREE
7915|GIRDWOOD
7916|GIRTY
7917|GIRVIN
7918|GISELA
7919|GLACIER
7920|GLAD VALLEY
7921|GLADBROOK
7922|GLADDEN
7923|GLADE
7924|GLADE MILLS
7925|GLADE SPRING
7926|GLADEVIEW
7927|GLADEVILLE
7928|GLADEWATER
7929|GLADIOLA
7930|GLADSTONE
7931|GLADWIN
7932|GLADWYNE
7933|GLADY
7934|GLADYS
7935|GLAMIS
7936|GLANCY
7937|GLANDORF
7938|GLASCO
7939|GLASFORD
7940|GLASGOW
7941|GLASGOW VILLAGE
7942|GLASS
7943|GLASSBORO
7944|GLASSMANOR
7945|GLASSPORT
7946|GLASTONBURY CENTER
7947|GLAZIER
7948|GLEASON
7949|GLEASONDALE
7950|GLEED
7951|GLEESON
7952|GLEN
7953|GLEN ALLAN
7954|GLEN ALLEN
7955|GLEN ALPINE
7956|GLEN ARBOR
7957|GLEN ARM
7958|GLEN AUBREY
7959|GLEN AVON
7960|GLEN BURNIE
7961|GLEN CAMPBELL
7962|GLEN CARBON
7963|GLEN COVE
7964|GLEN DEAN
7965|GLEN ECHO
7966|GLEN ECHO PARK
7967|GLEN ELDER
7968|GLEN ELLEN
7969|GLEN ELLYN
7970|GLEN ESTE
7971|GLEN FERRIS
7972|GLEN FLORA
7973|GLEN FORK
7974|GLEN GARDNER
7975|GLEN HAVEN
7976|GLEN HEAD
7977|GLEN HOPE
7978|GLEN JEAN
7979|GLEN LYN
7980|GLEN LYON
7981|GLEN PARK
7982|GLEN RAVEN
7983|GLEN RIDDLE
7984|GLEN RIDGE
7985|GLEN ROCK
7986|GLEN ROGERS
7987|GLEN ROSE
7988|GLEN SAINT MARY
7989|GLEN ULLIN
7990|GLEN WHITE
7991|GLEN WILTON
7992|GLENAIRE
7993|GLENALLEN
7994|GLENARDEN
7995|GLENBAR
7996|GLENBEULAH
7997|GLENBROOK
7998|GLENBURN
7999|GLENCOE
8000|GLENCROSS
8001|GLENDALE
8002|GLENDALE HEIGHTS
8003|GLENDALE SPRINGS
8004|GLENDEVEY
8005|GLENDIVE
8006|GLENDO
8007|GLENDON
8008|GLENDORA
8009|GLENEAGLE
8010|GLENFIELD
8011|GLENFORD
8012|GLENHAM
8013|GLENLOCH
8014|GLENMONT
8015|GLENMOOR
8016|GLENMOORE
8017|GLENMORA
8018|GLENN
8019|GLENN DALE
8020|GLENN HEIGHTS
8021|GLENNALLEN
8022|GLENNIE
8023|GLENNS FERRY
8024|GLENNVILLE
8025|GLENOLDEN
8026|GLENOMA
8027|GLENPOOL
8028|GLENRIDGE
8029|GLENROCK
8030|GLENS
8031|GLENS FALLS
8032|GLENSHAW
8033|GLENSIDE
8034|GLENTANA
8035|GLENVAR
8036|GLENVAR HEIGHTS
8037|GLENVIEW
8038|GLENVIEW HILLS
8039|GLENVIEW MANOR
8040|GLENVIL
8041|GLENVILLE
8042|GLENWILLARD
8043|GLENWILLOW
8044|GLENWOOD
8045|GLENWOOD CITY
8046|GLENWOOD LANDING
8047|GLENWOOD SPRINGS
8048|GLIDDEN
8049|GLIDE
8050|GLOBE
8051|GLORIA GLENS PARK
8052|GLORIETA
8053|GLOSTER
8054|GLOUCESTER
8055|GLOUCESTER CITY
8056|GLOUCESTER COURTHOUSE
8057|GLOUCESTER POINT
8058|GLOUSTER
8059|GLOVER
8060|GLOVERSVILLE
8061|GLOVERVILLE
8062|GLUCK
8063|GLUEK
8064|GLYNDON
8065|GLYNN
8066|GNADENHUTTEN
8067|GOBER
8068|GOBLER
8069|GOBLES
8070|GODDARD
8071|GODFREY
8072|GODLEY
8073|GODWIN
8074|GODWINSVILLE
8075|GOEHNER
8076|GOESSEL
8077|GOFF
8078|GOFFS
8079|GOFFSTOWN
8080|GOLCONDA
8081|GOLD
8082|GOLD ACRES
8083|GOLD BAR
8084|GOLD BEACH
8085|GOLD CANYON
8086|GOLD HILL
8087|GOLD KEY LAKE
8088|GOLD POINT
8089|GOLD RIVER
8090|GOLDCREEK
8091|GOLDEN
8092|GOLDEN BEACH
8093|GOLDEN CITY
8094|GOLDEN EAGLE
8095|GOLDEN GATE
8096|GOLDEN GLADES
8097|GOLDEN GROVE
8098|GOLDEN HILLS
8099|GOLDEN MEADOW
8100|GOLDEN TRIANGLE
8101|GOLDEN VALLEY
8102|GOLDENDALE
8103|GOLDENROD
8104|GOLDENS BRIDGE
8105|GOLDFIELD
8106|GOLDMAN
8107|GOLDONNA
8108|GOLDSBORO
8109|GOLDSBY
8110|GOLDSMITH
8111|GOLDSTON
8112|GOLDTHWAITE
8113|GOLDVEIN
8114|GOLDVILLE
8115|GOLETA
8116|GOLF
8117|GOLF MANOR
8118|GOLF VIEW
8119|GOLIAD
8120|GOLINDA
8121|GOLOVIN
8122|GOLTRY
8123|GOLVA
8124|GOMEZ
8125|GONVICK
8126|GONZALES
8127|GONZALEZ
8128|GOOBER HILL
8129|GOOCHLAND
8130|GOOD HART
8131|GOOD HOPE
8132|GOOD THUNDER
8133|GOODE
8134|GOODELL
8135|GOODENOW
8136|GOODFIELD
8137|GOODHUE
8138|GOODING
8139|GOODINGS GROVE
8140|GOODLAND
8141|GOODLETT
8142|GOODLETTSVILLE
8143|GOODLOW PARK
8144|GOODMAN
8145|GOODNEWS BAY
8146|GOODNIGHT
8147|GOODNO
8148|GOODNOE HILLS
8149|GOODRICH
8150|GOODRIDGE
8151|GOODSPRINGS
8152|GOODVIEW
8153|GOODVILLE
8154|GOODWATER
8155|GOODWELL
8156|GOODWILL
8157|GOODWIN
8158|GOODWINE
8159|GOODYEAR
8160|GOODYEARS BAR
8161|GOOFY RIDGE
8162|GOOSE CREEK
8163|GOOSE LAKE
8164|GOOSE PRAIRIE
8165|GOOSPORT
8166|GORDO
8167|GORDON
8168|GORDON HEIGHTS
8169|GORDONSVILLE
8170|GORDONVILLE
8171|GORDY
8172|GORE
8173|GOREE
8174|GOREVILLE
8175|GORGAS
8176|GORHAM
8177|GORIN
8178|GORMAN
8179|GORST
8180|GORUM
8181|GOSHEN
8182|GOSHENVILLE
8183|GOSHUTE
8184|GOSNELL
8185|GOSPORT
8186|GOSS
8187|GOST CREEK
8188|GOTEBO
8189|GOTHA
8190|GOTHAM
8191|GOTHENBURG
8192|GOUDEAU
8193|GOUGH
8194|GOUGLERSVILLE
8195|GOULD
8196|GOULD CITY
8197|GOULDING
8198|GOULDS
8199|GOULDSBORO
8200|GOUVERNEUR
8201|GOVAN
8202|GOVE
8203|GOVERNMENT CAMP
8204|GOWAN
8205|GOWANDA
8206|GOWEN
8207|GOWER
8208|GOWRIE
8209|GRABALL
8210|GRABILL
8211|GRACE
8212|GRACE CITY
8213|GRACEMONT
8214|GRACETON
8215|GRACEVILLE
8216|GRACEWOOD
8217|GRACEY
8218|GRADY
8219|GRADYVILLE
8220|GRAEAGLE
8221|GRAETTINGER
8222|GRAF
8223|GRAFORD
8224|GRAFTON
8225|GRAHAM
8226|GRAHAMTOWN
8227|GRAIN VALLEY
8228|GRAINFIELD
8229|GRAINOLA
8230|GRAINTON
8231|GRAMA
8232|GRAMBLING
8233|GRAMERCY
8234|GRAMLING
8235|GRAMPIAN
8236|GRAN QUIVIRA
8237|GRANADA
8238|GRANBURY
8239|GRANBY
8240|GRAND BAY
8241|GRAND BEACH
8242|GRAND BLANC
8243|GRAND CANE
8244|GRAND CANYON
8245|GRAND CHAIN
8246|GRAND CHENIER
8247|GRAND COTEAU
8248|GRAND COULEE
8249|GRAND DETOUR
8250|GRAND ECORE
8251|GRAND FALLS
8252|GRAND FALLS PLAZA
8253|GRAND FORKS
8254|GRAND GLAISE
8255|GRAND GULF
8256|GRAND HAVEN
8257|GRAND ISLAND
8258|GRAND ISLE
8259|GRAND JUNCTION
8260|GRAND LAKE
8261|GRAND LAKE TOWNE
8262|GRAND LEDGE
8263|GRAND MARAIS
8264|GRAND MARSH
8265|GRAND MEADOW
8266|GRAND MESA
8267|GRAND MOUND
8268|GRAND PASS
8269|GRAND POINT
8270|GRAND PORTAGE
8271|GRAND PRAIRIE
8272|GRAND RAPIDS
8273|GRAND RIDGE
8274|GRAND RIVER
8275|GRAND RIVERS
8276|GRAND RONDE
8277|GRAND SALINE
8278|GRAND TERRACE
8279|GRAND TOWER
8280|GRAND VIEW
8281|GRAND VIEW ESTATES
8282|GRAND VIEW-ON-HUDSON
8283|GRANDE
8284|GRANDFALLS
8285|GRANDFATHER
8286|GRANDFIELD
8287|GRANDIN
8288|GRANDVIEW
8289|GRANDVIEW HEIGHTS
8290|GRANDVIEW PLAZA
8291|GRANDVILLE
8292|GRANDWOOD PARK
8293|GRANDY
8294|GRANDYLE VILLAGE
8295|GRANGER
8296|GRANGEVILLE
8297|GRANITE
8298|GRANITE BAY
8299|GRANITE CITY
8300|GRANITE FALLS
8301|GRANITE HILLS
8302|GRANITE QUARRY
8303|GRANITE SHOALS
8304|GRANITE SPRINGS
8305|GRANITEVILLE
8306|GRANJENO
8307|GRANNIS
8308|GRANO
8309|GRANT
8310|GRANT CITY
8311|GRANT PARK
8312|GRANT TOWN
8313|GRANT-VALKARIA
8314|GRANTFORK
8315|GRANTLEY
8316|GRANTON
8317|GRANTS
8318|GRANTS PASS
8319|GRANTSBORO
8320|GRANTSBURG
8321|GRANTSDALE
8322|GRANTSVILLE
8323|GRANTVILLE
8324|GRANTWOOD VILLAGE
8325|GRANVILLE
8326|GRAPE CREEK
8327|GRAPELAND
8328|GRAPEVIEW
8329|GRAPEVILLE
8330|GRAPEVINE
8331|GRASMERE
8332|GRASONVILLE
8333|GRASS CREEK
8334|GRASS LAKE
8335|GRASS RANGE
8336|GRASS VALLEY
8337|GRASSFLAT
8338|GRASSTON
8339|GRASSY
8340|GRASSY BUTTE
8341|GRASSY CREEK
8342|GRATERFORD
8343|GRATIOT
8344|GRATIS
8345|GRATON
8346|GRATTON
8347|GRATZ
8348|GRAVELLY
8349|GRAVES
8350|GRAVETTE
8351|GRAVOIS MILLS
8352|GRAWN
8353|GRAY COURT
8354|GRAY HAWK
8355|GRAY HORSE
8356|GRAY MOUNTAIN
8357|GRAY SUMMIT
8358|GRAYBURG
8359|GRAYLAND
8360|GRAYLING
8361|GRAYMOOR-DEVONDALE
8362|GRAYRIDGE
8363|GRAYS
8364|GRAYS BRANCH
8365|GRAYS HILL
8366|GRAYS PRAIRIE
8367|GRAYS RIVER
8368|GRAYSLAKE
8369|GRAYSON
8370|GRAYSON VALLEY
8371|GRAYSVILLE
8372|GRAYVILLE
8373|GRAZIERVILLE
8374|GREASEWOOD
8375|GREASY
8376|GREAT BARRINGTON
8377|GREAT BEND
8378|GREAT CACAPON
8379|GREAT FALLS
8380|GREAT MEADOWS
8381|GREAT NECK
8382|GREAT NECK ESTATES
8383|GREAT NECK GARDENS
8384|GREAT NECK PLAZA
8385|GREAT RIVER
8386|GREATWOOD
8387|GREECE
8388|GREELEY
8389|GREELEY HILL
8390|GREELEYVILLE
8391|GREEN ACRES
8392|GREEN BANK
8393|GREEN BAY
8394|GREEN BLUFF
8395|GREEN BRIER
8396|GREEN CAMP
8397|GREEN CASTLE
8398|GREEN CITY
8399|GREEN COVE SPRINGS
8400|GREEN FOREST
8401|GREEN GRASS
8402|GREEN GROVE
8403|GREEN HARBOR
8404|GREEN HILL
8405|GREEN HILLS
8406|GREEN ISLAND
8407|GREEN ISLE
8408|GREEN KNOLL
8409|GREEN LAKE
8410|GREEN LANE
8411|GREEN LEVEL
8412|GREEN MEADOWS
8413|GREEN MOUNTAIN
8414|GREEN MOUNTAIN FALLS
8415|GREEN OAKS
8416|GREEN PARK
8417|GREEN POND
8418|GREEN RIDGE
8419|GREEN RIVER
8420|GREEN ROCK
8421|GREEN SPRING
8422|GREEN SPRINGS
8423|GREEN TREE
8424|GREEN VALLEY
8425|GREEN VALLEY FARMS
8426|GREEN VALLEY LAKE
8427|GREEN VILLAGE
8428|GREENACRES
8429|GREENACRES CITY
8430|GREENBACK
8431|GREENBACKVILLE
8432|GREENBANK
8433|GREENBELT
8434|GREENBRAE
8435|GREENBRIAR
8436|GREENBRIER
8437|GREENBUSH
8438|GREENCASTLE
8439|GREENDALE
8440|GREENE
8441|GREENEVERS
8442|GREENEVILLE
8443|GREENFIELD
8444|GREENFIELD HILL
8445|GREENFIELDS
8446|GREENFORD
8447|GREENHILLS
8448|GREENHORN
8449|GREENLAND
8450|GREENLAWN
8451|GREENLEAF
8452|GREENLEAFTON
8453|GREENOCK
8454|GREENOUGH
8455|GREENPORT
8456|GREENS FARMS
8457|GREENS FORK
8458|GREENSBORO
8459|GREENSBORO BEND
8460|GREENSBURG
8461|GREENTOP
8462|GREENTOWN
8463|GREENTREE
8464|GREENUP
8465|GREENVALE
8466|GREENVIEW
8467|GREENVILLE
8468|GREENWALD
8469|GREENWATER
8470|GREENWAY
8471|GREENWICH
8472|GREENWICH HEIGHTS
8473|GREENWOOD
8474|GREENWOOD LAKE
8475|GREENWOOD VILLAGE
8476|GREER
8477|GREERS FERRY
8478|GREGORY
8479|GREIGSVILLE
8480|GREILICKVILLE
8481|GRENADA
8482|GRENOLA
8483|GRENORA
8484|GRENVILLE
8485|GRESHAM
8486|GRESHAM PARK
8487|GRESSITT
8488|GRETNA
8489|GREY EAGLE
8490|GREY FOREST
8491|GREYBULL
8492|GREYCLIFF
8493|GREYSTONE
8494|GRIDER
8495|GRIDLEY
8496|GRIER CITY
8497|GRIFFIN
8498|GRIFFINS MILLS
8499|GRIFFITH
8500|GRIFFITHSVILLE
8501|GRIFFITHVILLE
8502|GRIFTON
8503|GRIGGSTOWN
8504|GRIGGSVILLE
8505|GRIGSTON
8506|GRILL
8507|GRIMES
8508|GRIMESLAND
8509|GRIMSLEY
8510|GRIND STONE CITY
8511|GRINDSTONE
8512|GRINGO
8513|GRINNELL
8514|GRISDALE
8515|GRISWOLD
8516|GRISWOLDVILLE
8517|GRIT
8518|GRIZZLY
8519|GROESBECK
8520|GROSSE POINTE
8521|GROSSE POINTE FARMS
8522|GROSSE POINTE PARK
8523|GROSSE POINTE SHORES
8524|GROSSE POINTE WOODS
8525|GROSSE TETE
8526|GROSSMONT
8527|GROTON
8528|GROTON LONG POINT
8529|GROTTO
8530|GROTTOES
8531|GROUSE
8532|GROUSE CREEK
8533|GROVANIA
8534|GROVE
8535|GROVE CENTER
8536|GROVE CITY
8537|GROVE HILL
8538|GROVE LAKE
8539|GROVELAND
8540|GROVEPORT
8541|GROVER
8542|GROVER BEACH
8543|GROVER HILL
8544|GROVERTOWN
8545|GROVES
8546|GROVESPRING
8547|GROVETON
8548|GROVETOWN
8549|GROVEVILLE
8550|GROVONT
8551|GROWLER
8552|GRUBBS
8553|GRUENE
8554|GRUETLI-LAAGER
8555|GRUHLKEY
8556|GRUNDY
8557|GRUNDY CENTER
8558|GRUVER
8559|GRYGLA
8560|GU OIDAK
8561|GU-WIN
8562|GUADALUPE
8563|GUADALUPITA
8564|GUAGE
8565|GUALALA
8566|GUASTI
8567|GUAYABAL
8568|GUAYABAL COMUNIDAD
8569|GUAYAMA
8570|GUAYAMA ZONA URBANA
8571|GUAYANILLA
8572|GUAYANILLA ZONA URBANA
8573|GUAYNABO
8574|GUAYNABO ZONA URBANA
8575|GUERNEVILLE
8576|GUERNSEY
8577|GUERRA
8578|GUEYDAN
8579|GUFFEY
8580|GUIDE ROCK
8581|GUILFORD
8582|GUIN
8583|GUINDA
8584|GUINEA
8585|GUION
8586|GULF
8587|GULF BREEZE
8588|GULF GATE ESTATES
8589|GULF HAMMOCK
8590|GULF HILLS
8591|GULF PARK ESTATES
8592|GULF SHORES
8593|GULF STREAM
8594|GULFCREST
8595|GULFPORT
8596|GULKANA
8597|GULLETT
8598|GULLY
8599|GULNARE
8600|GUM BRANCH
8601|GUM SPRINGS
8602|GUMLOG
8603|GUN BARREL CITY
8604|GUN CLUB ESTATES
8605|GUNBARREL
8606|GUNDER
8607|GUNLOCK
8608|GUNN
8609|GUNN CITY
8610|GUNNISON
8611|GUNTER
8612|GUNTERSVILLE
8613|GUNTOWN
8614|GURABO
8615|GURABO ZONA URBANA
8616|GURDON
8617|GURLEY
8618|GURNEE
8619|GUSTAVUS
8620|GUSTINE
8621|GUSTON
8622|GUTHRIE
8623|GUTHRIE CENTER
8624|GUTHRIESVILLE
8625|GUTTENBERG
8626|GUY
8627|GUYMON
8628|GUYS
8629|GUYS MILLS
8630|GUYTON
8631|GUÁNICA
8632|GUÁNICA ZONA URBANA
8633|GWENFORD
8634|GWINN
8635|GWINNER
8636|GWYNEDD VALLEY
8637|GWYNN
8638|GWYNN OAK
8639|GYPSUM
8640|GYPSY
8641|H. RIVERA COLON
8642|H. RIVERA COLÓN COMUNIDAD
8643|HAASWOOD
8644|HABERSHAM
8645|HACHITA
8646|HACIENDA HEIGHTS
8647|HACIENDA SAN JOSÉ COMUNIDAD
8648|HACIENDA VILLAGE
8649|HACKAMORE
8650|HACKBERRY
8651|HACKENSACK
8652|HACKER VALLEY
8653|HACKETT
8654|HACKETTSTOWN
8655|HACKLEBURG
8656|HACKNEY
8657|HACKNEYVILLE
8658|HACODA
8659|HADAR
8660|HADDAM
8661|HADDOCK
8662|HADDON HEIGHTS
8663|HADDONFIELD
8664|HADLEY
8665|HAGAMAN
8666|HAGAN
8667|HAGARVILLE
8668|HAGEMAN
8669|HAGER CITY
8670|HAGERHILL
8671|HAGERMAN
8672|HAGERSTOWN
8673|HAGEWOOD
8674|HAGUE
8675|HAHIRA
8676|HAHNTOWN
8677|HAHNVILLE
8678|HAIG
8679|HAIGLER
8680|HAILE
8681|HAILESBORO
8682|HAILEY
8683|HAILEYVILLE
8684|HAINES
8685|HAINES CITY
8686|HAINESBURG
8687|HAINESPORT
8688|HAINESVILLE
8689|HAIVANA NAKYA
8690|HAIWEE
8691|HALAʻULA
8692|HALBUR
8693|HALCHITA
8694|HALDANE
8695|HALDEMAN
8696|HALE
8697|HALE CENTER
8698|HALEBURG
8699|HALEDON
8700|HALES CORNERS
8701|HALESITE
8702|HALETHORPE
8703|HALEY
8704|HALEYVILLE
8705|HALEʻIWA
8706|HALF DAY
8707|HALF MOON
8708|HALF MOON BAY
8709|HALFA
8710|HALFMOON LANDING
8711|HALFWAY
8712|HALFWAY HOUSE
8713|HALIBUT COVE
8714|HALIFAX
8715|HALL
8716|HALL SUMMIT
8717|HALLAM
8718|HALLANDALE BEACH
8719|HALLECK
8720|HALLETT
8721|HALLETTSVILLE
8722|HALLEY
8723|HALLIDAY
8724|HALLOCK
8725|HALLOWELL
8726|HALLS
8727|HALLS CROSSING
8728|HALLS CROSSROADS
8729|HALLS GAP
8730|HALLS SUMMIT
8731|HALLSBORO
8732|HALLSBURG
8733|HALLSTEAD
8734|HALLSVILLE
8735|HALLTOWN
8736|HALLWOOD
8737|HALMA
8738|HALSEY
8739|HALSTAD
8740|HALSTEAD
8741|HALTOM CITY
8742|HAM LAKE
8743|HAMBERG
8744|HAMBLETON
8745|HAMBURG
8746|HAMDEN
8747|HAMEL
8748|HAMER
8749|HAMERSVILLE
8750|HAMILL
8751|HAMILTON
8752|HAMILTON BRANCH
8753|HAMILTON CITY
8754|HAMILTON DOME
8755|HAMILTON SQUARE
8756|HAMILTONS FORT
8757|HAMLER
8758|HAMLET
8759|HAMLETSBURG
8760|HAMLIN
8761|HAMMERSLEY FORK
8762|HAMMETT
8763|HAMMON
8764|HAMMOND
8765|HAMMONDSPORT
8766|HAMMONDVILLE
8767|HAMMONTON
8768|HAMORTON
8769|HAMPDEN
8770|HAMPDEN HIGHLANDS
8771|HAMPDEN SYDNEY
8772|HAMPSHIRE
8773|HAMPSTEAD
8774|HAMPTON
8775|HAMPTON BAYS
8776|HAMPTON BEACH
8777|HAMPTON MANOR
8778|HAMPTON SPRINGS
8779|HAMTRAMCK
8780|HANAHAN
8781|HANALEI
8782|HANAMĀʻULU
8783|HANAPĒPĒ
8784|HANCEVILLE
8785|HANCOCK
8786|HANCOCKS BRIDGE
8787|HANDLEY
8788|HANDSHOE
8789|HANFORD
8790|HANGING LIMB
8791|HANGING ROCK
8792|HANKAMER
8793|HANKINSON
8794|HANKSVILLE
8795|HANLEY FALLS
8796|HANLEY HILLS
8797|HANLONTOWN
8798|HANNA
8799|HANNA CITY
8800|HANNAFORD
8801|HANNAH
8802|HANNAHS MILL
8803|HANNASTOWN
8804|HANNASVILLE
8805|HANNAWA FALLS
8806|HANNIBAL
8807|HANNOVER
8808|HANOVER
8809|HANOVER CENTER
8810|HANOVER PARK
8811|HANOVERTON
8812|HANSBORO
8813|HANSELL
8814|HANSEN
8815|HANSKA
8816|HANSON
8817|HANSTON
8818|HANSVILLE
8819|HAPEVILLE
8820|HAPPY
8821|HAPPY CAMP
8822|HAPPY JACK
8823|HAPPY VALLEY
8824|HAPPYS INN
8825|HARAHAN
8826|HARALSON
8827|HARBERT
8828|HARBINE
8829|HARBISON CANYON
8830|HARBOR
8831|HARBOR BEACH
8832|HARBOR BLUFFS
8833|HARBOR HILLS
8834|HARBOR ISLE
8835|HARBOR SPRINGS
8836|HARBOR VIEW
8837|HARBORTON
8838|HARBOUR HEIGHTS
8839|HARBOUR POINTE
8840|HARCOURT
8841|HARCUVAR
8842|HARDAWAY
8843|HARDEEVILLE
8844|HARDESTY
8845|HARDIN
8846|HARDING
8847|HARDING LAKE
8848|HARDINSBURG
8849|HARDTNER
8850|HARDWICK
8851|HARDY
8852|HARDYVILLE
8853|HARGILL
8854|HARGIS
8855|HARING
8856|HARKER HEIGHTS
8857|HARKERS ISLAND
8858|HARKEYVILLE
8859|HARLAN
8860|HARLEIGH
8861|HARLEM
8862|HARLEM HEIGHTS
8863|HARLEM SPRINGS
8864|HARLETON
8865|HARLEYSVILLE
8866|HARLEYVILLE
8867|HARLINGEN
8868|HARLOW
8869|HARLOWTON
8870|HARMAN
8871|HARMANS
8872|HARMAR HEIGHTS
8873|HARMARVILLE
8874|HARMON
8875|HARMONSBURG
8876|HARMONY
8877|HARNEY
8878|HAROLD
8879|HARPER
8880|HARPER WOODS
8881|HARPERS FERRY
8882|HARPERSVILLE
8883|HARPERVILLE
8884|HARPSTER
8885|HARRAH
8886|HARRELL
8887|HARRELLS
8888|HARRELLSVILLE
8889|HARRIET
8890|HARRIETTA
8891|HARRIETTSVILLE
8892|HARRIMAN
8893|HARRINGTON
8894|HARRINGTON PARK
8895|HARRIS
8896|HARRIS HILL
8897|HARRISBURG
8898|HARRISON
8899|HARRISON CITY
8900|HARRISON GROVE
8901|HARRISON TOWNSHIP
8902|HARRISON VALLEY
8903|HARRISONBURG
8904|HARRISONVILLE
8905|HARRISTON
8906|HARRISTOWN
8907|HARRISVILLE
8908|HARROD
8909|HARRODSBURG
8910|HARROGATE
8911|HARROLD
8912|HARSHAW
8913|HART
8914|HARTFIELD
8915|HARTFORD
8916|HARTFORD CITY
8917|HARTINGTON
8918|HARTLAND
8919|HARTLETON
8920|HARTLEY
8921|HARTLINE
8922|HARTLY
8923|HARTMAN
8924|HARTRANDT
8925|HARTS
8926|HARTSBURG
8927|HARTSDALE
8928|HARTSEL
8929|HARTSELLE
8930|HARTSHORN
8931|HARTSHORNE
8932|HARTSTOWN
8933|HARTSVILLE
8934|HARTVILLE
8935|HARTWELL
8936|HARTWICK
8937|HARVARD
8938|HARVEL
8939|HARVEST
8940|HARVEY
8941|HARVEY CEDARS
8942|HARVEYS LAKE
8943|HARVEYSBURG
8944|HARVEYVILLE
8945|HARVIELL
8946|HARWICH PORT
8947|HARWICK
8948|HARWOOD
8949|HARWOOD HEIGHTS
8950|HASBROUCK HEIGHTS
8951|HASKELL
8952|HASKINS
8953|HASLET
8954|HASLETT
8955|HASSE
8956|HASSELL
8957|HASSMAN
8958|HASSON HEIGHTS
8959|HASTINGS
8960|HASTINGS-ON-HUDSON
8961|HASTY
8962|HASWELL
8963|HAT CREEK
8964|HATBORO
8965|HATCH
8966|HATCHBEND
8967|HATCHECHUBBEE
8968|HATCHEL
8969|HATFIELD
8970|HATHAWAY
8971|HATILLO
8972|HATILLO ZONA URBANA
8973|HATLEY
8974|HATO ARRIBA
8975|HATO ARRIBA COMUNIDAD
8976|HATO CANDAL
8977|HATO CANDAL COMUNIDAD
8978|HATTERAS
8979|HATTIESBURG
8980|HATTIEVILLE
8981|HATTON
8982|HAUBSTADT
8983|HAUGAN
8984|HAUGEN
8985|HAUGHTON
8986|HAUPPAUGE
8987|HAUSER
8988|HAUʻULA
8989|HAVANA
8990|HAVELOCK
8991|HAVEN
8992|HAVENSVILLE
8993|HAVERFORD
8994|HAVERHILL
8995|HAVERSTRAW
8996|HAVERTOWN
8997|HAVILAND
8998|HAVRE
8999|HAVRE DE GRACE
9000|HAW RIVER
9001|HAWAIIAN ACRES
9002|HAWAIIAN BEACHES
9003|HAWAIIAN GARDENS
9004|HAWAIIAN OCEAN VIEW
9005|HAWAIIAN PARADISE PARK
9006|HAWARDEN
9007|HAWESVILLE
9008|HAWICK
9009|HAWK COVE
9010|HAWK INLET
9011|HAWK POINT
9012|HAWK RUN
9013|HAWK SPRINGS
9014|HAWKEYE
9015|HAWKINS
9016|HAWKINSVILLE
9017|HAWKS
9018|HAWLEY
9019|HAWORTH
9020|HAWTHORN
9021|HAWTHORN WOODS
9022|HAWTHORNE
9023|HAXTUN
9024|HAY
9025|HAY CREEK
9026|HAY SPRINGS
9027|HAYCOCK
9028|HAYDEN
9029|HAYDEN LAKE
9030|HAYDEN ROW
9031|HAYDENVILLE
9032|HAYES
9033|HAYES CENTER
9034|HAYESVILLE
9035|HAYFIELD
9036|HAYFORD
9037|HAYFORK
9038|HAYLOW
9039|HAYMARKET
9040|HAYNES
9041|HAYNESVILLE
9042|HAYNEVILLE
9043|HAYS
9044|HAYSI
9045|HAYSVILLE
9046|HAYTI
9047|HAYTI HEIGHTS
9048|HAYWARD
9049|HAYWOOD
9050|HAYWOOD CITY
9051|HAZARD
9052|HAZARDVILLE
9053|HAZEL
9054|HAZEL CREST
9055|HAZEL DELL
9056|HAZEL GREEN
9057|HAZEL HURST
9058|HAZEL PARK
9059|HAZEL RUN
9060|HAZELTON
9061|HAZELWOOD
9062|HAZEN
9063|HAZLEHURST
9064|HAZLET
9065|HAZLETON
9066|HEAD OF THE HARBOR
9067|HEADLAND
9068|HEADQUARTERS
9069|HEADRICK
9070|HEADS
9071|HEAFFORD JUNCTION
9072|HEALDSBURG
9073|HEALDTON
9074|HEALING SPRINGS
9075|HEALY
9076|HEALY LAKE
9077|HEARNE
9078|HEART BUTTE
9079|HEARTWELL
9080|HEATH
9081|HEATH SPRINGS
9082|HEATHCOTE
9083|HEATHROW
9084|HEATHSVILLE
9085|HEATON
9086|HEAVENER
9087|HEBARDVILLE
9088|HEBBARDSVILLE
9089|HEBBRONVILLE
9090|HEBBVILLE
9091|HEBER
9092|HEBER CITY
9093|HEBER SPRINGS
9094|HEBO
9095|HEBRON
9096|HEBRON ESTATES
9097|HECKER
9098|HECKSCHERVILLE
9099|HECKVILLE
9100|HECLA
9101|HECTOR
9102|HEDGESVILLE
9103|HEDLEY
9104|HEDRICK
9105|HEDVILLE
9106|HEDWIG VILLAGE
9107|HEDWIGS HILL
9108|HEENEY
9109|HEFLIN
9110|HEGINS
9111|HEGLAR
9112|HEIBERGER
9113|HEIDELBERG
9114|HEIDLERSBURG
9115|HEIDRICK
9116|HEIL
9117|HEILWOOD
9118|HEIMDAL
9119|HEIZER
9120|HELEN
9121|HELENA
9122|HELENA-WEST HELENA
9123|HELENDALE
9124|HELENVILLE
9125|HELENWOOD
9126|HELIX
9127|HELLERTOWN
9128|HELM
9129|HELMER
9130|HELMETTA
9131|HELMVILLE
9132|HELOTES
9133|HELPER
9134|HELTON
9135|HELTONVILLE
9136|HELVETIA
9137|HEMATITE
9138|HEMBY BRIDGE
9139|HEMET
9140|HEMINGFORD
9141|HEMINGWAY
9142|HEMLOCK
9143|HEMLOCK FARMS
9144|HEMPHILL
9145|HEMPSTEAD
9146|HENAGAR
9147|HENDERSON
9148|HENDERSON POINT
9149|HENDERSONVILLE
9150|HENDLEY
9151|HENDRICKS
9152|HENDRIX
9153|HENDRON
9154|HENDRUM
9155|HENEFER
9156|HENLAWSON
9157|HENLEY
9158|HENLOPEN ACRES
9159|HENLY
9160|HENNEPIN
9161|HENNESSEY
9162|HENNIKER
9163|HENNING
9164|HENRICO
9165|HENRIETTA
9166|HENRIETTE
9167|HENRIEVILLE
9168|HENRY
9169|HENRY FORK
9170|HENRYETTA
9171|HENRYVILLE
9172|HENSEL
9173|HENSHAW
9174|HENSLER
9175|HENSLEY
9176|HEPBURN
9177|HEPHZIBAH
9178|HEPLER
9179|HEPPNER
9180|HEPZIBAH
9181|HERALD
9182|HERALD HARBOR
9183|HERBST
9184|HERBSTER
9185|HERCULANEUM
9186|HERCULES
9187|HERD
9188|HEREFORD
9189|HERENDEEN BAY
9190|HERINGTON
9191|HERITAGE CREEK
9192|HERITAGE HILLS
9193|HERITAGE LAKE
9194|HERITAGE VILLAGE
9195|HERKIMER
9196|HERLONG
9197|HERMAN
9198|HERMANN
9199|HERMANSVILLE
9200|HERMANTOWN
9201|HERMANVILLE
9202|HERMINIE
9203|HERMISTON
9204|HERMITAGE
9205|HERMITAGE SPRINGS
9206|HERMLEIGH
9207|HERMON
9208|HERMOSA
9209|HERMOSA BEACH
9210|HERNANDEZ
9211|HERNANDO
9212|HERNANDO BEACH
9213|HERNDON
9214|HERNSHAW
9215|HEROD
9216|HERON
9217|HERON BAY
9218|HERON LAKE
9219|HERREID
9220|HERRICK
9221|HERRICKS
9222|HERRIMAN
9223|HERRIN
9224|HERRING
9225|HERRINGS
9226|HERRON
9227|HERSCHER
9228|HERSEY
9229|HERSHEY
9230|HERTEL
9231|HERTFORD
9232|HERTY
9233|HERZMAN MESA
9234|HESLER
9235|HESPERIA
9236|HESPERUS
9237|HESS
9238|HESSEL
9239|HESSMER
9240|HESSTON
9241|HESSVILLE
9242|HESTER
9243|HETLAND
9244|HETTICK
9245|HETTINGER
9246|HEUVELTON
9247|HEWINS
9248|HEWITT
9249|HEWLETT
9250|HEWLETT BAY PARK
9251|HEWLETT HARBOR
9252|HEWLETT NECK
9253|HEXT
9254|HEYBURN
9255|HEYWORTH
9256|HEʻEIA
9257|HI-NELLA
9258|HIALEAH
9259|HIALEAH GARDENS
9260|HIATTVILLE
9261|HIAWASSEE
9262|HIAWATHA
9263|HIBBARD
9264|HIBBING
9265|HIBERNIA
9266|HICKMAN
9267|HICKOK
9268|HICKORY
9269|HICKORY CORNERS
9270|HICKORY CREEK
9271|HICKORY FLAT
9272|HICKORY GROVE
9273|HICKORY HILL
9274|HICKORY HILLS
9275|HICKORY PLAINS
9276|HICKORY RIDGE
9277|HICKORY VALLEY
9278|HICKOX
9279|HICKS
9280|HICKSON
9281|HICKSVILLE
9282|HICO
9283|HIDALGO
9284|HIDDEN HILLS
9285|HIDDEN LAKE
9286|HIDDEN MEADOWS
9287|HIDDEN TIMBER
9288|HIDDEN VALLEY
9289|HIDDEN VALLEY LAKE
9290|HIDDENITE
9291|HIDE-A-WAY HILLS
9292|HIDE-A-WAY LAKE
9293|HIDEAWAY
9294|HIDEOUT
9295|HIGBEE
9296|HIGDEN
9297|HIGGANUM
9298|HIGGINS
9299|HIGGINSON
9300|HIGGINSPORT
9301|HIGGINSVILLE
9302|HIGGSTON
9303|HIGH AMANA
9304|HIGH BRIDGE
9305|HIGH FALLS
9306|HIGH HILL
9307|HIGH ISLAND
9308|HIGH LANDING
9309|HIGH POINT
9310|HIGH RIDGE
9311|HIGH ROCK
9312|HIGH ROLLS
9313|HIGH SHOALS
9314|HIGH SPRINGS
9315|HIGHBANK
9316|HIGHCLIFF
9317|HIGHFILL
9318|HIGHGROVE
9319|HIGHLAND
9320|HIGHLAND ACRES
9321|HIGHLAND BEACH
9322|HIGHLAND CENTER
9323|HIGHLAND CITY
9324|HIGHLAND FALLS
9325|HIGHLAND HAVEN
9326|HIGHLAND HEIGHTS
9327|HIGHLAND HILLS
9328|HIGHLAND HOLIDAY
9329|HIGHLAND HOME
9330|HIGHLAND LAKE
9331|HIGHLAND LAKES
9332|HIGHLAND MILLS
9333|HIGHLAND PARK
9334|HIGHLAND SPRINGS
9335|HIGHLAND VIEW
9336|HIGHLAND VILLAGE
9337|HIGHLANDS
9338|HIGHLANDS RANCH
9339|HIGHLANDVILLE
9340|HIGHMORE
9341|HIGHPOINT
9342|HIGHSPIRE
9343|HIGHTSTOWN
9344|HIGHTSVILLE
9345|HIGHWOOD
9346|HIGHWOODS
9347|HIGLEY
9348|HIKO
9349|HILAND
9350|HILBERT
9351|HILBURN
9352|HILDA
9353|HILDALE
9354|HILDEBRAN
9355|HILDEN
9356|HILDRETH
9357|HILGARD
9358|HILGER
9359|HILL 'N DALE
9360|HILL CITY
9361|HILL COUNTRY VILLAGE
9362|HILL TOP
9363|HILL VIEW HEIGHTS
9364|HILLAND
9365|HILLANDALE
9366|HILLBURN
9367|HILLCREST
9368|HILLCREST HEIGHTS
9369|HILLDALE
9370|HILLEMANN
9371|HILLER
9372|HILLHOUSE
9373|HILLIARD
9374|HILLIARDS
9375|HILLISTER
9376|HILLMAN
9377|HILLROSE
9378|HILLS
9379|HILLS AND DALES
9380|HILLS PRAIRIE
9381|HILLSBORO
9382|HILLSBORO BEACH
9383|HILLSBORO PINES
9384|HILLSBOROUGH
9385|HILLSDALE
9386|HILLSIDE
9387|HILLSIDE LAKE
9388|HILLSIDE MANOR
9389|HILLSVIEW
9390|HILLSVILLE
9391|HILLTOP
9392|HILLTOP COLONIA
9393|HILLTOP LAKES
9394|HILLVIEW
9395|HILMAR
9396|HILO
9397|HILSHIRE VILLAGE
9398|HILT
9399|HILTON
9400|HILTON HEAD ISLAND
9401|HILTONIA
9402|HINCHCLIFF
9403|HINCKLEY
9404|HINDMAN
9405|HINDSBORO
9406|HINDSVILLE
9407|HINES
9408|HINESBURG
9409|HINESTON
9410|HINESVILLE
9411|HINGHAM
9412|HINKLEY
9413|HINSDALE
9414|HINSON
9415|HINTON
9416|HIOUCHI
9417|HIRAM
9418|HISEVILLE
9419|HISLE
9420|HISSOP
9421|HITCHCOCK
9422|HITCHITA
9423|HITCHLAND
9424|HITEMAN
9425|HITSCHMANN
9426|HITTERDAL
9427|HIWANNEE
9428|HIWASSE
9429|HIWASSEE
9430|HIXSON
9431|HIXTON
9432|HO-HO-KUS
9433|HOADLY
9434|HOAGLAND
9435|HOBACK
9436|HOBAN
9437|HOBART
9438|HOBART BAY
9439|HOBBS
9440|HOBE SOUND
9441|HOBERG
9442|HOBERGS
9443|HOBGOOD
9444|HOBOKEN
9445|HOBSON
9446|HOBSON CITY
9447|HOBUCKEN
9448|HOCHHEIM
9449|HOCKESSIN
9450|HOCKINGPORT
9451|HOCKINSON
9452|HOCKLEY
9453|HODGE
9454|HODGENVILLE
9455|HODGES
9456|HODGESVILLE
9457|HODGKINS
9458|HOEHNE
9459|HOFFMAN
9460|HOFFMAN ESTATES
9461|HOGANSBURG
9462|HOGANSVILLE
9463|HOGATZA
9464|HOGELAND
9465|HOHENWALD
9466|HOISINGTON
9467|HOKAH
9468|HOKENDAUQUA
9469|HOKES BLUFF
9470|HOLABIRD
9471|HOLBROOK
9472|HOLCOMB
9473|HOLCOMBE
9474|HOLCUT
9475|HOLDEN
9476|HOLDEN BEACH
9477|HOLDEN HEIGHTS
9478|HOLDENVILLE
9479|HOLDER
9480|HOLDINGFORD
9481|HOLDREGE
9482|HOLGATE
9483|HOLIDAY
9484|HOLIDAY BEACH
9485|HOLIDAY CITY
9486|HOLIDAY HEIGHTS
9487|HOLIDAY HILLS
9488|HOLIDAY ISLAND
9489|HOLIDAY LAKE
9490|HOLIDAY LAKES
9491|HOLIDAY POCONO
9492|HOLIDAY SHORES
9493|HOLIDAY VALLEY
9494|HOLIKACHUK
9495|HOLLADAY
9496|HOLLAND
9497|HOLLAND PATENT
9498|HOLLANDALE
9499|HOLLANDSBURG
9500|HOLLANSBURG
9501|HOLLENBERG
9502|HOLLEY
9503|HOLLIDAY
9504|HOLLIDAYSBURG
9505|HOLLINS
9506|HOLLIS
9507|HOLLIS CROSSROADS
9508|HOLLISTER
9509|HOLLOW CREEK
9510|HOLLOW ROCK
9511|HOLLOWAY
9512|HOLLOWAY TERRACE
9513|HOLLOWAYVILLE
9514|HOLLY
9515|HOLLY BEACH
9516|HOLLY BLUFF
9517|HOLLY GROVE
9518|HOLLY HILL
9519|HOLLY HILLS
9520|HOLLY OAK
9521|HOLLY POND
9522|HOLLY RIDGE
9523|HOLLY SPRINGS
9524|HOLLYHILL
9525|HOLLYMEAD
9526|HOLLYVILLA
9527|HOLLYWOOD
9528|HOLLYWOOD HEIGHTS
9529|HOLLYWOOD PARK
9530|HOLMAN
9531|HOLMDEL
9532|HOLMEN
9533|HOLMES BEACH
9534|HOLMES CITY
9535|HOLMESVILLE
9536|HOLOPAW
9537|HOLSTEIN
9538|HOLT
9539|HOLTON
9540|HOLTS CORNER
9541|HOLTS SUMMIT
9542|HOLTSVILLE
9543|HOLTVILLE
9544|HOLTWOOD
9545|HOLY CROSS
9546|HOLYOKE
9547|HOLYROOD
9548|HOMA HILLS
9549|HOME GARDEN
9550|HOME GARDENS
9551|HOMEACRE
9552|HOMECROFT
9553|HOMEDALE
9554|HOMELAND
9555|HOMELAND PARK
9556|HOMER
9557|HOMER CITY
9558|HOMER GLEN
9559|HOMERVILLE
9560|HOMESTEAD
9561|HOMESTEAD PARK
9562|HOMESTOWN
9563|HOMETOWN
9564|HOMEVILLE
9565|HOMEWOOD
9566|HOMEWORTH
9567|HOMINY
9568|HOMOSASSA
9569|HOMOSASSA SPRINGS
9570|HON
9571|HONAKER
9572|HONALO
9573|HONCUT
9574|HONDA
9575|HONDO
9576|HONEA PATH
9577|HONEOYE
9578|HONEOYE FALLS
9579|HONESDALE
9580|HONEY BROOK
9581|HONEY GROVE
9582|HONEY ISLAND
9583|HONEYDEW
9584|HONEYVILLE
9585|HONOBIA
9586|HONOKAHUA
9587|HONOKAʻA
9588|HONOLULU
9589|HONOMU
9590|HONOR
9591|HONORAVILLE
9592|HONUʻAPO
9593|HOOD
9594|HOOD RIVER
9595|HOODSPORT
9596|HOOKDALE
9597|HOOKER
9598|HOOKERTON
9599|HOOKS
9600|HOOKSETT
9601|HOOKSTOWN
9602|HOONAH
9603|HOOPA
9604|HOOPER
9605|HOOPER BAY
9606|HOOPERS CREEK
9607|HOOPERSVILLE
9608|HOOPESTON
9609|HOOPLE
9610|HOOPPOLE
9611|HOOSICK FALLS
9612|HOOT OWL
9613|HOOVEN
9614|HOOVER
9615|HOOVERSON HEIGHTS
9616|HOOVERSVILLE
9617|HOP BOTTOM
9618|HOPATCONG
9619|HOPE
9620|HOPE MILLS
9621|HOPE VALLEY
9622|HOPEDALE
9623|HOPEFUL HEIGHTS
9624|HOPELAND
9625|HOPETON
9626|HOPEWELL
9627|HOPEWELL JUNCTION
9628|HOPKINS
9629|HOPKINS PARK
9630|HOPKINSVILLE
9631|HOPKINTON
9632|HOPLAND
9633|HOPPER
9634|HOPWOOD
9635|HOQUIAM
9636|HORACE
9637|HORATIO
9638|HORATIO GARDENS
9639|HORD
9640|HORDVILLE
9641|HORICON
9642|HORINE
9643|HORIZON CITY
9644|HORMIGUEROS
9645|HORMIGUEROS ZONA URBANA
9646|HORN HILL
9647|HORN LAKE
9648|HORNBEAK
9649|HORNBECK
9650|HORNBROOK
9651|HORNELL
9652|HORNERSTOWN
9653|HORNERSVILLE
9654|HORNICK
9655|HORNITOS
9656|HORNS
9657|HORNSBY
9658|HORNSBY BEND
9659|HORNTOWN
9660|HORREL HILL
9661|HORSE BRANCH
9662|HORSE CAVE
9663|HORSE CREEK
9664|HORSE PASTURE
9665|HORSE SHOE
9666|HORSEHEAD
9667|HORSEHEADS
9668|HORSESHOE BAY
9669|HORSESHOE BEACH
9670|HORSESHOE BEND
9671|HORSESHOE LAKE
9672|HORSHAM
9673|HORTENSE
9674|HORTON
9675|HORTON BAY
9676|HORTONVILLE
9677|HOSCHTON
9678|HOSFORD
9679|HOSKINS
9680|HOSKINSTON
9681|HOSMER
9682|HOSPERS
9683|HOSSTON
9684|HOSTETTER
9685|HOT SPRINGS
9686|HOT SPRINGS LANDING
9687|HOT SPRINGS VILLAGE
9688|HOT SULPHUR SPRINGS
9689|HOTCHKISS
9690|HOTEVILLA
9691|HOTEVILLA-BACAVI
9692|HOUCK
9693|HOUGH
9694|HOUGHTON
9695|HOUGHTON LAKE
9696|HOULKA
9697|HOULTON
9698|HOUMA
9699|HOUMONT PARK
9700|HOUSATONIC
9701|HOUSE SPRINGS
9702|HOUSERVILLE
9703|HOUSTON
9704|HOUSTON ACRES
9705|HOUSTON LAKE
9706|HOUSTONIA
9707|HOUTZDALE
9708|HOVEN
9709|HOVLAND
9710|HOWARD
9711|HOWARD CITY
9712|HOWARD LAKE
9713|HOWARDS GROVE
9714|HOWARDSTOWN
9715|HOWARDVILLE
9716|HOWARDWICK
9717|HOWE
9718|HOWELL
9719|HOWELLS
9720|HOWES
9721|HOWES MILL
9722|HOWESVILLE
9723|HOWIE IN THE HILLS
9724|HOWISON
9725|HOWLAND
9726|HOWLAND CENTER
9727|HOXIE
9728|HOYLETON
9729|HOYT
9730|HOYT LAKES
9731|HOYTSVILLE
9732|HOYTVILLE
9733|HOʻOLEHUA
9734|HUACHUCA CITY
9735|HUBBARD
9736|HUBBARD LAKE
9737|HUBBARDSTON
9738|HUBBELL
9739|HUBER
9740|HUBER HEIGHTS
9741|HUBER RIDGE
9742|HUBLERSBURG
9743|HUCKABAY
9744|HUDSON
9745|HUDSON BEND
9746|HUDSON FALLS
9747|HUDSON LAKE
9748|HUDSON OAKS
9749|HUDSONVILLE
9750|HUETTER
9751|HUEY
9752|HUEYTOWN
9753|HUFFMAN
9754|HUGH
9755|HUGHES
9756|HUGHES SPRINGS
9757|HUGHESTOWN
9758|HUGHESVILLE
9759|HUGHSON
9760|HUGO
9761|HUGOTON
9762|HUGULEY
9763|HULAH
9764|HULBERT
9765|HULETT
9766|HULL
9767|HULMEVILLE
9768|HUMACAO
9769|HUMACAO ZONA URBANA
9770|HUMANSVILLE
9771|HUMAROCK
9772|HUMBIRD
9773|HUMBLE
9774|HUMBLE CITY
9775|HUMBOLDT
9776|HUMBOLDT HILL
9777|HUME
9778|HUMESTON
9779|HUMMELS WHARF
9780|HUMMELSTOWN
9781|HUMNOKE
9782|HUMPHREY
9783|HUMPHREYS
9784|HUMPTULIPS
9785|HUNDRED
9786|HUNGERFORD
9787|HUNGRY HORSE
9788|HUNKER
9789|HUNNEWELL
9790|HUNT
9791|HUNTER
9792|HUNTERDON
9793|HUNTERS
9794|HUNTERS CREEK
9795|HUNTERS CREEK VILLAGE
9796|HUNTERS HOLLOW
9797|HUNTERSTOWN
9798|HUNTERSVILLE
9799|HUNTERTOWN
9800|HUNTING VALLEY
9801|HUNTINGBURG
9802|HUNTINGDON
9803|HUNTINGTON
9804|HUNTINGTON BAY
9805|HUNTINGTON BEACH
9806|HUNTINGTON PARK
9807|HUNTINGTON STATION
9808|HUNTINGTON WOODS
9809|HUNTINGTOWN
9810|HUNTLAND
9811|HUNTLEIGH
9812|HUNTLEY
9813|HUNTOON
9814|HUNTS POINT
9815|HUNTSDALE
9816|HUNTSVILLE
9817|HURDLAND
9818|HURDLE MILLS
9819|HURDSFIELD
9820|HURDTOWN
9821|HURFFVILLE
9822|HURLEY
9823|HURLOCK
9824|HURON
9825|HURON BEACH
9826|HURRICANE
9827|HURST
9828|HURSTBOURNE
9829|HURSTBOURNE ACRES
9830|HURSTVILLE
9831|HURT
9832|HURTSBORO
9833|HUSCHER
9834|HUSHPUCKENA
9835|HUSLIA
9836|HUSON
9837|HUSSER
9838|HUSTISFORD
9839|HUSTLER
9840|HUSTON
9841|HUSTONVILLE
9842|HUSUM
9843|HUTCHINS
9844|HUTCHINSON
9845|HUTSONVILLE
9846|HUTTIG
9847|HUTTO
9848|HUTTON
9849|HUTTONSVILLE
9850|HUXFORD
9851|HUXLEY
9852|HYAK
9853|HYAMPOM
9854|HYANNIS
9855|HYATTSVILLE
9856|HYATTVILLE
9857|HYBART
9858|HYBLA VALLEY
9859|HYDABURG
9860|HYDE
9861|HYDE PARK
9862|HYDEN
9863|HYDER
9864|HYDESVILLE
9865|HYDETOWN
9866|HYDRO
9867|HYE
9868|HYGIENE
9869|HYMER
9870|HYMERA
9871|HYNDMAN
9872|HYPOLUXO
9873|HYRUM
9874|HYSHAM
9875|HYTOP
9876|HĀLAWA
9877|HĀLIʻIMAILE
9878|HĀNA
9879|HĀWĪ
9880|HĀʻENA
9881|HŌLUALOA
9882|IAEGER
9883|IAGO
9884|IATAN
9885|IBAPAH
9886|IBERIA
9887|IBERVILLE
9888|ICARD
9889|ICKESBURG
9890|ICONIUM
9891|IDA
9892|IDA GROVE
9893|IDA MAY
9894|IDABEL
9895|IDAHO CITY
9896|IDAHO FALLS
9897|IDAHO SPRINGS
9898|IDALIA
9899|IDALOU
9900|IDAMAY
9901|IDANA
9902|IDANHA
9903|IDAVILLE
9904|IDER
9905|IDLEDALE
9906|IDLEWILD
9907|IDLEYLD PARK
9908|IDMON
9909|IDRIA
9910|IDYLLWILD
9911|IDYLSIDE
9912|IDYLWOOD
9913|IGIUGIG
9914|IGLOO
9915|IGNACIO
9916|IGO
9917|IHLEN
9918|IKATAN
9919|ILA
9920|ILCHESTER
9921|ILIAD
9922|ILIAMNA
9923|ILIFF
9924|ILION
9925|ILLINOIS CITY
9926|ILLIOPOLIS
9927|ILLMO
9928|ILWACO
9929|IMBERY
9930|IMBLER
9931|IMBODEN
9932|IMBS
9933|IMBÉRY COMUNIDAD
9934|IMLAY
9935|IMLAY CITY
9936|IMLAYSTOWN
9937|IMMOKALEE
9938|IMOGENE
9939|IMPACT
9940|IMPERIAL
9941|IMPERIAL BEACH
9942|INA
9943|INADALE
9944|INAVALE
9945|INCHELIUM
9946|INCLINE VILLAGE
9947|INDEPENDENCE
9948|INDEPENDENCE CORNER
9949|INDEPENDENCE HILL
9950|INDEPENDENT HILL
9951|INDEX
9952|INDIA
9953|INDIA HOOK
9954|INDIAHOMA
9955|INDIALANTIC
9956|INDIAN BEACH
9957|INDIAN CREEK
9958|INDIAN CREEK VILLAGE
9959|INDIAN FALLS
9960|INDIAN HARBOUR BEACH
9961|INDIAN HEAD
9962|INDIAN HEAD PARK
9963|INDIAN HEIGHTS
9964|INDIAN HILLS
9965|INDIAN LAKE
9966|INDIAN MOUND
9967|INDIAN MOUNTAIN LAKE
9968|INDIAN PASS
9969|INDIAN POINT
9970|INDIAN RIVER
9971|INDIAN RIVER CITY
9972|INDIAN RIVER ESTATES
9973|INDIAN RIVER SHORES
9974|INDIAN ROCKS BEACH
9975|INDIAN SHORES
9976|INDIAN SPRINGS
9977|INDIAN SPRINGS VILLAGE
9978|INDIAN TRAIL
9979|INDIAN VALLEY
9980|INDIAN VILLAGE
9981|INDIAN WELLS
9982|INDIANA
9983|INDIANAPOLIS
9984|INDIANOLA
9985|INDIANTOWN
9986|INDIO
9987|INDIO HILLS
9988|INDIOS
9989|INDIOS COMUNIDAD
9990|INDRIO
9991|INDUS
9992|INDUSTRY
9993|INEZ
9994|INGALLS
9995|INGALLS PARK
9996|INGENIO
9997|INGENIO COMUNIDAD
9998|INGER
9999|INGERSOLL
10000|INGLEFIELD
10001|INGLESIDE
10002|INGLESIDE ON-THE-BAY
10003|INGLEWOOD
10004|INGLIS
10005|INGOLD
10006|INGOMAR
10007|INGOT
10008|INGRAHAM
10009|INGRAM
10010|INGUADONA
10011|INKERMAN
10012|INKOM
10013|INKSTER
10014|INLAND
10015|INMAN
10016|INMAN MILLS
10017|INNIS
10018|INNISWOLD
10019|INNSBROOK
10020|INOLA
10021|INSTITUTE
10022|INTERCESSION CITY
10023|INTERIOR
10024|INTERLACHEN
10025|INTERLAKEN
10026|INTERLOCHEN
10027|INTERNATIONAL FALLS
10028|INTRACOASTAL CITY
10029|INVER GROVE HEIGHTS
10030|INVERNESS
10031|INWOOD
10032|INYOKERN
10033|IOLA
10034|IONA
10035|IONE
10036|IONIA
10037|IOTA
10038|IOWA
10039|IOWA CITY
10040|IOWA COLONY
10041|IOWA FALLS
10042|IOWA PARK
10043|IOWA POINT
10044|IPAVA
10045|IPSWICH
10046|IRA
10047|IRAAN
10048|IRASBURG
10049|IRBY
10050|IREDELL
10051|IRELAND
10052|IRENA
10053|IRENE
10054|IRETON
10055|IRMA
10056|IRMO
10057|IRON BELT
10058|IRON CITY
10059|IRON GATE
10060|IRON GATES
10061|IRON HILL
10062|IRON HORSE
10063|IRON JUNCTION
10064|IRON LIGHTNING
10065|IRON MOUNTAIN
10066|IRON MOUNTAIN LAKE
10067|IRON POST
10068|IRON RIDGE
10069|IRON RIVER
10070|IRON SPRINGS
10071|IRON STATION
10072|IRONATON
10073|IRONDALE
10074|IRONDEQUOIT
10075|IRONIA
10076|IRONSIDE
10077|IRONTON
10078|IRONVILLE
10079|IRONWOOD
10080|IROQUOIS
10081|IROQUOIS POINT
10082|IRRIGON
10083|IRVINE
10084|IRVING
10085|IRVINGTON
10086|IRVONA
10087|IRWIN
10088|IRWINDALE
10089|IRWINTON
10090|IRWINVILLE
10091|ISABEL
10092|ISABELA
10093|ISABELA ZONA URBANA
10094|ISABELLA
10095|ISANTI
10096|ISBELL
10097|ISELIN
10098|ISHPEMING
10099|ISLA
10100|ISLA VISTA
10101|ISLAMORADA
10102|ISLAND
10103|ISLAND CITY
10104|ISLAND GROVE
10105|ISLAND HEIGHTS
10106|ISLAND LAKE
10107|ISLAND MOUNTAIN
10108|ISLAND PARK
10109|ISLAND POND
10110|ISLAND VIEW
10111|ISLANDIA
10112|ISLANDTON
10113|ISLE
10114|ISLE AU HAUT
10115|ISLE OF HOPE
10116|ISLE OF PALMS
10117|ISLE OF WIGHT
10118|ISLEN
10119|ISLETA
10120|ISLETON
10121|ISLINGTON
10122|ISLIP
10123|ISLIP TERRACE
10124|ISMAY
10125|ISOLA
10126|ISSAQUAH
10127|ISTACHATTA
10128|ITALIA
10129|ITALY
10130|ITASCA
10131|ITHACA
10132|ITMANN
10133|ITTA BENA
10134|IUKA
10135|IVA
10136|IVALEE
10137|IVAN
10138|IVANHOE
10139|IVANOF BAY
10140|IVANPAH
10141|IVES ESTATES
10142|IVESDALE
10143|IVEY
10144|IVINS
10145|IVOR
10146|IVYDALE
10147|IVYLAND
10148|IXL
10149|IXONIA
10150|IZAGORA
10151|IZEE
10152|JAARS
10153|JACINTO CITY
10154|JACKPOT
10155|JACKSBORO
10156|JACKSON
10157|JACKSON CENTER
10158|JACKSON HEIGHTS
10159|JACKSON JUNCTION
10160|JACKSONBORO
10161|JACKSONBURG
10162|JACKSONPORT
10163|JACKSONS GAP
10164|JACKSONS MILLS
10165|JACKSONTOWN
10166|JACKSONVILLE
10167|JACKSONVILLE BEACH
10168|JACKSONWALD
10169|JACKSTOWN
10170|JACOB LAKE
10171|JACOBS
10172|JACOBSBURG
10173|JACOBSON
10174|JACOBSVILLE
10175|JACOBUS
10176|JACONA
10177|JACONITA
10178|JACUMBA HOT SPRINGS
10179|JAFFREY
10180|JAGUAL
10181|JAGUAL COMUNIDAD
10182|JAKES CORNER
10183|JAKIN
10184|JAKOLOF BAY
10185|JAL
10186|JALAPA
10187|JAMACHA JUNCTION
10188|JAMAICA
10189|JAMAICA BEACH
10190|JAMES
10191|JAMES CITY
10192|JAMES TOWN
10193|JAMESBURG
10194|JAMESON
10195|JAMESPORT
10196|JAMESTOWN
10197|JAMESVILLE
10198|JAMIESON
10199|JAMISON
10200|JAMISON CITY
10201|JAMUL
10202|JAN-PHYL VILLAGE
10203|JANE
10204|JANE LEW
10205|JANESVILLE
10206|JANNEY
10207|JANSEN
10208|JAPTON
10209|JARALES
10210|JARBIDGE
10211|JARDINE
10212|JAROSO
10213|JARRATT
10214|JARREAU
10215|JARRELL
10216|JARRETTSVILLE
10217|JARVISBURG
10218|JASMINE ESTATES
10219|JASONVILLE
10220|JASPER
10221|JAUCA
10222|JAUCA COMUNIDAD
10223|JAVA
10224|JAY
10225|JAYTON
10226|JAYUYA
10227|JAYUYA ZONA URBANA
10228|JEAN
10229|JEAN LAFITTE
10230|JEANERETTE
10231|JEANNETTE
10232|JEDDITO
10233|JEDDO
10234|JEFF
10235|JEFFERS
10236|JEFFERSON
10237|JEFFERSON CITY
10238|JEFFERSON HEIGHTS
10239|JEFFERSON HILLS
10240|JEFFERSON ISLAND
10241|JEFFERSON VALLEY
10242|JEFFERSONTON
10243|JEFFERSONTOWN
10244|JEFFERSONVILLE
10245|JEFFREY
10246|JEFFREY CITY
10247|JEISYVILLE
10248|JELLICO
10249|JELLOWAY
10250|JELM
10251|JEMEZ PUEBLO
10252|JEMEZ SPRINGS
10253|JEMISON
10254|JENA
10255|JENERA
10256|JENIFER
10257|JENISON
10258|JENKINJONES
10259|JENKINS
10260|JENKINSBURG
10261|JENKINSVILLE
10262|JENKINTOWN
10263|JENKS
10264|JENNER
10265|JENNERS
10266|JENNERSTOWN
10267|JENNERSVILLE
10268|JENNETTE
10269|JENNIE
10270|JENNINGS
10271|JENNINGS LODGE
10272|JENSEN
10273|JENSEN BEACH
10274|JERICHO
10275|JERICO
10276|JERICO SPRINGS
10277|JERMYN
10278|JEROME
10279|JEROMESVILLE
10280|JERRY CITY
10281|JERRYVILLE
10282|JERSEY
10283|JERSEY CITY
10284|JERSEY SHORE
10285|JERSEY VILLAGE
10286|JERSEYTOWN
10287|JERSEYVILLE
10288|JERUSALEM
10289|JESMOND DENE
10290|JESSIE
10291|JESSIETOWN
10292|JESSIEVILLE
10293|JESSUP
10294|JESTERVILLE
10295|JESUP
10296|JET
10297|JETERSVILLE
10298|JETMORE
10299|JETTE
10300|JEWELL
10301|JEWELL RIDGE
10302|JEWELL VALLEY
10303|JEWETT
10304|JEWETT CITY
10305|JEWETTVILLE
10306|JIGGER
10307|JIM FALLS
10308|JIM THORPE
10309|JINGO
10310|JOANNA
10311|JOAQUIN
10312|JOBOS
10313|JOBOS COMUNIDAD
10314|JOBSTOWN
10315|JOEL
10316|JOES
10317|JOFFRE
10318|JOHANNESBURG
10319|JOHN DAY
10320|JOHNETTA
10321|JOHNFARRIS
10322|JOHNS
10323|JOHNS CREEK
10324|JOHNS ISLAND
10325|JOHNSBURG
10326|JOHNSON
10327|JOHNSON CITY
10328|JOHNSON CORNER
10329|JOHNSON CREEK
10330|JOHNSON LANE
10331|JOHNSON SIDING
10332|JOHNSON VILLAGE
10333|JOHNSONBURG
10334|JOHNSONDALE
10335|JOHNSONS STATION
10336|JOHNSONVILLE
10337|JOHNSTON
10338|JOHNSTON CITY
10339|JOHNSTONE
10340|JOHNSTONVILLE
10341|JOHNSTOWN
10342|JOHNSTOWN CENTER
10343|JOHNSVILLE
10344|JOHNTOWN
10345|JOICE
10346|JOINER
10347|JOLIET
10348|JOLIVUE
10349|JOLLEY
10350|JOLLY
10351|JOLLYVILLE
10352|JONAH
10353|JONANCY
10354|JONES CHAPEL
10355|JONES CREEK
10356|JONES MILLS
10357|JONES POINT
10358|JONESBORO
10359|JONESBOROUGH
10360|JONESBURG
10361|JONESTOWN
10362|JONESVILLE
10363|JOPLIN
10364|JOPPA
10365|JOPPATOWNE
10366|JORDAN
10367|JORDAN HILL
10368|JORDAN VALLEY
10369|JOSEPH
10370|JOSEPH CITY
10371|JOSEPHINE
10372|JOSEPHVILLE
10373|JOSHUA
10374|JOSHUA TREE
10375|JOSLIN
10376|JOURDANTON
10377|JOY
10378|JOYCE
10379|JUANA DÍAZ
10380|JUANA DÍAZ ZONA URBANA
10381|JUANITA
10382|JUBILEE SPRINGS
10383|JUD
10384|JUDA
10385|JUDITH GAP
10386|JUDSON
10387|JUDSONIA
10388|JUDYVILLE
10389|JUGTOWN
10390|JUILLIARD
10391|JULESBURG
10392|JULIAETTA
10393|JULIAN
10394|JULIETTE
10395|JULIFF
10396|JULIUSTOWN
10397|JUMP RIVER
10398|JUMPERTOWN
10399|JUNCAL
10400|JUNCAL COMUNIDAD
10401|JUNCOS
10402|JUNCOS ZONA URBANA
10403|JUNCTION CITY
10404|JUNE LAKE
10405|JUNE PARK
10406|JUNEAU
10407|JUNIATA
10408|JUNIATA TERRACE
10409|JUNIOR
10410|JUNIPER
10411|JUNIUS
10412|JUNO
10413|JUNO BEACH
10414|JUNO RIDGE
10415|JUNTURA
10416|JUPITER
10417|JUPITER INLET BEACH COLONY
10418|JUPITER ISLAND
10419|JUSTICE
10420|JUSTICEBURG
10421|JUSTIN
10422|JUSTUS
10423|K I SAWYER
10424|K-BAR RANCH
10425|KACHEMAK CITY
10426|KACHINA VILLAGE
10427|KACKLEY
10428|KADANE CORNER
10429|KADOKA
10430|KAFFIR
10431|KAHAKULOA
10432|KAHALUʻU
10433|KAHLOTUS
10434|KAHOKA
10435|KAHUKU
10436|KAHULUI
10437|KAIBAB
10438|KAIBITO
10439|KAILUA
10440|KAKA
10441|KAKE
10442|KAKTOVIK
10443|KALALOCH
10444|KALAMA
10445|KALAMAZOO
10446|KALAOA
10447|KALAUPAPA
10448|KALEVA
10449|KALIDA
10450|KALIFORNSKY
10451|KALIHI WAI
10452|KALISPELL
10453|KALKASKA
10454|KALONA
10455|KALSKAG
10456|KALTAG
10457|KALUAʻAHA
10458|KALVESTA
10459|KALĀHEO
10460|KAMALŌ
10461|KAMAS
10462|KAMEY
10463|KAMIAH
10464|KAMPSVILLE
10465|KAMRAR
10466|KANAB
10467|KANARANZI
10468|KANARRAVILLE
10469|KANASKAT
10470|KANAUGA
10471|KANAWHA
10472|KANDIYOHI
10473|KANE
10474|KANEVILLE
10475|KANGLEY
10476|KANKAKEE
10477|KANNAPOLIS
10478|KANOPOLIS
10479|KANORADO
10480|KANOSH
10481|KANSAS
10482|KANSAS CITY
10483|KAOLIN
10484|KAPALUA
10485|KAPAʻA
10486|KAPAʻAU
10487|KAPLAN
10488|KAPOLEI
10489|KAPOWSIN
10490|KAPP HEIGHTS
10491|KAPPA
10492|KARLSRUHE
10493|KARLSTAD
10494|KARLUK
10495|KARNACK
10496|KARNAK
10497|KARNES CITY
10498|KARNS
10499|KARNS CITY
10500|KARTHAUS
10501|KARVAL
10502|KASAAN
10503|KASER
10504|KASHEGELOK
10505|KASIGLUK
10506|KASILOF
10507|KASKASKIA
10508|KASOTA
10509|KASSON
10510|KATALLA
10511|KATEMCY
10512|KATHERINE
10513|KATHLEEN
10514|KATHRYN
10515|KATIE
10516|KATONAH
10517|KATY
10518|KAUFMAN
10519|KAUKAUNA
10520|KAUMAKANI
10521|KAUMALAPAU
10522|KAUNAKAKAI
10523|KAW CITY
10524|KAWAIHAE
10525|KAWEAH
10526|KAWELA BAY
10527|KAWKAWLIN
10528|KAYCEE
10529|KAYENTA
10530|KAYLOR
10531|KAYSVILLE
10532|KAʻAʻAWA
10533|KEALAKEKUA
10534|KEAMS CANYON
10535|KEANSBURG
10536|KEARNEY
10537|KEARNEY PARK
10538|KEARNEYSVILLE
10539|KEARNS
10540|KEARNY
10541|KEATCHIE
10542|KEATING
10543|KEATS
10544|KEAUHOU
10545|KEAVY
10546|KEAʻAU
10547|KECHI
10548|KEDDIE
10549|KEDRON
10550|KEEDYSVILLE
10551|KEEFTON
10552|KEEGO HARBOR
10553|KEELER
10554|KEELINE
10555|KEENAN
10556|KEENE
10557|KEENER
10558|KEENES
10559|KEENESBURG
10560|KEENEYVILLE
10561|KEENSBURG
10562|KEESEVILLE
10563|KEEWATIN
10564|KEISER
10565|KEITHSBURG
10566|KEITHVILLE
10567|KEIZER
10568|KEKAHA
10569|KEKOSKEE
10570|KELAYRES
10571|KELFORD
10572|KELL
10573|KELLER
10574|KELLERTON
10575|KELLERVILLE
10576|KELLEY
10577|KELLEYS ISLAND
10578|KELLIHER
10579|KELLNER
10580|KELLNERSVILLE
10581|KELLOGG
10582|KELLOGGSVILLE
10583|KELLY
10584|KELLY LAKE
10585|KELLYTON
10586|KELLYVILLE
10587|KELSAY
10588|KELSEY
10589|KELSEYVILLE
10590|KELSO
10591|KELTON
10592|KELTYS
10593|KELVIN
10594|KEMAH
10595|KEMBLESVILLE
10596|KEMMERER
10597|KEMP
10598|KEMP MILL
10599|KEMPNER
10600|KEMPSTER
10601|KEMPTON
10602|KEN CARYL
10603|KENAI
10604|KENANSVILLE
10605|KENBRIDGE
10606|KENDALE LAKES
10607|KENDALL
10608|KENDALL PARK
10609|KENDALLVILLE
10610|KENDLETON
10611|KENDRICK
10612|KENEDY
10613|KENEFIC
10614|KENEFICK
10615|KENEL
10616|KENESAW
10617|KENHORST
10618|KENILWORTH
10619|KENLY
10620|KENMAR
10621|KENMARE
10622|KENMAWR
10623|KENMORE
10624|KENNA
10625|KENNAN
10626|KENNARD
10627|KENNARD CORNER
10628|KENNEBEC
10629|KENNEBUNK
10630|KENNEBUNKPORT
10631|KENNEDALE
10632|KENNEDY
10633|KENNEDYVILLE
10634|KENNER
10635|KENNERDELL
10636|KENNESAW
10637|KENNETH
10638|KENNETH CITY
10639|KENNETT
10640|KENNETT SQUARE
10641|KENNEWICK
10642|KENNEY
10643|KENNY LAKE
10644|KENNYDALE
10645|KENO
10646|KENOSHA
10647|KENOVA
10648|KENSAL
10649|KENSETT
10650|KENSINGTON
10651|KENSINGTON PARK
10652|KENT
10653|KENT ACRES
10654|KENT CITY
10655|KENT NARROWS
10656|KENT PARK
10657|KENTFIELD
10658|KENTLAND
10659|KENTMORE PARK
10660|KENTON
10661|KENTON VALE
10662|KENTWOOD
10663|KENVIL
10664|KENVIR
10665|KENWOOD
10666|KENYON
10667|KEO
10668|KEOKEE
10669|KEOKUK
10670|KEOMAH VILLAGE
10671|KEOSAUQUA
10672|KEOTA
10673|KERBY
10674|KERENS
10675|KERHONKSON
10676|KERKHOVEN
10677|KERMAN
10678|KERMIT
10679|KERNERSVILLE
10680|KERNVILLE
10681|KERR
10682|KERRICK
10683|KERRTOWN
10684|KERRVILLE
10685|KERSEY
10686|KERSHAW
10687|KESHENA
10688|KESLEY
10689|KESWICK
10690|KETCHIKAN
10691|KETCHUM
10692|KETRON
10693|KETTERING
10694|KETTLE FALLS
10695|KETTLE RIVER
10696|KETTLEMAN CITY
10697|KETTLERSVILLE
10698|KEUKA
10699|KEUKA PARK
10700|KEVIL
10701|KEVIN
10702|KEWA
10703|KEWANEE
10704|KEWANNA
10705|KEWASKUM
10706|KEWAUNEE
10707|KEWEENAW BAY
10708|KEY
10709|KEY BISCAYNE
10710|KEY CENTER
10711|KEY COLONY BEACH
10712|KEY LARGO
10713|KEY WEST
10714|KEYAPAHA
10715|KEYES
10716|KEYES SUMMIT
10717|KEYESPORT
10718|KEYPORT
10719|KEYS
10720|KEYSER
10721|KEYSTONE
10722|KEYSTONE HEIGHTS
10723|KEYSVILLE
10724|KEYTESVILLE
10725|KEZAR FALLS
10726|KIAHSVILLE
10727|KIANA
10728|KIAWAH ISLAND
10729|KIBLAH
10730|KIBLER
10731|KICKING HORSE
10732|KIDDER
10733|KIDRON
10734|KIEF
10735|KIEFER
10736|KIEL
10737|KIELER
10738|KIESTER
10739|KILA
10740|KILBOURNE
10741|KILDARE
10742|KILDEER
10743|KILGORE
10744|KILKARE WOODS
10745|KILKENNY
10746|KILL DEVIL HILLS
10747|KILLBUCK
10748|KILLDEER
10749|KILLDUFF
10750|KILLEEN
10751|KILLEN
10752|KILLIAN
10753|KILLONA
10754|KILMARNOCK
10755|KILMICHAEL
10756|KILN
10757|KIM
10758|KIMBALL
10759|KIMBALLTON
10760|KIMBERLING CITY
10761|KIMBERLY
10762|KIMBERTON
10763|KIMBOLTON
10764|KIMBROUGH
10765|KIMMELL
10766|KIMMINS
10767|KIMMSWICK
10768|KIMPER
10769|KINARD
10770|KINARDS
10771|KINBRAE
10772|KINCAID
10773|KINDE
10774|KINDER
10775|KINDERHOOK
10776|KINDERLOU
10777|KINDRED
10778|KING
10779|KING AND QUEEN COURT HOUSE
10780|KING ARTHUR PARK
10781|KING CITY
10782|KING COVE
10783|KING GEORGE
10784|KING HILL
10785|KING LAKE
10786|KING OF PRUSSIA
10787|KING SALMON
10788|KING WILLIAM
10789|KINGDOM CITY
10790|KINGFISHER
10791|KINGMAN
10792|KINGS
10793|KINGS BEACH
10794|KINGS CANYON
10795|KINGS GRANT
10796|KINGS MILLS
10797|KINGS MOUNTAIN
10798|KINGS PARK
10799|KINGS POINT
10800|KINGS VALLEY
10801|KINGSBURG
10802|KINGSBURY
10803|KINGSDALE
10804|KINGSDOWN
10805|KINGSFORD
10806|KINGSFORD HEIGHTS
10807|KINGSLAND
10808|KINGSLEY
10809|KINGSMILL
10810|KINGSPORT
10811|KINGSTON
10812|KINGSTON ESTATES
10813|KINGSTON MINES
10814|KINGSTON SPRINGS
10815|KINGSTOWN
10816|KINGSTREE
10817|KINGSVILLE
10818|KINGVALE
10819|KINGWOOD
10820|KINLOCH
10821|KINMUNDY
10822|KINNEAR
10823|KINNELON
10824|KINNEY
10825|KINO SPRINGS
10826|KINROSS
10827|KINSALE
10828|KINSEY
10829|KINSLEY
10830|KINSMAN
10831|KINSTON
10832|KINTA
10833|KINTER
10834|KINTYRE
10835|KINWOOD
10836|KIOWA
10837|KIPLING
10838|KIPNUK
10839|KIPP
10840|KIPTON
10841|KIRBY
10842|KIRBYVILLE
10843|KIRE
10844|KIRK
10845|KIRKERSVILLE
10846|KIRKLAND
10847|KIRKLAND JUNCTION
10848|KIRKLIN
10849|KIRKMAN
10850|KIRKMANSVILLE
10851|KIRKPATRICK
10852|KIRKSEY
10853|KIRKSVILLE
10854|KIRKVILLE
10855|KIRKWOOD
10856|KIRLEY
10857|KIRON
10858|KIRTLAND
10859|KIRTLAND HILLS
10860|KIRVIN
10861|KIRWIN
10862|KIRYAS JOEL
10863|KISATCHIE
10864|KISKIMERE
10865|KISMET
10866|KISSEE MILLS
10867|KISSIMMEE
10868|KISTLER
10869|KIT CARSON
10870|KITALOU
10871|KITE
10872|KITSAP LAKE
10873|KITTANNING
10874|KITTERY
10875|KITTERY POINT
10876|KITTITAS
10877|KITTREDGE
10878|KITTRELL
10879|KITTS HILL
10880|KITTY HAWK
10881|KITZMILLER
10882|KIVALINA
10883|KIWALIK
10884|KLAGETOH
10885|KLAMATH
10886|KLAMATH AGENCY
10887|KLAMATH FALLS
10888|KLAMATH RIVER
10889|KLAWOCK
10890|KLEIN
10891|KLEMME
10892|KLICKITAT
10893|KLINE
10894|KLINGERSTOWN
10895|KLONDIKE
10896|KLOSSNER
10897|KLUKWAN
10898|KNAPP
10899|KNAPPA
10900|KNAUERTOWN
10901|KNEELAND
10902|KNIERIM
10903|KNIFE RIVER
10904|KNIFLEY
10905|KNIGHT
10906|KNIGHTDALE
10907|KNIGHTS
10908|KNIGHTS LANDING
10909|KNIGHTSEN
10910|KNIGHTSTOWN
10911|KNIGHTSVILLE
10912|KNIK
10913|KNIMAN
10914|KNIPPA
10915|KNOB LICK
10916|KNOB NOSTER
10917|KNOBEL
10918|KNOKE
10919|KNOLLS
10920|KNOLLWOOD
10921|KNOTTS ISLAND
10922|KNOWLES
10923|KNOWLTON
10924|KNOX
10925|KNOX CITY
10926|KNOXVILLE
10927|KO VAYA
10928|KOBUK
10929|KODIAK
10930|KOEHLER
10931|KOFA
10932|KOGGIUNG
10933|KOHATK
10934|KOHLER
10935|KOHLS RANCH
10936|KOHRVILLE
10937|KOKADJO
10938|KOKHANOK
10939|KOKOMO
10940|KOKRINES
10941|KOLEEN
10942|KOLIGANEK
10943|KOLIN
10944|KOLOLA SPRINGS
10945|KOMALTY
10946|KOMANDORSKI VILLAGE
10947|KOMATKE
10948|KONAWA
10949|KONGIGANAK
10950|KONNAROCK
10951|KOONTZ LAKE
10952|KOONTZVILLE
10953|KOOSHAREM
10954|KOOSKIA
10955|KOOTENAI
10956|KOPPEL
10957|KOPPERL
10958|KOPPERSTON
10959|KORBEL
10960|KORONA
10961|KOSCIUSKO
10962|KOSHKONONG
10963|KOSSE
10964|KOSSUTH
10965|KOSZTA
10966|KOTLIK
10967|KOTZEBUE
10968|KOUNTZE
10969|KOUTS
10970|KOYUK
10971|KOYUKUK
10972|KRAEMER
10973|KRAGNES
10974|KRAKOW
10975|KRAMER
10976|KRAMER JUNCTION
10977|KRANZBURG
10978|KRATZERVILLE
10979|KREAMER
10980|KREBS
10981|KREMLIN
10982|KREMMLING
10983|KREOLE
10984|KRESS
10985|KRESSON
10986|KRIDER
10987|KRONBORG
10988|KRONENWETTER
10989|KROTZ SPRINGS
10990|KRUGERVILLE
10991|KRUM
10992|KUALAPUʻU
10993|KUKUIHAELE
10994|KULM
10995|KULPMONT
10996|KULPSVILLE
10997|KUMMER
10998|KUNA
10999|KUNKLE
11000|KUNKLETOWN
11001|KUPREANOF
11002|KURE BEACH
11003|KURTEN
11004|KURTHWOOD
11005|KURTISTOWN
11006|KURTZ
11007|KUSTATAN
11008|KUTTAWA
11009|KUTZTOWN
11010|KVICHAK
11011|KWETHLUK
11012|KWIGILLINGOK
11013|KYBURZ
11014|KYKOTSMOVI VILLAGE
11015|KYLE
11016|KYLERTOWN
11017|KYSORVILLE
11018|KĀNEʻOHE
11019|KĀʻANAPALI
11020|KĒŌKEA
11021|KĪHEI
11022|KĪLAUEA
11023|KĪPAHULU
11024|KŌLOA
11025|L'ANSE
11026|LA ALIANZA
11027|LA ALIANZA COMUNIDAD
11028|LA BARGE
11029|LA BELLE
11030|LA BLANCA
11031|LA CASITA
11032|LA CAÑADA FLINTRIDGE
11033|LA CENTER
11034|LA CIENEGA
11035|LA CLEDE
11036|LA CONNER
11037|LA COSTE
11038|LA CRESCENT
11039|LA CRESCENTA
11040|LA CROFT
11041|LA CROSSE
11042|LA CUEVA
11043|LA CYGNE
11044|LA DOLORES
11045|LA DOLORES COMUNIDAD
11046|LA DUE
11047|LA FARGE
11048|LA FARGEVILLE
11049|LA FERIA
11050|LA FERMINA
11051|LA FERMINA COMUNIDAD
11052|LA FONTAINE
11053|LA GARITA
11054|LA GRANDE
11055|LA GRANGE
11056|LA GRANGE PARK
11057|LA GRULLA
11058|LA HABRA
11059|LA HABRA HEIGHTS
11060|LA HARPE
11061|LA HOMA
11062|LA HONDA
11063|LA HUERTA
11064|LA JARA
11065|LA JOYA
11066|LA JUNTA
11067|LA JUNTA GARDENS
11068|LA LIGA COMUNIDAD
11069|LA LUISA
11070|LA LUISA COMUNIDAD
11071|LA LUZ
11072|LA MADERA
11073|LA MARQUE
11074|LA MESA
11075|LA MESILLA
11076|LA MIRADA
11077|LA MOILLE
11078|LA MONTE
11079|LA MOTTE
11080|LA PALMA
11081|LA PALOMA
11082|LA PALOMA ADDITION COLONIA
11083|LA PARGUERA
11084|LA PARGUERA COMUNIDAD
11085|LA PAZ
11086|LA PAZ VALLEY
11087|LA PINE
11088|LA PLANT
11089|LA PLATA
11090|LA PLATTE
11091|LA PLAYA
11092|LA PLAYA COMUNIDAD
11093|LA PLENA
11094|LA PLENA COMUNIDAD
11095|LA PORTE
11096|LA PORTE CITY
11097|LA PRAIRIE
11098|LA PRESA
11099|LA PRYOR
11100|LA PUEBLA
11101|LA PUENTE
11102|LA PUERTA
11103|LA PUSH
11104|LA QUINTA
11105|LA REFORMA
11106|LA RIVIERA
11107|LA ROSE
11108|LA ROSITA
11109|LA RUE
11110|LA RUSSELL
11111|LA SAL
11112|LA SALLE
11113|LA SELVA BEACH
11114|LA TINA RANCH
11115|LA UNION
11116|LA VALE
11117|LA VALLE
11118|LA VERGNE
11119|LA VERNE
11120|LA VERNIA
11121|LA VETA
11122|LA VICTORIA
11123|LA VILLA
11124|LA VILLITA
11125|LA VINA
11126|LA VISTA
11127|LA WARD
11128|LA YUCA COMUNIDAD
11129|LABADIE
11130|LABADIEVILLE
11131|LABELLE
11132|LABETTE
11133|LABISH VILLAGE
11134|LABOLT
11135|LAC DU FLAMBEAU
11136|LAC LA BELLE
11137|LACASSINE
11138|LACEY
11139|LACEYVILLE
11140|LACHINE
11141|LACKAWANNA
11142|LACKEY
11143|LACKMANS
11144|LACLEDE
11145|LACOMB
11146|LACOMBE
11147|LACON
11148|LACONA
11149|LACONIA
11150|LACOOCHEE
11151|LACY-LAKEVIEW
11152|LADD
11153|LADDONIA
11154|LADELLE
11155|LADENTOWN
11156|LADERA
11157|LADERA HEIGHTS
11158|LADERA RANCH
11159|LADNER
11160|LADOGA
11161|LADONIA
11162|LADORA
11163|LADSON
11164|LADUE
11165|LADY LAKE
11166|LADYSMITH
11167|LAFAYETTE
11168|LAFE
11169|LAFFERTY
11170|LAFITTE
11171|LAFLIN
11172|LAFOLLETTE
11173|LAFONTAINE
11174|LAFOURCHE
11175|LAGO
11176|LAGO VISTA
11177|LAGRANGE
11178|LAGRO
11179|LAGUNA
11180|LAGUNA BEACH
11181|LAGUNA HEIGHTS
11182|LAGUNA HILLS
11183|LAGUNA NIGUEL
11184|LAGUNA PARK
11185|LAGUNA SECA
11186|LAGUNA VISTA
11187|LAGUNA WOODS
11188|LAGUNITAS
11189|LAHAINA
11190|LAHOMA
11191|LAINGSBURG
11192|LAIR
11193|LAIRD
11194|LAIRD HILL
11195|LAJAS
11196|LAJAS ZONA URBANA
11197|LAJITAS
11198|LAKE
11199|LAKE ALFRED
11200|LAKE ALMANOR COUNTRY CLUB
11201|LAKE ALMANOR PENINSULA
11202|LAKE ALMANOR WEST
11203|LAKE ALUMA
11204|LAKE ANDES
11205|LAKE ANGELUS
11206|LAKE ANN
11207|LAKE ANNETTE
11208|LAKE ARBOR
11209|LAKE ARIEL
11210|LAKE ARROWHEAD
11211|LAKE ARTHUR
11212|LAKE ARTHUR ESTATES
11213|LAKE BARCROFT
11214|LAKE BARRINGTON
11215|LAKE BELVEDERE ESTATES
11216|LAKE BENTON
11217|LAKE BEULAH
11218|LAKE BLUFF
11219|LAKE BOSWORTH
11220|LAKE BRIDGEPORT
11221|LAKE BRONSON
11222|LAKE BROWNWOOD
11223|LAKE BUENA VISTA
11224|LAKE BUTLER
11225|LAKE CAMELOT
11226|LAKE CARMEL
11227|LAKE CATHERINE
11228|LAKE CAVANAUGH
11229|LAKE CHARLES
11230|LAKE CITY
11231|LAKE CLARKE SHORES
11232|LAKE CLEAR
11233|LAKE COMO
11234|LAKE CREEK
11235|LAKE CRYSTAL
11236|LAKE DALECARLIA
11237|LAKE DALLAS
11238|LAKE DARBY
11239|LAKE DAVIS
11240|LAKE DELTON
11241|LAKE DUNLAP
11242|LAKE ELMO
11243|LAKE ELSINORE
11244|LAKE END
11245|LAKE ERIE BEACH
11246|LAKE FENTON
11247|LAKE FIVE
11248|LAKE FOREST
11249|LAKE FOREST PARK
11250|LAKE FORK
11251|LAKE GENEVA
11252|LAKE GEORGE
11253|LAKE GOODWIN
11254|LAKE GROVE
11255|LAKE HALLIE
11256|LAKE HAMILTON
11257|LAKE HARBOR
11258|LAKE HART
11259|LAKE HAVASU CITY
11260|LAKE HELEN
11261|LAKE HENRY
11262|LAKE HERITAGE
11263|LAKE HIAWATHA
11264|LAKE HILLS
11265|LAKE HOLIDAY
11266|LAKE HUGHES
11267|LAKE IN THE HILLS
11268|LAKE ISABELLA
11269|LAKE ITASCA
11270|LAKE JACKSON
11271|LAKE JUNALUSKA
11272|LAKE KA-HO
11273|LAKE KATHRYN
11274|LAKE KATRINE
11275|LAKE KETCHUM
11276|LAKE KIOWA
11277|LAKE KOSHKONONG
11278|LAKE LAFAYETTE
11279|LAKE LAKENGREN
11280|LAKE LATONKA
11281|LAKE LEELANAU
11282|LAKE LILLIAN
11283|LAKE LINDEN
11284|LAKE LINDSEY
11285|LAKE LORRAINE
11286|LAKE LOS ANGELES
11287|LAKE LOTAWANA
11288|LAKE LOUISE
11289|LAKE LURE
11290|LAKE LUZERNE
11291|LAKE MAGDALENE
11292|LAKE MARY
11293|LAKE MARY RONAN
11294|LAKE MCDONALD
11295|LAKE MCMURRAY
11296|LAKE MEADE
11297|LAKE MICHIGAN BEACH
11298|LAKE MILLS
11299|LAKE MILTON
11300|LAKE MINCHUMINA
11301|LAKE MOHAWK
11302|LAKE MOHEGAN
11303|LAKE MONROE
11304|LAKE MONTEZUMA
11305|LAKE MONTICELLO
11306|LAKE MYKEE TOWN
11307|LAKE NACIMIENTO
11308|LAKE NEBAGAMON
11309|LAKE NORDEN
11310|LAKE ODESSA
11311|LAKE OF THE PINES
11312|LAKE OF THE WOODS
11313|LAKE ORION
11314|LAKE OSWEGO
11315|LAKE OZARK
11316|LAKE PANASOFFKEE
11317|LAKE PANORAMA
11318|LAKE PARK
11319|LAKE PETERSBURG
11320|LAKE PINE
11321|LAKE PLACID
11322|LAKE POCOTOPAUG
11323|LAKE PRESTON
11324|LAKE PROVIDENCE
11325|LAKE QUIVIRA
11326|LAKE RIDGE
11327|LAKE RIPLEY
11328|LAKE ROESIGER
11329|LAKE RONKONKOMA
11330|LAKE SAINT CROIX BEACH
11331|LAKE SAINT LOUIS
11332|LAKE SAN MARCOS
11333|LAKE SANTEETLAH
11334|LAKE SARASOTA
11335|LAKE SECESSION
11336|LAKE SENECA
11337|LAKE SHANGRILA
11338|LAKE SHORE
11339|LAKE SPRING
11340|LAKE STATION
11341|LAKE STEVENS
11342|LAKE STICKNEY
11343|LAKE SUCCESS
11344|LAKE SUMMERSET
11345|LAKE SUMNER
11346|LAKE TANGLEWOOD
11347|LAKE TANSI
11348|LAKE TAPAWINGO
11349|LAKE TELEMARK
11350|LAKE TOMAHAWK
11351|LAKE TOXAWAY
11352|LAKE VALLEY
11353|LAKE VIEW
11354|LAKE VILLA
11355|LAKE VILLAGE
11356|LAKE WACCAMAW
11357|LAKE WALES
11358|LAKE WAUKOMIS
11359|LAKE WAZEECHA
11360|LAKE WILDWOOD
11361|LAKE WILSON
11362|LAKE WINNEBAGO
11363|LAKE WINOLA
11364|LAKE WISCONSIN
11365|LAKE WISSOTA
11366|LAKE WORTH
11367|LAKE WYLIE
11368|LAKE WYNONAH
11369|LAKE ZURICH
11370|LAKEBAY
11371|LAKEFIELD
11372|LAKEHEAD
11373|LAKEHILLS
11374|LAKEHURST
11375|LAKELAND
11376|LAKELAND HEIGHTS
11377|LAKELAND HIGHLANDS
11378|LAKELAND SHORES
11379|LAKELAND VILLAGE
11380|LAKELINE
11381|LAKEMONT
11382|LAKEMOOR
11383|LAKEMORE
11384|LAKEPORT
11385|LAKERIDGE
11386|LAKES OF THE FOUR SEASONS
11387|LAKESHIRE
11388|LAKESHORE
11389|LAKESIDE
11390|LAKESIDE CITY
11391|LAKESIDE PARK
11392|LAKESITE
11393|LAKETON
11394|LAKETOWN
11395|LAKEVIEW
11396|LAKEVIEW ESTATES
11397|LAKEVIEW HEIGHTS
11398|LAKEVILLE
11399|LAKEWAY
11400|LAKEWOOD
11401|LAKEWOOD CLUB
11402|LAKEWOOD HEIGHTS
11403|LAKEWOOD PARK
11404|LAKEWOOD SHORES
11405|LAKEWOOD VILLAGE
11406|LAKIN
11407|LAKOTA
11408|LAMAR
11409|LAMAR HEIGHTS
11410|LAMASCO
11411|LAMBERT
11412|LAMBERTON
11413|LAMBERTVILLE
11414|LAMBOGLIA
11415|LAMBOGLIA COMUNIDAD
11416|LAMBROOK
11417|LAMBS GROVE
11418|LAME DEER
11419|LAMESA
11420|LAMINE
11421|LAMINGTON
11422|LAMISON
11423|LAMKIN
11424|LAMOILLE
11425|LAMOINE
11426|LAMONA
11427|LAMONI
11428|LAMONT
11429|LAMOURE
11430|LAMOURIE
11431|LAMPASAS
11432|LAMPETER
11433|LAMPSON
11434|LAMY
11435|LANAGAN
11436|LANARE
11437|LANARK
11438|LANARK VILLAGE
11439|LANCASTER
11440|LANCE CREEK
11441|LANCING
11442|LAND
11443|LAND O' LAKES
11444|LAND OF PINES
11445|LANDA
11446|LANDEN
11447|LANDENBERG
11448|LANDER
11449|LANDERSVILLE
11450|LANDESS
11451|LANDFALL
11452|LANDING
11453|LANDINGVILLE
11454|LANDIS
11455|LANDISBURG
11456|LANDISVILLE
11457|LANDMARK
11458|LANDO
11459|LANDOVER
11460|LANDOVER HILLS
11461|LANDRUM
11462|LANDUSKY
11463|LANE
11464|LANE CITY
11465|LANEBURG
11466|LANESBORO
11467|LANESVILLE
11468|LANETT
11469|LANEVILLE
11470|LANGDON
11471|LANGDON PLACE
11472|LANGELOTH
11473|LANGES CORNERS
11474|LANGFORD
11475|LANGHORNE
11476|LANGHORNE MANOR
11477|LANGLEY
11478|LANGLEY PARK
11479|LANGLEYVILLE
11480|LANGLOIS
11481|LANGSTON
11482|LANGTRY
11483|LANGWORTHY
11484|LANHAM
11485|LANKIN
11486|LANNON
11487|LANSDALE
11488|LANSDOWNE
11489|LANSFORD
11490|LANSING
11491|LANTANA
11492|LANTON
11493|LANTRY
11494|LANYON
11495|LAONA
11496|LAOTTO
11497|LAPEER
11498|LAPEL
11499|LAPLACE
11500|LAPOINT
11501|LAPORTE
11502|LAPWAI
11503|LARAMIE
11504|LARCHMONT
11505|LARCHWOOD
11506|LAREDO
11507|LAREDO RANCHETTES
11508|LARES
11509|LARES ZONA URBANA
11510|LARGO
11511|LARIAT
11512|LARIMER
11513|LARIMERS CORNER
11514|LARIMORE
11515|LARK
11516|LARKSPUR
11517|LARKSVILLE
11518|LARNED
11519|LAROSE
11520|LARRABEE
11521|LARSEN
11522|LARSEN BAY
11523|LARSLAN
11524|LARSMONT
11525|LARSON
11526|LARTO
11527|LARUE
11528|LARWILL
11529|LAS ANIMAS
11530|LAS CAROLINAS
11531|LAS CAROLINAS COMUNIDAD
11532|LAS CROABAS
11533|LAS CROABAS COMUNIDAD
11534|LAS CRUCES
11535|LAS FLORES
11536|LAS LOMAS
11537|LAS LOMITAS
11538|LAS MARAVILLAS
11539|LAS MARIAS
11540|LAS MARÍAS COMUNIDAD
11541|LAS MARÍAS ZONA URBANA
11542|LAS NUTRIAS
11543|LAS OCHENTA
11544|LAS OCHENTA COMUNIDAD
11545|LAS OLLAS
11546|LAS OLLAS COMUNIDAD
11547|LAS PALMAS
11548|LAS PALOMAS
11549|LAS PIEDRAS
11550|LAS PIEDRAS ZONA URBANA
11551|LAS QUINTAS FRONTERIZAS
11552|LAS QUINTAS FRONTERIZAS COLONIA
11553|LAS VEGAS
11554|LASANA
11555|LASARA
11556|LASHMEET
11557|LASKER
11558|LASSATER
11559|LAST CHANCE
11560|LASTRUP
11561|LATAH
11562|LATEXO
11563|LATHAM
11564|LATHAM PARK
11565|LATHROP
11566|LATHRUP VILLAGE
11567|LATIMER
11568|LATON
11569|LATOUR
11570|LATROBE
11571|LATTA
11572|LATTASBURG
11573|LATTIMER
11574|LATTIMORE
11575|LATTINGTOWN
11576|LATTY
11577|LAUADA
11578|LAUD
11579|LAUDERDALE
11580|LAUDERDALE LAKES
11581|LAUDERDALE-BY-THE-SEA
11582|LAUDERHILL
11583|LAUGHLIN
11584|LAUNIUPOKO
11585|LAUPĀHOEHOE
11586|LAURA
11587|LAUREL
11588|LAUREL BAY
11589|LAUREL GARDENS
11590|LAUREL GROVE
11591|LAUREL HILL
11592|LAUREL HOLLOW
11593|LAUREL LAKE
11594|LAUREL MOUNTAIN PARK
11595|LAUREL PARK
11596|LAUREL RUN
11597|LAUREL SPRINGS
11598|LAURELDALE
11599|LAURELES
11600|LAURELTON
11601|LAURELVILLE
11602|LAURENCE HARBOR
11603|LAURENS
11604|LAURIE
11605|LAURIER
11606|LAURINBURG
11607|LAURIUM
11608|LAURYS STATION
11609|LAUTZ
11610|LAVA HOT SPRINGS
11611|LAVACA
11612|LAVALETTE
11613|LAVALLETTE
11614|LAVEEN
11615|LAVELLE
11616|LAVERKIN
11617|LAVERNE
11618|LAVINA
11619|LAVINIA
11620|LAVON
11621|LAVONIA
11622|LAWEN
11623|LAWLER
11624|LAWLEY
11625|LAWN
11626|LAWNDALE
11627|LAWNSIDE
11628|LAWNTON
11629|LAWRENCE
11630|LAWRENCE CREEK
11631|LAWRENCE PARK
11632|LAWRENCEBURG
11633|LAWRENCEVILLE
11634|LAWS
11635|LAWSON
11636|LAWSON HEIGHTS
11637|LAWSONIA
11638|LAWTELL
11639|LAWTEY
11640|LAWTON
11641|LAXON
11642|LAY
11643|LAYHIGH
11644|LAYHILL
11645|LAYMANTOWN
11646|LAYTON
11647|LAYTONSVILLE
11648|LAYTONVILLE
11649|LAZARE
11650|LAZEAR
11651|LAZY ACRES
11652|LAZY LAKE
11653|LAZY MOUNTAIN
11654|LE CENTER
11655|LE CLAIRE
11656|LE GRAND
11657|LE LOUP
11658|LE MARS
11659|LE MOYEN
11660|LE RAYSVILLE
11661|LE ROY
11662|LE SOURDSVILLE
11663|LE SUEUR
11664|LEABURG
11665|LEACH
11666|LEACHVILLE
11667|LEACOCK
11668|LEAD HILL
11669|LEADER
11670|LEADINGTON
11671|LEADORE
11672|LEADPOINT
11673|LEADVILLE
11674|LEADWOOD
11675|LEAF RIVER
11676|LEAGUE CITY
11677|LEAKESVILLE
11678|LEAKEY
11679|LEAL
11680|LEALMAN
11681|LEAMINGTON
11682|LEANDER
11683|LEANDO
11684|LEARY
11685|LEASBURG
11686|LEATHERSVILLE
11687|LEATHERWOOD
11688|LEAVENWORTH
11689|LEAVITTSBURG
11690|LEAWOOD
11691|LEBAM
11692|LEBANON
11693|LEBANON CHURCH
11694|LEBANON JUNCTION
11695|LEBEAU
11696|LEBEC
11697|LEBO
11698|LECANTO
11699|LECHEE
11700|LECOMPTE
11701|LECOMPTON
11702|LEDBETTER
11703|LEDFORD
11704|LEDGER
11705|LEDGEWOOD
11706|LEDOUX
11707|LEDYARD
11708|LEE ACRES
11709|LEE BAYOU
11710|LEE CENTER
11711|LEE CITY
11712|LEE CREEK
11713|LEE MONT
11714|LEE VINING
11715|LEECHBURG
11716|LEEDEY
11717|LEEDS
11718|LEEDY
11719|LEEPER
11720|LEES CAMP
11721|LEES SUMMIT
11722|LEESBURG
11723|LEESPORT
11724|LEESVILLE
11725|LEETON
11726|LEETONIA
11727|LEETSDALE
11728|LEEVILLE
11729|LEEWOOD
11730|LEFLORE
11731|LEFOR
11732|LEFORS
11733|LEGEND LAKE
11734|LEGGETT
11735|LEHI
11736|LEHIGH
11737|LEHIGH ACRES
11738|LEHIGHTON
11739|LEHMAN
11740|LEHR
11741|LEICESTER
11742|LEIGH
11743|LEIGHTON
11744|LEILANI ESTATES
11745|LEIPERS FORK
11746|LEIPSIC
11747|LEISURE CITY
11748|LEISURE KNOLL
11749|LEISURE VILLAGE
11750|LEISURE VILLAGE EAST
11751|LEISURE VILLAGE WEST
11752|LEISURETOWNE
11753|LEITCH
11754|LEITCHFIELD
11755|LEITER
11756|LEITERSBURG
11757|LEITH
11758|LELA
11759|LELAND
11760|LELAND GROVE
11761|LELIA LAKE
11762|LELY
11763|LELY RESORT
11764|LEMANNVILLE
11765|LEMAY
11766|LEMETA
11767|LEMHI
11768|LEMING
11769|LEMITAR
11770|LEMMON
11771|LEMMON VALLEY
11772|LEMON GROVE
11773|LEMON HEIGHTS
11774|LEMONCOVE
11775|LEMONT
11776|LEMONT FURNACE
11777|LEMOORE
11778|LEMOYNE
11779|LENAPAH
11780|LENAPE
11781|LENAPE HEIGHTS
11782|LENEXA
11783|LENGBY
11784|LENHARTSVILLE
11785|LENKERVILLE
11786|LENNEP
11787|LENNON
11788|LENNOX
11789|LENOIR
11790|LENOIR CITY
11791|LENOLA
11792|LENORA
11793|LENORAH
11794|LENORE
11795|LENOX
11796|LENOXBURG
11797|LENWOOD
11798|LENZ
11799|LENZBURG
11800|LEO-CEDARVILLE
11801|LEOLA
11802|LEOMA
11803|LEOMINSTER
11804|LEON
11805|LEON JUNCTION
11806|LEON VALLEY
11807|LEONA
11808|LEONA VALLEY
11809|LEONARD
11810|LEONARDO
11811|LEONARDSVILLE
11812|LEONARDTOWN
11813|LEONARDVILLE
11814|LEONIA
11815|LEONIDAS
11816|LEONORE
11817|LEONVILLE
11818|LEOPOLD
11819|LEOPOLIS
11820|LEOTA
11821|LEOTI
11822|LEOVILLE
11823|LEPANTO
11824|LEQUIRE
11825|LERNA
11826|LERNERVILLE
11827|LEROY
11828|LESAGE
11829|LESHARA
11830|LESLEY
11831|LESLIE
11832|LESSLEY
11833|LESSLIE
11834|LESTER
11835|LESTER PRAIRIE
11836|LESTERVILLE
11837|LETART FALLS
11838|LETCHER
11839|LETHA
11840|LETOHATCHEE
11841|LETONA
11842|LETTS
11843|LETTSWORTH
11844|LEUCADIA
11845|LEUPP
11846|LEUPP CORNER
11847|LEVAN
11848|LEVANT
11849|LEVASY
11850|LEVEL GREEN
11851|LEVEL PARK
11852|LEVEL PLAINS
11853|LEVELLAND
11854|LEVELOCK
11855|LEVERING
11856|LEVITTOWN
11857|LEVITTOWN COMUNIDAD
11858|LEVY
11859|LEWELLEN
11860|LEWES
11861|LEWIS
11862|LEWIS AND CLARK VILLAGE
11863|LEWIS CENTER
11864|LEWIS RUN
11865|LEWIS SPRINGS
11866|LEWISBERRY
11867|LEWISBURG
11868|LEWISETTA
11869|LEWISPORT
11870|LEWISTON
11871|LEWISTON ORCHARDS
11872|LEWISTON WOODVILLE
11873|LEWISTOWN
11874|LEWISTOWN HEIGHTS
11875|LEWISVILLE
11876|LEXA
11877|LEXIE
11878|LEXINGTON
11879|LEXINGTON HEIGHTS
11880|LEXINGTON HILLS
11881|LEXINGTON PARK
11882|LEYDEN
11883|LEYNER
11884|LIBBY
11885|LIBBYVILLE
11886|LIBERTY CENTER
11887|LIBERTY CITY
11888|LIBERTY CORNER
11889|LIBERTY GROVE
11890|LIBERTY HILL
11891|LIBERTY LAKE
11892|LIBERTY PARK
11893|LIBERTY PLAIN
11894|LIBERTY POLE
11895|LIBERTYTOWN
11896|LIBERTYVILLE
11897|LIBORIO NEGRON TORRES
11898|LIBORIO NEGRÓN TORRES COMUNIDAD
11899|LIBUSE
11900|LICKING
11901|LIDA
11902|LIDDERDALE
11903|LIDDIEVILLE
11904|LIDGERWOOD
11905|LIDO BEACH
11906|LIEBENTHAL
11907|LIGHT OAK
11908|LIGHT STREET
11909|LIGHTHOUSE POINT
11910|LIGNITE
11911|LIGNUM
11912|LIGON
11913|LIGONIER
11914|LIGURTA
11915|LIKELY
11916|LILBERT
11917|LILBOURN
11918|LILBURN
11919|LILESVILLE
11920|LILITA
11921|LILLE
11922|LILLIAN
11923|LILLIE
11924|LILLINGTON
11925|LILLIWAUP
11926|LILLY
11927|LILY
11928|LILY CACHE
11929|LILY LAKE
11930|LILYDALE
11931|LILYMOOR
11932|LIM ROCK
11933|LIMA
11934|LIMAVILLE
11935|LIME CITY
11936|LIME CREEK
11937|LIME LAKE
11938|LIME RIDGE
11939|LIME SPRINGS
11940|LIME VILLAGE
11941|LIMERICK
11942|LIMESTONE
11943|LIMESTONE CREEK
11944|LIMON
11945|LINBY
11946|LINCH
11947|LINCOLN
11948|LINCOLN ACRES
11949|LINCOLN BEACH
11950|LINCOLN CITY
11951|LINCOLN ESTATES
11952|LINCOLN HEIGHTS
11953|LINCOLN HILLS
11954|LINCOLN PARK
11955|LINCOLN VILLAGE
11956|LINCOLNDALE
11957|LINCOLNIA
11958|LINCOLNSHIRE
11959|LINCOLNTON
11960|LINCOLNVILLE
11961|LINCOLNWOOD
11962|LINCROFT
11963|LIND
11964|LINDA
11965|LINDALE
11966|LINDBERG
11967|LINDCOVE
11968|LINDEN
11969|LINDENAU
11970|LINDENHURST
11971|LINDENWOLD
11972|LINDENWOOD
11973|LINDISFARNE
11974|LINDON
11975|LINDSAY
11976|LINDSBORG
11977|LINDSEY
11978|LINDSEYVILLE
11979|LINDSIDE
11980|LINDSTROM
11981|LINDY
11982|LINESVILLE
11983|LINEVILLE
11984|LINFIELD
11985|LINGANORE
11986|LINGLE
11987|LINGLESTOWN
11988|LINN
11989|LINN CREEK
11990|LINN GROVE
11991|LINN VALLEY
11992|LINNDALE
11993|LINNEUS
11994|LINNTOWN
11995|LINO LAKES
11996|LINTHICUM
11997|LINTON
11998|LINTON HALL
11999|LINVILLE
12000|LINWOOD
12001|LIONVILLE
12002|LIPAN
12003|LIPSCOMB
12004|LISABEULA
12005|LISBON
12006|LISBON FALLS
12007|LISCO
12008|LISCOMB
12009|LISLE
12010|LISMAN
12011|LISMORE
12012|LISSIE
12013|LITCHFIELD
12014|LITCHFIELD PARK
12015|LITCHVILLE
12016|LITERBERRY
12017|LITHIA SPRINGS
12018|LITHIUM
12019|LITHONIA
12020|LITHOPOLIS
12021|LITITZ
12022|LITROE
12023|LITTIG
12024|LITTLE AMERICA
12025|LITTLE BRITAIN
12026|LITTLE CANADA
12027|LITTLE CEDAR
12028|LITTLE CHUTE
12029|LITTLE CREEK
12030|LITTLE CYPRESS
12031|LITTLE EAGLE
12032|LITTLE ELM
12033|LITTLE FALLS
12034|LITTLE FERRY
12035|LITTLE FLOCK
12036|LITTLE GRASS VALLEY
12037|LITTLE HOCKING
12038|LITTLE LAKE
12039|LITTLE MARAIS
12040|LITTLE MEADOWS
12041|LITTLE MOUNTAIN
12042|LITTLE ORLEANS
12043|LITTLE RAPIDS
12044|LITTLE RIVER
12045|LITTLE RIVER-ACADEMY
12046|LITTLE ROCK
12047|LITTLE ROUND LAKE
12048|LITTLE SAUK
12049|LITTLE SILVER
12050|LITTLE SIOUX
12051|LITTLE STURGEON
12052|LITTLE VALLEY
12053|LITTLE YORK
12054|LITTLEFIELD
12055|LITTLEFORK
12056|LITTLEJOHN ISLAND
12057|LITTLEPORT
12058|LITTLEROCK
12059|LITTLESTOWN
12060|LITTLETON
12061|LITTLETON COMMON
12062|LITTLETOWN
12063|LITTLEVILLE
12064|LIVE OAK
12065|LIVE OAK SPRINGS
12066|LIVELY
12067|LIVENGOOD
12068|LIVERMORE
12069|LIVERMORE FALLS
12070|LIVERPOOL
12071|LIVIA
12072|LIVINGSTON
12073|LIVINGSTON MANOR
12074|LIVONA
12075|LIVONIA
12076|LIVONIA CENTER
12077|LIZELLA
12078|LIZEMORES
12079|LIZTON
12080|LLANO
12081|LLANO DEL MEDIO
12082|LLANO GRANDE
12083|LLOYD
12084|LLOYD HARBOR
12085|LLOYDELL
12086|LLUVERAS
12087|LLUVERAS COMUNIDAD
12088|LOA
12089|LOACHAPOKA
12090|LOAG
12091|LOAMI
12092|LOBECO
12093|LOBELVILLE
12094|LOBO
12095|LOCH ARBOUR
12096|LOCH LLOYD
12097|LOCH LOMOND
12098|LOCH LYNN HEIGHTS
12099|LOCH SHELDRAKE
12100|LOCHBUIE
12101|LOCHEARN
12102|LOCHIEL
12103|LOCHLOOSA
12104|LOCHMOOR WATERWAY ESTATES
12105|LOCHSLOY
12106|LOCK HAVEN
12107|LOCK SPRINGS
12108|LOCKBOURNE
12109|LOCKEFORD
12110|LOCKESBURG
12111|LOCKETT
12112|LOCKHART
12113|LOCKINGTON
12114|LOCKLAND
12115|LOCKNEY
12116|LOCKPORT
12117|LOCKPORT HEIGHTS
12118|LOCKRIDGE
12119|LOCKWOOD
12120|LOCO
12121|LOCO HILLS
12122|LOCUST
12123|LOCUST CORNER
12124|LOCUST FORK
12125|LOCUST GROVE
12126|LOCUST LAKE
12127|LOCUST VALLEY
12128|LOCUSTDALE
12129|LODA
12130|LODGE
12131|LODGE GRASS
12132|LODGE POLE
12133|LODGEPOLE
12134|LODI
12135|LODOGA
12136|LOEB
12137|LOFALL
12138|LOFGREEN
12139|LOG CABIN
12140|LOG LANE VILLAGE
12141|LOGAN
12142|LOGAN ELM VILLAGE
12143|LOGANDALE
12144|LOGANSPORT
12145|LOGANTON
12146|LOGANVILLE
12147|LOGHILL VILLAGE
12148|LOGSDEN
12149|LOHMAN
12150|LOHRVILLE
12151|LOLA
12152|LOLETA
12153|LOLITA
12154|LOLO
12155|LOLO HOT SPRINGS
12156|LOMA
12157|LOMA ALTA
12158|LOMA GRANDE COLONIA
12159|LOMA LINDA
12160|LOMA LINDA COLONIA
12161|LOMA LINDA EAST COLONIA
12162|LOMA MAR
12163|LOMA RICA
12164|LOMA VISTA COLONIA
12165|LOMAN
12166|LOMAS
12167|LOMAS COMUNIDAD
12168|LOMAX
12169|LOMBARD
12170|LOMETA
12171|LOMIRA
12172|LOMITA
12173|LOMPICO
12174|LOMPOC
12175|LONACONING
12176|LONDON
12177|LONDON MILLS
12178|LONDONDERRY
12179|LONE ELM
12180|LONE GROVE
12181|LONE JACK
12182|LONE MOUNTAIN
12183|LONE OAK
12184|LONE PINE
12185|LONE ROCK
12186|LONE STAR
12187|LONE TREE
12188|LONE WOLF
12189|LONEDELL
12190|LONELYVILLE
12191|LONEPINE
12192|LONEROCK
12193|LONETREE
12194|LONG BARN
12195|LONG BEACH
12196|LONG BRANCH
12197|LONG BRIDGE
12198|LONG CREEK
12199|LONG GROVE
12200|LONG HILL
12201|LONG ISLAND
12202|LONG LAKE
12203|LONG MEADOW
12204|LONG MOTT
12205|LONG NECK
12206|LONG PINE
12207|LONG POINT
12208|LONG POND
12209|LONG PRAIRIE
12210|LONG RIDGE
12211|LONG VALLEY
12212|LONGBOAT KEY
12213|LONGBRANCH
12214|LONGDALE
12215|LONGFELLOW
12216|LONGFORD
12217|LONGHURST
12218|LONGMEADOW
12219|LONGMIRE
12220|LONGMONT
12221|LONGPORT
12222|LONGRUN
12223|LONGS
12224|LONGSTREET
12225|LONGTON
12226|LONGTOWN
12227|LONGVIEW
12228|LONGVIEW HEIGHTS
12229|LONGVILLE
12230|LONGWOOD
12231|LONGWOODS
12232|LONGWORTH
12233|LONO
12234|LONOKE
12235|LONSDALE
12236|LOOGOOTEE
12237|LOOKEBA
12238|LOOKINGGLASS
12239|LOOKOUT
12240|LOOKOUT MOUNTAIN
12241|LOOMIS
12242|LOON LAKE
12243|LOOSE CREEK
12244|LOPEZVILLE
12245|LOPEÑO
12246|LORAIN
12247|LORAINE
12248|LORANE
12249|LORANGER
12250|LORD
12251|LORDSBURG
12252|LORDSTOWN
12253|LORE CITY
12254|LOREAUVILLE
12255|LORENA
12256|LORENTZ
12257|LORENZ PARK
12258|LORENZO
12259|LORETTA
12260|LORETTO
12261|LORIDA
12262|LORIMOR
12263|LORING
12264|LORIS
12265|LORMAN
12266|LORRAINE
12267|LORTON
12268|LOS ALAMITOS
12269|LOS ALAMOS
12270|LOS ALTOS
12271|LOS ALTOS COLONIA
12272|LOS ALTOS HILLS
12273|LOS ALVAREZ
12274|LOS ANGELES
12275|LOS BANOS
12276|LOS BARRERAS
12277|LOS BERROS
12278|LOS CHAVEZ
12279|LOS EBANOS
12280|LOS EBANOS COLONIA
12281|LOS FRESNOS
12282|LOS GATOS
12283|LOS INDIOS
12284|LOS LLANOS
12285|LOS LLANOS COMUNIDAD
12286|LOS LUCEROS
12287|LOS LUNAS
12288|LOS MEDANOS
12289|LOS MOLINOS
12290|LOS NIETOS
12291|LOS OJOS
12292|LOS OLIVOS
12293|LOS OSOS
12294|LOS PADILLAS
12295|LOS PANES COMUNIDAD
12296|LOS PINOS
12297|LOS PRADOS COMUNIDAD
12298|LOS RANCHOS DE ALBUQUERQUE
12299|LOS SERRANOS
12300|LOS TRANCOS WOODS
12301|LOS TRUJILLOS
12302|LOS VILLAREALES
12303|LOS YBANEZ
12304|LOSANTVILLE
12305|LOST BRIDGE VILLAGE
12306|LOST CABIN
12307|LOST CITY
12308|LOST CREEK
12309|LOST HILLS
12310|LOST LAKE WOODS
12311|LOST NATION
12312|LOST RIVER
12313|LOST SPRINGS
12314|LOSTANT
12315|LOSTINE
12316|LOSTWOOD
12317|LOTHAIR
12318|LOTSEE
12319|LOTT
12320|LOTTAVILLE
12321|LOTUS WOODS
12322|LOUANN
12323|LOUDON
12324|LOUDONVILLE
12325|LOUGHMAN
12326|LOUIN
12327|LOUISA
12328|LOUISBURG
12329|LOUISE
12330|LOUISIANA
12331|LOUISVILLE
12332|LOUP CITY
12333|LOURDES
12334|LOUVALE
12335|LOUVIERS
12336|LOVE VALLEY
12337|LOVEJOY
12338|LOVELACEVILLE
12339|LOVELADY
12340|LOVELAND
12341|LOVELAND PARK
12342|LOVELL
12343|LOVELLS
12344|LOVELOCK
12345|LOVES PARK
12346|LOVETT
12347|LOVETTSVILLE
12348|LOVEWELL
12349|LOVILIA
12350|LOVING
12351|LOVINGSTON
12352|LOVINGTON
12353|LOW MOOR
12354|LOW MOUNTAIN
12355|LOWDEN
12356|LOWELL
12357|LOWELL POINT
12358|LOWELLTOWN
12359|LOWELLVILLE
12360|LOWEMONT
12361|LOWER ALLEN
12362|LOWER BRULE
12363|LOWER BURRELL
12364|LOWER GRAND LAGOON
12365|LOWER KALSKAG
12366|LOWER LAKE
12367|LOWER MARLBORO
12368|LOWER SALEM
12369|LOWER SQUANKUM
12370|LOWER TONSINA
12371|LOWES
12372|LOWES ISLAND
12373|LOWESVILLE
12374|LOWGAP
12375|LOWLAND
12376|LOWMAN
12377|LOWNDESBORO
12378|LOWNDESVILLE
12379|LOWRY
12380|LOWRY CITY
12381|LOWRY CROSSING
12382|LOWRYS
12383|LOWSVILLE
12384|LOWVILLE
12385|LOXA
12386|LOXAHATCHEE
12387|LOXAHATCHEE GROVES
12388|LOXLEY
12389|LOYAL
12390|LOYAL VALLEY
12391|LOYALHANNA
12392|LOYALL
12393|LOYALTON
12394|LOYD
12395|LOYOLA
12396|LOYSBURG
12397|LOYSVILLE
12398|LOZANO
12399|LOZEAU
12400|LOÍZA
12401|LOÍZA ZONA URBANA
12402|LU VERNE
12403|LUANA
12404|LUBBOCK
12405|LUBEC
12406|LUBECK
12407|LUBLIN
12408|LUCAMA
12409|LUCAN
12410|LUCAS
12411|LUCAS VALLEY
12412|LUCASVILLE
12413|LUCCA
12414|LUCE
12415|LUCEDALE
12416|LUCERNE
12417|LUCERNE MINES
12418|LUCERNE VALLEY
12419|LUCERO
12420|LUCIEN
12421|LUCILE
12422|LUCIN
12423|LUCINDA
12424|LUCK
12425|LUCKEY
12426|LUCKY
12427|LUCY
12428|LUDDEN
12429|LUDELL
12430|LUDINGTON
12431|LUDLAM
12432|LUDLOW
12433|LUDLOW FALLS
12434|LUDLOWVILLE
12435|LUDOWICI
12436|LUDWIGS CORNER
12437|LUEDERS
12438|LUELLA
12439|LUFKIN
12440|LUGERT
12441|LUGOFF
12442|LUHRIG
12443|LUIS LLORENS TORRES
12444|LUIS LLORÉNS TORRES COMUNIDAD
12445|LUIS LOPEZ
12446|LUIS M. CINTRON
12447|LUIS M. CINTRÓN COMUNIDAD
12448|LUKACHUKAI
12449|LUKE
12450|LUKEVILLE
12451|LULA
12452|LULING
12453|LULU
12454|LUM
12455|LUMBER BRIDGE
12456|LUMBER CITY
12457|LUMBERPORT
12458|LUMBERTON
12459|LUMPKIN
12460|LUMS CHAPEL
12461|LUNA
12462|LUNA PIER
12463|LUND
12464|LUNDELL
12465|LUNDS
12466|LUNDY
12467|LUNENBURG
12468|LUNING
12469|LUPTON
12470|LUPUS
12471|LUQUILLO
12472|LUQUILLO ZONA URBANA
12473|LURAVILLE
12474|LURAY
12475|LURTON
12476|LUSBY
12477|LUSHTON
12478|LUSK
12479|LUSTRE
12480|LUTAK
12481|LUTCHER
12482|LUTHER
12483|LUTHERSBURG
12484|LUTHERSVILLE
12485|LUTHERVILLE
12486|LUTIE
12487|LUTON
12488|LUTSEN
12489|LUTTRELL
12490|LUTTS
12491|LUTZ
12492|LUVERNE
12493|LUXEMBURG
12494|LUXOR
12495|LUXORA
12496|LUYANDO
12497|LUYANDO COMUNIDAD
12498|LUZERNE
12499|LYCAN
12500|LYDEN
12501|LYDIA
12502|LYDICK
12503|LYERLY
12504|LYFORD
12505|LYKENS
12506|LYLE
12507|LYLES
12508|LYMAN
12509|LYNBROOK
12510|LYNCH
12511|LYNCH STATION
12512|LYNCHBURG
12513|LYNCOURT
12514|LYND
12515|LYNDELL
12516|LYNDEN
12517|LYNDHURST
12518|LYNDON
12519|LYNDON STATION
12520|LYNDONVILLE
12521|LYNDORA
12522|LYNN
12523|LYNN GARDEN
12524|LYNN GROVE
12525|LYNN HAVEN
12526|LYNNDYL
12527|LYNNE
12528|LYNNFIELD
12529|LYNNVIEW
12530|LYNNVILLE
12531|LYNNWOOD
12532|LYNWOOD
12533|LYNWOOD HILLS
12534|LYNXVILLE
12535|LYON
12536|LYON MOUNTAIN
12537|LYONS
12538|LYONS FALLS
12539|LYONS PLAIN
12540|LYSITE
12541|LYTLE
12542|LYTLE CREEK
12543|LYTTON
12544|LĀNAʻI CITY
12545|LĀWAʻI
12546|LĀʻIE
12547|LĪHUʻE
12548|MABANA
12549|MABANK
12550|MABEL
12551|MABELLE
12552|MABELVALE
12553|MABEN
12554|MABIE
12555|MABLETON
12556|MABSCOTT
12557|MABTON
12558|MACARTHUR
12559|MACCLENNY
12560|MACCLESFIELD
12561|MACDOEL
12562|MACDONA
12563|MACEDON
12564|MACEDONIA
12565|MACEO
12566|MACHENS
12567|MACHESNEY PARK
12568|MACHIAS
12569|MACHOVEC
12570|MACK
12571|MACKAY
12572|MACKENZIE
12573|MACKEY
12574|MACKEYS
12575|MACKINAC ISLAND
12576|MACKINAW
12577|MACKINAW CITY
12578|MACKS CREEK
12579|MACKSBURG
12580|MACKSVILLE
12581|MACKVILLE
12582|MACLAND
12583|MACOMB
12584|MACON
12585|MACOPIN
12586|MACUNGIE
12587|MACWAHOC
12588|MACY
12589|MAD RIVER
12590|MADAKET
12591|MADAWASKA
12592|MADDEN
12593|MADDOCK
12594|MADEIRA
12595|MADEIRA BEACH
12596|MADELIA
12597|MADELINE
12598|MADERA
12599|MADERA ACRES
12600|MADILL
12601|MADISON
12602|MADISON HEIGHTS
12603|MADISON LAKE
12604|MADISON MILLS
12605|MADISON PARK
12606|MADISONBURG
12607|MADISONVILLE
12608|MADOC
12609|MADONNA
12610|MADRAS
12611|MADRID
12612|MADRONE
12613|MAESER
12614|MAEYSTOWN
12615|MAGALIA
12616|MAGAS ARRIBA
12617|MAGAS ARRIBA COMUNIDAD
12618|MAGASCO
12619|MAGAZINE
12620|MAGDALENA
12621|MAGEE
12622|MAGGIE VALLEY
12623|MAGMA
12624|MAGNA
12625|MAGNESS
12626|MAGNET
12627|MAGNET COVE
12628|MAGNETIC SPRINGS
12629|MAGNOLIA
12630|MAGNOLIA BEACH
12631|MAGNOLIA GARDENS
12632|MAGNOLIA SPRINGS
12633|MAGOUN
12634|MAGUAYO
12635|MAGUAYO COMUNIDAD
12636|MAGWALT
12637|MAHAFFEY
12638|MAHANOY CITY
12639|MAHARISHI VEDIC CITY
12640|MAHASKA
12641|MAHNOMEN
12642|MAHOMET
12643|MAHOPAC
12644|MAHTOMEDI
12645|MAHTOWA
12646|MAHWAH
12647|MAIDA
12648|MAIDEN
12649|MAIDEN ROCK
12650|MAINE
12651|MAINEVILLE
12652|MAINVILLE
12653|MAISH VAYA
12654|MAITLAND
12655|MAIZE
12656|MAJENICA
12657|MAJESTIC
12658|MAKAKILO CITY
12659|MAKANDA
12660|MAKAWAO
12661|MAKEMIE PARK
12662|MAKINEN
12663|MAKOTI
12664|MALABAR
12665|MALAD CITY
12666|MALAGA
12667|MALAKOFF
12668|MALCOLM
12669|MALCOM
12670|MALDEN
12671|MALDEN-ON-HUDSON
12672|MALESUS
12673|MALIBU
12674|MALIN
12675|MALINTA
12676|MALJAMAR
12677|MALLARD
12678|MALLORY
12679|MALMO
12680|MALO
12681|MALONE
12682|MALOTT
12683|MALOY
12684|MALTA
12685|MALTA BEND
12686|MALTBY
12687|MALVADO
12688|MALVERN
12689|MALVERNE
12690|MALVERNE PARK OAKS
12691|MAMARONECK
12692|MAMERS
12693|MAMMOTH
12694|MAMMOTH CAVE
12695|MAMMOTH LAKES
12696|MAMMOTH SPRING
12697|MAMONT
12698|MAMOU
12699|MANACK
12700|MANAHAWKIN
12701|MANAKIN
12702|MANALAPAN
12703|MANANNAH
12704|MANASOTA KEY
12705|MANASQUAN
12706|MANASSA
12707|MANASSAS
12708|MANASSAS PARK
12709|MANATEE ROAD
12710|MANATÍ
12711|MANATÍ ZONA URBANA
12712|MANAWA
12713|MANCELONA
12714|MANCHAC
12715|MANCHACA
12716|MANCHESTER
12717|MANCHESTER CENTER
12718|MANCHESTER TOWNSHIP
12719|MANCHESTER-BY-THE-SEA
12720|MANCOS
12721|MANDAN
12722|MANDAREE
12723|MANDERFIELD
12724|MANDERSON
12725|MANDEVILLE
12726|MANES
12727|MANGHAM
12728|MANGO
12729|MANGONIA PARK
12730|MANGUM
12731|MANHASSET
12732|MANHASSET HILLS
12733|MANHATTAN
12734|MANHATTAN BEACH
12735|MANHEIM
12736|MANIFEST
12737|MANIFOLD
12738|MANILA
12739|MANILLA
12740|MANISTEE
12741|MANISTIQUE
12742|MANITO
12743|MANITOU
12744|MANITOU BEACH
12745|MANITOU SPRINGS
12746|MANITOWISH
12747|MANITOWOC
12748|MANKATO
12749|MANKINS
12750|MANLEY
12751|MANLEY HOT SPRINGS
12752|MANLIUS
12753|MANLY
12754|MANNFORD
12755|MANNING
12756|MANNINGTON
12757|MANNS CHOICE
12758|MANNS HARBOR
12759|MANNSVILLE
12760|MANOKOTAK
12761|MANOR
12762|MANOR CREEK
12763|MANORHAVEN
12764|MANORVILLE
12765|MANSFIELD
12766|MANSFIELD CENTER
12767|MANSON
12768|MANSURA
12769|MANTACHIE
12770|MANTADOR
12771|MANTECA
12772|MANTEE
12773|MANTENO
12774|MANTEO
12775|MANTER
12776|MANTI
12777|MANTOLOKING
12778|MANTON
12779|MANTORVILLE
12780|MANTUA
12781|MANUELITO
12782|MANVEL
12783|MANVILLE
12784|MANY
12785|MANY FARMS
12786|MANZANITA
12787|MANZANO
12788|MANZANO SPRINGS
12789|MANZANOLA
12790|MAPLE BAY
12791|MAPLE BLUFF
12792|MAPLE CITY
12793|MAPLE FALLS
12794|MAPLE GLEN
12795|MAPLE GROVE
12796|MAPLE HEIGHTS
12797|MAPLE HILL
12798|MAPLE LAKE
12799|MAPLE PARK
12800|MAPLE PLAIN
12801|MAPLE RAPIDS
12802|MAPLE RIDGE
12803|MAPLE SHADE
12804|MAPLE VALLEY
12805|MAPLESVILLE
12806|MAPLETON
12807|MAPLETOWN
12808|MAPLEVIEW
12809|MAPLEVILLE
12810|MAPLEWOOD
12811|MAPLEWOOD PARK
12812|MAPPSBURG
12813|MAPPSVILLE
12814|MAQUOKETA
12815|MAQUON
12816|MAR-MAC
12817|MARAMEC
12818|MARANA
12819|MARATHON
12820|MARATHON SHORES
12821|MARBLE
12822|MARBLE CANYON
12823|MARBLE CITY
12824|MARBLE CLIFF
12825|MARBLE FALLS
12826|MARBLE HILL
12827|MARBLE ROCK
12828|MARBLEDALE
12829|MARBLEHEAD
12830|MARBLEMOUNT
12831|MARBLETON
12832|MARBURY
12833|MARCELINE
12834|MARCELL
12835|MARCELLA
12836|MARCELLUS
12837|MARCHE
12838|MARCO
12839|MARCOLA
12840|MARCUS
12841|MARCUS HOOK
12842|MARDELA SPRINGS
12843|MARENGO
12844|MARENISCO
12845|MARFA
12846|MARGARET
12847|MARGARETVILLE
12848|MARGATE
12849|MARGATE CITY
12850|MARGIE
12851|MARGUERITE
12852|MARIA ANTONIA
12853|MARIANNA
12854|MARIANNE
12855|MARIANO COLÓN
12856|MARIANO COLÓN COMUNIDAD
12857|MARIAVILLE LAKE
12858|MARIBA
12859|MARIBEL
12860|MARICAO
12861|MARICAO ZONA URBANA
12862|MARICOPA
12863|MARIE
12864|MARIEMONT
12865|MARIENTHAL
12866|MARIENVILLE
12867|MARIETTA
12868|MARIN CITY
12869|MARINA
12870|MARINA DEL REY
12871|MARINE
12872|MARINE CITY
12873|MARINE ON SAINT CROIX
12874|MARINELAND
12875|MARINETTE
12876|MARINGOUIN
12877|MARINWOOD
12878|MARION
12879|MARION CENTER
12880|MARION HEIGHTS
12881|MARION HILL
12882|MARION JUNCTION
12883|MARIONVILLE
12884|MARIPOSA
12885|MARISSA
12886|MARK
12887|MARKED TREE
12888|MARKESAN
12889|MARKHAM
12890|MARKLE
12891|MARKLEEVILLE
12892|MARKLESBURG
12893|MARKLEVILLE
12894|MARKLEYSBURG
12895|MARKS
12896|MARKSBORO
12897|MARKSVILLE
12898|MARKVILLE
12899|MARLAND
12900|MARLBORO
12901|MARLBORO MEADOWS
12902|MARLBOROUGH
12903|MARLETTE
12904|MARLEY
12905|MARLIN
12906|MARLINTON
12907|MARLOW
12908|MARLOW HEIGHTS
12909|MARLTON
12910|MARMADUKE
12911|MARMARTH
12912|MARMET
12913|MARNE
12914|MAROA
12915|MARQUAND
12916|MARQUETTE
12917|MARQUETTE HEIGHTS
12918|MARQUEZ
12919|MARRERO
12920|MARRIOTT-SLATERVILLE
12921|MARROWBONE
12922|MARROWSTONE
12923|MARS
12924|MARS HILL
12925|MARSEILLES
12926|MARSH
12927|MARSHALL
12928|MARSHALLBERG
12929|MARSHALLTON
12930|MARSHALLTOWN
12931|MARSHALLVILLE
12932|MARSHDALE
12933|MARSHFIELD
12934|MARSHFIELD CENTER
12935|MARSHFIELD HILLS
12936|MARSHVILLE
12937|MARSING
12938|MARSLAND
12939|MARSTON
12940|MARSTONS MILLS
12941|MART
12942|MARTEL
12943|MARTELL
12944|MARTELLE
12945|MARTENSDALE
12946|MARTHA
12947|MARTHA LAKE
12948|MARTHASVILLE
12949|MARTHAVILLE
12950|MARTIN
12951|MARTIN BLUFF
12952|MARTIN CITY
12953|MARTIN LAKE
12954|MARTINDALE
12955|MARTINEZ
12956|MARTINS ADDITIONS
12957|MARTINS CREEK
12958|MARTINS FERRY
12959|MARTINS MILL
12960|MARTINSBURG
12961|MARTINSDALE
12962|MARTINSVILLE
12963|MARTINTON
12964|MARTINVILLE
12965|MARTORELL
12966|MARTORELL COMUNIDAD
12967|MARTY
12968|MARUEÑO
12969|MARUEÑO COMUNIDAD
12970|MARVEL
12971|MARVELL
12972|MARVIN
12973|MARY ESTHER
12974|MARYDEL
12975|MARYHILL
12976|MARYHILL ESTATES
12977|MARYLAND CITY
12978|MARYLAND HEIGHTS
12979|MARYNEAL
12980|MARYS CORNER
12981|MARYS HOME
12982|MARYSVALE
12983|MARYSVILLE
12984|MARYVILLE
12985|MARÍA ANTONIA COMUNIDAD
12986|MASARYKTOWN
12987|MASCOT
12988|MASCOTTE
12989|MASCOUTAH
12990|MASHPEE NECK
12991|MASHULAVILLE
12992|MASKELL
12993|MASON
12994|MASON CITY
12995|MASONTOWN
12996|MASONVILLE
12997|MASPETH
12998|MASSAC
12999|MASSADONA
13000|MASSANETTA SPRINGS
13001|MASSANUTTEN
13002|MASSAPEQUA
13003|MASSAPEQUA PARK
13004|MASSENA
13005|MASSIES MILL
13006|MASSIEVILLE
13007|MASSILLON
13008|MASTERS
13009|MASTERSON
13010|MASTHOPE
13011|MASTIC
13012|MASTIC BEACH
13013|MASURY
13014|MATADOR
13015|MATAGORDA
13016|MATAMORAS
13017|MATANUSKA
13018|MATAWAN
13019|MATEWAN
13020|MATFIELD GREEN
13021|MATHENY
13022|MATHER
13023|MATHERVILLE
13024|MATHESON
13025|MATHEWS
13026|MATHIAS
13027|MATHIS
13028|MATHISTON
13029|MATINECOCK
13030|MATLACHA
13031|MATLOCK
13032|MATOACA
13033|MATOAKA
13034|MATTAPEX
13035|MATTAWA
13036|MATTAWAN
13037|MATTAWANA
13038|MATTAWOMAN
13039|MATTESE
13040|MATTESON
13041|MATTHEWS
13042|MATTITUCK
13043|MATTOON
13044|MATTOXTOWN
13045|MATTSON
13046|MATTYDALE
13047|MAUCKPORT
13048|MAUD
13049|MAUDLOW
13050|MAUGANSVILLE
13051|MAULDIN
13052|MAUMEE
13053|MAUMELLE
13054|MAUNABO
13055|MAUNABO ZONA URBANA
13056|MAUNALOA
13057|MAUNAWILI
13058|MAUNIE
13059|MAUPIN
13060|MAURERTOWN
13061|MAURICE
13062|MAURICEVILLE
13063|MAURINE
13064|MAURY
13065|MAURY CITY
13066|MAUSDALE
13067|MAUSTON
13068|MAUSTOWN
13069|MAVERICK
13070|MAVISDALE
13071|MAX
13072|MAX MEADOWS
13073|MAXBASS
13074|MAXEYS
13075|MAXIE
13076|MAXIMO
13077|MAXTON
13078|MAXVILLE
13079|MAXWELL
13080|MAXWELTON
13081|MAY CITY
13082|MAY CREEK
13083|MAYAGÜEZ
13084|MAYAGÜEZ ZONA URBANA
13085|MAYBEE
13086|MAYBELL
13087|MAYBEURY
13088|MAYBROOK
13089|MAYDAY
13090|MAYDELLE
13091|MAYER
13092|MAYERSVILLE
13093|MAYESVILLE
13094|MAYETTA
13095|MAYFIELD
13096|MAYFIELD HEIGHTS
13097|MAYFLOWER
13098|MAYFLOWER VILLAGE
13099|MAYHEW
13100|MAYHILL
13101|MAYKING
13102|MAYLENE
13103|MAYNA
13104|MAYNARD
13105|MAYNARDVILLE
13106|MAYO
13107|MAYODAN
13108|MAYOWORTH
13109|MAYPEARL
13110|MAYPENS
13111|MAYS
13112|MAYS CHAPEL
13113|MAYS LANDING
13114|MAYS LICK
13115|MAYSFIELD
13116|MAYSVILLE
13117|MAYTOWN
13118|MAYVIEW
13119|MAYVILLE
13120|MAYWOOD
13121|MAYWOOD PARK
13122|MAZAMA
13123|MAZEPPA
13124|MAZIE
13125|MAZOMANIE
13126|MAZON
13127|MC LEAN
13128|MCADAMS
13129|MCADENVILLE
13130|MCADOO
13131|MCAFEE
13132|MCALESTER
13133|MCALISTER
13134|MCALISTERVILLE
13135|MCALLEN
13136|MCALLISTER
13137|MCALMONT
13138|MCALPIN
13139|MCARTHUR
13140|MCBAIN
13141|MCBAINE
13142|MCBEAN
13143|MCBEE
13144|MCBRIDE
13145|MCCABE
13146|MCCALL
13147|MCCALL CREEK
13148|MCCALLSBURG
13149|MCCALLUM
13150|MCCAMEY
13151|MCCAMMON
13152|MCCARR
13153|MCCARTHY
13154|MCCARTYS
13155|MCCASKILL
13156|MCCAULLEY
13157|MCCAUSLAND
13158|MCCAYSVILLE
13159|MCCLAVE
13160|MCCLEARY
13161|MCCLELLAND
13162|MCCLELLANVILLE
13163|MCCLOUD
13164|MCCLURE
13165|MCCLUSKY
13166|MCCOLL
13167|MCCOMB
13168|MCCONNELL
13169|MCCONNELLS
13170|MCCONNELLSBURG
13171|MCCONNELLSTOWN
13172|MCCONNELSVILLE
13173|MCCONNICO
13174|MCCOOK
13175|MCCOOL
13176|MCCOOL JUNCTION
13177|MCCOOLE
13178|MCCORD
13179|MCCORD BEND
13180|MCCORDSVILLE
13181|MCCORMICK
13182|MCCOY
13183|MCCOYS CORNER
13184|MCCRACKEN
13185|MCCREDIE SPRINGS
13186|MCCRORY
13187|MCCULLOM LAKE
13188|MCCUNE
13189|MCCUNEVILLE
13190|MCCURTAIN
13191|MCCUTCHENVILLE
13192|MCDADE
13193|MCDANIEL
13194|MCDANIELS
13195|MCDAVID
13196|MCDERMITT
13197|MCDERMOTT
13198|MCDONALD
13199|MCDONALD CHAPEL
13200|MCDONOUGH
13201|MCDOUGAL
13202|MCDOWELL
13203|MCELHATTAN
13204|MCEWEN
13205|MCEWENSVILLE
13206|MCFADDEN
13207|MCFADDIN
13208|MCFALL
13209|MCFARLAN
13210|MCFARLAND
13211|MCGEE
13212|MCGEHEE
13213|MCGILL
13214|MCGONIGLE
13215|MCGOVERN
13216|MCGRADY
13217|MCGRATH
13218|MCGRAW
13219|MCGREGOR
13220|MCGREW
13221|MCGUFFEY
13222|MCHENRY
13223|MCINTIRE
13224|MCINTOSH
13225|MCINTYRE
13226|MCKAMIE
13227|MCKEANSBURG
13228|MCKEE
13229|MCKEES ROCKS
13230|MCKEESPORT
13231|MCKENNA
13232|MCKENNEY
13233|MCKENZIE
13234|MCKENZIE BRIDGE
13235|MCKIBBEN
13236|MCKINLEY
13237|MCKINLEY HEIGHTS
13238|MCKINLEYVILLE
13239|MCKINNEY
13240|MCKINNEY ACRES
13241|MCKINNON
13242|MCKITTRICK
13243|MCKNIGHT
13244|MCKNIGHTSTOWN
13245|MCLAIN
13246|MCLAUGHLIN
13247|MCLAURIN
13248|MCLEAN
13249|MCLEANSBORO
13250|MCLEANSVILLE
13251|MCLEMORESVILLE
13252|MCLENDON-CHISHOLM
13253|MCLEOD
13254|MCLOUD
13255|MCLOUTH
13256|MCMANUS
13257|MCMECHEN
13258|MCMILLAN
13259|MCMILLIN
13260|MCMINNVILLE
13261|MCMULLEN
13262|MCMULLIN
13263|MCMURRAY
13264|MCNAB
13265|MCNABB
13266|MCNAIR
13267|MCNARY
13268|MCNAUGHTON
13269|MCNEAL
13270|MCNEIL
13271|MCNEILL
13272|MCPHERSON
13273|MCQUADY
13274|MCQUEEN
13275|MCQUEENEY
13276|MCRAE
13277|MCROBERTS
13278|MCSHERRYSTOWN
13279|MCVEIGH
13280|MCVEYTOWN
13281|MCVILLE
13282|MCWHORTER
13283|MCWILLIAMS
13284|MCWILLIE
13285|MEACHAM
13286|MEAD
13287|MEAD VALLEY
13288|MEADE
13289|MEADOW
13290|MEADOW ACRES
13291|MEADOW BRIDGE
13292|MEADOW CREEK
13293|MEADOW GLADE
13294|MEADOW GROVE
13295|MEADOW LAKE
13296|MEADOW LAKES
13297|MEADOW LANDS
13298|MEADOW VALE
13299|MEADOW VALLEY
13300|MEADOW VIEW ADDITION
13301|MEADOW VISTA
13302|MEADOW WOODS
13303|MEADOWBROOK
13304|MEADOWBROOK FARM
13305|MEADOWBROOK TERRACE
13306|MEADOWDALE
13307|MEADOWLAKES
13308|MEADOWLANDS
13309|MEADOWOOD
13310|MEADOWS
13311|MEADOWS PLACE
13312|MEADOWVIEW
13313|MEADOWVIEW ESTATES
13314|MEADVIEW
13315|MEADVILLE
13316|MEANSVILLE
13317|MEAUX
13318|MEBANE
13319|MECCA
13320|MECHANIC FALLS
13321|MECHANICSBURG
13322|MECHANICSTOWN
13323|MECHANICSVILLE
13324|MECHANICVILLE
13325|MECKLING
13326|MECOSTA
13327|MEDANALES
13328|MEDART
13329|MEDARYVILLE
13330|MEDFIELD
13331|MEDFORD
13332|MEDFORD LAKES
13333|MEDFRA
13334|MEDIA
13335|MEDIAPOLIS
13336|MEDICAL LAKE
13337|MEDICINE BOW
13338|MEDICINE LAKE
13339|MEDICINE LODGE
13340|MEDICINE MOUND
13341|MEDICINE PARK
13342|MEDINA
13343|MEDINAH
13344|MEDLEY
13345|MEDON
13346|MEDORA
13347|MEDULLA
13348|MEEKER
13349|MEEKS BAY
13350|MEERS
13351|MEETEETSE
13352|MEGARGEL
13353|MEGGETT
13354|MEGLER
13355|MEHAMA
13356|MEHERRIN
13357|MEHLVILLE
13358|MEIGS
13359|MEINERS OAKS
13360|MEINHARD
13361|MEIRE GROVE
13362|MEKINOCK
13363|MEKORYUK
13364|MELBA
13365|MELBETA
13366|MELBOURNE
13367|MELBOURNE BEACH
13368|MELBOURNE VILLAGE
13369|MELBY
13370|MELCHER-DALLAS
13371|MELDER
13372|MELDRUM
13373|MELFA
13374|MELISSA
13375|MELITOTA
13376|MELLEN
13377|MELLETTE
13378|MELLIN
13379|MELLOTT
13380|MELMORE
13381|MELODY HILL
13382|MELODY HILLS
13383|MELROSE
13384|MELROSE PARK
13385|MELRUDE
13386|MELSTONE
13387|MELSTRAND
13388|MELVERN
13389|MELVILLE
13390|MELVIN
13391|MELVIN VILLAGE
13392|MELVINA
13393|MELVINDALE
13394|MEMPHIS
13395|MEMPHIS JUNCTION
13396|MENA
13397|MENAHGA
13398|MENAN
13399|MENANDS
13400|MENARD
13401|MENASHA
13402|MENCHALVILLE
13403|MENDELTNA
13404|MENDENHALL
13405|MENDES
13406|MENDHAM
13407|MENDOCINO
13408|MENDON
13409|MENDOTA
13410|MENDOTA HEIGHTS
13411|MENDOZA
13412|MENFRO
13413|MENIFEE
13414|MENLO
13415|MENLO PARK
13416|MENNO
13417|MENO
13418|MENOKEN
13419|MENOMINEE
13420|MENOMONEE FALLS
13421|MENTASTA LAKE
13422|MENTMORE
13423|MENTONE
13424|MENTOR
13425|MENTOR-ON-THE-LAKE
13426|MEPPEN
13427|MEQUON
13428|MER ROUGE
13429|MERAUX
13430|MERCED
13431|MERCEDES
13432|MERCER
13433|MERCER ISLAND
13434|MERCERSBURG
13435|MERCERSVILLE
13436|MERCERVILLE
13437|MERCHANTVILLE
13438|MERCURY
13439|MEREDITH
13440|MEREDOSIA
13441|MERIDEAN
13442|MERIDEN
13443|MERIDIAN
13444|MERIDIAN HILLS
13445|MERIDIANVILLE
13446|MERIGOLD
13447|MERINO
13448|MERIT
13449|MERIWETHER
13450|MERKEL
13451|MERLIN
13452|MERMENTAU
13453|MERNA
13454|MEROM
13455|MERRIAM
13456|MERRIAM WOODS
13457|MERRICK
13458|MERRIFIELD
13459|MERRILL
13460|MERRILLAN
13461|MERRILLVILLE
13462|MERRIMAC
13463|MERRIMAN
13464|MERRIMON
13465|MERRIONETTE PARK
13466|MERRITT
13467|MERRITT ISLAND
13468|MERRYDALE
13469|MERRYVILLE
13470|MERSHON
13471|MERTENS
13472|MERTON
13473|MERTZON
13474|MERTZTOWN
13475|MERWIN
13476|MESA
13477|MESA DEL CABALLO
13478|MESA GRANDE
13479|MESA VERDE
13480|MESA VISTA
13481|MESCAL
13482|MESCALERO
13483|MESERVEY
13484|MESHOPPEN
13485|MESIC
13486|MESICK
13487|MESILLA
13488|MESITA
13489|MESQUITE
13490|MESQUITE CREEK
13491|META
13492|METAIRIE
13493|METALINE
13494|METALINE FALLS
13495|METAMORA
13496|METCALF
13497|METCALF GAP
13498|METCALFE
13499|METEA
13500|METHOW
13501|METHUEN
13502|METLAKATLA
13503|METOLIUS
13504|METOMPKIN
13505|METROPOLIS
13506|METTAWA
13507|METTER
13508|METTLER
13509|METUCHEN
13510|METZ
13511|METZGER
13512|MEXIA
13513|MEXICAN COLONY
13514|MEXICAN HAT
13515|MEXICAN WATER
13516|MEXICO
13517|MEXICO BEACH
13518|MEYER
13519|MEYERS
13520|MEYERS CHUCK
13521|MEYERS LAKE
13522|MEYERSDALE
13523|MI-WUK VILLAGE
13524|MIAMI
13525|MIAMI BEACH
13526|MIAMI GARDENS
13527|MIAMI HEIGHTS
13528|MIAMI LAKES
13529|MIAMI SHORES
13530|MIAMI SPRINGS
13531|MIAMISBURG
13532|MIAMITOWN
13533|MIAMIVILLE
13534|MICANOPY
13535|MICAVILLE
13536|MICCO
13537|MICCOSUKEE
13538|MICHIANA
13539|MICHIANA SHORES
13540|MICHIE
13541|MICHIGAMME
13542|MICHIGAN
13543|MICHIGAN CENTER
13544|MICHIGAN CITY
13545|MICHIGANTOWN
13546|MICKLETON
13547|MIDAS
13548|MIDDLE AMANA
13549|MIDDLE GROVE
13550|MIDDLE ISLAND
13551|MIDDLE POINT
13552|MIDDLE RIVER
13553|MIDDLE VALLEY
13554|MIDDLE VILLAGE
13555|MIDDLE WATER
13556|MIDDLEBERG
13557|MIDDLEBORO
13558|MIDDLEBOURNE
13559|MIDDLEBROOK
13560|MIDDLEBURG
13561|MIDDLEBURG HEIGHTS
13562|MIDDLEBURGH
13563|MIDDLEBURY
13564|MIDDLEBUSH
13565|MIDDLEFIELD
13566|MIDDLEPORT
13567|MIDDLESBORO
13568|MIDDLESEX
13569|MIDDLETON
13570|MIDDLETOWN
13571|MIDDLEVILLE
13572|MIDDLEWAY
13573|MIDFIELD
13574|MIDLAND
13575|MIDLAND CITY
13576|MIDLAND PARK
13577|MIDLOTHIAN
13578|MIDNIGHT
13579|MIDPINES
13580|MIDTOWN
13581|MIDVALE
13582|MIDVALE CORNER
13583|MIDVILLE
13584|MIDWAY
13585|MIDWAY CITY
13586|MIDWAY PARK
13587|MIDWEST
13588|MIDWEST CITY
13589|MIER
13590|MIESVILLE
13591|MIFFLIN
13592|MIFFLINBURG
13593|MIFFLINTOWN
13594|MIFFLINVILLE
13595|MIGNON
13596|MIKADO
13597|MIKKALO
13598|MILA DOCE
13599|MILACA
13600|MILAM
13601|MILAN
13602|MILANO
13603|MILBANK
13604|MILBURN
13605|MILDRED
13606|MILES
13607|MILES CITY
13608|MILESBURG
13609|MILESVILLE
13610|MILEY
13611|MILFORD
13612|MILFORD CENTER
13613|MILFORD CROSSROADS
13614|MILFORD MILL
13615|MILFORD SQUARE
13616|MILILANI TOWN
13617|MILL BROOK
13618|MILL CITY
13619|MILL CREEK
13620|MILL GROVE
13621|MILL HALL
13622|MILL IRON
13623|MILL NECK
13624|MILL SHOALS
13625|MILL SPRING
13626|MILL VALLEY
13627|MILL VILLAGE
13628|MILLADORE
13629|MILLARD
13630|MILLBORO
13631|MILLBOURNE
13632|MILLBRAE
13633|MILLBROOK
13634|MILLBURN
13635|MILLBURY
13636|MILLCREEK
13637|MILLEDGEVILLE
13638|MILLEN
13639|MILLER
13640|MILLER CITY
13641|MILLER HOUSE
13642|MILLER PLACE
13643|MILLERS COVE
13644|MILLERS CREEK
13645|MILLERS FALLS
13646|MILLERS FERRY
13647|MILLERS LANDING
13648|MILLERSBURG
13649|MILLERSPORT
13650|MILLERSTOWN
13651|MILLERSVIEW
13652|MILLERSVILLE
13653|MILLERTON
13654|MILLERVILLE
13655|MILLETT
13656|MILLEVILLE BEACH
13657|MILLFIELD
13658|MILLGROVE
13659|MILLHAVEN
13660|MILLHEIM
13661|MILLHOUSEN
13662|MILLHURST
13663|MILLICAN
13664|MILLIGAN
13665|MILLIGANTOWN
13666|MILLIKEN
13667|MILLIKIN
13668|MILLINGPORT
13669|MILLINGTON
13670|MILLINOCKET
13671|MILLPORT
13672|MILLRY
13673|MILLS
13674|MILLS RIVER
13675|MILLSAP
13676|MILLSBORO
13677|MILLSTADT
13678|MILLSTON
13679|MILLSTONE
13680|MILLTOWN
13681|MILLVALE
13682|MILLVILLE
13683|MILLWOOD
13684|MILNER
13685|MILNESAND
13686|MILNOR
13687|MILO
13688|MILOLIʻI
13689|MILPITAS
13690|MILROY
13691|MILSTEAD
13692|MILTON
13693|MILTON CENTER
13694|MILTON MILLS
13695|MILTON-FREEWATER
13696|MILTONA
13697|MILTONSBURG
13698|MILTONVALE
13699|MILTONVILLE
13700|MILWAUKEE
13701|MILWAUKIE
13702|MIMBRES
13703|MIMOSA PARK
13704|MIMS
13705|MINA
13706|MINAM
13707|MINATARE
13708|MINBURN
13709|MINCO
13710|MINDEN
13711|MINDEN CITY
13712|MINDENMINES
13713|MINDORO
13714|MINE HILL
13715|MINE LA MOTTE
13716|MINEOLA
13717|MINER
13718|MINERAL
13719|MINERAL BLUFF
13720|MINERAL CITY
13721|MINERAL HILLS
13722|MINERAL HOT SPRINGS
13723|MINERAL POINT
13724|MINERAL RIDGE
13725|MINERAL SPRINGS
13726|MINERAL WELLS
13727|MINERSVILLE
13728|MINERVA
13729|MINERVA PARK
13730|MINETTO
13731|MINEVILLE
13732|MINFORD
13733|MINGO
13734|MINGO JUNCTION
13735|MINGOVILLE
13736|MINGUS
13737|MINIDOKA
13738|MINIER
13739|MINK CREEK
13740|MINKLER
13741|MINNEAPOLIS
13742|MINNEHAHA
13743|MINNEHAHA SPRINGS
13744|MINNEISKA
13745|MINNEOLA
13746|MINNEOTA
13747|MINNESOTA CITY
13748|MINNESOTA LAKE
13749|MINNESOTT BEACH
13750|MINNETONKA
13751|MINNETONKA BEACH
13752|MINNETRISTA
13753|MINNEWAUKAN
13754|MINOA
13755|MINOCQUA
13756|MINONG
13757|MINONK
13758|MINOOKA
13759|MINOR HILL
13760|MINORCA
13761|MINOT
13762|MINQUADALE
13763|MINSTER
13764|MINT HILL
13765|MINTER
13766|MINTER CITY
13767|MINTERS CHAPEL
13768|MINTLE
13769|MINTO
13770|MINTURN
13771|MIO
13772|MIRA
13773|MIRA LOMA
13774|MIRA MONTE
13775|MIRACLE HOT SPRINGS
13776|MIRACLE VALLEY
13777|MIRAMAR
13778|MIRAMAR BEACH
13779|MIRAMIGUOA PARK
13780|MIRANDA
13781|MIRANDA COMUNIDAD
13782|MIRANDO CITY
13783|MIRRORMONT
13784|MISENHEIMER
13785|MISHAWAKA
13786|MISHICOT
13787|MISQUAMICUT
13788|MISSION
13789|MISSION BEND
13790|MISSION CANYON
13791|MISSION HILL
13792|MISSION HILLS
13793|MISSION RIDGE
13794|MISSION VIEJO
13795|MISSION WOODS
13796|MISSOULA
13797|MISSOURI CITY
13798|MISSOURI VALLEY
13799|MIST
13800|MITCHELL
13801|MITCHELL HEIGHTS
13802|MITCHELLSBURG
13803|MITCHELLSVILLE
13804|MITCHELLTOWN
13805|MITCHELLVILLE
13806|MITIWANGA
13807|MITTIE
13808|MIXERSVILLE
13809|MIZE
13810|MIZPAH
13811|MOAB
13812|MOAPA
13813|MOAPA TOWN
13814|MOAPA VALLEY
13815|MOARK
13816|MOBEETIE
13817|MOBERLY
13818|MOBILE
13819|MOBILE CITY
13820|MOBRIDGE
13821|MOCA
13822|MOCA ZONA URBANA
13823|MOCANAQUA
13824|MOCANE
13825|MOCCASIN
13826|MOCKINGBIRD VALLEY
13827|MOCKSVILLE
13828|MOCLIPS
13829|MODALE
13830|MODDERSVILLE
13831|MODEL
13832|MODEL CITY
13833|MODENA
13834|MODEST TOWN
13835|MODESTE
13836|MODESTO
13837|MODOC
13838|MOENKOPI
13839|MOFFAT
13840|MOFFETT
13841|MOFFIT
13842|MOGADORE
13843|MOGOTE
13844|MOGUL
13845|MOHALL
13846|MOHAVE VALLEY
13847|MOHAWK
13848|MOHAWK VISTA
13849|MOHLER
13850|MOHNTON
13851|MOHRSVILLE
13852|MOIESE
13853|MOINGONA
13854|MOJAVE
13855|MOJAVE RANCH ESTATES
13856|MOKANE
13857|MOKELUMNE HILL
13858|MOKENA
13859|MOKULĒʻIA
13860|MOLALLA
13861|MOLE LAKE
13862|MOLENA
13863|MOLINA
13864|MOLINE
13865|MOLINE ACRES
13866|MOLINO
13867|MOLLUSK
13868|MOLSON
13869|MOLT
13870|MOLYNEAUX CORNERS
13871|MOMENCE
13872|MOMEYER
13873|MONA
13874|MONACA
13875|MONAHANS
13876|MONANGO
13877|MONARCH
13878|MONAVILLE
13879|MONCHES
13880|MONCKS CORNER
13881|MONCURE
13882|MONDAMIN
13883|MONDOVI
13884|MONEE
13885|MONELL
13886|MONERO
13887|MONESSEN
13888|MONETA
13889|MONETT
13890|MONETTA
13891|MONETTE
13892|MONEY
13893|MONEY CREEK
13894|MONFORT HEIGHTS
13895|MONIAC
13896|MONIDA
13897|MONINGER
13898|MONKSTOWN
13899|MONKTON
13900|MONMOUTH
13901|MONMOUTH BEACH
13902|MONMOUTH JUNCTION
13903|MONO CITY
13904|MONO VISTA
13905|MONOLITH
13906|MONOMOSCOY ISLAND
13907|MONON
13908|MONONA
13909|MONONGAH
13910|MONONGAHELA
13911|MONOWI
13912|MONROE
13913|MONROE CENTER
13914|MONROE CITY
13915|MONROETON
13916|MONROEVILLE
13917|MONROVIA
13918|MONSE
13919|MONSERRATE
13920|MONSERRATE COMUNIDAD
13921|MONSEY
13922|MONSON
13923|MONT ALTO
13924|MONT BELVIEU
13925|MONT CLARE
13926|MONT IDA
13927|MONTA VISTA
13928|MONTAGUE
13929|MONTALBA
13930|MONTALVIN
13931|MONTALVO
13932|MONTANA
13933|MONTANA CITY
13934|MONTANDON
13935|MONTARA
13936|MONTAUK
13937|MONTBROOK
13938|MONTCALM
13939|MONTCHANIN
13940|MONTCLAIR
13941|MONTE ALTO
13942|MONTE GRANDE
13943|MONTE GRANDE COMUNIDAD
13944|MONTE RIO
13945|MONTE SERENO
13946|MONTE VERDE COMUNIDAD
13947|MONTE VISTA
13948|MONTEAGLE
13949|MONTEBELLO
13950|MONTECITO
13951|MONTEGUT
13952|MONTEITH
13953|MONTELLO
13954|MONTEREY
13955|MONTEREY PARK
13956|MONTESANO
13957|MONTEVALLO
13958|MONTEVIDEO
13959|MONTEVIEW
13960|MONTEZUMA
13961|MONTEZUMA CREEK
13962|MONTFORT
13963|MONTGOMERY
13964|MONTGOMERY CITY
13965|MONTGOMERY CREEK
13966|MONTGOMERY VILLAGE
13967|MONTGOMERYVILLE
13968|MONTICELLO
13969|MONTIER
13970|MONTMORENCI
13971|MONTOUR
13972|MONTOUR FALLS
13973|MONTOURSVILLE
13974|MONTOYA
13975|MONTPELIER
13976|MONTREAL
13977|MONTREAT
13978|MONTROSE
13979|MONTROSE HILL
13980|MONTROSE MANOR
13981|MONTROSS
13982|MONTVALE
13983|MONTVERDE
13984|MONTVILLE
13985|MONTZ
13986|MONUMENT
13987|MONUMENT BEACH
13988|MOODUS
13989|MOODY
13990|MOODYS
13991|MOOERS
13992|MOOLEYVILLE
13993|MOON
13994|MOON RUN
13995|MOONACHIE
13996|MOONSHINE HILL
13997|MOONSTONE
13998|MOORCROFT
13999|MOORE
14000|MOORE HAVEN
14001|MOORE STATION
14002|MOOREFIELD
14003|MOORELAND
14004|MOORES BRIDGE
14005|MOORES HILL
14006|MOORES MILL
14007|MOORESBORO
14008|MOORESBURG
14009|MOORESTOWN
14010|MOORESVILLE
14011|MOORETON
14012|MOOREVILLE
14013|MOOREWOOD
14014|MOORHEAD
14015|MOORING
14016|MOORINGSPORT
14017|MOORLAND
14018|MOORPARK
14019|MOOSE
14020|MOOSE CREEK
14021|MOOSE LAKE
14022|MOOSE PASS
14023|MOOSE WILSON ROAD
14024|MOOSIC
14025|MOOSUP
14026|MOQUAH
14027|MOQUINO
14028|MORA
14029|MORA COMUNIDAD
14030|MORADA
14031|MORAGA
14032|MORAINE
14033|MORALES
14034|MORAN
14035|MORAVIA
14036|MORAVIAN FALLS
14037|MOREAUVILLE
14038|MOREHEAD
14039|MOREHEAD CITY
14040|MOREHOUSE
14041|MORELAND
14042|MORELAND HILLS
14043|MORENCI
14044|MORENO
14045|MORENO VALLEY
14046|MORGAN
14047|MORGAN CITY
14048|MORGAN FARM COLONIA
14049|MORGAN HILL
14050|MORGAN MILL
14051|MORGANA
14052|MORGANDALE
14053|MORGANFIELD
14054|MORGANS POINT
14055|MORGANS POINT RESORT
14056|MORGANTON
14057|MORGANTOWN
14058|MORGANVILLE
14059|MORGANZA
14060|MORGNEC
14061|MORIARTY
14062|MORICHES
14063|MORITA
14064|MORLAND
14065|MORLEY
14066|MORMON LAKE
14067|MORNING GLORY
14068|MORNING SUN
14069|MORNINGSIDE
14070|MORO
14071|MORO BAY
14072|MOROCCO
14073|MORONGO VALLEY
14074|MORONI
14075|MOROVIS
14076|MOROVIS ZONA URBANA
14077|MORRAL
14078|MORRICE
14079|MORRILL
14080|MORRILTON
14081|MORRIS
14082|MORRIS PLAINS
14083|MORRIS RANCH
14084|MORRISDALE
14085|MORRISON
14086|MORRISON BLUFF
14087|MORRISON CROSSROAD
14088|MORRISONVILLE
14089|MORRISTON
14090|MORRISTOWN
14091|MORRISVILLE
14092|MORRO BAY
14093|MORROW
14094|MORROWVILLE
14095|MORSE
14096|MORSE BLUFF
14097|MORSE JUNCTION
14098|MORSTEIN
14099|MORTMAR
14100|MORTON
14101|MORTON GROVE
14102|MORTON MILLS
14103|MORTON VALLEY
14104|MORTONS GAP
14105|MORTONSVILLE
14106|MORVEN
14107|MORZHOVOI
14108|MOSBY
14109|MOSCA
14110|MOSCOW
14111|MOSCOW MILLS
14112|MOSELEY
14113|MOSELLE
14114|MOSES LAKE
14115|MOSHANNON
14116|MOSHEIM
14117|MOSHER
14118|MOSIER
14119|MOSINEE
14120|MOSQUERO
14121|MOSQUITO LAKE
14122|MOSS
14123|MOSS BEACH
14124|MOSS BLUFF
14125|MOSS HILL
14126|MOSS LANDING
14127|MOSS POINT
14128|MOSSES
14129|MOSSVILLE
14130|MOSSY HEAD
14131|MOSSYROCK
14132|MOTLEY
14133|MOTT
14134|MOULTON
14135|MOULTON HEIGHTS
14136|MOULTRIE
14137|MOUND
14138|MOUND BAYOU
14139|MOUND CITY
14140|MOUND VALLEY
14141|MOUNDRIDGE
14142|MOUNDS
14143|MOUNDS VIEW
14144|MOUNDSVILLE
14145|MOUNDVILLE
14146|MOUNT AETNA
14147|MOUNT AIRY
14148|MOUNT ANDREW
14149|MOUNT ANGEL
14150|MOUNT ARLINGTON
14151|MOUNT AUBURN
14152|MOUNT AYR
14153|MOUNT BALDY
14154|MOUNT BETHEL
14155|MOUNT BLANCHARD
14156|MOUNT BRIAR
14157|MOUNT CALM
14158|MOUNT CALVARY
14159|MOUNT CARBON
14160|MOUNT CARMEL
14161|MOUNT CARROLL
14162|MOUNT CHARLESTON
14163|MOUNT CLARE
14164|MOUNT CLEMENS
14165|MOUNT COBB
14166|MOUNT CORY
14167|MOUNT CRAWFORD
14168|MOUNT CRESTED BUTTE
14169|MOUNT CROGHAN
14170|MOUNT DORA
14171|MOUNT EAGLE
14172|MOUNT EATON
14173|MOUNT EDEN
14174|MOUNT ENTERPRISE
14175|MOUNT EPHRAIM
14176|MOUNT ERIE
14177|MOUNT ETNA
14178|MOUNT FERN
14179|MOUNT FREEDOM
14180|MOUNT GILEAD
14181|MOUNT GRETNA
14182|MOUNT GRETNA HEIGHTS
14183|MOUNT HAMILL
14184|MOUNT HARMONY
14185|MOUNT HEALTHY
14186|MOUNT HEALTHY HEIGHTS
14187|MOUNT HEBRON
14188|MOUNT HERMON
14189|MOUNT HOLLY
14190|MOUNT HOLLY SPRINGS
14191|MOUNT HOOD
14192|MOUNT HOOD VILLAGE
14193|MOUNT HOPE
14194|MOUNT HOREB
14195|MOUNT HOUSTON
14196|MOUNT IDA
14197|MOUNT IVY
14198|MOUNT JACKSON
14199|MOUNT JEWETT
14200|MOUNT JOY
14201|MOUNT JUDEA
14202|MOUNT JULIET
14203|MOUNT KISCO
14204|MOUNT LAGUNA
14205|MOUNT LAUREL
14206|MOUNT LEBANON
14207|MOUNT LENA
14208|MOUNT LEONARD
14209|MOUNT LIBERTY
14210|MOUNT MONTGOMERY
14211|MOUNT MORIAH
14212|MOUNT MORRIS
14213|MOUNT NEBO
14214|MOUNT OLIVE
14215|MOUNT OLIVER
14216|MOUNT OLIVET
14217|MOUNT ORAB
14218|MOUNT PENN
14219|MOUNT PLEASANT
14220|MOUNT PLEASANT MILLS
14221|MOUNT PLYMOUTH
14222|MOUNT POCONO
14223|MOUNT PROSPECT
14224|MOUNT PULASKI
14225|MOUNT RAINIER
14226|MOUNT REPOSE
14227|MOUNT ROSE
14228|MOUNT ROYAL
14229|MOUNT SAVAGE
14230|MOUNT SELMAN
14231|MOUNT SHASTA
14232|MOUNT SIDNEY
14233|MOUNT SINAI
14234|MOUNT SOLON
14235|MOUNT STERLING
14236|MOUNT STORM
14237|MOUNT SUMMIT
14238|MOUNT TABOR
14239|MOUNT TRUMBULL
14240|MOUNT UNION
14241|MOUNT UPTON
14242|MOUNT VERNON
14243|MOUNT VICTORY
14244|MOUNT VISTA
14245|MOUNT WASHINGTON
14246|MOUNT WOLF
14247|MOUNT ZION
14248|MOUNTAIN
14249|MOUNTAIN BROOK
14250|MOUNTAIN CENTER
14251|MOUNTAIN CITY
14252|MOUNTAIN CREEK
14253|MOUNTAIN GATE
14254|MOUNTAIN GREEN
14255|MOUNTAIN GROVE
14256|MOUNTAIN HOME
14257|MOUNTAIN HOUSE
14258|MOUNTAIN IRON
14259|MOUNTAIN LAKE
14260|MOUNTAIN LAKE PARK
14261|MOUNTAIN LAKES
14262|MOUNTAIN LODGE PARK
14263|MOUNTAIN MEADOWS
14264|MOUNTAIN MESA
14265|MOUNTAIN PARK
14266|MOUNTAIN PINE
14267|MOUNTAIN RANCH
14268|MOUNTAIN ROAD
14269|MOUNTAIN TOP
14270|MOUNTAIN VALLEY
14271|MOUNTAIN VIEW
14272|MOUNTAIN VIEW ACRES
14273|MOUNTAIN VILLAGE
14274|MOUNTAINAIR
14275|MOUNTAINAIRE
14276|MOUNTAINBURG
14277|MOUNTAINHOME
14278|MOUNTAINSIDE
14279|MOUNTLAKE TERRACE
14280|MOUNTVILLE
14281|MOUSER
14282|MOUSIE
14283|MOUTH OF WILSON
14284|MOVICO
14285|MOVILLE
14286|MOWEAQUA
14287|MOWRYSTOWN
14288|MOXAHALA
14289|MOXEE CITY
14290|MOXLEY
14291|MOYERS
14292|MOYIE SPRINGS
14293|MOYLAN
14294|MOYOCK
14295|MOZELLE
14296|MUCARABONES
14297|MUCARABONES COMUNIDAD
14298|MUD BAY
14299|MUD BUTTE
14300|MUD LAKE
14301|MUDDY
14302|MUDDY GAP
14303|MUENSTER
14304|MUHLENBERG PARK
14305|MUIR
14306|MUIR BEACH
14307|MUKILTEO
14308|MUKWONAGO
14309|MULAT
14310|MULBERRY
14311|MULBERRY GROVE
14312|MULDOON
14313|MULDRAUGH
14314|MULDROW
14315|MULE CREEK
14316|MULESHOE
14317|MULFORD
14318|MULGA
14319|MULHALL
14320|MULINO
14321|MULKEYTOWN
14322|MULLAN
14323|MULLEN
14324|MULLENS
14325|MULLICA HILL
14326|MULLIKEN
14327|MULLIN
14328|MULLINS
14329|MULLINVILLE
14330|MULVANE
14331|MUMFORD
14332|MUNCIE
14333|MUNCY
14334|MUNDAY
14335|MUNDELEIN
14336|MUNDEN
14337|MUNDS PARK
14338|MUNDYS CORNER
14339|MUNFORD
14340|MUNFORDVILLE
14341|MUNGER
14342|MUNHALL
14343|MUNICH
14344|MUNISING
14345|MUNIZ
14346|MUNJOR
14347|MUNNERLYN
14348|MUNNSVILLE
14349|MUNROE FALLS
14350|MUNSEY PARK
14351|MUNSON
14352|MUNSONS CORNERS
14353|MUNSTER
14354|MURCHISON
14355|MURDO
14356|MURDOCK
14357|MURFREESBORO
14358|MURILLO COLONIA
14359|MURPHY
14360|MURPHY CITY
14361|MURPHYS
14362|MURPHYS CORNER
14363|MURPHYS ESTATES
14364|MURPHYSBORO
14365|MURPHYTOWN
14366|MURRAY
14367|MURRAY CITY
14368|MURRAY HILL
14369|MURRAYSVILLE
14370|MURRAYVILLE
14371|MURRELLS INLET
14372|MURRIETA
14373|MURRY HILL
14374|MURRYSVILLE
14375|MURTAUGH
14376|MUSCATINE
14377|MUSCLE SHOALS
14378|MUSCODA
14379|MUSCOTAH
14380|MUSCOY
14381|MUSE
14382|MUSELLA
14383|MUSICKS FERRY
14384|MUSKEGO
14385|MUSKEGON
14386|MUSKEGON HEIGHTS
14387|MUSKOGEE
14388|MUSSELSHELL
14389|MUSTANG
14390|MUSTANG RIDGE
14391|MUSTOE
14392|MUTTONTOWN
14393|MUTUAL
14394|MYAKKA CITY
14395|MYERS
14396|MYERS CORNER
14397|MYERS FLAT
14398|MYERSTOWN
14399|MYERSVILLE
14400|MYLO
14401|MYNARD
14402|MYOMA
14403|MYRA
14404|MYRICK
14405|MYRON
14406|MYRTLE
14407|MYRTLE BEACH
14408|MYRTLE CREEK
14409|MYRTLE GROVE
14410|MYRTLE POINT
14411|MYRTLE SPRINGS
14412|MYRTLETOWN
14413|MYRTLEWOOD
14414|MYSTIC
14415|MYSTIC ISLAND
14416|MYTON
14417|MĀHUKONA
14418|MĀKAHA
14419|MĀKAHA VALLEY
14420|MĀKENA
14421|MĀNĀ
14422|MĀʻALAEA
14423|MĀʻILI
14424|NABB
14425|NABESNA
14426|NABNASSET
14427|NABORTON
14428|NACHES
14429|NACO
14430|NACOGDOCHES
14431|NADA
14432|NADINE
14433|NAGEEZI
14434|NAGS HEAD
14435|NAGUABO
14436|NAGUABO ZONA URBANA
14437|NAHANT
14438|NAHMA
14439|NAHUNTA
14440|NAIRN
14441|NAKAIBITO
14442|NAKNEK
14443|NALLEN
14444|NAMBE
14445|NAMEKAGON
14446|NAMPA
14447|NANAFALIA
14448|NANCES CREEK
14449|NANCY
14450|NANKIN
14451|NANSON
14452|NANTICOKE
14453|NANTICOKE ACRES
14454|NANTUCKET
14455|NANTY GLO
14456|NANUET
14457|NANWALEK
14458|NAOMI
14459|NAPA
14460|NAPAKIAK
14461|NAPANOCH
14462|NAPASKIAK
14463|NAPAVINE
14464|NAPEAGUE
14465|NAPER
14466|NAPERVILLE
14467|NAPIER FIELD
14468|NAPLATE
14469|NAPLES
14470|NAPLES MANOR
14471|NAPLES PARK
14472|NAPOLEON
14473|NAPOLEONVILLE
14474|NAPONEE
14475|NAPPANEE
14476|NARA VISA
14477|NARANJA
14478|NARANJITO
14479|NARANJITO ZONA URBANA
14480|NARBERTH
14481|NARCISSA
14482|NARCISSO
14483|NARCOOSSEE
14484|NARDIN
14485|NARKA
14486|NAROD
14487|NARRAGANSETT PIER
14488|NARROWS
14489|NARROWSBURG
14490|NARUNA
14491|NASCHITTI
14492|NASELLE
14493|NASH
14494|NASHOBA
14495|NASHOTAH
14496|NASHUA
14497|NASHVILLE
14498|NASHWAUK
14499|NASON
14500|NASONVILLE
14501|NASSAU
14502|NASSAU BAY
14503|NASSAU SHORES
14504|NASSAWADOX
14505|NATALBANY
14506|NATALIA
14507|NATCHEZ
14508|NATCHITOCHES
14509|NATHALIE
14510|NATHAN
14511|NATIONAL
14512|NATIONAL CITY
14513|NATIONAL MINE
14514|NATIONAL PARK
14515|NATOMA
14516|NATRONA
14517|NATRONA HEIGHTS
14518|NATURAL BRIDGE
14519|NATURAL BRIDGE STATION
14520|NATURAL DAM
14521|NATURAL STEPS
14522|NATURITA
14523|NATWICK
14524|NAUBINWAY
14525|NAUGATUCK
14526|NAUKATI BAY
14527|NAUVOO
14528|NAVAJO
14529|NAVAJO DAM
14530|NAVAJO MOUNTAIN
14531|NAVARINO
14532|NAVARRE
14533|NAVARRO
14534|NAVASOTA
14535|NAVASSA
14536|NAVESINK
14537|NAVY YARD CITY
14538|NAYLOR
14539|NAYTAHWAUSH
14540|NAZARETH
14541|NAZLINI
14542|NEAH BAY
14543|NEAHKAHNIE
14544|NEAL
14545|NEAME
14546|NEAPOLIS
14547|NEAVITT
14548|NEBO
14549|NEBRASKA CITY
14550|NECEDAH
14551|NECHE
14552|NECHES
14553|NECK CITY
14554|NECTAR
14555|NEDERLAND
14556|NEDROW
14557|NEEDHAM
14558|NEEDLES
14559|NEEDMORE
14560|NEEDVILLE
14561|NEELY
14562|NEELYS LANDING
14563|NEELYVILLE
14564|NEENAH
14565|NEESES
14566|NEFFS
14567|NEGAUNEE
14568|NEGLEY
14569|NEGRA
14570|NEGREET
14571|NEHALEM
14572|NEHAWKA
14573|NEIBERT
14574|NEIHART
14575|NEILLSVILLE
14576|NEILTON
14577|NEKOMA
14578|NEKOOSA
14579|NELAGONEY
14580|NELCHINA
14581|NELIGH
14582|NELLIE
14583|NELLIEBURG
14584|NELLISTON
14585|NELLYSFORD
14586|NELSON
14587|NELSON LAGOON
14588|NELSONIA
14589|NELSONVILLE
14590|NEMACOLIN
14591|NEMAH
14592|NEMAHA
14593|NEMO
14594|NENAHNEZAD
14595|NENANA
14596|NENZEL
14597|NEODESHA
14598|NEOGA
14599|NEOLA
14600|NEOPIT
14601|NEOSHO
14602|NEOSHO FALLS
14603|NEOSHO RAPIDS
14604|NEPHI
14605|NEPONSET
14606|NEPTUNE
14607|NEPTUNE BEACH
14608|NEPTUNE CITY
14609|NERSTRAND
14610|NESBIT
14611|NESBITT
14612|NESCATUNGA
14613|NESCO
14614|NESCONSET
14615|NESCOPECK
14616|NESHAMINY
14617|NESHANIC STATION
14618|NESHKORO
14619|NESHOBA
14620|NESIKA BEACH
14621|NESKOWIN
14622|NESMITH
14623|NESPELEM
14624|NESQUEHONING
14625|NESS CITY
14626|NESSEN CITY
14627|NESTORIA
14628|NESTORVILLE
14629|NETARTS
14630|NETAWAKA
14631|NETCONG
14632|NETHERS
14633|NETT LAKE
14634|NETTIE
14635|NETTLE LAKE
14636|NETTLETON
14637|NEUBERT
14638|NEUSE
14639|NEUSE FOREST
14640|NEUVILLE
14641|NEVADA
14642|NEVADA CITY
14643|NEVILLE
14644|NEVINVILLE
14645|NEVIS
14646|NEW ALBANY
14647|NEW ALBIN
14648|NEW ALEXANDRIA
14649|NEW ALMELO
14650|NEW AMSTERDAM
14651|NEW ATHENS
14652|NEW AUBURN
14653|NEW AUGUSTA
14654|NEW BADEN
14655|NEW BALTIMORE
14656|NEW BAVARIA
14657|NEW BEAVER
14658|NEW BEDFORD
14659|NEW BERLIN
14660|NEW BERLINVILLE
14661|NEW BERN
14662|NEW BETHLEHEM
14663|NEW BLAINE
14664|NEW BLOOMFIELD
14665|NEW BLOOMINGTON
14666|NEW BOSTON
14667|NEW BRAUNFELS
14668|NEW BREMEN
14669|NEW BRIGHTON
14670|NEW BRITAIN
14671|NEW BROCKTON
14672|NEW BRUNSWICK
14673|NEW BUFFALO
14674|NEW BURLINGTON
14675|NEW BURNSIDE
14676|NEW CALIFORNIA
14677|NEW CAMBRIA
14678|NEW CANEY
14679|NEW CANTON
14680|NEW CARLISLE
14681|NEW CARROLLTON
14682|NEW CASSEL
14683|NEW CASTLE
14684|NEW CENTERVILLE
14685|NEW CHAPEL HILL
14686|NEW CHICAGO
14687|NEW CHURCH
14688|NEW CITY
14689|NEW COLUMBIA
14690|NEW COLUMBUS
14691|NEW CONCORD
14692|NEW COURT VILLAGE
14693|NEW CREEK
14694|NEW CUMBERLAND
14695|NEW CUYAMA
14696|NEW DEAL
14697|NEW DOUGLAS
14698|NEW EAGLE
14699|NEW EDINBURG
14700|NEW EFFINGTON
14701|NEW EGYPT
14702|NEW ELLENTON
14703|NEW ELLIOTT
14704|NEW ENGLAND
14705|NEW ERA
14706|NEW FAIRVIEW
14707|NEW FALCON
14708|NEW FLORENCE
14709|NEW FRANKEN
14710|NEW FRANKLIN
14711|NEW FREEDOM
14712|NEW FREEPORT
14713|NEW GALILEE
14714|NEW GERMANY
14715|NEW GLARUS
14716|NEW GOSHEN
14717|NEW GRAND CHAIN
14718|NEW HAMILTON
14719|NEW HAMPSHIRE
14720|NEW HAMPTON
14721|NEW HARMONY
14722|NEW HARTFORD
14723|NEW HAVEN
14724|NEW HEBRON
14725|NEW HEMPSTEAD
14726|NEW HOLLAND
14727|NEW HOLSTEIN
14728|NEW HOME
14729|NEW HOPE
14730|NEW HRADEC
14731|NEW HUDSON
14732|NEW HYDE PARK
14733|NEW IBERIA
14734|NEW JERUSALEM
14735|NEW JOHNSONVILLE
14736|NEW KENSINGTON
14737|NEW KENT
14738|NEW KINGSTOWN
14739|NEW KNOXVILLE
14740|NEW LAGUNA
14741|NEW LANCASTER
14742|NEW LEBANON
14743|NEW LEIPZIG
14744|NEW LENOX
14745|NEW LEXINGTON
14746|NEW LIBERTY
14747|NEW LISBON
14748|NEW LLANO
14749|NEW LONDON
14750|NEW LOTHROP
14751|NEW LYME STATION
14752|NEW MADISON
14753|NEW MADRID
14754|NEW MARKET
14755|NEW MARSHFIELD
14756|NEW MARTINSVILLE
14757|NEW MATAMORAS
14758|NEW MEADOWS
14759|NEW MELLE
14760|NEW MIAMI
14761|NEW MIDDLETOWN
14762|NEW MILFORD
14763|NEW MILTON
14764|NEW MINDEN
14765|NEW MORGAN
14766|NEW MUNICH
14767|NEW MUNSTER
14768|NEW ORLEANS
14769|NEW OXFORD
14770|NEW PALESTINE
14771|NEW PALTZ
14772|NEW PARIS
14773|NEW PEKIN
14774|NEW PETERSBURG
14775|NEW PHILADELPHIA
14776|NEW PINE CREEK
14777|NEW PITTSBURG
14778|NEW PLYMOUTH
14779|NEW POINT
14780|NEW PORT RICHEY
14781|NEW POST
14782|NEW PRAGUE
14783|NEW PRESTON
14784|NEW PROVIDENCE
14785|NEW RAYMER
14786|NEW RICHLAND
14787|NEW RICHMOND
14788|NEW RIEGEL
14789|NEW RINGGOLD
14790|NEW RIVER
14791|NEW ROADS
14792|NEW ROCHELLE
14793|NEW ROCKFORD
14794|NEW ROME
14795|NEW ROSS
14796|NEW SALEM
14797|NEW SALISBURY
14798|NEW SARPY
14799|NEW SEABURY
14800|NEW SHARON
14801|NEW SHEFFIELD
14802|NEW SITE
14803|NEW SMYRNA BEACH
14804|NEW SQUARE
14805|NEW STANTON
14806|NEW STRAITSVILLE
14807|NEW STRAWN
14808|NEW STUYAHOK
14809|NEW SUFFOLK
14810|NEW SUMMERFIELD
14811|NEW TAITON
14812|NEW TAZEWELL
14813|NEW TERRITORY
14814|NEW TOKEEN
14815|NEW TOWN
14816|NEW TRENTON
14817|NEW TRIER
14818|NEW TRIPOLI
14819|NEW TROY
14820|NEW ULM
14821|NEW UNDERWOOD
14822|NEW UNION
14823|NEW VERNON
14824|NEW VIENNA
14825|NEW VILLAGE
14826|NEW VIRGINIA
14827|NEW WASHINGTON
14828|NEW WASHOE CITY
14829|NEW WATERFORD
14830|NEW WAVERLY
14831|NEW WESTON
14832|NEW WHITELAND
14833|NEW WILLARD
14834|NEW WILMINGTON
14835|NEW WINDSOR
14836|NEW WOODSTOCK
14837|NEW WOODVILLE
14838|NEW YORK
14839|NEW YORK MILLS
14840|NEW ZION
14841|NEWALD
14842|NEWARK
14843|NEWARK VALLEY
14844|NEWAUKUM
14845|NEWAYGO
14846|NEWBERG
14847|NEWBERN
14848|NEWBERRY
14849|NEWBERRY SPRINGS
14850|NEWBORN
14851|NEWBURG
14852|NEWBURGH
14853|NEWBURGH HEIGHTS
14854|NEWBURN
14855|NEWBURY
14856|NEWBURYPORT
14857|NEWCASTLE
14858|NEWCOMB
14859|NEWCOMERSTOWN
14860|NEWDALE
14861|NEWELL
14862|NEWELLTON
14863|NEWFANE
14864|NEWFIELD
14865|NEWFIELDS
14866|NEWFOLDEN
14867|NEWFOUNDLAND
14868|NEWHALEM
14869|NEWHALEN
14870|NEWHALL
14871|NEWHOPE
14872|NEWINGTON
14873|NEWKIRK
14874|NEWLAND
14875|NEWLIN
14876|NEWLONSBURG
14877|NEWMAN
14878|NEWMAN GROVE
14879|NEWMAN LAKE
14880|NEWMANSTOWN
14881|NEWMARKET
14882|NEWNAN
14883|NEWPORT
14884|NEWPORT BEACH
14885|NEWPORT CENTER
14886|NEWPORT HILLS
14887|NEWPORT NEWS
14888|NEWPORTVILLE TERRACE
14889|NEWRY
14890|NEWSOME
14891|NEWSOMS
14892|NEWTOK
14893|NEWTON
14894|NEWTON FALLS
14895|NEWTON GROVE
14896|NEWTON HAMILTON
14897|NEWTONIA
14898|NEWTONSVILLE
14899|NEWTONVILLE
14900|NEWTOWN
14901|NEWTOWN GRANT
14902|NEWTOWN SQUARE
14903|NEWVILLE
14904|NEY
14905|NEYLANDVILLE
14906|NEZPERCE
14907|NIAGARA
14908|NIAGARA FALLS
14909|NIANGUA
14910|NIANTIC
14911|NIARADA
14912|NIBLEY
14913|NICASIO
14914|NICE
14915|NICEVILLE
14916|NICHOLASVILLE
14917|NICHOLLS
14918|NICHOLS
14919|NICHOLS HILLS
14920|NICHOLSON
14921|NICHOLVILLE
14922|NICKEL CREEK STATION
14923|NICKELSVILLE
14924|NICKERSON
14925|NICKSVILLE
14926|NICODEMUS
14927|NICOLAUS
14928|NICOLLET
14929|NICOMA PARK
14930|NICUT
14931|NIEDERWALD
14932|NIELSVILLE
14933|NIGHTHAWK
14934|NIGHTMUTE
14935|NIKEP
14936|NIKISKI
14937|NIKOLAEVSK
14938|NIKOLAI
14939|NIKOLSKI
14940|NILAND
14941|NILE
14942|NILES
14943|NILWOOD
14944|NIMMONS
14945|NIMROD
14946|NINA
14947|NINAVIEW
14948|NINE MILE FALLS
14949|NINETY SIX
14950|NINILCHIK
14951|NINNEKAH
14952|NINOCK
14953|NIOBE
14954|NIOBRARA
14955|NIOTA
14956|NIOTAZE
14957|NIPINNAWASEE
14958|NIPOMO
14959|NIPTON
14960|NISKAYUNA
14961|NISLAND
14962|NISQUALLY
14963|NISSEQUOGUE
14964|NISSWA
14965|NITER
14966|NITRO
14967|NITTA YUMA
14968|NITTANY
14969|NIULIʻI
14970|NIVERTON
14971|NIVERVILLE
14972|NIWOT
14973|NIXA
14974|NIXON
14975|NIXONS CROSSROADS
14976|NO NAME
14977|NOANK
14978|NOATAK
14979|NOBLE
14980|NOBLESTOWN
14981|NOBLESVILLE
14982|NOBLETON
14983|NOCATEE
14984|NOCONA
14985|NOCONA HILLS
14986|NODAWAY
14987|NOEL
14988|NOELKE
14989|NOGAL
14990|NOGALES
14991|NOHLY
14992|NOKESVILLE
14993|NOKOMIS
14994|NOLANVILLE
14995|NOLENSVILLE
14996|NOLIC
14997|NOMA
14998|NOME
14999|NONDALTON
15000|NOOKSACK
15001|NOONAN
15002|NOONDAY
15003|NOORVIK
15004|NOPAL
15005|NORA
15006|NORA SPRINGS
15007|NORBECK
15008|NORBORNE
15009|NORBOURNE ESTATES
15010|NORCATUR
15011|NORCO
15012|NORCROSS
15013|NORD
15014|NORDEN
15015|NORDHEIM
15016|NORDLAND
15017|NORDMAN
15018|NORFLEET
15019|NORFOLK
15020|NORFORK
15021|NORGE
15022|NORIAS
15023|NORLINA
15024|NORMAN
15025|NORMAN PARK
15026|NORMANDY
15027|NORMANDY PARK
15028|NORMANGEE
15029|NORMANNA
15030|NORMANS
15031|NORMANTOWN
15032|NORPHLET
15033|NORRIDGE
15034|NORRIDGEWOCK
15035|NORRIE
15036|NORRIS
15037|NORRIS CITY
15038|NORRISTOWN
15039|NORSELAND
15040|NORSHOR JUNCTION
15041|NORTH
15042|NORTH ABINGTON
15043|NORTH ACOMITA VILLAGE
15044|NORTH ADAMS
15045|NORTH ALAMO
15046|NORTH ALBANY
15047|NORTH AMHERST
15048|NORTH AMITY
15049|NORTH AMITYVILLE
15050|NORTH ANDOVER
15051|NORTH APOLLO
15052|NORTH ARLINGTON
15053|NORTH ATLANTA
15054|NORTH ATTLEBORO
15055|NORTH AUBURN
15056|NORTH AUGUSTA
15057|NORTH AURORA
15058|NORTH BABYLON
15059|NORTH BALTIMORE
15060|NORTH BARRINGTON
15061|NORTH BAY
15062|NORTH BAY SHORE
15063|NORTH BAY VILLAGE
15064|NORTH BEACH
15065|NORTH BEACH HAVEN
15066|NORTH BELLE VERNON
15067|NORTH BELLINGHAM
15068|NORTH BELLMORE
15069|NORTH BELLPORT
15070|NORTH BEND
15071|NORTH BENNINGTON
15072|NORTH BERGEN
15073|NORTH BERWICK
15074|NORTH BETHESDA
15075|NORTH BIBB
15076|NORTH BILLERICA
15077|NORTH BLOOMFIELD
15078|NORTH BONNEVILLE
15079|NORTH BOSTON
15080|NORTH BRADDOCK
15081|NORTH BRANCH
15082|NORTH BRENTWOOD
15083|NORTH BROOKFIELD
15084|NORTH BROOKSVILLE
15085|NORTH BROWNING
15086|NORTH BUENA VISTA
15087|NORTH BUFFALO
15088|NORTH CALDWELL
15089|NORTH CANTON
15090|NORTH CAPE
15091|NORTH CAPE MAY
15092|NORTH CARROLLTON
15093|NORTH CATASAUQUA
15094|NORTH CHARLEROI
15095|NORTH CHARLESTON
15096|NORTH CHELMSFORD
15097|NORTH CHEVY CHASE
15098|NORTH CHICAGO
15099|NORTH CHILI
15100|NORTH CITY
15101|NORTH CLEVELAND
15102|NORTH COHASSET
15103|NORTH COLLEGE HILL
15104|NORTH COLLINS
15105|NORTH CONWAY
15106|NORTH CORBIN
15107|NORTH COURTLAND
15108|NORTH COWDEN
15109|NORTH CREEK
15110|NORTH CROSSETT
15111|NORTH CROWS NEST
15112|NORTH DECATUR
15113|NORTH DELAND
15114|NORTH DRUID HILLS
15115|NORTH EAGLE BUTTE
15116|NORTH EAST
15117|NORTH EAST CARRY
15118|NORTH EASTHAM
15119|NORTH EATON
15120|NORTH EDWARDS
15121|NORTH EL MONTE
15122|NORTH ENGLISH
15123|NORTH ENID
15124|NORTH EPWORTH
15125|NORTH ESCOBARES
15126|NORTH EVANS
15127|NORTH FAIR OAKS
15128|NORTH FAIRFIELD
15129|NORTH FALMOUTH
15130|NORTH FOND DU LAC
15131|NORTH FORK
15132|NORTH FORT MYERS
15133|NORTH FOSTER
15134|NORTH FREEDOM
15135|NORTH GATES
15136|NORTH GLEN ELLYN
15137|NORTH GRANBY
15138|NORTH GREAT RIVER
15139|NORTH GROSVENOR DALE
15140|NORTH HALEDON
15141|NORTH HAMPTON
15142|NORTH HANOVER
15143|NORTH HARTLAND
15144|NORTH HARTSVILLE
15145|NORTH HAVEN
15146|NORTH HAVERHILL
15147|NORTH HENDERSON
15148|NORTH HIGH SHOALS
15149|NORTH HIGHLANDS
15150|NORTH HILL
15151|NORTH HILLS
15152|NORTH HODGE
15153|NORTH HORNELL
15154|NORTH HOUSTON
15155|NORTH HUDSON
15156|NORTH HURLEY
15157|NORTH INDUSTRY
15158|NORTH IRWIN
15159|NORTH JOHNS
15160|NORTH JUDSON
15161|NORTH KANSAS CITY
15162|NORTH KENSINGTON
15163|NORTH KEY LARGO
15164|NORTH KINGSVILLE
15165|NORTH KOMELIK
15166|NORTH LA JUNTA
15167|NORTH LAKEVILLE
15168|NORTH LAS VEGAS
15169|NORTH LAUDERDALE
15170|NORTH LAUREL
15171|NORTH LAWRENCE
15172|NORTH LEWISBURG
15173|NORTH LIBERTY
15174|NORTH LILBOURN
15175|NORTH LIMA
15176|NORTH LINDENHURST
15177|NORTH LITTLE ROCK
15178|NORTH LOGAN
15179|NORTH LOUP
15180|NORTH LYNBROOK
15181|NORTH LYNNWOOD
15182|NORTH MADISON
15183|NORTH MANCHESTER
15184|NORTH MANITOU
15185|NORTH MANKATO
15186|NORTH MARSHFIELD
15187|NORTH MARYSVILLE
15188|NORTH MASSAPEQUA
15189|NORTH MERRICK
15190|NORTH MIAMI
15191|NORTH MIAMI BEACH
15192|NORTH MIDDLETOWN
15193|NORTH MUSKEGON
15194|NORTH MYRTLE BEACH
15195|NORTH NAPLES
15196|NORTH NEW HYDE PARK
15197|NORTH NEWTON
15198|NORTH OAKS
15199|NORTH OGDEN
15200|NORTH OLMSTED
15201|NORTH OMAK
15202|NORTH PALM BEACH
15203|NORTH PARK
15204|NORTH PATCHOGUE
15205|NORTH PEARSALL
15206|NORTH PEKIN
15207|NORTH PEMBROKE
15208|NORTH PERRY
15209|NORTH PHILIPSBURG
15210|NORTH PLAINFIELD
15211|NORTH PLAINS
15212|NORTH PLATTE
15213|NORTH PLYMOUTH
15214|NORTH POLE
15215|NORTH PORT
15216|NORTH POTOMAC
15217|NORTH POWDER
15218|NORTH PRAIRIE
15219|NORTH PUYALLUP
15220|NORTH RANDALL
15221|NORTH REDINGTON BEACH
15222|NORTH REDWOOD
15223|NORTH RICHLAND HILLS
15224|NORTH RICHMOND
15225|NORTH RIDGE
15226|NORTH RIDGEVILLE
15227|NORTH RIM
15228|NORTH RIVER
15229|NORTH RIVER SHORES
15230|NORTH RIVERSIDE
15231|NORTH ROBINSON
15232|NORTH ROBY
15233|NORTH ROCK SPRINGS
15234|NORTH ROSE
15235|NORTH ROYALTON
15236|NORTH SAINT PAUL
15237|NORTH SALEM
15238|NORTH SALT LAKE
15239|NORTH SAN JUAN
15240|NORTH SAN PEDRO
15241|NORTH SAN YSIDRO
15242|NORTH SARASOTA
15243|NORTH SCITUATE
15244|NORTH SEA
15245|NORTH SEEKONK
15246|NORTH SHORE
15247|NORTH SIOUX CITY
15248|NORTH SPRINGFIELD
15249|NORTH STRATFORD
15250|NORTH SUDBURY
15251|NORTH SULTAN
15252|NORTH SUTTON
15253|NORTH SYRACUSE
15254|NORTH TERRE HAUTE
15255|NORTH TEWKSBURY
15256|NORTH TONAWANDA
15257|NORTH TOPSAIL BEACH
15258|NORTH TROY
15259|NORTH TRURO
15260|NORTH TUNICA
15261|NORTH TUSTIN
15262|NORTH VACHERIE
15263|NORTH VALLEY
15264|NORTH VALLEY STREAM
15265|NORTH VANDERGRIFT
15266|NORTH VERNON
15267|NORTH WALES
15268|NORTH WALPOLE
15269|NORTH WANTAGH
15270|NORTH WARREN
15271|NORTH WASHINGTON
15272|NORTH WATERFORD
15273|NORTH WEBSTER
15274|NORTH WESTMINSTER
15275|NORTH WESTPORT
15276|NORTH WHITE PLAINS
15277|NORTH WILDWOOD
15278|NORTH WILKESBORO
15279|NORTH WILMINGTON
15280|NORTH WINDHAM
15281|NORTH WOLCOTT
15282|NORTH WOODSTOCK
15283|NORTH YELM
15284|NORTH YORK
15285|NORTH ZANESVILLE
15286|NORTH ZULCH
15287|NORTHAMPTON
15288|NORTHBORO
15289|NORTHBOROUGH
15290|NORTHBRANCH
15291|NORTHBROOK
15292|NORTHCOTE
15293|NORTHCREST
15294|NORTHDALE
15295|NORTHERN CAMBRIA
15296|NORTHFIELD
15297|NORTHFIELD CENTER
15298|NORTHFORK
15299|NORTHGATE
15300|NORTHGLENN
15301|NORTHLAKE
15302|NORTHLAKES
15303|NORTHLAND
15304|NORTHMOOR
15305|NORTHOME
15306|NORTHPORT
15307|NORTHRIDGE
15308|NORTHROP
15309|NORTHUMBERLAND
15310|NORTHVALE
15311|NORTHVIEW
15312|NORTHVILLE
15313|NORTHVUE
15314|NORTHWAY
15315|NORTHWAY JUNCTION
15316|NORTHWAY VILLAGE
15317|NORTHWEST
15318|NORTHWEST HARBOR
15319|NORTHWOOD
15320|NORTHWOODS
15321|NORTHWOODS BEACH
15322|NORTHWYE
15323|NORTON
15324|NORTON SHORES
15325|NORTONVILLE
15326|NORVELT
15327|NORWALK
15328|NORWAY
15329|NORWICH
15330|NORWOOD
15331|NORWOOD COURT
15332|NORWOOD YOUNG AMERICA
15333|NOTASULGA
15334|NOTCHIETOWN
15335|NOTIECHTOWN
15336|NOTREES
15337|NOTTOWAY COURT HOUSE
15338|NOTUS
15339|NOUGH
15340|NOUNAN
15341|NOVA
15342|NOVATO
15343|NOVELTY
15344|NOVI
15345|NOVICE
15346|NOVINGER
15347|NOWATA
15348|NOWLIN
15349|NOWTHEN
15350|NOXAPATER
15351|NOXEN
15352|NOXON
15353|NOYACK
15354|NOYES
15355|NUANGOLA
15356|NUBIEBER
15357|NUCLA
15358|NUEVO
15359|NUIQSUT
15360|NULATO
15361|NUMA
15362|NUMIDIA
15363|NUNAKA VALLEY
15364|NUNAM IQUA
15365|NUNAPITCHUK
15366|NUNDA
15367|NUNEZ
15368|NUNN
15369|NUNNELLY
15370|NUREMBERG
15371|NUSHAGAK
15372|NUTLEY
15373|NUTRIOSO
15374|NUTT
15375|NUTTER FORT
15376|NUTTING LAKE
15377|NUYAKA
15378|NYAC
15379|NYACK
15380|NYE
15381|NYSSA
15382|NĀNĀKULI
15383|NĀNĀWALE ESTATES
15384|NĀʻĀLEHU
15385|O'BRIEN
15386|O'DONNELL
15387|O'FALLON
15388|O'KEAN
15389|O'NEALS
15390|O'NEILL
15391|OACOMA
15392|OAK
15393|OAK BEACH
15394|OAK BROOK
15395|OAK CITY
15396|OAK CREEK
15397|OAK FOREST
15398|OAK GLEN
15399|OAK GROVE
15400|OAK GROVE HEIGHTS
15401|OAK GROVE VILLAGE
15402|OAK HALL
15403|OAK HARBOR
15404|OAK HILL
15405|OAK HILLS
15406|OAK HILLS PLACE
15407|OAK ISLAND
15408|OAK LAWN
15409|OAK LEAF
15410|OAK LEVEL
15411|OAK PARK
15412|OAK PARK HEIGHTS
15413|OAK POINT
15414|OAK RIDGE
15415|OAK RIDGE NORTH
15416|OAK RUN
15417|OAK SPRINGS
15418|OAK TRAIL SHORES
15419|OAK VALE
15420|OAK VALLEY
15421|OAK VIEW
15422|OAKBORO
15423|OAKBROOK
15424|OAKBROOK TERRACE
15425|OAKDALE
15426|OAKES
15427|OAKESDALE
15428|OAKFIELD
15429|OAKFORD
15430|OAKGROVE
15431|OAKHAVEN
15432|OAKHURST
15433|OAKLAND
15434|OAKLAND ACRES
15435|OAKLAND CITY
15436|OAKLAND HEIGHTS
15437|OAKLAND PARK
15438|OAKLEY
15439|OAKLEY PARK
15440|OAKLYN
15441|OAKMAN
15442|OAKMONT
15443|OAKPARK
15444|OAKRIDGE
15445|OAKS
15446|OAKSHADE
15447|OAKTON
15448|OAKTOWN
15449|OAKVALE
15450|OAKVIEW
15451|OAKVILLE
15452|OAKWOOD
15453|OAKWOOD HILLS
15454|OAKWOOD MANOR
15455|OAKWOOD PARK
15456|OARK
15457|OASIS
15458|OATFIELD
15459|OATMAN
15460|OBAR
15461|OBERLIN
15462|OBERON
15463|OBERT
15464|OBETZ
15465|OBION
15466|OBLONG
15467|OCALA
15468|OCATE
15469|OCCIDENTAL
15470|OCCOQUAN
15471|OCEAN
15472|OCEAN ACRES
15473|OCEAN BEACH
15474|OCEAN BLUFF
15475|OCEAN BREEZE PARK
15476|OCEAN CITY
15477|OCEAN GATE
15478|OCEAN GROVE
15479|OCEAN ISLE BEACH
15480|OCEAN PARK
15481|OCEAN PINES
15482|OCEAN RIDGE
15483|OCEAN SHORES
15484|OCEAN SPRINGS
15485|OCEAN VIEW
15486|OCEANA
15487|OCEANO
15488|OCEANPORT
15489|OCEANSIDE
15490|OCEE
15491|OCEOLA
15492|OCHELATA
15493|OCHEYEDAN
15494|OCHLOCKNEE
15495|OCHOA
15496|OCHOPEE
15497|OCILLA
15498|OCOEE
15499|OCONEE
15500|OCONOMOWOC
15501|OCONOMOWOC LAKE
15502|OCONTO
15503|OCONTO FALLS
15504|OCOTILLO
15505|OCRACOKE
15506|OCTA
15507|OCTAVIA
15508|ODANAH
15509|ODEBOLT
15510|ODELL
15511|ODEM
15512|ODEN
15513|ODENTON
15514|ODENVILLE
15515|ODESSA
15516|ODESSADALE
15517|ODIN
15518|ODON
15519|ODUM
15520|OELRICHS
15521|OELWEIN
15522|OFFERLE
15523|OFFERMAN
15524|OGALLAH
15525|OGALLALA
15526|OGDEN
15527|OGDEN DUNES
15528|OGDENSBURG
15529|OGEMA
15530|OGEMAW
15531|OGG
15532|OGILBY
15533|OGILVIE
15534|OGLALA
15535|OGLESBY
15536|OGLETHORPE
15537|OGLETOWN
15538|OHATCHEE
15539|OHIO
15540|OHIO CITY
15541|OHIOPYLE
15542|OHIOVILLE
15543|OHIOWA
15544|OHLMAN
15545|OHOOPEE
15546|OHOP
15547|OIL CITY
15548|OIL TROUGH
15549|OILDALE
15550|OILMONT
15551|OILTON
15552|OJAI
15553|OJO AMARILLO
15554|OJO CALIENTE
15555|OJO FELIZ
15556|OJO SARCO
15557|OJUS
15558|OKABENA
15559|OKAHUMPKA
15560|OKANOGAN
15561|OKARCHE
15562|OKATON
15563|OKAUCHEE
15564|OKAUCHEE LAKE
15565|OKAWVILLE
15566|OKEANA
15567|OKEECHOBEE
15568|OKEELANTA
15569|OKEENE
15570|OKEMAH
15571|OKEMOS
15572|OKETO
15573|OKLAHOMA
15574|OKLAHOMA CITY
15575|OKLAUNION
15576|OKLEE
15577|OKMULGEE
15578|OKOBOJI
15579|OKOLONA
15580|OKREEK
15581|OKTAHA
15582|OLA
15583|OLALLA
15584|OLAMON
15585|OLANCHA
15586|OLANTA
15587|OLAR
15588|OLATHE
15589|OLATON
15590|OLBERG
15591|OLCOTT
15592|OLD AGENCY
15593|OLD APPLETON
15594|OLD BENNINGTON
15595|OLD BETHPAGE
15596|OLD BRIDGE
15597|OLD BROOKVILLE
15598|OLD BROWNSBORO PLACE
15599|OLD EUCHA
15600|OLD FIELD
15601|OLD FIELDS
15602|OLD FORGE
15603|OLD FORT
15604|OLD GLORY
15605|OLD GREENWICH
15606|OLD HARBOR
15607|OLD HUNDRED
15608|OLD JEFFERSON
15609|OLD LEXINGTON
15610|OLD MILL CREEK
15611|OLD MINES
15612|OLD MINTO
15613|OLD MONROE
15614|OLD MYSTIC
15615|OLD OCEAN
15616|OLD ORCHARD
15617|OLD ORCHARD BEACH
15618|OLD RIPLEY
15619|OLD RIVER-WINFREE
15620|OLD SHAWNEETOWN
15621|OLD STATION
15622|OLD TAPPAN
15623|OLD TOWN
15624|OLD WASHINGTON
15625|OLD WESTBURY
15626|OLDE WEST CHESTER
15627|OLDEN
15628|OLDENBURG
15629|OLDHAM
15630|OLDS
15631|OLDSMAR
15632|OLDTOWN
15633|OLEAN
15634|OLENA
15635|OLENE
15636|OLEX
15637|OLEY
15638|OLGA
15639|OLIMPO
15640|OLIMPO COMUNIDAD
15641|OLIN
15642|OLIVAREZ
15643|OLIVE
15644|OLIVE BRANCH
15645|OLIVE HILL
15646|OLIVEHURST
15647|OLIVER
15648|OLIVER SPRINGS
15649|OLIVET
15650|OLIVETTE
15651|OLIVIA
15652|OLLA
15653|OLLIE
15654|OLMITO
15655|OLMITZ
15656|OLMOS PARK
15657|OLMSTEAD
15658|OLMSTED
15659|OLMSTED FALLS
15660|OLNES
15661|OLNEY
15662|OLNEY SPRINGS
15663|OLOWALU
15664|OLPE
15665|OLSBURG
15666|OLSONVILLE
15667|OLTON
15668|OLUSTEE
15669|OLVEY
15670|OLYMPIA
15671|OLYMPIA FIELDS
15672|OLYMPIA HEIGHTS
15673|OLYMPIAN VILLAGE
15674|OLYMPIC VIEW
15675|OLYPHANT
15676|OMA
15677|OMAHA
15678|OMAK
15679|OMAR
15680|OMEGA
15681|OMEMEE
15682|OMENA
15683|OMER
15684|OMO RANCH
15685|OMRO
15686|ONA
15687|ONAGA
15688|ONAKA
15689|ONALASKA
15690|ONAMIA
15691|ONANCOCK
15692|ONARGA
15693|ONAVA
15694|ONAWA
15695|ONAWAY
15696|ONEGO
15697|ONEIDA
15698|ONEIDA CASTLE
15699|ONEKAMA
15700|ONEONTA
15701|ONG
15702|ONIDA
15703|ONLEY
15704|ONO
15705|ONSET
15706|ONSLOW
15707|ONSTED
15708|ONTARIO
15709|ONTON
15710|ONTONAGON
15711|ONWARD
15712|ONYCHA
15713|ONYX
15714|OOLITIC
15715|OOLOGAH
15716|OOLTEWAH
15717|OOSTBURG
15718|OPA LOCKA
15719|OPA-LOCKA
15720|OPAL
15721|OPAL CLIFFS
15722|OPDYKE
15723|OPDYKE WEST
15724|OPELIKA
15725|OPELOUSAS
15726|OPHEIM
15727|OPHIR
15728|OPIHIKAO
15729|OPOLIS
15730|OPP
15731|OPPELO
15732|OPTIMO
15733|OQUAWKA
15734|OQUOSSOC
15735|ORACLE
15736|ORACLE JUNCTION
15737|ORADELL
15738|ORAIBI
15739|ORAN
15740|ORANGE
15741|ORANGE BEACH
15742|ORANGE CITY
15743|ORANGE COVE
15744|ORANGE GROVE
15745|ORANGE HEIGHTS
15746|ORANGE LAKE
15747|ORANGE PARK
15748|ORANGE PARK ACRES
15749|ORANGEBURG
15750|ORANGETREE
15751|ORANGEVALE
15752|ORANGEVILLE
15753|ORASON ACRES COLONIA
15754|ORBISONIA
15755|ORCAS
15756|ORCHARD
15757|ORCHARD BEACH
15758|ORCHARD CITY
15759|ORCHARD FARM
15760|ORCHARD GRASS HILLS
15761|ORCHARD HILL
15762|ORCHARD HILLS
15763|ORCHARD HOMES
15764|ORCHARD LAKE
15765|ORCHARD MESA
15766|ORCHARD PARK
15767|ORCHARD VALLEY
15768|ORCHARDS
15769|ORCHID
15770|ORCHIDLANDS ESTATES
15771|ORCUTT
15772|ORD
15773|ORDERVILLE
15774|ORDWAY
15775|ORE CITY
15776|OREANA
15777|OREGON
15778|OREGON CITY
15779|OREGONIA
15780|ORELAND
15781|OREM
15782|ORESTES
15783|ORETTA
15784|ORFORDVILLE
15785|ORGAN
15786|ORICK
15787|ORIENT
15788|ORIENT PARK
15789|ORIENTA
15790|ORIENTAL
15791|ORIN
15792|ORINDA
15793|ORIOLE BEACH
15794|ORION
15795|ORISKA
15796|ORISKANY
15797|ORISKANY FALLS
15798|ORLA
15799|ORLAND
15800|ORLAND HILLS
15801|ORLAND PARK
15802|ORLANDO
15803|ORLEANS
15804|ORLINDA
15805|ORLOVISTA
15806|ORME
15807|ORMOND BEACH
15808|ORMOND-BY-THE-SEA
15809|ORMSBY
15810|ORO GRANDE
15811|ORO VALLEY
15812|OROCOVIS
15813|OROCOVIS ZONA URBANA
15814|OROFINO
15815|OROGRANDE
15816|ORONO
15817|ORONOCO
15818|ORONOGO
15819|OROSI
15820|OROVADA
15821|OROVILLE
15822|ORPHA
15823|ORR
15824|ORRICK
15825|ORRIN
15826|ORRSTOWN
15827|ORRTANNA
15828|ORRUM
15829|ORRVILLE
15830|ORSON
15831|ORTING
15832|ORTLEY
15833|ORTONVILLE
15834|ORVISTON
15835|ORWELL
15836|ORWIGSBURG
15837|ORWIN
15838|OSAGE
15839|OSAGE BEACH
15840|OSAGE CITY
15841|OSAKIS
15842|OSAWATOMIE
15843|OSBORN
15844|OSBORNE
15845|OSBURN
15846|OSCARVILLE
15847|OSCEOLA
15848|OSCEOLA MILLS
15849|OSCODA
15850|OSCURA
15851|OSGOOD
15852|OSHKOSH
15853|OSHOTO
15854|OSIERFIELD
15855|OSINO
15856|OSKALOOSA
15857|OSKAWALIK
15858|OSLO
15859|OSMAN
15860|OSMOND
15861|OSNABROCK
15862|OSO
15863|OSPREY
15864|OSSEO
15865|OSSIAN
15866|OSSINEKE
15867|OSSINING
15868|OSSIPEE
15869|OSSUN
15870|OSTEEN
15871|OSTERDOCK
15872|OSTERVILLE
15873|OSTRANDER
15874|OSWAYO
15875|OSWEGO
15876|OSYKA
15877|OTAY
15878|OTEGO
15879|OTHELLO
15880|OTHO
15881|OTIS
15882|OTIS ORCHARDS
15883|OTISCO
15884|OTISVILLE
15885|OTLEY
15886|OTO
15887|OTOE
15888|OTRANTO
15889|OTSEGO
15890|OTSEGO LAKE
15891|OTTAWA
15892|OTTAWA HILLS
15893|OTTER
15894|OTTER CREEK
15895|OTTER LAKE
15896|OTTERBEIN
15897|OTTERTAIL
15898|OTTERVILLE
15899|OTTO
15900|OTTOSEN
15901|OTTOVILLE
15902|OTTUMWA
15903|OTTUSVILLE
15904|OTWAY
15905|OTWELL
15906|OUACHITA
15907|OUR TOWN
15908|OURAY
15909|OUTING
15910|OUTLOOK
15911|OUZINKIE
15912|OVAL
15913|OVALO
15914|OVANDO
15915|OVERBROOK
15916|OVERGAARD
15917|OVERLAND
15918|OVERLAND PARK
15919|OVERLEA
15920|OVERLY
15921|OVERPECK
15922|OVERTON
15923|OVETT
15924|OVID
15925|OVIEDO
15926|OVILLA
15927|OWANECO
15928|OWANKA
15929|OWASA
15930|OWASSO
15931|OWATONNA
15932|OWEGO
15933|OWENDALE
15934|OWENS
15935|OWENS CROSS ROADS
15936|OWENSBORO
15937|OWENSBURG
15938|OWENSVILLE
15939|OWENTON
15940|OWENTOWN
15941|OWENYO
15942|OWINGS
15943|OWINGS MILLS
15944|OWINGSVILLE
15945|OWL CREEK
15946|OWL RANCH
15947|OWOSSO
15948|OWYHEE
15949|OXBOW
15950|OXBOW ESTATES
15951|OXFORD
15952|OXFORD JUNCTION
15953|OXLY
15954|OXNARD
15955|OXON HILL
15956|OYEHUT
15957|OYENS
15958|OYLEN
15959|OYSTER BAY
15960|OYSTER BAY COVE
15961|OYSTER CREEK
15962|OYSTERVILLE
15963|OZAN
15964|OZARK
15965|OZAWKIE
15966|OZONA
15967|OZONE
15968|OZORA
15969|PABLO
15970|PACE
15971|PACHECO
15972|PACHUTA
15973|PACIFIC BEACH
15974|PACIFIC CITY
15975|PACIFIC GROVE
15976|PACIFIC JUNCTION
15977|PACIFICA
15978|PACKARD
15979|PACKWAUKEE
15980|PACKWOOD
15981|PACOLET
15982|PACOLET MILLS
15983|PADDOCK LAKE
15984|PADEN
15985|PADEN CITY
15986|PADERBORN
15987|PADONIA
15988|PADRONI
15989|PADUCAH
15990|PAGE
15991|PAGE CITY
15992|PAGE MANOR
15993|PAGE PARK
15994|PAGEDALE
15995|PAGELAND
15996|PAGETON
15997|PAGOSA JUNCTION
15998|PAGOSA SPRINGS
15999|PAGUATE
16000|PAHOKEE
16001|PAHRUMP
16002|PAICINES
16003|PAIGE
16004|PAINCOURTVILLE
16005|PAINESDALE
16006|PAINESVILLE
16007|PAINT
16008|PAINT BANK
16009|PAINT CREEK
16010|PAINT LICK
16011|PAINT ROCK
16012|PAINTED HILLS
16013|PAINTED POST
16014|PAINTER
16015|PAINTERSVILLE
16016|PAINTERTOWN
16017|PAINTSVILLE
16018|PAISANO PARK COLONIA
16019|PAISLEY
16020|PAJARITO
16021|PAJARO
16022|PAJONAL
16023|PAJONAL COMUNIDAD
16024|PALA
16025|PALACIOS
16026|PALATINE
16027|PALATINE BRIDGE
16028|PALATKA
16029|PALCO
16030|PALENVILLE
16031|PALERMO
16032|PALESTINE
16033|PALISADE
16034|PALISADES
16035|PALISADES PARK
16036|PALITO BLANCO
16037|PALM BAY
16038|PALM BEACH
16039|PALM BEACH GARDENS
16040|PALM BEACH SHORES
16041|PALM CITY
16042|PALM COAST
16043|PALM DESERT
16044|PALM DESERT COUNTRY
16045|PALM HARBOR
16046|PALM RIVER
16047|PALM SHORES
16048|PALM SPRINGS
16049|PALM VALLEY
16050|PALMAREJO
16051|PALMAREJO COMUNIDAD
16052|PALMAS
16053|PALMAS COMUNIDAD
16054|PALMAS DEL MAR
16055|PALMAS DEL MAR COMUNIDAD
16056|PALMDALE
16057|PALMER
16058|PALMER COMUNIDAD
16059|PALMER HEIGHTS
16060|PALMER LAKE
16061|PALMER PARK
16062|PALMERS CROSSING
16063|PALMERSVILLE
16064|PALMERTON
16065|PALMETTO
16066|PALMETTO BAY
16067|PALMETTO ESTATES
16068|PALMHURST
16069|PALMONA PARK
16070|PALMVIEW
16071|PALMYRA
16072|PALO
16073|PALO ALTO
16074|PALO CEDRO
16075|PALO PINTO
16076|PALO SECO
16077|PALO SECO COMUNIDAD
16078|PALO VERDE
16079|PALOMAR PARK
16080|PALOMAS
16081|PALOMAS COMUNIDAD
16082|PALOMINAS
16083|PALOS HEIGHTS
16084|PALOS HILLS
16085|PALOS PARK
16086|PALOS VERDES ESTATES
16087|PALOS VERDES PENINSULA
16088|PALOUSE
16089|PAMELIA CENTER
16090|PAMLICO BEACH
16091|PAMPA
16092|PAMPLICO
16093|PAMPLIN
16094|PANA
16095|PANACA
16096|PANACEA
16097|PANAMA
16098|PANAMA CITY
16099|PANAMA CITY BEACH
16100|PANCO
16101|PANCOASTBURG
16102|PANDORA
16103|PANGBURN
16104|PANGUITCH
16105|PANHANDLE
16106|PANOLA
16107|PANORA
16108|PANORAMA HEIGHTS
16109|PANORAMA PARK
16110|PANORAMA VILLAGE
16111|PANTANO
16112|PANTEGO
16113|PANTHER
16114|PANTHERSVILLE
16115|PANTOPS
16116|PAOLA
16117|PAOLI
16118|PAONIA
16119|PAPALOTE
16120|PAPILLION
16121|PAPINEAU
16122|PARACHUTE
16123|PARADE
16124|PARADIS
16125|PARADISE
16126|PARADISE BEACH
16127|PARADISE HEIGHTS
16128|PARADISE HILL
16129|PARADISE HILLS
16130|PARADISE PARK
16131|PARADISE VALLEY
16132|PARAGON
16133|PARAGON ESTATES
16134|PARAGONAH
16135|PARAGOULD
16136|PARAJE
16137|PARALOMA
16138|PARAMOUNT
16139|PARAMUS
16140|PARC
16141|PARCELAS DE NAVARRO COMUNIDAD
16142|PARCELAS LA MILAGROSA
16143|PARCELAS LA MILAGROSA COMUNIDAD
16144|PARCELAS MANDRY COMUNIDAD
16145|PARCELAS NUEVAS
16146|PARCELAS NUEVAS COMUNIDAD
16147|PARCELAS PEÑUELAS
16148|PARCELAS PEÑUELAS COMUNIDAD
16149|PARCELAS VIEJAS BORINQUEN COMUNIDAD
16150|PARCHMENT
16151|PARCOAL
16152|PARDEESVILLE
16153|PARDEEVILLE
16154|PARHAMS
16155|PARIS
16156|PARIS CROSSING
16157|PARISH
16158|PARISHVILLE
16159|PARK
16160|PARK CITY
16161|PARK CREST
16162|PARK FALLS
16163|PARK FOREST
16164|PARK FOREST VILLAGE
16165|PARK GROVE
16166|PARK HILL
16167|PARK HILLS
16168|PARK LAYNE
16169|PARK RAPIDS
16170|PARK RIDGE
16171|PARK RIVER
16172|PARK VALLEY
16173|PARK VIEW
16174|PARKDALE
16175|PARKER
16176|PARKER CITY
16177|PARKER CROSSROADS
16178|PARKER FORD
16179|PARKER SCHOOL
16180|PARKER STRIP
16181|PARKERFIELD
16182|PARKERS
16183|PARKERS PRAIRIE
16184|PARKERS SETTLEMENT
16185|PARKERSBURG
16186|PARKERTON
16187|PARKERTOWN
16188|PARKERVILLE
16189|PARKESBURG
16190|PARKFIELD
16191|PARKIN
16192|PARKLAND
16193|PARKLINE
16194|PARKMAN
16195|PARKS
16196|PARKSDALE
16197|PARKSIDE
16198|PARKSLEY
16199|PARKSTON
16200|PARKSVILLE
16201|PARKTON
16202|PARKVILLE
16203|PARKWAY
16204|PARKWAY VILLAGE
16205|PARKWOOD
16206|PARLIER
16207|PARLIN
16208|PARMA
16209|PARMA HEIGHTS
16210|PARMALEE
16211|PARMELE
16212|PARMELEE
16213|PARMERTON
16214|PARNELL
16215|PAROLE
16216|PARON
16217|PAROWAN
16218|PARRAL
16219|PARRAN
16220|PARRISH
16221|PARROTT
16222|PARROTTSVILLE
16223|PARRYVILLE
16224|PARSHALL
16225|PARSIPPANY
16226|PARSONS
16227|PARSONSBURG
16228|PARTHENON
16229|PARTRIDGE
16230|PASADENA
16231|PASADENA HILLS
16232|PASADENA PARK
16233|PASATIEMPO
16234|PASCAGOULA
16235|PASCO
16236|PASCOAG
16237|PASCOLA
16238|PASKENTA
16239|PASO ROBLES
16240|PASS CHRISTIAN
16241|PASSAIC
16242|PASSAPATANZY
16243|PASTORIA
16244|PASTOS
16245|PASTOS COMUNIDAD
16246|PASTURA
16247|PATAGONIA
16248|PATAHA
16249|PATASKALA
16250|PATCH GROVE
16251|PATCHOGUE
16252|PATEROS
16253|PATERSON
16254|PATESVILLE
16255|PATETOWN
16256|PATHFORK
16257|PATILLAS
16258|PATILLAS ZONA URBANA
16259|PATMOS
16260|PATOKA
16261|PATON
16262|PATRICIA
16263|PATRICK
16264|PATRICK SPRINGS
16265|PATRICKSBURG
16266|PATRIOT
16267|PATROON
16268|PATSVILLE
16269|PATTERSON
16270|PATTERSON HEIGHTS
16271|PATTERSON SPRINGS
16272|PATTISON
16273|PATTON
16274|PATTON VILLAGE
16275|PATTONSBURG
16276|PATTONVILLE
16277|PATZAU
16278|PAUKAA
16279|PAUL
16280|PAUL SMITHS
16281|PAUL SPUR
16282|PAULDEN
16283|PAULDING
16284|PAULETTE
16285|PAULINA
16286|PAULINE
16287|PAULLINA
16288|PAULS CROSSROADS
16289|PAULS VALLEY
16290|PAULSBORO
16291|PAULTON
16292|PAVILION
16293|PAVILLION
16294|PAVO
16295|PAW CREEK
16296|PAW PAW
16297|PAW PAW LAKE
16298|PAWCATUCK
16299|PAWHUSKA
16300|PAWLEYS ISLAND
16301|PAWLING
16302|PAWNEE
16303|PAWNEE CITY
16304|PAWNEE ROCK
16305|PAWNEE STATION
16306|PAWTUCKET
16307|PAX
16308|PAXICO
16309|PAXSON
16310|PAXTANG
16311|PAXTON
16312|PAXTONIA
16313|PAXTONVILLE
16314|PAXVILLE
16315|PAYETTE
16316|PAYNE
16317|PAYNE GAP
16318|PAYNE SPRINGS
16319|PAYNES
16320|PAYNES CREEK
16321|PAYNESVILLE
16322|PAYSON
16323|PAYTES
16324|PAʻAUILO
16325|PE ELL
16326|PEA RIDGE
16327|PEABODY
16328|PEACEFUL VALLEY
16329|PEACH CREEK
16330|PEACH LAKE
16331|PEACH ORCHARD
16332|PEACH SPRINGS
16333|PEACHBURG
16334|PEACHLAND
16335|PEACHTREE CITY
16336|PEACHTREE CORNERS
16337|PEACOCK
16338|PEAK
16339|PEAKS MILL
16340|PEAPACK
16341|PEARBLOSSOM
16342|PEARCE
16343|PEARCY
16344|PEARISBURG
16345|PEARL
16346|PEARL BEACH
16347|PEARL CITY
16348|PEARL RIVER
16349|PEARLAND
16350|PEARLINGTON
16351|PEARSALL
16352|PEARSON
16353|PEARSONVILLE
16354|PEASE
16355|PEASTER
16356|PEAVINE
16357|PEBBLE BEACH
16358|PEBBLE CREEK
16359|PECAN ACRES
16360|PECAN GAP
16361|PECAN GROVE
16362|PECAN HILL
16363|PECAN PLANTATION
16364|PECATONICA
16365|PECK
16366|PECKHAM
16367|PECKTONVILLE
16368|PECONIC
16369|PECOS
16370|PECULIAR
16371|PEDEN
16372|PEDERNAL
16373|PEDLEY
16374|PEDRICKTOWN
16375|PEDRO
16376|PEDRO BAY
16377|PEE DEE
16378|PEEBLES
16379|PEEKSKILL
16380|PEEL
16381|PEEPLES VALLEY
16382|PEERLESS
16383|PEETZ
16384|PEEVER
16385|PEGGS
16386|PEGRAM
16387|PEKIN
16388|PELAHATCHIE
16389|PELETIER
16390|PELHAM
16391|PELHAM MANOR
16392|PELICAN
16393|PELICAN BAY
16394|PELICAN LAKE
16395|PELICAN RAPIDS
16396|PELION
16397|PELKIE
16398|PELL CITY
16399|PELL LAKE
16400|PELLA
16401|PELLAND
16402|PELLETTOWN
16403|PELLSTON
16404|PELLVILLE
16405|PELZER
16406|PEMBERTON
16407|PEMBERTON HEIGHTS
16408|PEMBERVILLE
16409|PEMBERWICK
16410|PEMBINA
16411|PEMBINE
16412|PEMBROKE
16413|PEMBROKE PARK
16414|PEMBROKE PINES
16415|PEN ARGYL
16416|PEN MAR
16417|PENALOSA
16418|PENBROOK
16419|PENCE
16420|PENCER
16421|PENDER
16422|PENDERGRASS
16423|PENDLETON
16424|PENDLETON CENTER
16425|PENDROY
16426|PENELOPE
16427|PENERMON
16428|PENFIELD
16429|PENGILLY
16430|PENHOOK
16431|PENINSULA
16432|PENITAS
16433|PENN
16434|PENN ESTATES
16435|PENN LAKE PARK
16436|PENN VALLEY
16437|PENN WYNNE
16438|PENN YAN
16439|PENNDEL
16440|PENNEY FARMS
16441|PENNGROVE
16442|PENNINGTON
16443|PENNINGTON GAP
16444|PENNOCK
16445|PENNS CREEK
16446|PENNS GROVE
16447|PENNS NECK
16448|PENNSBORO
16449|PENNSBURG
16450|PENNSBURY VILLAGE
16451|PENNSIDE
16452|PENNSUCO
16453|PENNSVILLE
16454|PENNVILLE
16455|PENNWYN
16456|PENROSE
16457|PENRYN
16458|PENSACOLA
16459|PENTON
16460|PENTRESS
16461|PENTWATER
16462|PENWELL
16463|PENZANCE
16464|PEOA
16465|PEORIA
16466|PEORIA HEIGHTS
16467|PEOSTA
16468|PEOTONE
16469|PEP
16470|PEPEʻEKEO
16471|PEPIN
16472|PEPPER PIKE
16473|PEPPERELL
16474|PEPPERMILL VILLAGE
16475|PEQUANNOCK
16476|PEQUOP
16477|PEQUOT LAKES
16478|PERALTA
16479|PERCILLA
16480|PERCIVAL
16481|PERCLE
16482|PERCY
16483|PERDIDO
16484|PERDIDO BEACH
16485|PEREZ
16486|PEREZVILLE
16487|PERHAM
16488|PERIDOT
16489|PERINTOWN
16490|PERKASIE
16491|PERKINS
16492|PERKINSTON
16493|PERKINSVILLE
16494|PERLA
16495|PERLEY
16496|PERMA
16497|PERNELL
16498|PEROTE
16499|PERRIN
16500|PERRINE
16501|PERRINTON
16502|PERRIS
16503|PERRY
16504|PERRY HALL
16505|PERRY HEIGHTS
16506|PERRY PARK
16507|PERRYDALE
16508|PERRYMAN
16509|PERRYOPOLIS
16510|PERRYSBURG
16511|PERRYSVILLE
16512|PERRYTON
16513|PERRYTOWN
16514|PERRYVILLE
16515|PERSIA
16516|PERTH
16517|PERTH AMBOY
16518|PERU
16519|PESCADERO
16520|PESHASTIN
16521|PESHAWBESTOWN
16522|PESHTIGO
16523|PESOTUM
16524|PETAL
16525|PETALUMA
16526|PETERBOROUGH
16527|PETERMAN
16528|PETERS
16529|PETERSBURG
16530|PETERSHAM
16531|PETERSON
16532|PETERSTOWN
16533|PETERSVILLE
16534|PETOSKEY
16535|PETREY
16536|PETROLEUM
16537|PETROLIA
16538|PETRONILA
16539|PETROS
16540|PETTIBONE
16541|PETTIGREW
16542|PETTISVILLE
16543|PETTIT
16544|PETTRY
16545|PETTUS
16546|PETTY
16547|PEVELY
16548|PEWAMO
16549|PEWAUKEE
16550|PEWEE VALLEY
16551|PEYTON
16552|PEÑA BLANCA
16553|PEÑA POBRE
16554|PEÑA POBRE COMUNIDAD
16555|PEÑASCO
16556|PEÑUELAS
16557|PEÑUELAS ZONA URBANA
16558|PFEIFER
16559|PFLUGERVILLE
16560|PHARR
16561|PHEBA
16562|PHELAN
16563|PHELPS
16564|PHELPS CITY
16565|PHENIX
16566|PHENIX CITY
16567|PHIL CAMPBELL
16568|PHILADELPHIA
16569|PHILBROOK
16570|PHILIP
16571|PHILIPP
16572|PHILIPPI
16573|PHILIPSBURG
16574|PHILLIPS
16575|PHILLIPSBURG
16576|PHILLIPSTOWN
16577|PHILLIPSVILLE
16578|PHILMONT
16579|PHILO
16580|PHILOMATH
16581|PHIPPSBURG
16582|PHLOX
16583|PHOENICIA
16584|PHOENIX
16585|PHOENIX LAKE
16586|PHOENIXVILLE
16587|PICA
16588|PICABO
16589|PICACHO
16590|PICAYUNE
16591|PICK CITY
16592|PICKENS
16593|PICKENSVILLE
16594|PICKERING
16595|PICKERINGTON
16596|PICKETT
16597|PICKFORD
16598|PICKRELL
16599|PICKSTOWN
16600|PICKTON
16601|PICNIC POINT
16602|PICO RIVERA
16603|PICTURE ROCKS
16604|PICURIS PUEBLO
16605|PIDCOKE
16606|PIE TOWN
16607|PIEDMONT
16608|PIEDRA
16609|PIEDRA AGUZA COMUNIDAD
16610|PIEDRA GORDA
16611|PIEDRA GORDA COMUNIDAD
16612|PIERCE
16613|PIERCE CITY
16614|PIERCETON
16615|PIERCEVILLE
16616|PIERCY
16617|PIERMONT
16618|PIERPONT
16619|PIERRE
16620|PIERRE PART
16621|PIERREPONT MANOR
16622|PIERRON
16623|PIERSON
16624|PIERZ
16625|PIFFARD
16626|PIGEON
16627|PIGEON COVE
16628|PIGEON CREEK
16629|PIGEON FALLS
16630|PIGEON FORGE
16631|PIGEON RIVER
16632|PIGGOTT
16633|PIKE
16634|PIKE CITY
16635|PIKE CREEK
16636|PIKE CREEK VALLEY
16637|PIKE ROAD
16638|PIKE VIEW
16639|PIKES CREEK
16640|PIKESVILLE
16641|PIKETON
16642|PIKEVIEW
16643|PIKEVILLE
16644|PILAR
16645|PILGER
16646|PILGRIM
16647|PILLAGER
16648|PILLOW
16649|PILLSBURY
16650|PILOT GROVE
16651|PILOT HILL
16652|PILOT KNOB
16653|PILOT MOUND
16654|PILOT MOUNTAIN
16655|PILOT POINT
16656|PILOT ROCK
16657|PILOT STATION
16658|PILOTTOWN
16659|PILSEN
16660|PILTZVILLE
16661|PIMA
16662|PIMACO TWO
16663|PIMENTO
16664|PIMMIT HILLS
16665|PIN OAK ACRES
16666|PINAL
16667|PINARDVILLE
16668|PINCH
16669|PINCKARD
16670|PINCKNEY
16671|PINCKNEYVILLE
16672|PINCONNING
16673|PINDALL
16674|PINE
16675|PINE AIRE
16676|PINE APPLE
16677|PINE BARREN
16678|PINE BEACH
16679|PINE BEND
16680|PINE BLUFF
16681|PINE BLUFFS
16682|PINE BROOK
16683|PINE BROOK HILL
16684|PINE BUSH
16685|PINE CASTLE
16686|PINE CENTER
16687|PINE CITY
16688|PINE COVE
16689|PINE CREST
16690|PINE FLAT
16691|PINE FOREST
16692|PINE GLEN
16693|PINE GROVE
16694|PINE GROVE MILLS
16695|PINE HALL
16696|PINE HAVEN
16697|PINE HILL
16698|PINE HILLS
16699|PINE HOLLOW
16700|PINE ISLAND
16701|PINE ISLAND CENTER
16702|PINE ISLAND RIDGE
16703|PINE KNOLL SHORES
16704|PINE KNOT
16705|PINE LAKE
16706|PINE LAKE PARK
16707|PINE LAKES
16708|PINE LAKES ADDITION
16709|PINE LAWN
16710|PINE LEVEL
16711|PINE LOG
16712|PINE MANOR
16713|PINE MOUNTAIN
16714|PINE MOUNTAIN CLUB
16715|PINE MOUNTAIN VALLEY
16716|PINE ORCHARD
16717|PINE PARK
16718|PINE PLAINS
16719|PINE POINT
16720|PINE PRAIRIE
16721|PINE REST
16722|PINE RIDGE
16723|PINE RIDGE AT CRESTWOOD
16724|PINE RIVER
16725|PINE SPRINGS
16726|PINE VALLEY
16727|PINE VILLAGE
16728|PINEBLUFF
16729|PINECLIFFE
16730|PINECREEK
16731|PINECREST
16732|PINEDA
16733|PINEDALE
16734|PINEHILL
16735|PINEHURST
16736|PINELAND
16737|PINELLAS PARK
16738|PINEOLA
16739|PINEORA
16740|PINERIDGE
16741|PINESBURG
16742|PINESDALE
16743|PINETOP-LAKESIDE
16744|PINETOPS
16745|PINETOWN
16746|PINETTA
16747|PINEVIEW
16748|PINEVILLE
16749|PINEWOOD
16750|PINEWOOD ESTATES
16751|PINEY
16752|PINEY FORK
16753|PINEY GREEN
16754|PINEY PARK
16755|PINEY POINT
16756|PINEY POINT VILLAGE
16757|PINEY RIVER
16758|PINEY VIEW
16759|PINEY WOODS
16760|PINGREE
16761|PINGREE GROVE
16762|PINHOOK
16763|PINHOOK CORNER
16764|PINK
16765|PINK HILL
16766|PINKSTAFF
16767|PINLAND
16768|PINNACLE
16769|PINOLA
16770|PINOLE
16771|PINON
16772|PINOPOLIS
16773|PINOS ALTOS
16774|PINSON
16775|PINTA
16776|PINTO
16777|PINTURA
16778|PIOCHE
16779|PIONEER
16780|PIONEER JUNCTION
16781|PIONEER VILLAGE
16782|PIPE
16783|PIPE CREEK
16784|PIPER
16785|PIPER CITY
16786|PIPERTON
16787|PIPESTONE
16788|PIPPA PASSES
16789|PIQUA
16790|PIRTLEVILLE
16791|PIRU
16792|PISCATAWAY
16793|PISEK
16794|PISGAH
16795|PISGAH FOREST
16796|PISINEMO
16797|PISMO BEACH
16798|PISTAKEE HIGHLANDS
16799|PISTOL RIVER
16800|PITCAIRN
16801|PITKAS POINT
16802|PITKIN
16803|PITMAN
16804|PITSBURG
16805|PITTMAN
16806|PITTMAN CENTER
16807|PITTS
16808|PITTSBORO
16809|PITTSBURG
16810|PITTSBURGH
16811|PITTSFIELD
16812|PITTSFORD
16813|PITTSTON
16814|PITTSVIEW
16815|PITTSVILLE
16816|PITTWOOD
16817|PIXLEY
16818|PIÑON
16819|PIÑON HILLS
16820|PLACEDO
16821|PLACENTIA
16822|PLACER
16823|PLACERVILLE
16824|PLACID
16825|PLACIDA
16826|PLACITAS
16827|PLAIN CITY
16828|PLAIN DEALING
16829|PLAIN VIEW
16830|PLAINEDGE
16831|PLAINFIELD
16832|PLAINS
16833|PLAINSBORO
16834|PLAINSBORO CENTER
16835|PLAINVIEW
16836|PLAINVILLE
16837|PLAINWELL
16838|PLANADA
16839|PLANDOME
16840|PLANDOME HEIGHTS
16841|PLANDOME MANOR
16842|PLANKINTON
16843|PLANO
16844|PLANT CITY
16845|PLANTATION
16846|PLANTATION ISLAND
16847|PLANTATION KEY
16848|PLANTATION MOBILE HOME PARK
16849|PLANTERSVILLE
16850|PLANTSVILLE
16851|PLAQUEMINE
16852|PLASKA
16853|PLASTER CITY
16854|PLAT
16855|PLATA
16856|PLATEA
16857|PLATINA
16858|PLATINUM
16859|PLATNER
16860|PLATO
16861|PLATO CENTER
16862|PLATTE
16863|PLATTE CENTER
16864|PLATTE CITY
16865|PLATTE WOODS
16866|PLATTEKILL
16867|PLATTER
16868|PLATTEVILLE
16869|PLATTSBURG
16870|PLATTSBURGH
16871|PLATTSMOUTH
16872|PLATTVILLE
16873|PLAUCHEVILLE
16874|PLAYA FORTUNA
16875|PLAYA FORTUNA COMUNIDAD
16876|PLAYAS
16877|PLAYITA
16878|PLAYITA COMUNIDAD
16879|PLAYITA CORTADA
16880|PLAYITA CORTADA COMUNIDAD
16881|PLAZA
16882|PLEAK
16883|PLEASANT CITY
16884|PLEASANT DALE
16885|PLEASANT GAP
16886|PLEASANT GARDEN
16887|PLEASANT GREEN
16888|PLEASANT GROVE
16889|PLEASANT HILL
16890|PLEASANT HILLS
16891|PLEASANT HOPE
16892|PLEASANT LAKE
16893|PLEASANT MOUND
16894|PLEASANT PLAIN
16895|PLEASANT PLAINS
16896|PLEASANT PRAIRIE
16897|PLEASANT RIDGE
16898|PLEASANT RUN
16899|PLEASANT RUN FARM
16900|PLEASANT SITE
16901|PLEASANT UNITY
16902|PLEASANT VALLEY
16903|PLEASANT VIEW
16904|PLEASANTON
16905|PLEASANTVILLE
16906|PLEASUREVILLE
16907|PLEDGER
16908|PLENTYWOOD
16909|PLESSIS
16910|PLETCHER
16911|PLETTENBERG
16912|PLEVNA
16913|PLOVER
16914|PLUCKEMIN
16915|PLUM
16916|PLUM BRANCH
16917|PLUM CITY
16918|PLUM CREEK
16919|PLUM GROVE
16920|PLUM SPRINGS
16921|PLUMAS EUREKA
16922|PLUMAS LAKE
16923|PLUMBSOCK
16924|PLUMERVILLE
16925|PLUMMER
16926|PLUMSTEADVILLE
16927|PLUMVILLE
16928|PLUMWOOD
16929|PLUSH
16930|PLYMOUTH
16931|PLYMOUTH MEETING
16932|PLYMPTONVILLE
16933|POAG
16934|POCA
16935|POCAHONTAS
16936|POCALLA SPRINGS
16937|POCASSET
16938|POCATALICO
16939|POCATELLO
16940|POCOLA
16941|POCOMOKE CITY
16942|POCONO MOUNTAIN LAKE ESTATES
16943|POCONO PINES
16944|POCONO RANCH LANDS
16945|POCONO SPRINGS
16946|POCOPSON
16947|POESTENKILL
16948|POHICK
16949|POINCIANA
16950|POINDEXTER
16951|POINT ARENA
16952|POINT BAKER
16953|POINT BLUE
16954|POINT CEDAR
16955|POINT CLEAR
16956|POINT COMFORT
16957|POINT HARBOR
16958|POINT HOPE
16959|POINT ISABEL
16960|POINT LAY
16961|POINT LOOKOUT
16962|POINT MACKENZIE
16963|POINT MARION
16964|POINT OF ROCKS
16965|POINT PLACE
16966|POINT PLEASANT
16967|POINT PLEASANT BEACH
16968|POINT REYES STATION
16969|POINT ROBERTS
16970|POINT VENTURE
16971|POINTE AUX PINS
16972|POINTE À LA HACHE
16973|POJOAQUE
16974|POLACCA
16975|POLAND
16976|POLARIS
16977|POLE OJEA
16978|POLE OJEA COMUNIDAD
16979|POLEBRIDGE
16980|POLK
16981|POLK CITY
16982|POLKTON
16983|POLKVILLE
16984|POLLARD
16985|POLLOCK
16986|POLLOCK PINES
16987|POLLOCKSVILLE
16988|POLLOK
16989|POLO
16990|POLONIA
16991|POLSON
16992|POLVADERA
16993|POMARIA
16994|POMEROY
16995|POMFRET
16996|POMONA
16997|POMONA HEIGHTS
16998|POMONA PARK
16999|POMONKEY
17000|POMPANO BEACH
17001|POMPANO PARK
17002|POMPEYS PILLAR
17003|POMPTON LAKES
17004|POMPTON PLAINS
17005|PONCA
17006|PONCA CITY
17007|PONCE
17008|PONCE DE LEON
17009|PONCE INLET
17010|PONCE ZONA URBANA
17011|PONCHA SPRINGS
17012|PONCHATOULA
17013|POND
17014|POND CREEK
17015|POND EDDY
17016|PONDER
17017|PONDERAY
17018|PONDEROSA
17019|PONDEROSA PARK
17020|PONDEROSA PINE
17021|PONDOSA
17022|PONDSVILLE
17023|PONEMAH
17024|PONETO
17025|PONSFORD
17026|PONSHEWAING
17027|PONTE VEDRA BEACH
17028|PONTIAC
17029|PONTOON BEACH
17030|PONTOOSUC
17031|PONTOTOC
17032|PONY
17033|POOLE
17034|POOLER
17035|POOLESVILLE
17036|POPE
17037|POPE VALLEY
17038|POPEJOY
17039|POPES CREEK
17040|POPLAR
17041|POPLAR BLUFF
17042|POPLAR BRANCH
17043|POPLAR CREEK
17044|POPLAR GROVE
17045|POPLAR HILLS
17046|POPLAR PLAINS
17047|POPLARVILLE
17048|POPPONESSET
17049|POPPONESSET ISLAND
17050|POQUONOCK BRIDGE
17051|POQUOSON
17052|POQUOTT
17053|PORCUPINE
17054|PORT ALEXANDER
17055|PORT ALLEGANY
17056|PORT ALLEN
17057|PORT ALSWORTH
17058|PORT ALTO
17059|PORT ANGELES
17060|PORT ARANSAS
17061|PORT ARMSTRONG
17062|PORT ARTHUR
17063|PORT ASHTON
17064|PORT AUSTIN
17065|PORT BARRE
17066|PORT BARRINGTON
17067|PORT BLAKELY
17068|PORT BOLIVAR
17069|PORT BYRON
17070|PORT CARBON
17071|PORT CHARLOTTE
17072|PORT CHESTER
17073|PORT CHILKOOT
17074|PORT CLARENCE
17075|PORT CLINTON
17076|PORT CLYDE
17077|PORT COLDEN
17078|PORT COSTA
17079|PORT DEPOSIT
17080|PORT DICKINSON
17081|PORT EDWARDS
17082|PORT EWEN
17083|PORT GAMBLE
17084|PORT GIBSON
17085|PORT GRAHAM
17086|PORT HADLOCK
17087|PORT HEIDEN
17088|PORT HENRY
17089|PORT HOPE
17090|PORT HUDSON
17091|PORT HUENEME
17092|PORT HURON
17093|PORT ISABEL
17094|PORT JEFFERSON
17095|PORT JEFFERSON STATION
17096|PORT JERVIS
17097|PORT KENT
17098|PORT LABELLE
17099|PORT LAVACA
17100|PORT LEYDEN
17101|PORT LIONS
17102|PORT LUDLOW
17103|PORT MADISON
17104|PORT MANSFIELD
17105|PORT MATILDA
17106|PORT MAYACA
17107|PORT MOLLER
17108|PORT MONMOUTH
17109|PORT MURRAY
17110|PORT NECHES
17111|PORT NORRIS
17112|PORT O'BRIEN
17113|PORT O'CONNOR
17114|PORT ORANGE
17115|PORT ORCHARD
17116|PORT ORFORD
17117|PORT PROTECTION
17118|PORT READING
17119|PORT REPUBLIC
17120|PORT RICHEY
17121|PORT ROYAL
17122|PORT SAINT JOE
17123|PORT SAINT JOHN
17124|PORT SAINT LUCIE
17125|PORT SALERNO
17126|PORT SANILAC
17127|PORT SEWALL
17128|PORT SULPHUR
17129|PORT TOBACCO
17130|PORT TOWNSEND
17131|PORT TREVORTON
17132|PORT UNION
17133|PORT VINCENT
17134|PORT VUE
17135|PORT WAKEFIELD
17136|PORT WASHINGTON
17137|PORT WASHINGTON NORTH
17138|PORT WENTWORTH
17139|PORT WILLIAM
17140|PORT WING
17141|PORTAGE
17142|PORTAGE CREEK
17143|PORTAGE DES SIOUX
17144|PORTAGE LAKES
17145|PORTAGEVILLE
17146|PORTAL
17147|PORTALES
17148|PORTER
17149|PORTER CENTER
17150|PORTER HEIGHTS
17151|PORTERDALE
17152|PORTERSVILLE
17153|PORTERVILLE
17154|PORTHILL
17155|PORTIA
17156|PORTIS
17157|PORTLAND
17158|PORTLAND MILLS
17159|PORTOLA
17160|PORTOLA VALLEY
17161|PORTSMOUTH
17162|PORTVILLE
17163|PORUM
17164|POSEN
17165|POSEY
17166|POSEYVILLE
17167|POSO PARK
17168|POSSESSION
17169|POST CREEK
17170|POST FALLS
17171|POST LAKE
17172|POST OAK
17173|POST OAK BEND CITY
17174|POSTELLE
17175|POSTON
17176|POSTVILLE
17177|POTALA PASTILLO
17178|POTALA PASTILLO COMUNIDAD
17179|POTATO CREEK
17180|POTEAU
17181|POTEET
17182|POTH
17183|POTLATCH
17184|POTOMAC
17185|POTOMAC HEIGHTS
17186|POTOMAC MILLS
17187|POTOMAC PARK
17188|POTOSI
17189|POTRERO
17190|POTSDAM
17191|POTTAWATTAMIE PARK
17192|POTTER
17193|POTTER LAKE
17194|POTTER VALLEY
17195|POTTERS HILL
17196|POTTERSVILLE
17197|POTTERVILLE
17198|POTTERY ADDITION
17199|POTTS CAMP
17200|POTTSBORO
17201|POTTSGROVE
17202|POTTSTOWN
17203|POTTSVILLE
17204|POTWIN
17205|POUDRE PARK
17206|POUGHKEEPSIE
17207|POULAN
17208|POULSBO
17209|POULTNEY
17210|POWAY
17211|POWDER RIVER
17212|POWDER SPRINGS
17213|POWDER WASH
17214|POWDERHORN
17215|POWDERLY
17216|POWDERSVILLE
17217|POWDERVILLE
17218|POWELL
17219|POWELL BUTTE
17220|POWELLHURST
17221|POWELLS CROSSROADS
17222|POWELLSVILLE
17223|POWELLTON
17224|POWELLVILLE
17225|POWELTON
17226|POWERS LAKE
17227|POWERSVILLE
17228|POWHATAN
17229|POWHATAN POINT
17230|POWHATTAN
17231|POY SIPPI
17232|POYDRAS
17233|POYEN
17234|POYNETTE
17235|POYNOR
17236|POʻIPŪ
17237|PRADO VERDE
17238|PRAGUE
17239|PRAIRIE
17240|PRAIRIE CITY
17241|PRAIRIE CREEK
17242|PRAIRIE DU CHIEN
17243|PRAIRIE DU ROCHER
17244|PRAIRIE DU SAC
17245|PRAIRIE FARM
17246|PRAIRIE GROVE
17247|PRAIRIE HILL
17248|PRAIRIE HOME
17249|PRAIRIE POINT
17250|PRAIRIE RIDGE
17251|PRAIRIE ROSE
17252|PRAIRIE VIEW
17253|PRAIRIE VILLAGE
17254|PRAIRIEBURG
17255|PRAIRIEVILLE
17256|PRATHERSVILLE
17257|PRATTS
17258|PRATTSBURGH
17259|PRATTSVILLE
17260|PRATTVILLE
17261|PREMONT
17262|PRENTICE
17263|PRENTISS
17264|PRESCOTT
17265|PRESCOTT VALLEY
17266|PRESHO
17267|PRESIDENTIAL LAKES ESTATES
17268|PRESIDIO
17269|PRESQUE ISLE
17270|PRESQUILLE
17271|PRESTBURY
17272|PRESTO
17273|PRESTON
17274|PRESTON HEIGHTS
17275|PRESTONSBURG
17276|PRESTONVILLE
17277|PRETTY BAYOU
17278|PRETTY PRAIRIE
17279|PREWITT
17280|PRICE
17281|PRICEDALE
17282|PRICES FORK
17283|PRICEVILLE
17284|PRICHARD
17285|PRIDDY
17286|PRIDE
17287|PRIDGEN
17288|PRIEN
17289|PRIEST RIVER
17290|PRIM
17291|PRIMERA
17292|PRIMGHAR
17293|PRIMROSE
17294|PRINCE
17295|PRINCE FREDERICK
17296|PRINCE GEORGE
17297|PRINCES LAKES
17298|PRINCESS ANNE
17299|PRINCETON
17300|PRINCETON JUNCTION
17301|PRINCETON MEADOWS
17302|PRINCEVILLE
17303|PRINEVILLE
17304|PRINGLE
17305|PRINSBURG
17306|PRIOR LAKE
17307|PRISMATIC
17308|PRITCHETT
17309|PRIVATEER
17310|PROBERTA
17311|PROCTOR
17312|PROCTORSVILLE
17313|PROCTORVILLE
17314|PROGRESO
17315|PROGRESO LAKES
17316|PROGRESS
17317|PROGRESS VILLAGE
17318|PROMISE CITY
17319|PROMISED LAND
17320|PROMPTON
17321|PRONTO
17322|PROPHETSTOWN
17323|PROSIT
17324|PROSPECT
17325|PROSPECT HEIGHTS
17326|PROSPECT PARK
17327|PROSPECT PLAINS
17328|PROSPECT VALLEY
17329|PROSPECTVILLE
17330|PROSPER
17331|PROSPERITY
17332|PROSSER
17333|PROTEM
17334|PROTIVIN
17335|PROVENCAL
17336|PROVIDENCE
17337|PROVIDENCE FORGE
17338|PROVINCETOWN
17339|PROVO
17340|PRUDENVILLE
17341|PRUDHOE BAY
17342|PRUE
17343|PRUNEDALE
17344|PRUNTYTOWN
17345|PRYOR
17346|PRYORSBURG
17347|PUAKŌ
17348|PUCKETT
17349|PUEBLITO
17350|PUEBLITO DEL CARMEN COMUNIDAD
17351|PUEBLITO DEL RIO
17352|PUEBLITO DEL RÍO COMUNIDAD
17353|PUEBLITOS
17354|PUEBLO
17355|PUEBLO NUEVO
17356|PUEBLO NUEVO COLONIA
17357|PUEBLO OF SANDIA VILLAGE
17358|PUEBLO PINTADO
17359|PUEBLO WEST
17360|PUENTE
17361|PUERTO DE LUNA
17362|PUERTO REAL
17363|PUERTO REAL COMUNIDAD
17364|PUHI
17365|PUKALANI
17366|PUKWANA
17367|PULASKI
17368|PULCIFER
17369|PULLMAN
17370|PULTNEYVILLE
17371|PUMPKIN CENTER
17372|PUMPVILLE
17373|PUNALUʻU
17374|PUNGOTEAGUE
17375|PUNTA GORDA
17376|PUNTA RASSA
17377|PUNTA SANTIAGO
17378|PUNTA SANTIAGO COMUNIDAD
17379|PUNXSUTAWNEY
17380|PURCELL
17381|PURCELLVILLE
17382|PURCHASE
17383|PURDIN
17384|PURDON
17385|PURDUM
17386|PURDY
17387|PURLEY
17388|PURPLE SAGE
17389|PURVES
17390|PURVIS
17391|PURYEAR
17392|PUT-IN-BAY
17393|PUTNAM
17394|PUTNAM HALL
17395|PUTNAM LAKE
17396|PUTNAMVILLE
17397|PUTNEY
17398|PUXICO
17399|PUYALLUP
17400|PUʻUWAI
17401|PYATT
17402|PYATTS
17403|PYLESVILLE
17404|PYOTE
17405|PYRAMID
17406|PYRITON
17407|PÁJAROS
17408|PÁJAROS COMUNIDAD
17409|PĀHALA
17410|PĀHOA
17411|PĀKALĀ VILLAGE
17412|PĀPAʻALOA
17413|PĀPAʻIKOU
17414|PĀʻIA
17415|PŪPŪKEA
17416|QUAIL
17417|QUAIL CREEK
17418|QUAKER CITY
17419|QUAKERTOWN
17420|QUAMBA
17421|QUANAH
17422|QUANTICO
17423|QUAPAW
17424|QUARRY
17425|QUARRYVILLE
17426|QUARTZ HILL
17427|QUARTZSITE
17428|QUASQUETON
17429|QUEALY
17430|QUEBEC
17431|QUEBECK
17432|QUEBRADA
17433|QUEBRADA COMUNIDAD
17434|QUEBRADA DEL AGUA COMUNIDAD
17435|QUEBRADILLAS
17436|QUEBRADILLAS ZONA URBANA
17437|QUECHEE
17438|QUEEN
17439|QUEEN ANNE
17440|QUEEN CITY
17441|QUEEN CREEK
17442|QUEEN VALLEY
17443|QUEENS
17444|QUEENSLAND
17445|QUEENSTOWN
17446|QUEETS
17447|QUEMADO
17448|QUENEMO
17449|QUENTIN
17450|QUESTA
17451|QUICK CITY
17452|QUIETUS
17453|QUIJOTOA
17454|QUILCENE
17455|QUIMBY
17456|QUINAULT
17457|QUINBY
17458|QUINCY
17459|QUINEBAUG
17460|QUINHAGAK
17461|QUINLAN
17462|QUINN
17463|QUINNESEC
17464|QUINNIMONT
17465|QUINTANA
17466|QUINTER
17467|QUINTETTE
17468|QUINTON
17469|QUINWOOD
17470|QUIOGUE
17471|QUITAQUE
17472|QUITMAN
17473|QUITO
17474|QUIVERO
17475|QULIN
17476|QUOGUE
17477|QUONOCHONTAUG
17478|RABBIT HASH
17479|RACELAND
17480|RACHAL
17481|RACHEL
17482|RACINE
17483|RADCLIFF
17484|RADCLIFFE
17485|RADERSBURG
17486|RADFORD
17487|RADISSON
17488|RADIUM
17489|RADIUM SPRINGS
17490|RADNOR
17491|RADOM
17492|RAEFORD
17493|RAEMON
17494|RAEVILLE
17495|RAFAEL CAPO
17496|RAFAEL CAPÓ COMUNIDAD
17497|RAFAEL GONZALEZ
17498|RAFAEL GONZÁLEZ COMUNIDAD
17499|RAFAEL HERNANDEZ
17500|RAFAEL HERNÁNDEZ COMUNIDAD
17501|RAFTER J RANCH
17502|RAGAN
17503|RAGLAND
17504|RAGLESVILLE
17505|RAGLEY
17506|RAGO
17507|RAGSDALE
17508|RAHWAY
17509|RAIFORD
17510|RAIL ROAD FLAT
17511|RAILROAD
17512|RAINBOW
17513|RAINBOW CITY
17514|RAINELLE
17515|RAINES
17516|RAINIER
17517|RAINS
17518|RAINSBURG
17519|RAINSVILLE
17520|RAISIN
17521|RAISIN CITY
17522|RAKE
17523|RALEIGH
17524|RALEIGH HILLS
17525|RALLS
17526|RALPH
17527|RALSTON
17528|RAMAH
17529|RAMBLEWOOD
17530|RAMER
17531|RAMEY
17532|RAMHURST
17533|RAMIRENO
17534|RAMIREZ
17535|RAMON
17536|RAMONA
17537|RAMOS
17538|RAMOS COMUNIDAD
17539|RAMPART
17540|RAMSAY
17541|RAMSEUR
17542|RAMSEY
17543|RAMTOWN
17544|RANBURNE
17545|RANCHESTER
17546|RANCHETTE ESTATES
17547|RANCHETTES
17548|RANCHITO
17549|RANCHITOS LAS LOMAS
17550|RANCHO ALEGRE
17551|RANCHO BANQUETE
17552|RANCHO CALAVERAS
17553|RANCHO CHICO
17554|RANCHO CORDOVA
17555|RANCHO CUCAMONGA
17556|RANCHO MIRAGE
17557|RANCHO MURIETA
17558|RANCHO PALOS VERDES
17559|RANCHO RINCONADA
17560|RANCHO SAN DIEGO
17561|RANCHO SANTA FE
17562|RANCHO SANTA MARGARITA
17563|RANCHO TEHAMA RESERVE
17564|RANCHO VIEJO
17565|RANCHOS DE TAOS
17566|RANCHOS PENITAS WEST
17567|RANCOCAS
17568|RANCOCAS WOODS
17569|RAND
17570|RANDADO
17571|RANDALIA
17572|RANDALL
17573|RANDALLSTOWN
17574|RANDLE
17575|RANDLE CLIFF BEACH
17576|RANDLEMAN
17577|RANDLETT
17578|RANDOLPH
17579|RANDOM LAKE
17580|RANDS
17581|RANDSBURG
17582|RANGELY
17583|RANGER
17584|RANGERVILLE
17585|RANIER
17586|RANKIN
17587|RANLO
17588|RANSHAW
17589|RANSOM
17590|RANSOM CANYON
17591|RANSOMVILLE
17592|RANSON
17593|RANTOUL
17594|RAOUL
17595|RAPELJE
17596|RAPID CITY
17597|RAPID VALLEY
17598|RAPIDS
17599|RAPIDS CITY
17600|RAQUETTE LAKE
17601|RARDEN
17602|RARDIN
17603|RARITAN
17604|RATAMOSA
17605|RATCLIFF
17606|RATHBUN
17607|RATHDRUM
17608|RATLIFF
17609|RATLIFF CITY
17610|RATON
17611|RATTAN
17612|RAUB
17613|RAUBSVILLE
17614|RAUCHTOWN
17615|RAVALLI
17616|RAVANNA
17617|RAVEN
17618|RAVENA
17619|RAVENDALE
17620|RAVENDEN
17621|RAVENDEN SPRINGS
17622|RAVENEL
17623|RAVENNA
17624|RAVENSDALE
17625|RAVENSWOOD
17626|RAVENSWORTH
17627|RAVENWOOD
17628|RAVIA
17629|RAVINE
17630|RAVINIA
17631|RAWLINGS
17632|RAWLINS
17633|RAWLS SPRINGS
17634|RAWSON
17635|RAWSONVILLE
17636|RAY
17637|RAY CITY
17638|RAYBURN
17639|RAYLAND
17640|RAYLE
17641|RAYMER
17642|RAYMOND
17643|RAYMONDVILLE
17644|RAYMORE
17645|RAYNE
17646|RAYNESFORD
17647|RAYNHAM
17648|RAYNHAM CENTER
17649|RAYSAL
17650|RAYTOWN
17651|RAYVILLE
17652|RAYWICK
17653|REA
17654|READER
17655|READING
17656|READINGTON
17657|READLAND
17658|READLYN
17659|READS LANDING
17660|READSBORO
17661|READSTOWN
17662|READSVILLE
17663|REAGAN
17664|REAGER
17665|REALITOS
17666|REAMSTOWN
17667|REARDAN
17668|REASNOR
17669|REBECCA
17670|REBERSBURG
17671|RECLUSE
17672|RECTOR
17673|RECTORVILLE
17674|RED ASH
17675|RED BANK
17676|RED BANKS
17677|RED BAY
17678|RED BIRD
17679|RED BLUFF
17680|RED BOILING SPRINGS
17681|RED BUD
17682|RED BUTTE
17683|RED BUTTES
17684|RED CHUTE
17685|RED CLIFF
17686|RED CLOUD
17687|RED CREEK
17688|RED CROSS
17689|RED DEVIL
17690|RED DOG MINE
17691|RED ELM
17692|RED FEATHER LAKES
17693|RED GATE
17694|RED HEAD
17695|RED HILL
17696|RED HOOK
17697|RED JACKET
17698|RED LAKE
17699|RED LAKE FALLS
17700|RED LEVEL
17701|RED LICK
17702|RED LION
17703|RED LODGE
17704|RED MESA
17705|RED MILLS
17706|RED MOUNTAIN
17707|RED OAK
17708|RED OAKS MILL
17709|RED RIVER
17710|RED RIVER HOT SPRINGS
17711|RED ROCK
17712|RED SHIRT
17713|RED SPRINGS
17714|RED STAR
17715|RED WING
17716|REDAN
17717|REDBANK
17718|REDBIRD
17719|REDBIRD SMITH
17720|REDBY
17721|REDCREST
17722|REDDELL
17723|REDDEN
17724|REDDICK
17725|REDDING
17726|REDFIELD
17727|REDFORD
17728|REDGRANITE
17729|REDIG
17730|REDINGS MILL
17731|REDINGTON
17732|REDINGTON BEACH
17733|REDINGTON SHORES
17734|REDKEY
17735|REDLAND
17736|REDLANDS
17737|REDMESA
17738|REDMON
17739|REDMOND
17740|REDONDO
17741|REDONDO BEACH
17742|REDOWL
17743|REDROCK
17744|REDSTONE
17745|REDVALE
17746|REDWATER
17747|REDWAY
17748|REDWOOD
17749|REDWOOD CITY
17750|REDWOOD FALLS
17751|REDWOOD TERRACE
17752|REDWOOD VALLEY
17753|REE HEIGHTS
17754|REECE
17755|REECE CITY
17756|REED
17757|REED CITY
17758|REED CREEK
17759|REED POINT
17760|REEDER
17761|REEDLEY
17762|REEDS
17763|REEDS SPRING
17764|REEDSBURG
17765|REEDSPORT
17766|REEDSVILLE
17767|REEDVILLE
17768|REEDY
17769|REELTOWN
17770|REESE
17771|REESEVILLE
17772|REEVES
17773|REEVESVILLE
17774|REFORM
17775|REFTON
17776|REFUGIO
17777|REGAL
17778|REGAN
17779|REGANTON
17780|REGENT
17781|REGGIO
17782|REGINA
17783|REGISTER
17784|REGO PARK
17785|REHOBETH
17786|REHOBOTH
17787|REHOBOTH BEACH
17788|REHRERSBURG
17789|REID
17790|REID HOPE KING COLONIA
17791|REIDLAND
17792|REIDSVILLE
17793|REIDVILLE
17794|REIFFTON
17795|REILES ACRES
17796|REILY
17797|REINBECK
17798|REINERSVILLE
17799|REINERTON
17800|REINHOLDS
17801|REISTERSTOWN
17802|REKLAW
17803|RELAMPAGO
17804|RELIANCE
17805|REMBERT
17806|REMBRANDT
17807|REMER
17808|REMERTON
17809|REMINDERVILLE
17810|REMINGTON
17811|REMSEN
17812|REMSENBURG
17813|REMY
17814|RENA
17815|RENDON
17816|RENDVILLE
17817|RENFROE
17818|RENFROW
17819|RENICK
17820|RENNER
17821|RENNER CORNER
17822|RENNERDALE
17823|RENNERT
17824|RENNINGERS
17825|RENO
17826|RENOVA
17827|RENOVO
17828|RENSSELAER
17829|RENSSELAER FALLS
17830|RENTCHLER
17831|RENTIESVILLE
17832|RENTON
17833|RENTZ
17834|RENVILLE
17835|RENWICK
17836|REPAUPO
17837|REPTON
17838|REPUBLIC
17839|REPUBLICAN CITY
17840|REQUA
17841|RERDELL
17842|RESACA
17843|RESERVE
17844|RESOTA BEACH
17845|REST HAVEN
17846|RESTON
17847|RETREAT
17848|RETROP
17849|RETSOF
17850|RETTA
17851|REUBENS
17852|REVA
17853|REVERE
17854|REVILLO
17855|REVLOC
17856|REW
17857|REWEY
17858|REX
17859|REXBURG
17860|REXFORD
17861|REXHAME
17862|REXTON
17863|REXVILLE
17864|REYDON
17865|REYNO
17866|REYNOLDS
17867|REYNOLDS HEIGHTS
17868|REYNOLDSBURG
17869|REYNOLDSVILLE
17870|RHAME
17871|RHEA
17872|RHEATOWN
17873|RHEEM
17874|RHEEMS
17875|RHINE
17876|RHINEBECK
17877|RHINECLIFF
17878|RHINELAND
17879|RHINELANDER
17880|RHODELL
17881|RHODES
17882|RHODHISS
17883|RHODODENDRON
17884|RHOME
17885|RIALTO
17886|RIB LAKE
17887|RIB MOUNTAIN
17888|RIBERA
17889|RICARDO
17890|RICE
17891|RICE LAKE
17892|RICEBORO
17893|RICES LANDING
17894|RICEVILLE
17895|RICH
17896|RICH CREEK
17897|RICH FOUNTAIN
17898|RICH HILL
17899|RICH POND
17900|RICH SQUARE
17901|RICH VALLEY
17902|RICHARDS
17903|RICHARDSON
17904|RICHARDSVILLE
17905|RICHARDTON
17906|RICHBORO
17907|RICHBURG
17908|RICHEY
17909|RICHFIELD
17910|RICHFIELD SPRINGS
17911|RICHFORD
17912|RICHGROVE
17913|RICHLAND
17914|RICHLAND CENTER
17915|RICHLAND HILLS
17916|RICHLAND SPRINGS
17917|RICHLANDS
17918|RICHLANDTOWN
17919|RICHLAWN
17920|RICHMOND
17921|RICHMOND BEACH
17922|RICHMOND DALE
17923|RICHMOND HEIGHTS
17924|RICHMOND HIGHLANDS
17925|RICHMOND HILL
17926|RICHMONDVILLE
17927|RICHTEX
17928|RICHTON
17929|RICHTON PARK
17930|RICHVALE
17931|RICHVIEW
17932|RICHVILLE
17933|RICHWOOD
17934|RICHWOODS
17935|RICKARDSVILLE
17936|RICKETTS
17937|RICKMAN
17938|RICKREALL
17939|RICO
17940|RIDDLE
17941|RIDDLESBURG
17942|RIDDLEVILLE
17943|RIDERWOOD
17944|RIDGE
17945|RIDGE FARM
17946|RIDGE MANOR
17947|RIDGE SPRING
17948|RIDGE WOOD HEIGHTS
17949|RIDGECREST
17950|RIDGEFIELD
17951|RIDGEFIELD PARK
17952|RIDGELAND
17953|RIDGELEY
17954|RIDGELY
17955|RIDGEMARK
17956|RIDGESIDE
17957|RIDGETOP
17958|RIDGEVIEW
17959|RIDGEVILLE
17960|RIDGEVILLE CORNERS
17961|RIDGEWAY
17962|RIDGEWOOD
17963|RIDGWAY
17964|RIDLEY PARK
17965|RIDOTT
17966|RIEGELSVILLE
17967|RIEGELWOOD
17968|RIENZI
17969|RIESEL
17970|RIETH
17971|RIFLE
17972|RIFTON
17973|RIGBY
17974|RIGGINS
17975|RILEY
17976|RILEYVILLE
17977|RILLITO
17978|RILLTON
17979|RIMERSBURG
17980|RIMFOREST
17981|RIMINI
17982|RINARD
17983|RINCON
17984|RINCÓN
17985|RINCÓN ZONA URBANA
17986|RINER
17987|RINEYVILLE
17988|RINGGOLD
17989|RINGLING
17990|RINGOLD
17991|RINGSTED
17992|RINGTON
17993|RINGTOWN
17994|RINGWOOD
17995|RIO
17996|RIO BLANCO
17997|RIO BRAVO
17998|RIO COMMUNITIES
17999|RIO CREEK
18000|RIO DEL MAR
18001|RIO DELL
18002|RIO EN MEDIO
18003|RIO GRANDE
18004|RIO GRANDE CITY
18005|RIO HONDO
18006|RIO LINDA
18007|RIO LUCIO
18008|RIO OSO
18009|RIO RANCHO
18010|RIO RICO
18011|RIO VERDE
18012|RIO VISTA
18013|RIOMEDINA
18014|RION
18015|RIOS
18016|RIPLEY
18017|RIPLINGER
18018|RIPON
18019|RIPPEY
18020|RIPPON
18021|RIRIE
18022|RISCO
18023|RISING CITY
18024|RISING FAWN
18025|RISING STAR
18026|RISING SUN
18027|RISINGSUN
18028|RISON
18029|RITCHEY
18030|RITCHIE
18031|RITTMAN
18032|RITZVILLE
18033|RIVA
18034|RIVANNA
18035|RIVER BEND
18036|RIVER BLUFF
18037|RIVER EDGE
18038|RIVER FALLS
18039|RIVER FOREST
18040|RIVER GROVE
18041|RIVER HEIGHTS
18042|RIVER HILLS
18043|RIVER OAKS
18044|RIVER PARK
18045|RIVER PINES
18046|RIVER RIDGE
18047|RIVER ROAD
18048|RIVER ROUGE
18049|RIVER SIOUX
18050|RIVER VIEW PARK
18051|RIVERA COLONIA
18052|RIVERBANK
18053|RIVERBEND
18054|RIVERDALE
18055|RIVERDALE PARK
18056|RIVERGROVE
18057|RIVERHEAD
18058|RIVERLAND
18059|RIVERLEA
18060|RIVERSIDE
18061|RIVERSIDE PARK
18062|RIVERTON
18063|RIVERVALE
18064|RIVERVIEW
18065|RIVERVIEW ESTATES
18066|RIVERVIEW FARMS
18067|RIVERWOOD
18068|RIVERWOODS
18069|RIVES
18070|RIVES JUNCTION
18071|RIVESVILLE
18072|RIVIERA
18073|RIVIERA BEACH
18074|RIXFORD
18075|ROACH
18076|ROACHDALE
18077|ROACHTOWN
18078|ROADS
18079|ROADS END
18080|ROAMING SHORES
18081|ROAN MOUNTAIN
18082|ROANE
18083|ROANN
18084|ROANOKE
18085|ROANOKE RAPIDS
18086|ROARING GAP
18087|ROARING SPRING
18088|ROARING SPRINGS
18089|ROBARDS
18090|ROBBIN
18091|ROBBINS
18092|ROBBINSDALE
18093|ROBBINSVILLE
18094|ROBBS
18095|ROBE
18096|ROBELINE
18097|ROBERSONVILLE
18098|ROBERT
18099|ROBERT LEE
18100|ROBERTA
18101|ROBERTA MILL
18102|ROBERTS
18103|ROBERTSBURG
18104|ROBERTSDALE
18105|ROBERTSON
18106|ROBERTSVILLE
18107|ROBESONIA
18108|ROBIN
18109|ROBINETTE
18110|ROBINS
18111|ROBINSON
18112|ROBINSONVILLE
18113|ROBINWOOD
18114|ROBSTOWN
18115|ROBY
18116|ROCA
18117|ROCHELLE
18118|ROCHEPORT
18119|ROCHERT
18120|ROCHESTER
18121|ROCHESTER HILLS
18122|ROCHFORD
18123|ROCK
18124|ROCK CAVE
18125|ROCK CITY
18126|ROCK CREEK
18127|ROCK CREEK PARK
18128|ROCK FALLS
18129|ROCK HALL
18130|ROCK HILL
18131|ROCK ISLAND
18132|ROCK LAKE
18133|ROCK MILLS
18134|ROCK POINT
18135|ROCK PORT
18136|ROCK RAPIDS
18137|ROCK RIVER
18138|ROCK SPRING
18139|ROCK SPRINGS
18140|ROCK VALLEY
18141|ROCKAWAY
18142|ROCKAWAY BEACH
18143|ROCKBRIDGE
18144|ROCKCREEK
18145|ROCKDALE
18146|ROCKDELL
18147|ROCKERVILLE
18148|ROCKFIELD
18149|ROCKFISH
18150|ROCKFORD
18151|ROCKFORD BAY
18152|ROCKHAM
18153|ROCKHILL
18154|ROCKHOLDS
18155|ROCKINGHAM
18156|ROCKLAND
18157|ROCKLEDGE
18158|ROCKLEIGH
18159|ROCKLIN
18160|ROCKMART
18161|ROCKPORT
18162|ROCKSPRINGS
18163|ROCKTON
18164|ROCKVALE
18165|ROCKVILLE
18166|ROCKVILLE CENTRE
18167|ROCKWALL
18168|ROCKWELL
18169|ROCKWELL CITY
18170|ROCKWOOD
18171|ROCKY
18172|ROCKY BOY'S AGENCY
18173|ROCKY COMFORT
18174|ROCKY FORD
18175|ROCKY FORK
18176|ROCKY FORK POINT
18177|ROCKY GAP
18178|ROCKY GROVE
18179|ROCKY HILL
18180|ROCKY MOUND
18181|ROCKY MOUNT
18182|ROCKY MOUNTAIN
18183|ROCKY POINT
18184|ROCKY RIDGE
18185|ROCKY RIDGE RANCH
18186|ROCKY RIPPLE
18187|ROCKY RIVER
18188|ROCKY TOP
18189|ROCKYPOINT
18190|RODANTHE
18191|RODARTE
18192|RODEO
18193|RODERFIELD
18194|RODESSA
18195|RODEY
18196|RODMAN
18197|RODNEY
18198|RODNEY VILLAGE
18199|RODRÍGUEZ HEVIA
18200|RODRÍGUEZ HEVIA COMUNIDAD
18201|ROE
18202|ROE PARK
18203|ROEBLING
18204|ROEBUCK
18205|ROELAND PARK
18206|ROELLEN
18207|ROESSLEVILLE
18208|ROEVILLE
18209|ROFF
18210|ROGANVILLE
18211|ROGERS
18212|ROGERS CITY
18213|ROGERSON
18214|ROGERSVILLE
18215|ROGGEN
18216|ROGUE RIVER
18217|ROHNERT PARK
18218|ROHNERVILLE
18219|ROHRERSVILLE
18220|ROHRSBURG
18221|ROHWER
18222|ROLAND
18223|ROLESVILLE
18224|ROLETTE
18225|ROLFE
18226|ROLINDA
18227|ROLL
18228|ROLLA
18229|ROLLING FIELDS
18230|ROLLING FORK
18231|ROLLING HILLS
18232|ROLLING HILLS ESTATES
18233|ROLLING MEADOWS
18234|ROLLING PRAIRIE
18235|ROLLINGBAY
18236|ROLLINGSTONE
18237|ROLLINGWOOD
18238|ROLLINS
18239|ROLLINSVILLE
18240|ROMA
18241|ROMA CREEK
18242|ROMA-LOS SAENZ
18243|ROMAN FOREST
18244|ROMANCOKE
18245|ROMAYOR
18246|ROMBAUER
18247|ROME
18248|ROME CITY
18249|ROMEO
18250|ROMEOVILLE
18251|ROMERO
18252|ROMEROVILLE
18253|ROMEVILLE
18254|ROMNEY
18255|ROMOLAND
18256|ROMULUS
18257|RONALD
18258|RONAN
18259|RONCEVERTE
18260|RONCO
18261|RONDA
18262|RONDO
18263|RONDOUT
18264|RONKONKOMA
18265|RONKS
18266|RONNEBY
18267|ROODHOUSE
18268|ROOPVILLE
18269|ROOSEVELT
18270|ROOSEVELT BEACH
18271|ROOSEVELT GARDENS
18272|ROOSEVELT PARK
18273|ROOSVILLE
18274|ROPER
18275|ROPESVILLE
18276|ROSA
18277|ROSA SANCHEZ
18278|ROSA SÁNCHEZ COMUNIDAD
18279|ROSALIA
18280|ROSALIE
18281|ROSAMOND
18282|ROSANKY
18283|ROSARIO
18284|ROSARYVILLE
18285|ROSATI
18286|ROSBORO
18287|ROSBURG
18288|ROSCOE
18289|ROSCOMMON
18290|ROSE
18291|ROSE BUD
18292|ROSE CITY
18293|ROSE CREEK
18294|ROSE FARM
18295|ROSE HAVEN
18296|ROSE HILL
18297|ROSE HILL ACRES
18298|ROSE HILL FARMS
18299|ROSE LAKE
18300|ROSE LODGE
18301|ROSE TREE
18302|ROSE VALLEY
18303|ROSEAU
18304|ROSEBORO
18305|ROSEBUD
18306|ROSEBURG
18307|ROSEBUSH
18308|ROSEDALE
18309|ROSEGLEN
18310|ROSELAND
18311|ROSELAWN
18312|ROSELLE
18313|ROSELLE PARK
18314|ROSEMARK
18315|ROSEMEAD
18316|ROSEMONT
18317|ROSEMOUNT
18318|ROSEN
18319|ROSENBERG
18320|ROSENDALE
18321|ROSENHAYN
18322|ROSEPINE
18323|ROSETO
18324|ROSETTA
18325|ROSETTE
18326|ROSEVILLE
18327|ROSEVILLE PARK
18328|ROSEWOOD
18329|ROSEWOOD HEIGHTS
18330|ROSEWORTH
18331|ROSHARON
18332|ROSHOLT
18333|ROSICLARE
18334|ROSIER
18335|ROSINE
18336|ROSITA
18337|ROSLYN
18338|ROSLYN ESTATES
18339|ROSLYN HARBOR
18340|ROSLYN HEIGHTS
18341|ROSMAN
18342|ROSS
18343|ROSS CORNER
18344|ROSS FORK
18345|ROSSBURG
18346|ROSSER
18347|ROSSFORD
18348|ROSSIE
18349|ROSSITER
18350|ROSSLYN FARMS
18351|ROSSMOOR
18352|ROSSMORE
18353|ROSSMOYNE
18354|ROSSTON
18355|ROSSVILLE
18356|ROSWELL
18357|ROTAN
18358|ROTE
18359|ROTHBURY
18360|ROTHSAY
18361|ROTHSCHILD
18362|ROTHSVILLE
18363|ROTHVILLE
18364|ROTONDA
18365|ROTTERDAM
18366|ROUGEMONT
18367|ROUGH AND READY
18368|ROUGH ROCK
18369|ROULETTE
18370|ROULO
18371|ROUND GROVE
18372|ROUND HILL
18373|ROUND LAKE
18374|ROUND LAKE BEACH
18375|ROUND LAKE HEIGHTS
18376|ROUND LAKE PARK
18377|ROUND MOUNTAIN
18378|ROUND OAK
18379|ROUND POND
18380|ROUND PRAIRIE
18381|ROUND ROCK
18382|ROUND TOP
18383|ROUND VALLEY
18384|ROUNDHEAD
18385|ROUNDUP
18386|ROUSES POINT
18387|ROUSEVILLE
18388|ROUZERVILLE
18389|ROVER
18390|ROWAN
18391|ROWDEN
18392|ROWE
18393|ROWENA
18394|ROWES RUN
18395|ROWESVILLE
18396|ROWLAND
18397|ROWLAND HEIGHTS
18398|ROWLESBURG
18399|ROWLETT
18400|ROWLEY
18401|ROWSBURG
18402|ROX
18403|ROXANA
18404|ROXBORO
18405|ROXBOROUGH PARK
18406|ROXBURY
18407|ROXIE
18408|ROXOBEL
18409|ROXTON
18410|ROY
18411|ROY LAKE
18412|ROYAL
18413|ROYAL CENTER
18414|ROYAL CITY
18415|ROYAL LAKES
18416|ROYAL OAK
18417|ROYAL PALM BEACH
18418|ROYAL PALM ESTATES
18419|ROYAL PINES
18420|ROYALTON
18421|ROYALTY
18422|ROYCE
18423|ROYERSFORD
18424|ROYSE CITY
18425|ROYSTON
18426|ROYVILLE
18427|ROZEL
18428|ROZELLVILLE
18429|ROZET
18430|RUBIDOUX
18431|RUBIO
18432|RUBONIA
18433|RUBY
18434|RUBY VALLEY
18435|RUCH
18436|RUCKER
18437|RUCKERSVILLE
18438|RUDD
18439|RUDEVILLE
18440|RUDOLPH
18441|RUDY
18442|RUDYARD
18443|RUETER
18444|RUFE
18445|RUFF
18446|RUFFIN
18447|RUFUS
18448|RUGBY
18449|RUIDOSA
18450|RUIDOSO
18451|RUIDOSO DOWNS
18452|RULEVILLE
18453|RULO
18454|RUMA
18455|RUMFORD
18456|RUMSON
18457|RUNAWAY BAY
18458|RUNGE
18459|RUNNELLS
18460|RUNNELSTOWN
18461|RUNNEMEDE
18462|RUNNING SPRINGS
18463|RUNNING WATER
18464|RUPERT
18465|RURAL HALL
18466|RURAL HILL
18467|RURAL RETREAT
18468|RURAL RIDGE
18469|RURAL VALLEY
18470|RUSH
18471|RUSH CENTER
18472|RUSH CITY
18473|RUSH HILL
18474|RUSH SPRINGS
18475|RUSH VALLEY
18476|RUSHFORD
18477|RUSHFORD VILLAGE
18478|RUSHMERE
18479|RUSHMORE
18480|RUSHSYLVANIA
18481|RUSHTON
18482|RUSHVILLE
18483|RUSK
18484|RUSKIN
18485|RUSO
18486|RUSSELL
18487|RUSSELL CITY
18488|RUSSELL GARDENS
18489|RUSSELL SPRINGS
18490|RUSSELLS POINT
18491|RUSSELLTON
18492|RUSSELLVILLE
18493|RUSSIA
18494|RUSSIAN MISSION
18495|RUSSIAVILLE
18496|RUSTAD
18497|RUSTBURG
18498|RUSTON
18499|RUTERSVILLE
18500|RUTH
18501|RUTHER GLEN
18502|RUTHERFORD
18503|RUTHERFORD COLLEGE
18504|RUTHERFORDTON
18505|RUTHERON
18506|RUTHSBURG
18507|RUTHTON
18508|RUTHVEN
18509|RUTHVILLE
18510|RUTLAND
18511|RUTLEDGE
18512|RYAN
18513|RYAN PARK
18514|RYDER
18515|RYDERWOOD
18516|RYE
18517|RYE BEACH
18518|RYE BROOK
18519|RYEGATE
18520|RYLAND
18521|RYLAND HEIGHTS
18522|RÍO BLANCO
18523|RÍO BLANCO COMUNIDAD
18524|RÍO CAÑAS ABAJO
18525|RÍO CAÑAS ABAJO COMUNIDAD
18526|RÍO GRANDE
18527|RÍO GRANDE ZONA URBANA
18528|RÍO LAJAS
18529|RÍO LAJAS COMUNIDAD
18530|SABANA
18531|SABANA COMUNIDAD
18532|SABANA ENEAS
18533|SABANA ENEAS COMUNIDAD
18534|SABANA GRANDE
18535|SABANA GRANDE ZONA URBANA
18536|SABANA HOYOS
18537|SABANA HOYOS COMUNIDAD
18538|SABANA SECA
18539|SABANA SECA COMUNIDAD
18540|SABATTIS
18541|SABETHA
18542|SABILLASVILLE
18543|SABIN
18544|SABINA
18545|SABINAL
18546|SABINE
18547|SABINE PASS
18548|SABINOSO
18549|SABINSVILLE
18550|SABULA
18551|SAC CITY
18552|SACATON
18553|SACHSE
18554|SACKETS HARBOR
18555|SACO
18556|SACRAMENTO
18557|SACRED HEART
18558|SADDLE BUTTE
18559|SADDLE RIVER
18560|SADDLE ROCK
18561|SADDLE ROCK ESTATES
18562|SADDLEBROOKE
18563|SADDLESTRING
18564|SADIEVILLE
18565|SADLER
18566|SADORUS
18567|SADSBURYVILLE
18568|SAEGERTOWN
18569|SAFETY HARBOR
18570|SAFFORD
18571|SAG HARBOR
18572|SAGAMORE
18573|SAGAMORE HILLS
18574|SAGAPONACK
18575|SAGE
18576|SAGERTON
18577|SAGEVILLE
18578|SAGINAW
18579|SAGUACHE
18580|SAHALEE
18581|SAHUARITA
18582|SAILOR SPRINGS
18583|SAINT ALBANS
18584|SAINT ANDREWS
18585|SAINT ANN
18586|SAINT ANN HIGHLANDS
18587|SAINT ANNE
18588|SAINT ANSGAR
18589|SAINT ANTHONY
18590|SAINT AUGUSTA
18591|SAINT AUGUSTINE
18592|SAINT AUGUSTINE BEACH
18593|SAINT AUGUSTINE SHORES
18594|SAINT AUGUSTINE SOUTH
18595|SAINT BENEDICT
18596|SAINT BERNARD
18597|SAINT BERNICE
18598|SAINT BETHLEHEM
18599|SAINT BONAVENTURE
18600|SAINT BONIFACIUS
18601|SAINT CATHERINE
18602|SAINT CHARLES
18603|SAINT CLAIR
18604|SAINT CLAIR HAVEN
18605|SAINT CLAIR SHORES
18606|SAINT CLAIRSVILLE
18607|SAINT CLEMENT
18608|SAINT CLOUD
18609|SAINT CROIX FALLS
18610|SAINT DAVID
18611|SAINT DONATUS
18612|SAINT EDWARD
18613|SAINT ELIZABETH
18614|SAINT ELMO
18615|SAINT FLORIAN
18616|SAINT FRANCIS
18617|SAINT FRANCISVILLE
18618|SAINT GABRIEL
18619|SAINT GEORGE
18620|SAINT GEORGE ISLAND
18621|SAINT GEORGES
18622|SAINT HEDWIG
18623|SAINT HELEN
18624|SAINT HELENA
18625|SAINT HELENS
18626|SAINT HENRY
18627|SAINT HILAIRE
18628|SAINT IGNACE
18629|SAINT IGNATIUS
18630|SAINT JACOB
18631|SAINT JAMES
18632|SAINT JAMES CITY
18633|SAINT JO
18634|SAINT JOE
18635|SAINT JOHN
18636|SAINT JOHNS
18637|SAINT JOHNSBURG
18638|SAINT JOHNSBURY
18639|SAINT JOHNSVILLE
18640|SAINT JOSEPH
18641|SAINT LANDRY
18642|SAINT LAWRENCE
18643|SAINT LEO
18644|SAINT LEON
18645|SAINT LEONARD
18646|SAINT LIBORY
18647|SAINT LOUIS
18648|SAINT LOUIS PARK
18649|SAINT LOUISVILLE
18650|SAINT LUCAS
18651|SAINT LUCIE
18652|SAINT MARIE
18653|SAINT MARIES
18654|SAINT MARKS
18655|SAINT MARTIN
18656|SAINT MARTINS
18657|SAINT MARTINVILLE
18658|SAINT MARY
18659|SAINT MARY-OF-THE-WOODS
18660|SAINT MARYS
18661|SAINT MARYS CITY
18662|SAINT MARYS POINT
18663|SAINT MATTHEWS
18664|SAINT MAURICE
18665|SAINT MEINRAD
18666|SAINT MICHAEL
18667|SAINT MICHAELS
18668|SAINT NAZIANZ
18669|SAINT NICHOLAS
18670|SAINT OLAF
18671|SAINT ONGE
18672|SAINT PARIS
18673|SAINT PAUL
18674|SAINT PAUL PARK
18675|SAINT PAULS
18676|SAINT PETE BEACH
18677|SAINT PETER
18678|SAINT PETERS
18679|SAINT PETERSBURG
18680|SAINT PIERRE
18681|SAINT REGIS
18682|SAINT REGIS FALLS
18683|SAINT REGIS PARK
18684|SAINT ROBERT
18685|SAINT ROSA
18686|SAINT ROSE
18687|SAINT SIMONS
18688|SAINT STEPHEN
18689|SAINT STEPHENS
18690|SAINT TERESA
18691|SAINT THOMAS
18692|SAINT VINCENT
18693|SAINT XAVIER
18694|SAINTE GENEVIEVE
18695|SAINTE MARIE
18696|SAKS
18697|SALADO
18698|SALAMANCA
18699|SALAMATOF
18700|SALAMONIA
18701|SALDURO
18702|SALE CITY
18703|SALE CREEK
18704|SALEM
18705|SALEM HEIGHTS
18706|SALEM LAKES
18707|SALEMBURG
18708|SALESVILLE
18709|SALIDA
18710|SALINA
18711|SALINAS
18712|SALINAS ZONA URBANA
18713|SALINEVILLE
18714|SALINEÑO
18715|SALISBURY
18716|SALISBURY MILLS
18717|SALITPA
18718|SALIX
18719|SALKUM
18720|SALLADASBURG
18721|SALLEY
18722|SALLIS
18723|SALLISAW
18724|SALLYARDS
18725|SALMON
18726|SALMON BROOK
18727|SALMON CREEK
18728|SALOL
18729|SALOME
18730|SALT CHUCK
18731|SALT CREEK
18732|SALT FLAT
18733|SALT FORK
18734|SALT GAP
18735|SALT LAKE CITY
18736|SALT LICK
18737|SALT POINT
18738|SALT ROCK
18739|SALT SPRINGS
18740|SALT WELLS
18741|SALTAIRE
18742|SALTER PATH
18743|SALTERS
18744|SALTESE
18745|SALTILLO
18746|SALTON CITY
18747|SALTON SEA BEACH
18748|SALTSBURG
18749|SALTVILLE
18750|SALUDA
18751|SALUNGA
18752|SALUS
18753|SALVISA
18754|SALVO
18755|SALYER
18756|SALYERSVILLE
18757|SAM RAYBURN
18758|SAMAK
18759|SAMANTHA
18760|SAMARIA
18761|SAMBURG
18762|SAMMAMISH
18763|SAMMONS POINT
18764|SAMNORWOOD
18765|SAMOA
18766|SAMOSET
18767|SAMPSON
18768|SAMSON
18769|SAMSULA
18770|SAMUELS
18771|SAN ACACIA
18772|SAN ACACIO
18773|SAN ANDREAS
18774|SAN ANGELO
18775|SAN ANSELMO
18776|SAN ANTONIO
18777|SAN ANTONIO COMUNIDAD
18778|SAN ANTONIO HEIGHTS
18779|SAN ANTONITO
18780|SAN ARDO
18781|SAN AUGUSTINE
18782|SAN BENITO
18783|SAN BERNARDINO
18784|SAN BRUNO
18785|SAN CARLOS
18786|SAN CARLOS NUMBER 1 COLONIA
18787|SAN CARLOS PARK
18788|SAN CLEMENTE
18789|SAN CRISTOBAL
18790|SAN DE FUCA
18791|SAN DIEGO
18792|SAN DIEGO COUNTRY ESTATES
18793|SAN DIMAS
18794|SAN ELIZARIO
18795|SAN FELIPE
18796|SAN FELIPE PUEBLO
18797|SAN FERNANDO
18798|SAN FIDEL
18799|SAN FRANCISCO
18800|SAN GABRIEL
18801|SAN GERMÁN
18802|SAN GERMÁN ZONA URBANA
18803|SAN GERONIMO
18804|SAN GREGORIO
18805|SAN IGNACIO
18806|SAN ILDEFONSO PUEBLO
18807|SAN ISIDRO
18808|SAN ISIDRO COMUNIDAD
18809|SAN JACINTO
18810|SAN JOAQUIN
18811|SAN JON
18812|SAN JOSE
18813|SAN JOSÉ
18814|SAN JOSÉ COMUNIDAD
18815|SAN JUAN
18816|SAN JUAN BAUTISTA
18817|SAN JUAN CAPISTRANO
18818|SAN JUAN COLONIA
18819|SAN JUAN HOT SPRINGS
18820|SAN JUAN PUEBLO
18821|SAN JUAN ZONA URBANA
18822|SAN LEANDRO
18823|SAN LEANNA
18824|SAN LEON
18825|SAN LORENZO
18826|SAN LORENZO ZONA URBANA
18827|SAN LUCAS
18828|SAN LUIS
18829|SAN LUIS OBISPO
18830|SAN LUIS REY
18831|SAN MANUEL
18832|SAN MAR
18833|SAN MARCIAL
18834|SAN MARCOS
18835|SAN MARINO
18836|SAN MARTIN
18837|SAN MATEO
18838|SAN MIGUEL
18839|SAN PABLO
18840|SAN PASQUAL
18841|SAN PATRICIO
18842|SAN PEDRO
18843|SAN PERLITA
18844|SAN PIERRE
18845|SAN QUENTIN
18846|SAN RAFAEL
18847|SAN RAMON
18848|SAN REMO
18849|SAN SABA
18850|SAN SEBASTIÁN
18851|SAN SEBASTIÁN ZONA URBANA
18852|SAN SIMEON
18853|SAN SIMON
18854|SAN TAN VALLEY
18855|SAN YGNACIO
18856|SAN YSIDRO
18857|SANAK
18858|SANATOGA
18859|SANATORIUM
18860|SANBORN
18861|SANBORNVILLE
18862|SANCTUARY
18863|SAND CITY
18864|SAND COULEE
18865|SAND CREEK
18866|SAND DRAW
18867|SAND FORK
18868|SAND HILL
18869|SAND LAKE
18870|SAND PASS
18871|SAND POINT
18872|SAND RIDGE
18873|SAND ROCK
18874|SAND SPRINGS
18875|SANDBORN
18876|SANDERS
18877|SANDERSON
18878|SANDERSVILLE
18879|SANDGAP
18880|SANDIA
18881|SANDIA HEIGHTS
18882|SANDIA KNOLLS
18883|SANDIA PARK
18884|SANDOVAL
18885|SANDOW
18886|SANDPOINT
18887|SANDS POINT
18888|SANDSTON
18889|SANDSTONE
18890|SANDUSKY
18891|SANDWICH
18892|SANDY
18893|SANDY BEACH
18894|SANDY BOTTOM
18895|SANDY CITY
18896|SANDY CREEK
18897|SANDY HOOK
18898|SANDY LAKE
18899|SANDY LEVEL
18900|SANDY OAKS
18901|SANDY PLAINS
18902|SANDY RIDGE
18903|SANDY SPRING
18904|SANDY SPRINGS
18905|SANDY VALLEY
18906|SANDYFIELD
18907|SANDYVILLE
18908|SANFORD
18909|SANGAREE
18910|SANGER
18911|SANGREY
18912|SANIBEL
18913|SANKERTOWN
18914|SANOSTEE
18915|SANS SOUCI
18916|SANSOM PARK
18917|SANTA
18918|SANTA ANA
18919|SANTA ANA HEIGHTS
18920|SANTA ANA PUEBLO
18921|SANTA ANNA
18922|SANTA BARBARA
18923|SANTA BÁRBARA COMUNIDAD
18924|SANTA CLARA
18925|SANTA CLARA COMUNIDAD
18926|SANTA CLARA PUEBLO
18927|SANTA CLARITA
18928|SANTA CLAUS
18929|SANTA CRUZ
18930|SANTA ELENA
18931|SANTA FE
18932|SANTA FE SPRINGS
18933|SANTA ISABEL
18934|SANTA ISABEL ZONA URBANA
18935|SANTA MARGARITA
18936|SANTA MARIA
18937|SANTA MONICA
18938|SANTA PAULA
18939|SANTA RITA
18940|SANTA ROSA
18941|SANTA ROSA BEACH
18942|SANTA ROSA COLONIA
18943|SANTA SUSANA
18944|SANTA TERESA
18945|SANTA VENETIA
18946|SANTA YNEZ
18947|SANTAQUIN
18948|SANTEE
18949|SANTIAGO
18950|SANTO
18951|SANTO DOMINGO
18952|SANTO DOMINGO COMUNIDAD
18953|SANTO DOMINGO PUEBLO
18954|SANTOS
18955|SAPELLO
18956|SAPELO ISLAND
18957|SAPPHO
18958|SAPPINGTON
18959|SAPULPA
18960|SARAGOSA
18961|SARAH
18962|SARAH ANN
18963|SARAHSVILLE
18964|SARALAND
18965|SARANAC
18966|SARANAC LAKE
18967|SARANAP
18968|SARASOTA
18969|SARASOTA SPRINGS
18970|SARATOGA
18971|SARATOGA SPRINGS
18972|SARBEN
18973|SARCOXIE
18974|SARDINIA
18975|SARDIS
18976|SARDIS CITY
18977|SAREPTA
18978|SARGEANT
18979|SARGENT
18980|SARGENTS
18981|SARITA
18982|SARLES
18983|SARONVILLE
18984|SARTELL
18985|SARVER
18986|SARVERSVILLE
18987|SASABE
18988|SASAKWA
18989|SASSER
18990|SATANTA
18991|SATARTIA
18992|SATELLITE BEACH
18993|SATICOY
18994|SATILLA
18995|SATIN
18996|SATOLAH
18997|SATSOP
18998|SATSUMA
18999|SATTLEY
19000|SATURN
19001|SAUCIER
19002|SAUGATUCK
19003|SAUGERTIES
19004|SAUGET
19005|SAUGUS
19006|SAUK CENTRE
19007|SAUK CITY
19008|SAUK RAPIDS
19009|SAUK VILLAGE
19010|SAUKVILLE
19011|SAULSBURY
19012|SAULT SAINTE MARIE
19013|SAUM
19014|SAUNDERS
19015|SAUNDERSTOWN
19016|SAUNEMIN
19017|SAUQUOIT
19018|SAUSALITO
19019|SAVAGE
19020|SAVAGE TOWN
19021|SAVAGEVILLE
19022|SAVANNA
19023|SAVANNAH
19024|SAVERY
19025|SAVONA
19026|SAVONBURG
19027|SAVOONGA
19028|SAVOY
19029|SAW CREEK
19030|SAWGRASS
19031|SAWMILL
19032|SAWMILLS
19033|SAWPIT
19034|SAWYER
19035|SAWYERS BAR
19036|SAWYERVILLE
19037|SAWYERWOOD
19038|SAXAPAHAW
19039|SAXE
19040|SAXIS
19041|SAXMAN
19042|SAXON
19043|SAXONBURG
19044|SAXTON
19045|SAXTONS RIVER
19046|SAYBROOK
19047|SAYBROOK MANOR
19048|SAYLORSBURG
19049|SAYLORVILLE
19050|SAYNER
19051|SAYRE
19052|SAYREVILLE
19053|SAYVILLE
19054|SCAGGSVILLE
19055|SCALES MOUND
19056|SCALLORN
19057|SCALP LEVEL
19058|SCALY MOUNTAIN
19059|SCAMMON
19060|SCAMMON BAY
19061|SCANDIA
19062|SCANDINAVIA
19063|SCANLON
19064|SCAPPOOSE
19065|SCARBORO
19066|SCARBOROUGH
19067|SCARBRO
19068|SCARLETS MILL
19069|SCARSDALE
19070|SCARVILLE
19071|SCENIC
19072|SCENIC OAKS
19073|SCHAAL
19074|SCHAEFFERSTOWN
19075|SCHAFFER
19076|SCHAGHTICOKE
19077|SCHALL CIRCLE
19078|SCHALLER
19079|SCHAUMBURG
19080|SCHELL CITY
19081|SCHELLSBURG
19082|SCHENECTADY
19083|SCHENEVUS
19084|SCHENLEY
19085|SCHERERVILLE
19086|SCHERR
19087|SCHERTZ
19088|SCHILLER PARK
19089|SCHLATER
19090|SCHLESWIG
19091|SCHLEY
19092|SCHLUSSER
19093|SCHNECKSVILLE
19094|SCHNEIDER
19095|SCHOENCHEN
19096|SCHOENECK
19097|SCHOFIELD
19098|SCHOHARIE
19099|SCHOLLE
19100|SCHOOLCRAFT
19101|SCHRAG
19102|SCHRAM CITY
19103|SCHRIEVER
19104|SCHROEDER
19105|SCHROON LAKE
19106|SCHUBERT
19107|SCHUCHK
19108|SCHULENBURG
19109|SCHULTE
19110|SCHULTER
19111|SCHULTZ
19112|SCHURZ
19113|SCHUYLER
19114|SCHUYLER LAKE
19115|SCHUYLERVILLE
19116|SCHUYLKILL HAVEN
19117|SCHWENKSVILLE
19118|SCIENCE HILL
19119|SCIO
19120|SCIOTA
19121|SCIOTO FURNACE
19122|SCIOTODALE
19123|SCIPIO
19124|SCITUATE
19125|SCOBEY
19126|SCOBEYVILLE
19127|SCOFIELD
19128|SCOOBA
19129|SCOTCHTOWN
19130|SCOTIA
19131|SCOTLAND
19132|SCOTLAND NECK
19133|SCOTLANDVILLE
19134|SCOTSDALE
19135|SCOTT CITY
19136|SCOTT DEPOT
19137|SCOTTDALE
19138|SCOTTS CORNERS
19139|SCOTTS HILL
19140|SCOTTS MILLS
19141|SCOTTS VALLEY
19142|SCOTTSBLUFF
19143|SCOTTSBORO
19144|SCOTTSBURG
19145|SCOTTSDALE
19146|SCOTTSMOOR
19147|SCOTTSVILLE
19148|SCOTTVILLE
19149|SCRANTON
19150|SCRAPER
19151|SCREVEN
19152|SCRIBNER
19153|SCURRY
19154|SEA BREEZE
19155|SEA BRIGHT
19156|SEA CLIFF
19157|SEA GIRT
19158|SEA ISLAND
19159|SEA ISLE CITY
19160|SEA RANCH
19161|SEA RANCH LAKES
19162|SEABECK
19163|SEABOARD
19164|SEABROOK
19165|SEABROOK BEACH
19166|SEABROOK FARMS
19167|SEABROOK ISLAND
19168|SEACLIFF
19169|SEADRIFT
19170|SEAFORD
19171|SEAFORTH
19172|SEAGOVILLE
19173|SEAGRAVES
19174|SEAGROVE
19175|SEAGROVE BEACH
19176|SEAHURST
19177|SEAL BEACH
19178|SEAL ROCK
19179|SEALE
19180|SEALEVEL
19181|SEALY
19182|SEAMA
19183|SEAMAN
19184|SEARCHLIGHT
19185|SEARCY
19186|SEARINGTOWN
19187|SEARLES
19188|SEARLES VALLEY
19189|SEARSBORO
19190|SEARSPORT
19191|SEASIDE
19192|SEASIDE HEIGHTS
19193|SEASIDE PARK
19194|SEAT PLEASANT
19195|SEATAC
19196|SEATON
19197|SEATONVILLE
19198|SEATTLE
19199|SEATTLE HEIGHTS
19200|SEBA DALKAI
19201|SEBASTIAN
19202|SEBASTOPOL
19203|SEBEKA
19204|SEBEWAING
19205|SEBOEIS
19206|SEBOYETA
19207|SEBREE
19208|SEBRELL
19209|SEBRING
19210|SECAUCUS
19211|SECO MINES
19212|SECOND MESA
19213|SECONSETT ISLAND
19214|SECOR
19215|SECRETARY
19216|SECTION
19217|SEDALIA
19218|SEDAN
19219|SEDGEFIELD
19220|SEDGEWICKVILLE
19221|SEDGWICK
19222|SEDILLO
19223|SEDLEY
19224|SEDONA
19225|SEDRO-WOOLLEY
19226|SEELEY
19227|SEELEY LAKE
19228|SEELYVILLE
19229|SEFFNER
19230|SEGNO
19231|SEGUIN
19232|SEGUNDO
19233|SEHILI
19234|SEIBERT
19235|SEILING
19236|SEKIU
19237|SELAH
19238|SELAWIK
19239|SELBY
19240|SELBYVILLE
19241|SELDEN
19242|SELDOVIA
19243|SELDOVIA VILLAGE
19244|SELFRIDGE
19245|SELIGMAN
19246|SELINSGROVE
19247|SELKIRK
19248|SELLECK
19249|SELLERS
19250|SELLERSBURG
19251|SELLERSVILLE
19252|SELLS
19253|SELMA
19254|SELMAN
19255|SELMAN CITY
19256|SELMER
19257|SELMONT
19258|SELTZER
19259|SELVIN
19260|SELZ
19261|SEMINARY
19262|SEMINOE DAM
19263|SEMINOLE
19264|SEMINOLE MANOR
19265|SEMMES
19266|SENA
19267|SENATH
19268|SENATOBIA
19269|SENECA
19270|SENECA FALLS
19271|SENECA GARDENS
19272|SENECA KNOLLS
19273|SENECAVILLE
19274|SENEY
19275|SENOIA
19276|SENTINEL
19277|SENTINEL BUTTE
19278|SEPAR
19279|SEQUIM
19280|SEQUNDO
19281|SEQUOYAH
19282|SERAFINA
19283|SERENA
19284|SERENADA
19285|SERGEANT BLUFF
19286|SERVIA
19287|SESPE
19288|SESSER
19289|SETAUKET
19290|SETH WARD
19291|SEVEN CORNERS
19292|SEVEN DEVILS
19293|SEVEN FIELDS
19294|SEVEN HILLS
19295|SEVEN LAKES
19296|SEVEN MILE
19297|SEVEN MILE FORD
19298|SEVEN OAKS
19299|SEVEN POINTS
19300|SEVEN SISTERS
19301|SEVEN SPRINGS
19302|SEVEN VALLEYS
19303|SEVENMILE
19304|SEVERANCE
19305|SEVERN
19306|SEVERNA PARK
19307|SEVERY
19308|SEVIER
19309|SEVIERVILLE
19310|SEVILLE
19311|SEWAL
19312|SEWALL'S POINT
19313|SEWANEE
19314|SEWARD
19315|SEWAREN
19316|SEWELL
19317|SEWICKLEY
19318|SEWICKLEY HEIGHTS
19319|SEWICKLEY HILLS
19320|SEXTON
19321|SEXTONVILLE
19322|SEYMOUR
19323|SEYMOURVILLE
19324|SHABBONA
19325|SHACKELFORD
19326|SHACKLE ISLAND
19327|SHADE
19328|SHADE GAP
19329|SHADEHILL
19330|SHADELAND
19331|SHADWELL
19332|SHADY
19333|SHADY COVE
19334|SHADY DALE
19335|SHADY GROVE
19336|SHADY HILLS
19337|SHADY HOLLOW
19338|SHADY POINT
19339|SHADY SHORES
19340|SHADY SIDE
19341|SHADY SPRING
19342|SHADYSIDE
19343|SHAFER
19344|SHAFTER
19345|SHAGELUK
19346|SHAKER HEIGHTS
19347|SHAKOPEE
19348|SHAKTOOLIK
19349|SHALIMAR
19350|SHALLOTTE
19351|SHALLOW WATER
19352|SHALLOWATER
19353|SHAMBAUGH
19354|SHAMOKIN
19355|SHAMOKIN DAM
19356|SHAMROCK
19357|SHAMROCK LAKES
19358|SHANDON
19359|SHANGHAI
19360|SHANIKO
19361|SHANKSVILLE
19362|SHANNON
19363|SHANNON CITY
19364|SHANNON HILLS
19365|SHANNONDALE
19366|SHARK RIVER HILLS
19367|SHARON
19368|SHARON HILL
19369|SHARON SPRINGS
19370|SHARONVILLE
19371|SHARPE
19372|SHARPES
19373|SHARPSBURG
19374|SHARPSVILLE
19375|SHARPTOWN
19376|SHARTLESVILLE
19377|SHASTA
19378|SHASTA LAKE
19379|SHATTUCK
19380|SHAUCK
19381|SHAVANO PARK
19382|SHAVER LAKE
19383|SHAVERTOWN
19384|SHAW
19385|SHAW HEIGHTS
19386|SHAW ISLAND
19387|SHAWAN
19388|SHAWANEE
19389|SHAWANO
19390|SHAWBORO
19391|SHAWHAN
19392|SHAWMUT
19393|SHAWNEE
19394|SHAWNEE HILLS
19395|SHAWNEE LAND
19396|SHAWNEETOWN
19397|SHAWSHEEN VILLAGE
19398|SHAWSVILLE
19399|SHAWVILLE
19400|SHAY
19401|SHEAKLEYVILLE
19402|SHEATOWN
19403|SHEBOYGAN
19404|SHEBOYGAN FALLS
19405|SHEDD
19406|SHEEP SPRINGS
19407|SHEFFIELD
19408|SHEFFIELD LAKE
19409|SHELBIANA
19410|SHELBINA
19411|SHELBURN
19412|SHELBURNE
19413|SHELBURNE FALLS
19414|SHELBY
19415|SHELBYVILLE
19416|SHELDAHL
19417|SHELDON
19418|SHELL
19419|SHELL BEACH
19420|SHELL KNOB
19421|SHELL LAKE
19422|SHELL POINT
19423|SHELL ROCK
19424|SHELL VALLEY
19425|SHELLEY
19426|SHELLMAN
19427|SHELLMAN BLUFF
19428|SHELLSBURG
19429|SHELLY
19430|SHELOCTA
19431|SHELTER COVE
19432|SHELTER ISLAND
19433|SHELTER ISLAND HEIGHTS
19434|SHELTON
19435|SHELTONS
19436|SHENANDOAH
19437|SHENANDOAH FARMS
19438|SHENANDOAH HEIGHTS
19439|SHENANDOAH JUNCTION
19440|SHENANDOAH RETREAT
19441|SHENANDOAH SHORES
19442|SHENOROCK
19443|SHEPARDSVILLE
19444|SHEPHERD
19445|SHEPHERDSTOWN
19446|SHEPHERDSVILLE
19447|SHEPPARD
19448|SHEPPERD
19449|SHEPPTON
19450|SHEPTON
19451|SHERACK
19452|SHERANDO
19453|SHERARD
19454|SHERBURN
19455|SHERBURNE
19456|SHERIDAN
19457|SHERIDAN BEACH
19458|SHERIDAN LAKE
19459|SHERMAN
19460|SHERMAN STATION
19461|SHERRARD
19462|SHERRELWOOD
19463|SHERRILL
19464|SHERRODSVILLE
19465|SHERWIN
19466|SHERWOOD
19467|SHERWOOD MANOR
19468|SHERWOOD SHORES
19469|SHESHEBEE
19470|SHEVLIN
19471|SHEYENNE
19472|SHICKLEY
19473|SHICKSHINNY
19474|SHIDLER
19475|SHIELDS
19476|SHILLINGTON
19477|SHILOH
19478|SHINDLER
19479|SHINER
19480|SHINGLE SPRINGS
19481|SHINGLEHOUSE
19482|SHINGLER
19483|SHINGLETON
19484|SHINGLETOWN
19485|SHINNECOCK HILLS
19486|SHINNSTON
19487|SHINROCK
19488|SHIOCTON
19489|SHIP BOTTOM
19490|SHIPLEY
19491|SHIPMAN
19492|SHIPPENSBURG
19493|SHIPPENVILLE
19494|SHIPPINGPORT
19495|SHIPROCK
19496|SHIPSHEWANA
19497|SHIREMANSTOWN
19498|SHIRLEY
19499|SHIRLEY MILLS
19500|SHIRLEYSBURG
19501|SHIRO
19502|SHISHMAREF
19503|SHIVELY
19504|SHIVERS
19505|SHIVWITS
19506|SHOAL CREEK DRIVE
19507|SHOAL CREEK ESTATES
19508|SHOALS
19509|SHOBONIER
19510|SHOEMAKERSVILLE
19511|SHOKAN
19512|SHOLES
19513|SHONGALOO
19514|SHONKIN
19515|SHONTO
19516|SHOOKS
19517|SHOP SPRINGS
19518|SHOPTON
19519|SHOPVILLE
19520|SHORE ACRES
19521|SHOREACRES
19522|SHOREHAM
19523|SHORELINE
19524|SHOREVIEW
19525|SHOREWOOD
19526|SHOREWOOD FOREST
19527|SHOREWOOD HILLS
19528|SHORT CREEK
19529|SHORT HILLS
19530|SHORT PUMP
19531|SHORTER
19532|SHORTERVILLE
19533|SHORTSVILLE
19534|SHOSHONE
19535|SHOSHONI
19536|SHOUNS
19537|SHOUP
19538|SHOVELTOWN
19539|SHOW LOW
19540|SHREVE
19541|SHREVEPORT
19542|SHREWSBURY
19543|SHRUB OAK
19544|SHUBERT
19545|SHUBUTA
19546|SHUEYVILLE
19547|SHULERVILLE
19548|SHULLSBURG
19549|SHUMWAY
19550|SHUNGNAK
19551|SHUQUALAK
19552|SIAM
19553|SIASCONSET
19554|SIBLEY
19555|SICARD
19556|SICILY ISLAND
19557|SICKLERVILLE
19558|SIDELL
19559|SIDMAN
19560|SIDNAW
19561|SIDNEY
19562|SIDNEY CENTER
19563|SIDON
19564|SIENNA PLANTATION
19565|SIEPER
19566|SIERRA BLANCA
19567|SIERRA BROOKS
19568|SIERRA CITY
19569|SIERRA MADRE
19570|SIERRA VIEW
19571|SIERRA VILLAGE
19572|SIERRA VISTA
19573|SIERRAVILLE
19574|SIESTA ACRES
19575|SIESTA KEY
19576|SIESTA SHORES
19577|SIGEL
19578|SIGLERVILLE
19579|SIGNAL HILL
19580|SIGNAL MOUNTAIN
19581|SIGOURNEY
19582|SIGSBEE
19583|SIGURD
19584|SIKES
19585|SIKESTON
19586|SIL NAKYA
19587|SILAS
19588|SILCO
19589|SILER CITY
19590|SILERTON
19591|SILESIA
19592|SILETZ
19593|SILEX
19594|SILICA
19595|SILIO
19596|SILK HOPE
19597|SILKWORTH
19598|SILO
19599|SILOAM
19600|SILOAM SPRINGS
19601|SILSBEE
19602|SILT
19603|SILTCOOS
19604|SILVA
19605|SILVANA
19606|SILVER
19607|SILVER BAY
19608|SILVER CITY
19609|SILVER CLIFF
19610|SILVER CREEK
19611|SILVER FIRS
19612|SILVER GATE
19613|SILVER GROVE
19614|SILVER HILL
19615|SILVER LAKE
19616|SILVER LAKES
19617|SILVER PEAK
19618|SILVER PLUME
19619|SILVER RIDGE
19620|SILVER SPRING
19621|SILVER SPRINGS
19622|SILVER SPRINGS SHORES
19623|SILVER STAR
19624|SILVER VALLEY
19625|SILVERADO
19626|SILVERDALE
19627|SILVERHILL
19628|SILVERSTREET
19629|SILVERTHORNE
19630|SILVERTIP
19631|SILVERTON
19632|SILVERVILLE
19633|SILVIES
19634|SILVIS
19635|SIMCOE
19636|SIMI VALLEY
19637|SIMILK BEACH
19638|SIMLA
19639|SIMMESPORT
19640|SIMMONS
19641|SIMMS
19642|SIMNASHO
19643|SIMONS
19644|SIMONTON
19645|SIMONTON LAKE
19646|SIMPSON
19647|SIMPSONS
19648|SIMPSONVILLE
19649|SIMS
19650|SIMS CHAPEL
19651|SIMSBORO
19652|SINAI
19653|SINCLAIR
19654|SINCLAIRVILLE
19655|SINGAC
19656|SINGER
19657|SINGLETON
19658|SINK CREEK
19659|SINKING SPRING
19660|SINTON
19661|SIOUX CENTER
19662|SIOUX CITY
19663|SIOUX FALLS
19664|SIOUX PASS
19665|SIOUX RAPIDS
19666|SIPSEY
19667|SIRACUSAVILLE
19668|SIREN
19669|SIRMANS
19670|SISCO HEIGHTS
19671|SISQUOC
19672|SISSETON
19673|SISSONVILLE
19674|SISTER BAY
19675|SISTER LAKES
19676|SISTERS
19677|SISTERSVILLE
19678|SITKA
19679|SIX MILE
19680|SIXES
19681|SIXTEEN
19682|SIXTEEN MILE STAND
19683|SKAGWAY
19684|SKAMOKAWA
19685|SKANEATELES
19686|SKEDEE
19687|SKELLYTOWN
19688|SKENE
19689|SKIATOOK
19690|SKIDAWAY ISLAND
19691|SKIDDY
19692|SKIDMORE
19693|SKIDWAY LAKE
19694|SKILLMAN
19695|SKIME
19696|SKIPPACK
19697|SKIPPERS CORNER
19698|SKIPPERTON
19699|SKIPTON
19700|SKOKIE
19701|SKOKOMISH
19702|SKOWHEGAN
19703|SKULL VALLEY
19704|SKWENTNA
19705|SKY LAKE
19706|SKY LONDA
19707|SKY VALLEY
19708|SKYFOREST
19709|SKYKOMISH
19710|SKYLAND
19711|SKYLAND ESTATES
19712|SKYLINE
19713|SKYLINE ACRES
19714|SKYLINE VIEW
19715|SKYWAY
19716|SLABTOWN
19717|SLACKWOODS
19718|SLADE
19719|SLAGLE
19720|SLANA
19721|SLANESVILLE
19722|SLAPOUT
19723|SLATE LICK
19724|SLATE SPRING
19725|SLATEDALE
19726|SLATER
19727|SLATERVILLE SPRINGS
19728|SLATINGTON
19729|SLATON
19730|SLATY FORK
19731|SLAUGHTER
19732|SLAUGHTER BEACH
19733|SLAUGHTERS
19734|SLAUGHTERVILLE
19735|SLAYDEN
19736|SLAYTON
19737|SLEDGE
19738|SLEEPER
19739|SLEEPY EYE
19740|SLEEPY HOLLOW
19741|SLEETMUTE
19742|SLEMP
19743|SLICK
19744|SLICKVILLE
19745|SLIDELL
19746|SLIGO
19747|SLINGER
19748|SLIPPERY ROCK
19749|SLOAN
19750|SLOAT
19751|SLOATSBURG
19752|SLOCOMB
19753|SLOCUM
19754|SLOVAN
19755|SMACKOVER
19756|SMALE
19757|SMALLEYTOWN
19758|SMALLWOOD
19759|SMARR
19760|SMARTSVILLE
19761|SMELTERTOWN
19762|SMELTERVILLE
19763|SMETHPORT
19764|SMICKSBURG
19765|SMILEY
19766|SMILEY PARK
19767|SMITH
19768|SMITH CENTER
19769|SMITH CORNER
19770|SMITH ISLAND
19771|SMITH MILLS
19772|SMITH POINT
19773|SMITH RIVER
19774|SMITH VILLAGE
19775|SMITHBORO
19776|SMITHBURG
19777|SMITHDALE
19778|SMITHERS
19779|SMITHFIELD
19780|SMITHLAND
19781|SMITHS CREEK
19782|SMITHS FERRY
19783|SMITHS GROVE
19784|SMITHS STATION
19785|SMITHSBURG
19786|SMITHTON
19787|SMITHTOWN
19788|SMITHVILLE
19789|SMITHVILLE FLATS
19790|SMITHWICK
19791|SMOAKS
19792|SMOCK
19793|SMOKE BEND
19794|SMOKE RISE
19795|SMOKETOWN
19796|SMOLAN
19797|SMOOT
19798|SMYER
19799|SMYRNA
19800|SMYRNA MILLS
19801|SNAKE CREEK
19802|SNAPFINGER
19803|SNEAD
19804|SNEADS
19805|SNEADS FERRY
19806|SNEEDVILLE
19807|SNELL
19808|SNELLING
19809|SNELLVILLE
19810|SNIDER
19811|SNOHOMISH
19812|SNOOK
19813|SNOQUALMIE
19814|SNOQUALMIE FALLS
19815|SNOQUALMIE PASS
19816|SNOVER
19817|SNOW HILL
19818|SNOW LAKE
19819|SNOW LAKE SHORES
19820|SNOW SHOE
19821|SNOWBALL
19822|SNOWDOUN
19823|SNOWFLAKE
19824|SNOWMASS
19825|SNOWMASS VILLAGE
19826|SNOWVILLE
19827|SNYDER
19828|SNYDERTOWN
19829|SNYDERVILLE
19830|SOAP LAKE
19831|SOBIESKI
19832|SOCASTEE
19833|SOCIAL CIRCLE
19834|SOCIAL HILL
19835|SOCIALVILLE
19836|SOCIETY HILL
19837|SOCORRO
19838|SODA BAY
19839|SODA SPRINGS
19840|SODAVILLE
19841|SODDY-DAISY
19842|SODERVILLE
19843|SODUS
19844|SODUS POINT
19845|SOFIA
19846|SOHAM
19847|SOLANA
19848|SOLANA BEACH
19849|SOLANO
19850|SOLDIER
19851|SOLDIER CREEK
19852|SOLDIER POND
19853|SOLDIER SUMMIT
19854|SOLDIERS GROVE
19855|SOLDOTNA
19856|SOLEDAD
19857|SOLEN
19858|SOLIS
19859|SOLITUDE
19860|SOLOMON
19861|SOLOMONS
19862|SOLON
19863|SOLON SPRINGS
19864|SOLROMAR
19865|SOLVANG
19866|SOLVAY
19867|SOLWAY
19868|SOMBRILLO
19869|SOMERDALE
19870|SOMERS
19871|SOMERS POINT
19872|SOMERSET
19873|SOMERSWORTH
19874|SOMERTON
19875|SOMERVILLE
19876|SOMES BAR
19877|SOMESVILLE
19878|SOMIS
19879|SOMONAUK
19880|SONDHEIMER
19881|SONESTOWN
19882|SONNETTE
19883|SONOITA
19884|SONOMA
19885|SONORA
19886|SONTAG
19887|SONTERRA
19888|SOPCHOPPY
19889|SOPER
19890|SOPERTON
19891|SOPHIA
19892|SOQUEL
19893|SORENTO
19894|SORREL
19895|SORRENTO
19896|SORUM
19897|SOSO
19898|SOUDAN
19899|SOUDERSBURG
19900|SOUDERTON
19901|SOULSBYVILLE
19902|SOUND BEACH
19903|SOUR LAKE
19904|SOURIS
19905|SOUTH ACTON
19906|SOUTH ALAMO
19907|SOUTH AMANA
19908|SOUTH AMBOY
19909|SOUTH AMHERST
19910|SOUTH APOPKA
19911|SOUTH ASHBURNHAM
19912|SOUTH BARRE
19913|SOUTH BARRINGTON
19914|SOUTH BAY
19915|SOUTH BEACH
19916|SOUTH BELOIT
19917|SOUTH BEND
19918|SOUTH BETHANY
19919|SOUTH BETHLEHEM
19920|SOUTH BLOOMFIELD
19921|SOUTH BLOOMING GROVE
19922|SOUTH BLOOMINGVILLE
19923|SOUTH BOARDMAN
19924|SOUTH BOSTON
19925|SOUTH BOUND BROOK
19926|SOUTH BRADENTON
19927|SOUTH BRANCH
19928|SOUTH BROADWAY
19929|SOUTH BROOKSVILLE
19930|SOUTH BROWNING
19931|SOUTH BURLINGTON
19932|SOUTH CANAL
19933|SOUTH CARROLLTON
19934|SOUTH CARTHAGE
19935|SOUTH CHARLESTON
19936|SOUTH CHELMSFORD
19937|SOUTH CHESCONESSEX
19938|SOUTH CHICAGO HEIGHTS
19939|SOUTH CHINA
19940|SOUTH CLE ELUM
19941|SOUTH CLEVELAND
19942|SOUTH COATESVILLE
19943|SOUTH COFFEYVILLE
19944|SOUTH COLTON
19945|SOUTH CONGAREE
19946|SOUTH CONNELLSVILLE
19947|SOUTH CORNING
19948|SOUTH COVENTRY
19949|SOUTH DARTMOUTH
19950|SOUTH DAYTON
19951|SOUTH DAYTONA
19952|SOUTH DEERFIELD
19953|SOUTH DENNIS
19954|SOUTH DOS PALOS
19955|SOUTH DUXBURY
19956|SOUTH EL MONTE
19957|SOUTH ELGIN
19958|SOUTH ELIOT
19959|SOUTH ENGLISH
19960|SOUTH EUCLID
19961|SOUTH FALLSBURG
19962|SOUTH FARMINGDALE
19963|SOUTH FLORAL PARK
19964|SOUTH FONTANA
19965|SOUTH FORK
19966|SOUTH FORK ESTATES
19967|SOUTH FULTON
19968|SOUTH GARCIA
19969|SOUTH GASTONIA
19970|SOUTH GATE
19971|SOUTH GATE RIDGE
19972|SOUTH GLASTONBURY
19973|SOUTH GLENS FALLS
19974|SOUTH GREELEY
19975|SOUTH GREENFIELD
19976|SOUTH GREENSBURG
19977|SOUTH GULL LAKE
19978|SOUTH HAVEN
19979|SOUTH HEART
19980|SOUTH HEIGHTS
19981|SOUTH HEMPSTEAD
19982|SOUTH HENDERSON
19983|SOUTH HIGHPOINT
19984|SOUTH HILL
19985|SOUTH HOLLAND
19986|SOUTH HOOKSETT
19987|SOUTH HOUSTON
19988|SOUTH HUNTINGTON
19989|SOUTH HUTCHINSON
19990|SOUTH JACKSONVILLE
19991|SOUTH JORDAN
19992|SOUTH KENSINGTON
19993|SOUTH KOMELIK
19994|SOUTH LAGRANGE
19995|SOUTH LAGUNA
19996|SOUTH LAKE
19997|SOUTH LAKE TAHOE
19998|SOUTH LANCASTER
19999|SOUTH LAUREL
20000|SOUTH LEAD HILL
20001|SOUTH LEBANON
20002|SOUTH LIMA
20003|SOUTH LINEVILLE
20004|SOUTH LOCKPORT
20005|SOUTH LYON
20006|SOUTH MANSFIELD
20007|SOUTH MIAMI
20008|SOUTH MIAMI HEIGHTS
20009|SOUTH MILLS
20010|SOUTH MILWAUKEE
20011|SOUTH MONROE
20012|SOUTH MONTROSE
20013|SOUTH MOUND
20014|SOUTH MOUNTAIN
20015|SOUTH NAKNEK
20016|SOUTH NEW BERLIN
20017|SOUTH NEW CASTLE
20018|SOUTH NEWPORT
20019|SOUTH NYACK
20020|SOUTH OGDEN
20021|SOUTH OROVILLE
20022|SOUTH OTSELIC
20023|SOUTH PADRE ISLAND
20024|SOUTH PALM BEACH
20025|SOUTH PARIS
20026|SOUTH PARK
20027|SOUTH PARK VIEW
20028|SOUTH PASADENA
20029|SOUTH PASS CITY
20030|SOUTH PATRICK SHORES
20031|SOUTH PEKIN
20032|SOUTH PERRY
20033|SOUTH PHILIPSBURG
20034|SOUTH PITTSBURG
20035|SOUTH PLAINFIELD
20036|SOUTH PLAINS
20037|SOUTH PLATTE
20038|SOUTH POINT
20039|SOUTH PONTE VEDRA BEACH
20040|SOUTH PORTLAND
20041|SOUTH POTTSTOWN
20042|SOUTH PRAIRIE
20043|SOUTH PUNTA GORDA HEIGHTS
20044|SOUTH RANGE
20045|SOUTH RENOVO
20046|SOUTH RICHMOND HILL
20047|SOUTH RIDING
20048|SOUTH RIVER
20049|SOUTH ROCKWOOD
20050|SOUTH ROSEMARY
20051|SOUTH ROXANA
20052|SOUTH ROYALTON
20053|SOUTH RUSSELL
20054|SOUTH SAINT PAUL
20055|SOUTH SALEM
20056|SOUTH SALT LAKE
20057|SOUTH SAN FRANCISCO
20058|SOUTH SAN GABRIEL
20059|SOUTH SAN JOSE HILLS
20060|SOUTH SANFORD
20061|SOUTH SARASOTA
20062|SOUTH SHAFTSBURY
20063|SOUTH SHORE
20064|SOUTH SIOUX CITY
20065|SOUTH SNOHOMISH
20066|SOUTH SOLON
20067|SOUTH SUMTER
20068|SOUTH SUPERIOR
20069|SOUTH TAFT
20070|SOUTH TEMPLE
20071|SOUTH TOLEDO BEND
20072|SOUTH TOMS RIVER
20073|SOUTH TORRINGTON
20074|SOUTH TUCSON
20075|SOUTH TUNNEL
20076|SOUTH UNIONTOWN
20077|SOUTH VACHERIE
20078|SOUTH VALLEY
20079|SOUTH VALLEY STREAM
20080|SOUTH VENICE
20081|SOUTH VIENNA
20082|SOUTH VINEMONT
20083|SOUTH WADESBORO
20084|SOUTH WALLINS
20085|SOUTH WALPOLE
20086|SOUTH WAVERLY
20087|SOUTH WAYNE
20088|SOUTH WEBER
20089|SOUTH WEBSTER
20090|SOUTH WELDON
20091|SOUTH WEST CITY
20092|SOUTH WESTPORT
20093|SOUTH WHITLEY
20094|SOUTH WHITTIER
20095|SOUTH WILLARD
20096|SOUTH WILLIAMSON
20097|SOUTH WILLIAMSPORT
20098|SOUTH WILMINGTON
20099|SOUTH WILSON
20100|SOUTH WINDHAM
20101|SOUTH WOODSTOCK
20102|SOUTH YARMOUTH
20103|SOUTH ZANESVILLE
20104|SOUTHAM
20105|SOUTHAMPTON
20106|SOUTHARD
20107|SOUTHAVEN
20108|SOUTHCHASE
20109|SOUTHDOWN
20110|SOUTHERN PINES
20111|SOUTHERN SHOPS
20112|SOUTHERN SHORES
20113|SOUTHERN VIEW
20114|SOUTHFIELD
20115|SOUTHFIELDS
20116|SOUTHGATE
20117|SOUTHINGTON
20118|SOUTHLAKE
20119|SOUTHLAND
20120|SOUTHMAYD
20121|SOUTHMONT
20122|SOUTHOLD
20123|SOUTHPORT
20124|SOUTHSIDE
20125|SOUTHSIDE PLACE
20126|SOUTHTON
20127|SOUTHVIEW
20128|SOUTHVILLE
20129|SOUTHWEST
20130|SOUTHWEST GREENSBURG
20131|SOUTHWEST HARBOR
20132|SOUTHWEST RANCHES
20133|SOUTHWOOD ACRES
20134|SOUTHWORTH
20135|SPACKENKILL
20136|SPADE
20137|SPALDING
20138|SPANAWAY
20139|SPANGLE
20140|SPANISH FORK
20141|SPANISH FORT
20142|SPANISH LAKE
20143|SPANISH SPRINGS
20144|SPANISH VALLEY
20145|SPARGURSVILLE
20146|SPARKILL
20147|SPARKMAN
20148|SPARKS
20149|SPARKSVILLE
20150|SPARLAND
20151|SPARLINGVILLE
20152|SPARR
20153|SPARTA
20154|SPARTANBURG
20155|SPARTANSBURG
20156|SPAULDING
20157|SPAVINAW
20158|SPEAKS
20159|SPEAR
20160|SPEARFISH
20161|SPEARMAN
20162|SPEARSVILLE
20163|SPEARVILLE
20164|SPECULATOR
20165|SPEEDWAY
20166|SPEER
20167|SPEERS
20168|SPEIGHT
20169|SPELTER
20170|SPENARD
20171|SPENCER MOUNTAIN
20172|SPENCERPORT
20173|SPENCERVILLE
20174|SPEONK
20175|SPERRY
20176|SPERRYVILLE
20177|SPICELAND
20178|SPICER
20179|SPICKARD
20180|SPILLERTOWN
20181|SPILLVILLE
20182|SPINDALE
20183|SPINK
20184|SPINNERSTOWN
20185|SPIRIT LAKE
20186|SPIRITWOOD
20187|SPIRITWOOD LAKE
20188|SPIRO
20189|SPIVEY
20190|SPIVEYS CORNER
20191|SPLENDORA
20192|SPOFFORD
20193|SPOKANE
20194|SPOKANE VALLEY
20195|SPOONER
20196|SPORTSMEN ACRES
20197|SPOTSWOOD
20198|SPOTSYLVANIA
20199|SPOTSYLVANIA COURTHOUSE
20200|SPOTTED HORSE
20201|SPOTTSVILLE
20202|SPRABERRY
20203|SPRAGUE
20204|SPRAGUE RIVER
20205|SPRAGUEVILLE
20206|SPREAD EAGLE
20207|SPRECKELS
20208|SPRING
20209|SPRING ARBOR
20210|SPRING BAY
20211|SPRING BRANCH
20212|SPRING BROOK
20213|SPRING CHURCH
20214|SPRING CITY
20215|SPRING CREEK
20216|SPRING GAP
20217|SPRING GARDEN
20218|SPRING GARDENS
20219|SPRING GLEN
20220|SPRING GREEN
20221|SPRING GROVE
20222|SPRING HILL
20223|SPRING HILLS
20224|SPRING HOPE
20225|SPRING HOUSE
20226|SPRING LAKE
20227|SPRING LAKE HEIGHTS
20228|SPRING LAKE PARK
20229|SPRING MILL
20230|SPRING MILLS
20231|SPRING MOUNT
20232|SPRING PARK
20233|SPRING PLACE
20234|SPRING RIDGE
20235|SPRING VALLEY
20236|SPRING VALLEY LAKE
20237|SPRINGBORO
20238|SPRINGBROOK
20239|SPRINGDALE
20240|SPRINGER
20241|SPRINGERTON
20242|SPRINGERVILLE
20243|SPRINGFIELD
20244|SPRINGFIELD GARDENS
20245|SPRINGHILL
20246|SPRINGLAKE
20247|SPRINGMONT
20248|SPRINGPORT
20249|SPRINGS
20250|SPRINGSIDE
20251|SPRINGTOWN
20252|SPRINGVALE
20253|SPRINGVIEW
20254|SPRINGVILLE
20255|SPROTT
20256|SPROUT
20257|SPRUCE PINE
20258|SPRY
20259|SPUR
20260|SPURGEON
20261|SPURGER
20262|SQUARE BUTTE
20263|SQUAW LAKE
20264|SQUAW VALLEY
20265|SQUIRE
20266|SQUIRES
20267|SQUIRREL MOUNTAIN VALLEY
20268|ST. JOHN
20269|STAATSBURG
20270|STACEY STREET
20271|STACY
20272|STACYVILLE
20273|STAFFORD
20274|STAFFORD SPRINGS
20275|STAGECOACH
20276|STAIRTOWN
20277|STALEY
20278|STALLINGS
20279|STALLION SPRINGS
20280|STALLO
20281|STALWART
20282|STAMFORD
20283|STAMPING GROUND
20284|STAMPLEY
20285|STANAFORD
20286|STANARDSVILLE
20287|STANBERRY
20288|STANCHFIELD
20289|STANDARD CITY
20290|STANDING PINE
20291|STANDING ROCK
20292|STANDISH
20293|STANDROD
20294|STANFIELD
20295|STANFORD
20296|STANHOPE
20297|STANLEY PARK
20298|STANLEYTOWN
20299|STANLEYVILLE
20300|STANNARDS
20301|STANSBURY PARK
20302|STANTON
20303|STANTONSBURG
20304|STANTONVILLE
20305|STANWOOD
20306|STAPLEHURST
20307|STAPLETON
20308|STAR CITY
20309|STAR CROSS
20310|STAR HARBOR
20311|STAR JUNCTION
20312|STAR LAKE
20313|STAR PRAIRIE
20314|STAR VALLEY
20315|STAR VALLEY RANCH
20316|STARBRICK
20317|STARBUCK
20318|STARK
20319|STARK CITY
20320|STARKE
20321|STARKEY
20322|STARKS
20323|STARKVILLE
20324|STARKWEATHER
20325|STARR
20326|STARR SCHOOL
20327|STARRS MILL
20328|STARRSVILLE
20329|STARRUCCA
20330|STARTEX
20331|STATE BRIDGE
20332|STATE CENTER
20333|STATE COLLEGE
20334|STATE LINE
20335|STATE LINE VILLAGE
20336|STATE PARK PLACE
20337|STATE ROAD
20338|STATEBURG
20339|STATELINE
20340|STATEN ISLAND
20341|STATENVILLE
20342|STATESBORO
20343|STATESVILLE
20344|STATHAM
20345|STAUNTON
20346|STAVES
20347|STAYTON
20348|STEAMBOAT
20349|STEAMBOAT ROCK
20350|STEAMBOAT SPRINGS
20351|STEARNS
20352|STEBBINS
20353|STECKER
20354|STEDMAN
20355|STEELE
20356|STEELE CITY
20357|STEELEVILLE
20358|STEELTON
20359|STEELVILLE
20360|STEEN
20361|STEENS
20362|STEEP FALLS
20363|STEGER
20364|STEHEKIN
20365|STEILACOOM
20366|STEINAUER
20367|STEINHATCHEE
20368|STELLA
20369|STELLA COMUNIDAD
20370|STELLA NIAGARA
20371|STENNETT
20372|STEPHAN
20373|STEPHEN
20374|STEPHEN CREEK
20375|STEPHENS
20376|STEPHENS CITY
20377|STEPHENSBURG
20378|STEPHENSON
20379|STEPHENVILLE
20380|STEPROCK
20381|STEPTOE
20382|STERLEY
20383|STERLING
20384|STERLING CITY
20385|STERLING FOREST
20386|STERLING HEIGHTS
20387|STERLING RUN
20388|STERLINGTON
20389|STERRETT
20390|STETSONVILLE
20391|STEUBEN
20392|STEUBENVILLE
20393|STEVENS CREEK
20394|STEVENS POINT
20395|STEVENS VILLAGE
20396|STEVENSON
20397|STEVENSTOWN
20398|STEVENSVILLE
20399|STEVINSON
20400|STEWARD
20401|STEWARDSON
20402|STEWART
20403|STEWART MANOR
20404|STEWARTSTOWN
20405|STEWARTSVILLE
20406|STEWARTVILLE
20407|STICKNEY
20408|STIDHAM
20409|STIGLER
20410|STILES
20411|STILESVILLE
20412|STILL POND
20413|STILL RIVER
20414|STILLINGS
20415|STILLMAN VALLEY
20416|STILLMORE
20417|STILLWATER
20418|STILLWELL
20419|STILSON
20420|STILWELL
20421|STINESVILLE
20422|STINNETT
20423|STINSON BEACH
20424|STIPPVILLE
20425|STIRLING
20426|STIRLING CITY
20427|STIRRAT
20428|STITES
20429|STITZER
20430|STOBO
20431|STOCK ISLAND
20432|STOCKBRIDGE
20433|STOCKDALE
20434|STOCKERTOWN
20435|STOCKETT
20436|STOCKHAM
20437|STOCKHOLM
20438|STOCKLAND
20439|STOCKMAN
20440|STOCKPORT
20441|STOCKTON
20442|STOCKVILLE
20443|STOCKWELL
20444|STODDARD
20445|STOKES
20446|STOKESDALE
20447|STOLLE
20448|STOLLINGS
20449|STONE CITY
20450|STONE CREEK
20451|STONE HARBOR
20452|STONE LAKE
20453|STONE MOUNTAIN
20454|STONE PARK
20455|STONE RIDGE
20456|STONEBANK
20457|STONEBORO
20458|STONEBURG
20459|STONECREST
20460|STONEFORT
20461|STONEGA
20462|STONEGATE
20463|STONEHAM
20464|STONER
20465|STONERSTOWN
20466|STONEVILLE
20467|STONEWALL
20468|STONEWALL GAP
20469|STONEWOOD
20470|STONEY POINT
20471|STONINGTON
20472|STONY BROOK
20473|STONY CREEK
20474|STONY CREEK MILLS
20475|STONY LAKE
20476|STONY POINT
20477|STONY PRAIRIE
20478|STONY RIDGE
20479|STONY RIVER
20480|STONYBROOK
20481|STONYFORD
20482|STORDEN
20483|STORLA
20484|STORM LAKE
20485|STORMSTOWN
20486|STORRIE
20487|STORRS
20488|STORY CITY
20489|STOTESBURY
20490|STOTTS CITY
20491|STOTTVILLE
20492|STOUCHSBURG
20493|STOUGHTON
20494|STOUTLAND
20495|STOUTSVILLE
20496|STOVALL
20497|STOVER
20498|STOW
20499|STOWE
20500|STOWELL
20501|STOY
20502|STOYSTOWN
20503|STRABANE
20504|STRAFFORD
20505|STRAHAN
20506|STRANDBURG
20507|STRANDELL
20508|STRANDQUIST
20509|STRANG
20510|STRANGE CREEK
20511|STRASBURG
20512|STRATFORD
20513|STRATHCONA
20514|STRATHMERE
20515|STRATHMOOR MANOR
20516|STRATHMOOR VILLAGE
20517|STRATHMORE
20518|STRATMOOR
20519|STRATTANVILLE
20520|STRATTON
20521|STRAUGHN
20522|STRAUSS
20523|STRAUSSTOWN
20524|STRAWBERRY
20525|STRAWBERRY PLAINS
20526|STRAWBERRY POINT
20527|STRAWN
20528|STREAMWOOD
20529|STREATOR
20530|STREETER
20531|STREETMAN
20532|STREETSBORO
20533|STREVELL
20534|STRING PRAIRIE
20535|STRINGER
20536|STRINGTOWN
20537|STRODES MILLS
20538|STROH
20539|STROMSBURG
20540|STRONACH
20541|STRONG CITY
20542|STRONGHURST
20543|STRONGSVILLE
20544|STROUD
20545|STROUDSBURG
20546|STRUBLE
20547|STRUM
20548|STRUTHERS
20549|STRYKER
20550|STRYKERSVILLE
20551|STUART
20552|STUARTS DRAFT
20553|STUCKEY
20554|STUDLEY
20555|STUDY BUTTE
20556|STULL
20557|STUMPY POINT
20558|STURBRIDGE
20559|STURGEON
20560|STURGEON BAY
20561|STURGEON LAKE
20562|STURGIS
20563|STURKIE
20564|STURTEVANT
20565|STUTTGART
20566|SUAMICO
20567|SUBIACO
20568|SUBLETT
20569|SUBLETTE
20570|SUBLIME
20571|SUBLIMITY
20572|SUCCASUNNA
20573|SUDAN
20574|SUDDEN VALLEY
20575|SUDLERSVILLE
20576|SUDLEY
20577|SUFFERN
20578|SUFFIELD DEPOT
20579|SUFFOLK
20580|SUGAR BUSH
20581|SUGAR BUSH KNOLLS
20582|SUGAR CITY
20583|SUGAR CREEK
20584|SUGAR GROVE
20585|SUGAR HILL
20586|SUGAR LAND
20587|SUGAR MOUNTAIN
20588|SUGAR NOTCH
20589|SUGAR TREE RIDGE
20590|SUGAR VALLEY
20591|SUGARCREEK
20592|SUGARLAND RUN
20593|SUGARLOAF
20594|SUGARLOAF MOUNTAIN PARK
20595|SUGARLOAF SAW MILL
20596|SUGARLOAF VILLAGE
20597|SUGARMILL WOODS
20598|SUGARTOWN
20599|SUGARVILLE
20600|SUGDEN
20601|SUISUN
20602|SUITLAND
20603|SULA
20604|SULLIGENT
20605|SULLIVAN
20606|SULLIVAN CITY
20607|SULLIVANS ISLAND
20608|SULLY
20609|SULPHUR
20610|SULPHUR BLUFF
20611|SULPHUR ROCK
20612|SULPHUR SPRINGS
20613|SULPHURDALE
20614|SULTAN
20615|SULTANA
20616|SUMAC
20617|SUMAS
20618|SUMATRA
20619|SUMIDERO
20620|SUMITON
20621|SUMMER HAVEN
20622|SUMMER LAKE
20623|SUMMER SHADE
20624|SUMMERDALE
20625|SUMMERFIELD
20626|SUMMERHAVEN
20627|SUMMERHILL
20628|SUMMERLAND
20629|SUMMERLAND KEY
20630|SUMMERS
20631|SUMMERSET
20632|SUMMERSIDE
20633|SUMMERSVILLE
20634|SUMMERTON
20635|SUMMERTOWN
20636|SUMMERVILLE
20637|SUMMIT
20638|SUMMIT CORNERS
20639|SUMMIT HILL
20640|SUMMIT LAKE
20641|SUMMIT PARK
20642|SUMMIT STATION
20643|SUMMITVIEW
20644|SUMMITVILLE
20645|SUMMUM
20646|SUMNER
20647|SUMPTER
20648|SUMRALL
20649|SUMTER
20650|SUMTERVILLE
20651|SUN CITY
20652|SUN CITY CENTER
20653|SUN CITY WEST
20654|SUN LAKES
20655|SUN PRAIRIE
20656|SUN RIVER
20657|SUN RIVER TERRACE
20658|SUN VALLEY
20659|SUNBEAM
20660|SUNBRIGHT
20661|SUNBURG
20662|SUNBURST
20663|SUNBURY
20664|SUNCOAST ESTATES
20665|SUNCOOK
20666|SUNCREST
20667|SUNDANCE
20668|SUNDERLAND
20669|SUNDOWN
20670|SUNFIELD
20671|SUNFISH LAKE
20672|SUNFLOWER
20673|SUNIZONA
20674|SUNLAND PARK
20675|SUNMAN
20676|SUNNILAND
20677|SUNNY CREST
20678|SUNNY ISLES BEACH
20679|SUNNY SIDE
20680|SUNNY SOUTH
20681|SUNNYBROOK
20682|SUNNYDALE
20683|SUNNYMEAD
20684|SUNNYSIDE
20685|SUNNYSLOPE
20686|SUNNYVALE
20687|SUNOL
20688|SUNRAY
20689|SUNRISE
20690|SUNRISE BEACH
20691|SUNRISE BEACH VILLAGE
20692|SUNRISE LAKE
20693|SUNRISE MANOR
20694|SUNRIVER
20695|SUNSET
20696|SUNSET ACRES COLONIA
20697|SUNSET BAY
20698|SUNSET BEACH
20699|SUNSET COLONIA
20700|SUNSET HILLS
20701|SUNSET VALLEY
20702|SUNSET VILLAGE
20703|SUNSHINE
20704|SUNTRANA
20705|SUPAI
20706|SUPERIOR
20707|SUPERIOR VILLAGE
20708|SUPREME
20709|SUQUALENA
20710|SUQUAMISH
20711|SURF CITY
20712|SURFSIDE
20713|SURFSIDE BEACH
20714|SURGOINSVILLE
20715|SURING
20716|SURPRISE
20717|SURRENCY
20718|SURREY
20719|SURRY
20720|SUSAN MOORE
20721|SUSANK
20722|SUSANVILLE
20723|SUSITNA
20724|SUSQUEHANNA
20725|SUSQUEHANNA TRAILS
20726|SUSSEX
20727|SUTCLIFFE
20728|SUTERSVILLE
20729|SUTHERLAND
20730|SUTHERLIN
20731|SUTTER
20732|SUTTER CREEK
20733|SUTTLE
20734|SUTTON
20735|SUTTONS BAY
20736|SUWANEE
20737|SUWANNEE
20738|SUÁREZ
20739|SUÁREZ COMUNIDAD
20740|SVEA
20741|SWAIN
20742|SWAINSBORO
20743|SWALEDALE
20744|SWAMPSCOTT
20745|SWAN LAKE
20746|SWAN RIVER
20747|SWAN VALLEY
20748|SWANDALE
20749|SWANLAKE
20750|SWANNANOA
20751|SWANQUARTER
20752|SWANSBORO
20753|SWANSEA
20754|SWANTON
20755|SWANVILLE
20756|SWANWICK
20757|SWARTHMORE
20758|SWARTZ
20759|SWARTZ CREEK
20760|SWARTZVILLE
20761|SWATARA
20762|SWAYZEE
20763|SWEA CITY
20764|SWEARINGEN
20765|SWEATMAN
20766|SWEDE HEAVEN
20767|SWEDEBORG
20768|SWEDEBURG
20769|SWEDEN
20770|SWEDEN VALLEY
20771|SWEDESBORO
20772|SWEDESBURG
20773|SWEENY
20774|SWEET AIR
20775|SWEET BRIAR STATION
20776|SWEET GRASS
20777|SWEET HOME
20778|SWEET SPRINGS
20779|SWEET VALLEY
20780|SWEET WATER
20781|SWEETSER
20782|SWEETWATER
20783|SWENSON
20784|SWEPSONVILLE
20785|SWIFT
20786|SWIFT FALLS
20787|SWIFT TRAIL JUNCTION
20788|SWIFTON
20789|SWIFTWATER
20790|SWINK
20791|SWINOMISH VILLAGE
20792|SWISHER
20793|SWISS ALP
20794|SWISSHOME
20795|SWISSVALE
20796|SWITZ CITY
20797|SWITZER
20798|SWORDS
20799|SWORMVILLE
20800|SWOYERSVILLE
20801|SYCAMORE
20802|SYCAMORE HILLS
20803|SYCAMORE VALLEY
20804|SYDNEY
20805|SYKESTON
20806|SYKESVILLE
20807|SYLACAUGA
20808|SYLVA
20809|SYLVAN BEACH
20810|SYLVAN GROVE
20811|SYLVAN HILLS
20812|SYLVAN LAKE
20813|SYLVAN SPRINGS
20814|SYLVANIA
20815|SYLVANITE
20816|SYLVARENA
20817|SYLVESTER
20818|SYLVIA
20819|SYMCO
20820|SYMERTON
20821|SYMSONIA
20822|SYNAREP
20823|SYOSSET
20824|SYRACUSE
20825|SYRIA
20826|TABERNACLE
20827|TABERNASH
20828|TABERVILLE
20829|TABIONA
20830|TABLE GROVE
20831|TABLE ROCK
20832|TABLER
20833|TABOR
20834|TABOR CITY
20835|TACNA
20836|TACOMA
20837|TACONIC SHORES
20838|TACONITE
20839|TACONITE HARBOR
20840|TAFT
20841|TAFT HEIGHTS
20842|TAFTON
20843|TAGG FLATS
20844|TAGUS
20845|TAHAWUS
20846|TAHLEQUAH
20847|TAHOE CITY
20848|TAHOE VISTA
20849|TAHOKA
20850|TAHOLAH
20851|TAHOMA
20852|TAHUYA
20853|TAIBAN
20854|TAINTER LAKE
20855|TAJIGUAS
20856|TAJIQUE
20857|TAKILMA
20858|TAKOMA PARK
20859|TAKOTNA
20860|TALALA
20861|TALBERT
20862|TALBOTT
20863|TALBOTTON
20864|TALCO
20865|TALENT
20866|TALIHINA
20867|TALISHEEK
20868|TALKEETNA
20869|TALKING ROCK
20870|TALL TIMBER
20871|TALL TIMBERS
20872|TALLABOA
20873|TALLABOA ALTA
20874|TALLABOA ALTA COMUNIDAD
20875|TALLABOA COMUNIDAD
20876|TALLADEGA
20877|TALLADEGA SPRINGS
20878|TALLAHASSEE
20879|TALLAPOOSA
20880|TALLASSEE
20881|TALLEVAST
20882|TALLEY CAVEY
20883|TALLEYVILLE
20884|TALLMADGE
20885|TALLMAN
20886|TALLULA
20887|TALLULAH
20888|TALLULAH FALLS
20889|TALMAGE
20890|TALMO
20891|TALOGA
20892|TALOWAH
20893|TALPA
20894|TALTY
20895|TAMA
20896|TAMAHA
20897|TAMAQUA
20898|TAMARAC
20899|TAMARACK
20900|TAMAROA
20901|TAMIAMI
20902|TAMINA
20903|TAMMS
20904|TAMO
20905|TAMOLA
20906|TAMORA
20907|TAMPA
20908|TAMPICO
20909|TANACROSS
20910|TANAINA
20911|TANANA
20912|TANEYTOWN
20913|TANEYVILLE
20914|TANGELO PARK
20915|TANGENT
20916|TANGERINE
20917|TANGIER
20918|TANGIPAHOA
20919|TANGLEWILDE
20920|TANGLEWOOD
20921|TANGLEWOOD FOREST
20922|TANKERSLEY
20923|TANNEHILL
20924|TANNER
20925|TANNERSVILLE
20926|TANQUE
20927|TANQUE VERDE
20928|TANSBORO
20929|TAOPI
20930|TAOS
20931|TAOS PUEBLO
20932|TAOS SKI VALLEY
20933|TAPPAHANNOCK
20934|TAPPAN
20935|TAPPEN
20936|TAR HEEL
20937|TARA
20938|TARA HILLS
20939|TARBORO
20940|TARENTUM
20941|TARIFFVILLE
20942|TARKIO
20943|TARLTON
20944|TARNOV
20945|TARPEY VILLAGE
20946|TARPON SPRINGS
20947|TARRANT
20948|TARRANTS
20949|TARRY
20950|TARRYALL
20951|TARRYTOWN
20952|TARVER
20953|TARZAN
20954|TASCO
20955|TASCOSA
20956|TASLEY
20957|TASSO
20958|TAT MOMOLI
20959|TATAMY
20960|TATE
20961|TATE CITY
20962|TATITLEK
20963|TATUM
20964|TATUMS
20965|TAUNTON
20966|TAVARES
20967|TAVERNIER
20968|TAVISTOCK
20969|TAWAS CITY
20970|TAYCHEEDAH
20971|TAYLOR
20972|TAYLOR CREEK
20973|TAYLOR LAKE VILLAGE
20974|TAYLOR LANDING
20975|TAYLOR MILL
20976|TAYLOR SPRINGS
20977|TAYLORS
20978|TAYLORS CREEK
20979|TAYLORS FALLS
20980|TAYLORS ISLAND
20981|TAYLORSPORT
20982|TAYLORSTOWN
20983|TAYLORSTOWN STATION
20984|TAYLORSVILLE
20985|TAYLORTOWN
20986|TAYLORVILLE
20987|TAZEWELL
20988|TAZLINA
20989|TCHULA
20990|TEACHEY
20991|TEAGUE
20992|TEASDALE
20993|TEATICKET
20994|TEAYS VALLEY
20995|TECATE
20996|TECOLOTE
20997|TECOLOTITO
20998|TECOPA
20999|TECUMSEH
21000|TEDROW
21001|TEE HARBOR
21002|TEEC NOS POS
21003|TEEDS GROVE
21004|TEES TOH
21005|TEGA CAY
21006|TEGARDEN
21007|TEHACHAPI
21008|TEHAMA
21009|TEHUACANA
21010|TEIGEN
21011|TEKAMAH
21012|TEKOA
21013|TEKONSHA
21014|TELEGRAPH
21015|TELEPHONE
21016|TELFERNER
21017|TELFORD
21018|TELIDA
21019|TELL CITY
21020|TELLER
21021|TELLICO PLAINS
21022|TELLURIDE
21023|TELMA
21024|TELOCASET
21025|TELOGIA
21026|TEMECULA
21027|TEMELEC
21028|TEMPE
21029|TEMPERANCE
21030|TEMPERANCEVILLE
21031|TEMPIUTE
21032|TEMPLE
21033|TEMPLE CITY
21034|TEMPLE HILL
21035|TEMPLE HILLS
21036|TEMPLE TERRACE
21037|TEMPLETON
21038|TEMPLEVILLE
21039|TEMVIK
21040|TEN BROECK
21041|TEN MILE
21042|TEN MILE RUN
21043|TEN SLEEP
21044|TENAFLY
21045|TENAHA
21046|TENAKEE SPRINGS
21047|TENDAL
21048|TENINO
21049|TENKILLER
21050|TENMILE
21051|TENNANT
21052|TENNENT
21053|TENNESSEE
21054|TENNESSEE CITY
21055|TENNESSEE COLONY
21056|TENNESSEE RIDGE
21057|TENNEY
21058|TENNILLE
21059|TENNYSON
21060|TENSAW
21061|TENSED
21062|TENSTRIKE
21063|TEQUESTA
21064|TERERRO
21065|TERESITA
21066|TERLINGUA
21067|TERLTON
21068|TERMINOUS
21069|TERMO
21070|TERRA ALTA
21071|TERRA BELLA
21072|TERRA LINDA
21073|TERRACE HEIGHTS
21074|TERRACE PARK
21075|TERRAL
21076|TERRAMUGGUS
21077|TERRE DU LAC
21078|TERRE HAUTE
21079|TERRE HILL
21080|TERREBONNE
21081|TERRELL
21082|TERRELL HILLS
21083|TERRETON
21084|TERRIL
21085|TERRY
21086|TERRYTOWN
21087|TERRYVILLE
21088|TESCO
21089|TESCOTT
21090|TESUQUE
21091|TESUQUE PUEBLO
21092|TETERBORO
21093|TETERVILLE
21094|TETLIN
21095|TETON
21096|TETON VILLAGE
21097|TETONIA
21098|TEUTOPOLIS
21099|TEXANNA
21100|TEXARKANA
21101|TEXAS CITY
21102|TEXAS CREEK
21103|TEXASVILLE
21104|TEXHOMA
21105|TEXICO
21106|TEXLINE
21107|TEXOLA
21108|TEXON
21109|THACH
21110|THACKERVILLE
21111|THALIA
21112|THALMANN
21113|THAMA
21114|THANE
21115|THATCHER
21116|THAWVILLE
21117|THAXTON
21118|THAYER
21119|THAYER JUNCTION
21120|THAYNE
21121|THE ACREAGE
21122|THE COLONY
21123|THE CROSSINGS
21124|THE DALLES
21125|THE GLEN
21126|THE GROVE
21127|THE HAMMOCKS
21128|THE HIDEOUT
21129|THE HILLS
21130|THE LAKES
21131|THE LANDING
21132|THE MEADOWS
21133|THE PINERY
21134|THE PLAINS
21135|THE ROCK
21136|THE VILLAGE
21137|THE VILLAGE OF INDIAN HILL
21138|THE VILLAGES
21139|THE WOODLANDS
21140|THEBA
21141|THEBES
21142|THEDFORD
21143|THEILMAN
21144|THELMA
21145|THENDARA
21146|THEODORE
21147|THEODOSIA
21148|THERESA
21149|THERESSA
21150|THERIOT
21151|THERMAL
21152|THERMALITO
21153|THERMOPOLIS
21154|THIBODAUX
21155|THIEF RIVER FALLS
21156|THIELLS
21157|THIENSVILLE
21158|THIRD LAKE
21159|THISTLE
21160|THOMAS
21161|THOMASBORO
21162|THOMASTON
21163|THOMASTOWN
21164|THOMASVILLE
21165|THOMPSON
21166|THOMPSON FALLS
21167|THOMPSON PLACE
21168|THOMPSON SPRINGS
21169|THOMPSON'S STATION
21170|THOMPSONS
21171|THOMPSONTOWN
21172|THOMPSONVILLE
21173|THOMSON
21174|THONOTOSASSA
21175|THOR
21176|THOREAU
21177|THORN
21178|THORNBURG
21179|THORNDALE
21180|THORNE
21181|THORNE BAY
21182|THORNFIELD
21183|THORNHILL
21184|THORNPORT
21185|THORNTON
21186|THORNTONVILLE
21187|THORNTOWN
21188|THORNVILLE
21189|THORNWOOD
21190|THOROFARE
21191|THORP
21192|THORSBY
21193|THOUSAND ISLAND PARK
21194|THOUSAND OAKS
21195|THOUSAND PALMS
21196|THOUSANDSTICKS
21197|THRALL
21198|THREE CREEK
21199|THREE CREEKS VILLAGE
21200|THREE FORKS
21201|THREE LAKES
21202|THREE MILE BAY
21203|THREE OAKS
21204|THREE POINTS
21205|THREE RIVERS
21206|THREE ROCKS
21207|THREE SPRINGS
21208|THREE WAY
21209|THREELINKS
21210|THROCKMORTON
21211|THROOP
21212|THUNDER BUTTE
21213|THUNDER HAWK
21214|THUNDERBOLT
21215|THURMAN
21216|THURMOND
21217|THURMONT
21218|THURSTON
21219|TIAWAH
21220|TIBBIE
21221|TIBES COMUNIDAD
21222|TIBURON
21223|TIBURONES
21224|TIBURONES COMUNIDAD
21225|TICE
21226|TICHIGAN
21227|TICHNOR
21228|TICKFAW
21229|TICONDEROGA
21230|TIDEWATER
21231|TIDIOUTE
21232|TIE PLANT
21233|TIE SIDING
21234|TIERRA AMARILLA
21235|TIERRA BONITA
21236|TIERRA GRANDE
21237|TIERRA VERDE
21238|TIERRAS NUEVAS PONIENTE
21239|TIERRAS NUEVAS PONIENTE COMUNIDAD
21240|TIETON
21241|TIFF CITY
21242|TIFFANY
21243|TIFFIN
21244|TIFTON
21245|TIGARD
21246|TIGER
21247|TIGER POINT
21248|TIGERTON
21249|TIGERVILLE
21250|TIGHTWAD
21251|TIGNALL
21252|TIJERAS
21253|TIKI ISLAND
21254|TILDEN
21255|TILDENVILLE
21256|TILFORD
21257|TILGHMAN
21258|TILGHMAN ISLAND
21259|TILGHMANTON
21260|TILINE
21261|TILLAMOOK
21262|TILLAR
21263|TILLATOBA
21264|TILLEDA
21265|TILLER
21266|TILLICUM
21267|TILLMAN
21268|TILLMANS CORNER
21269|TILLSON
21270|TILTON
21271|TILTONSVILLE
21272|TIMBER
21273|TIMBER HILLS
21274|TIMBER LAKE
21275|TIMBER LAKES
21276|TIMBER PINES
21277|TIMBERCREEK CANYON
21278|TIMBERLAKE
21279|TIMBERLANE
21280|TIMBERON
21281|TIMBERVILLE
21282|TIMBERWOOD PARK
21283|TIMBLIN
21284|TIMBO
21285|TIMEWELL
21286|TIMKEN
21287|TIMMONSVILLE
21288|TIMNATH
21289|TIMONIUM
21290|TIMPAS
21291|TIMPIE
21292|TIMPSON
21293|TIN CITY
21294|TINA
21295|TINAJA
21296|TINDALL
21297|TINGLEY
21298|TINLEY PARK
21299|TINSLEY
21300|TINSMAN
21301|TINTAH
21302|TINTON FALLS
21303|TIOGA
21304|TIONESTA
21305|TIPLERSVILLE
21306|TIPP CITY
21307|TIPPECANOE
21308|TIPPETT
21309|TIPTON
21310|TIPTONVILLE
21311|TIPTOP
21312|TIRA
21313|TIRO
21314|TISCH MILLS
21315|TISHOMINGO
21316|TISKILWA
21317|TITANIC
21318|TITICUS
21319|TITLEY
21320|TITONKA
21321|TITUSVILLE
21322|TIVERTON
21323|TIVOLI
21324|TOA ALTA
21325|TOA ALTA ZONA URBANA
21326|TOA BAJA
21327|TOA BAJA ZONA URBANA
21328|TOAD HOP
21329|TOANO
21330|TOAST
21331|TOBACCOVILLE
21332|TOBIAS
21333|TOBIN
21334|TOBIQUE
21335|TOBOSO
21336|TOBYHANNA
21337|TOCA
21338|TOCCOA
21339|TOCCOPOLA
21340|TOCITO
21341|TOCO
21342|TOCSIN
21343|TODD
21344|TODD CREEK
21345|TODD MISSION
21346|TODDVILLE
21347|TOETERVILLE
21348|TOFTE
21349|TOFTREES
21350|TOFTY
21351|TOGA
21352|TOGIAK
21353|TOGO
21354|TOHATCHI
21355|TOK
21356|TOKEEN
21357|TOKELAND
21358|TOKIO
21359|TOKSOOK BAY
21360|TOLANI LAKE
21361|TOLAR
21362|TOLBERT
21363|TOLCHESTER
21364|TOLCHESTER BEACH
21365|TOLEDO
21366|TOLLESON
21367|TOLLETTE
21368|TOLLEY
21369|TOLLHOUSE
21370|TOLNA
21371|TOLONO
21372|TOLSONA
21373|TOLSTOY
21374|TOLTEC
21375|TOLU
21376|TOLUCA
21377|TOM
21378|TOM BEAN
21379|TOMAH
21380|TOMAHAWK
21381|TOMALES
21382|TOMATO
21383|TOMBALL
21384|TOMBSTONE
21385|TOME
21386|TOMKINS COVE
21387|TOMNOLEN
21388|TOMPKINSVILLE
21389|TOMS BROOK
21390|TOMS PLACE
21391|TOMS RIVER
21392|TONALEA
21393|TONASKET
21394|TONAWANDA
21395|TONET
21396|TONGANOXIE
21397|TONICA
21398|TONKA BAY
21399|TONKAWA
21400|TONOPAH
21401|TONSINA
21402|TONTITOWN
21403|TONTO BASIN
21404|TONTO VILLAGE
21405|TONTOGANY
21406|TONY
21407|TONYVILLE
21408|TOOELE
21409|TOOMSBORO
21410|TOOMSUBA
21411|TOONE
21412|TOONERVILLE
21413|TOPANGA
21414|TOPAWA
21415|TOPAZ
21416|TOPAZ LAKE
21417|TOPEKA
21418|TOPEKA JUNCTION
21419|TOPINABEE
21420|TOPOCK
21421|TOPONAS
21422|TOPPENISH
21423|TOPSAIL BEACH
21424|TOPSFIELD
21425|TOPSHAM
21426|TOPSTONE
21427|TOPTON
21428|TOQUERVILLE
21429|TORBOY
21430|TORNILLO
21431|TORO
21432|TORO CANYON
21433|TORONTO
21434|TORRANCE
21435|TORREON
21436|TORREY
21437|TORRINGTON
21438|TORTILLA FLAT
21439|TOSTON
21440|TOTOWA
21441|TOUCHET
21442|TOUGALOO
21443|TOUGHKENAMON
21444|TOUHY
21445|TOULON
21446|TOVEY
21447|TOWACO
21448|TOWAMENSING TRAILS
21449|TOWANDA
21450|TOWAOC
21451|TOWER
21452|TOWER CITY
21453|TOWER HILL
21454|TOWER LAKE
21455|TOWERS CORNERS
21456|TOWN 'N' COUNTRY
21457|TOWN AND COUNTRY
21458|TOWN CREEK
21459|TOWN LINE
21460|TOWN OF PINES
21461|TOWN WEST
21462|TOWNER
21463|TOWNS
21464|TOWNSEND
21465|TOWNSVILLE
21466|TOWNVILLE
21467|TOWSON
21468|TOXEY
21469|TOYAH
21470|TOYAHVALE
21471|TOYEI
21472|TRABUCO CANYON
21473|TRABUCO HIGHLANDS
21474|TRACY
21475|TRACY CITY
21476|TRACYS LANDING
21477|TRACYTON
21478|TRADESVILLE
21479|TRADEWINDS
21480|TRAER
21481|TRAFALGAR
21482|TRAFFORD
21483|TRAIL
21484|TRAIL CITY
21485|TRAIL CREEK
21486|TRAINER
21487|TRAMMEL
21488|TRAMMELS
21489|TRAMWAY
21490|TRANQUILLITY
21491|TRANSYLVANIA
21492|TRAPPE
21493|TRAPPER CREEK
21494|TRASKWOOD
21495|TRAVELERS REST
21496|TRAVER
21497|TRAVERSE
21498|TRAVERSE CITY
21499|TRAVILAH
21500|TRAWICK
21501|TREASURE ISLAND
21502|TREASURE LAKE
21503|TREBLOC
21504|TREES MILLS
21505|TREGO
21506|TREMENTINA
21507|TREMONT
21508|TREMONT CITY
21509|TREMONTON
21510|TREMPEALEAU
21511|TRENARY
21512|TRENT
21513|TRENT WOODS
21514|TRENTON
21515|TRENTWOOD
21516|TRES PIEDRAS
21517|TRES PINOS
21518|TRESCKOW
21519|TREVESKYN
21520|TREVLAC
21521|TREVORTON
21522|TREVOSE
21523|TREXLERTOWN
21524|TREYNOR
21525|TREZEVANT
21526|TRI-CITY
21527|TRI-LAKES
21528|TRIADELPHIA
21529|TRIANA
21530|TRIBBEY
21531|TRIBES HILL
21532|TRIBUNE
21533|TRIDENT
21534|TRILBY
21535|TRIMBLE
21536|TRIMMER
21537|TRIMONT
21538|TRINCHERA
21539|TRINIDAD
21540|TRINITY
21541|TRINITY CENTER
21542|TRINITY VILLAGE
21543|TRINWAY
21544|TRION
21545|TRIPLET
21546|TRIPLETT
21547|TRIPOLI
21548|TRIPP
21549|TRIUMPH
21550|TROMMALD
21551|TRONA
21552|TROOPER
21553|TROPHY CLUB
21554|TROPIC
21555|TROSKY
21556|TROTTERS
21557|TROTWOOD
21558|TROUP
21559|TROUSDALE
21560|TROUT
21561|TROUT CREEK
21562|TROUT DALE
21563|TROUT LAKE
21564|TROUT RUN
21565|TROUT VALLEY
21566|TROUTDALE
21567|TROUTMAN
21568|TROUTVILLE
21569|TROWBRIDGE
21570|TROWBRIDGE PARK
21571|TROXELVILLE
21572|TROY
21573|TROY GROVE
21574|TROY HILLS
21575|TRUCHAS
21576|TRUCKEE
21577|TRUCKSVILLE
21578|TRUESDALE
21579|TRUFANT
21580|TRUJILLO
21581|TRUJILLO ALTO
21582|TRUJILLO ALTO ZONA URBANA
21583|TRUMAN
21584|TRUMANN
21585|TRUMANSBURG
21586|TRUMBAUERSVILLE
21587|TRUMBULL
21588|TRURO
21589|TRUSCOTT
21590|TRUSSVILLE
21591|TRUTH OR CONSEQUENCES
21592|TRUXALL
21593|TRUXTON
21594|TRYON
21595|TSCHETTER COLONY
21596|TSE BONITO
21597|TSELAKAI DEZZA
21598|TUALATIN
21599|TUBA CITY
21600|TUBAC
21601|TUCKAHOE
21602|TUCKER
21603|TUCKERMAN
21604|TUCKERS CROSSING
21605|TUCKERTON
21606|TUCSON
21607|TUCSON ESTATES
21608|TUCUMCARI
21609|TUKWILA
21610|TULA
21611|TULALIP
21612|TULARE
21613|TULAROSA
21614|TULELAKE
21615|TULETA
21616|TULIA
21617|TULIP
21618|TULL
21619|TULLAHASSEE
21620|TULLAHOMA
21621|TULLOS
21622|TULLY
21623|TULLYTOWN
21624|TULSA
21625|TULSITA
21626|TULUKSAK
21627|TUMACACORI
21628|TUMALO
21629|TUMBLING SHOALS
21630|TUMWATER
21631|TUNAS
21632|TUNDRA
21633|TUNICA
21634|TUNICA RESORTS
21635|TUNIS
21636|TUNIS MILLS
21637|TUNKHANNOCK
21638|TUNNEL CITY
21639|TUNNEL HILL
21640|TUNNEL SPRINGS
21641|TUNNELHILL
21642|TUNNELTON
21643|TUNTUTULIAK
21644|TUNUNAK
21645|TUOLUMNE
21646|TUOLUMNE CITY
21647|TUPELO
21648|TUPMAN
21649|TUPPER LAKE
21650|TUPPERS PLAINS
21651|TURAH
21652|TURBEVILLE
21653|TURBOTVILLE
21654|TURIN
21655|TURKEY
21656|TURKEY CREEK
21657|TURKEY CREEK MEADOWS
21658|TURLEY
21659|TURLOCK
21660|TURNBULL
21661|TURNER
21662|TURNER CORNER
21663|TURNERS FALLS
21664|TURNERSVILLE
21665|TURNERVILLE
21666|TURNEY
21667|TURON
21668|TURPIN
21669|TURPIN HILLS
21670|TURRELL
21671|TURTLE CREEK
21672|TURTLE LAKE
21673|TURTLE RIVER
21674|TURTON
21675|TUSAYAN
21676|TUSCALOOSA
21677|TUSCARAWAS
21678|TUSCARORA
21679|TUSCOLA
21680|TUSCULUM
21681|TUSCUMBIA
21682|TUSHKA
21683|TUSKAHOMA
21684|TUSKEGEE
21685|TUSTIN
21686|TUTHILL
21687|TUTTLE
21688|TUTTLETOWN
21689|TUTU
21690|TUTUILLA
21691|TUTWILER
21692|TUXEDO
21693|TUXEDO PARK
21694|TWAIN
21695|TWAIN HARTE
21696|TWENTYNINE PALMS
21697|TWICHELL
21698|TWILIGHT
21699|TWIN
21700|TWIN BRIDGES
21701|TWIN BROOKS
21702|TWIN CITY
21703|TWIN FALLS
21704|TWIN GROVE
21705|TWIN GROVES
21706|TWIN HILLS
21707|TWIN LAKE
21708|TWIN LAKES
21709|TWIN LAKES VILLAGE
21710|TWIN MOUNTAIN
21711|TWIN OAKS
21712|TWIN PEAKS
21713|TWIN RIVERS
21714|TWIN VALLEY
21715|TWINING
21716|TWINSBURG
21717|TWINSBURG HEIGHTS
21718|TWISP
21719|TWITTY
21720|TWO BUTTES
21721|TWO GUNS
21722|TWO HARBORS
21723|TWO INLETS
21724|TWO RIVERS
21725|TWO STRIKE
21726|TWODOT
21727|TY TY
21728|TYASKIN
21729|TYBEE ISLAND
21730|TYE
21731|TYGH VALLEY
21732|TYHEE
21733|TYLER
21734|TYLERSBURG
21735|TYLERSVILLE
21736|TYLERTOWN
21737|TYNAN
21738|TYNDALL
21739|TYNER
21740|TYNGSBORO
21741|TYONEK
21742|TYRO
21743|TYRONE
21744|TYRONZA
21745|TYSONS
21746|UALAPUʻE
21747|UBLY
21748|UCOLO
21749|UCON
21750|UDALL
21751|UDELL
21752|UEHLING
21753|UGASHIK
21754|UHLAND
21755|UHRICHSVILLE
21756|UINTAH
21757|UKIAH
21758|ULEN
21759|ULLIN
21760|ULM
21761|ULMER
21762|ULSTER
21763|ULUPALAKUA
21764|ULYSSES
21765|UMAPINE
21766|UMATILLA
21767|UMBARGER
21768|UMBER VIEW HEIGHTS
21769|UMIAT
21770|UMKUMIUTE
21771|UMPIRE
21772|UMPQUA
21773|UNADILLA
21774|UNALAKLEET
21775|UNALASKA
21776|UNCAS
21777|UNCASVILLE
21778|UNCERTAIN
21779|UNDERWOOD
21780|UNGA
21781|UNICOI
21782|UNIFIED GOVERNMENT OF GREELEY COUNTY (BALANCE)
21783|UNION
21784|UNION BEACH
21785|UNION BRIDGE
21786|UNION CENTER
21787|UNION CHURCH
21788|UNION CITY
21789|UNION CREEK
21790|UNION DALE
21791|UNION DEPOSIT
21792|UNION FURNACE
21793|UNION GAP
21794|UNION GROVE
21795|UNION HALL
21796|UNION HILL
21797|UNION LAKE
21798|UNION LEVEL
21799|UNION PARK
21800|UNION POINT
21801|UNION SPRINGS
21802|UNION STAR
21803|UNION VALLEY
21804|UNION VILLAGE
21805|UNIONDALE
21806|UNIONTOWN
21807|UNIONVALE
21808|UNIONVILLE
21809|UNIONVILLE CENTER
21810|UNIOPOLIS
21811|UNITED
21812|UNITY
21813|UNITY VILLAGE
21814|UNITYVILLE
21815|UNIVERSAL
21816|UNIVERSAL CITY
21817|UNIVERSITY
21818|UNIVERSITY CENTER
21819|UNIVERSITY CITY
21820|UNIVERSITY GARDENS
21821|UNIVERSITY HEIGHTS
21822|UNIVERSITY PARK
21823|UNIVERSITY PLACE
21824|UPALCO
21825|UPATOI
21826|UPHAM
21827|UPLAND
21828|UPLANDS PARK
21829|UPPER ARLINGTON
21830|UPPER BROOKVILLE
21831|UPPER CROSSROADS
21832|UPPER DARBY
21833|UPPER EXETER
21834|UPPER FRUITLAND
21835|UPPER GRAND LAGOON
21836|UPPER LAKE
21837|UPPER MARLBORO
21838|UPPER MILL
21839|UPPER MONTCLAIR
21840|UPPER NYACK
21841|UPPER PRESTON
21842|UPPER SADDLE RIVER
21843|UPPER SAINT CLAIR
21844|UPPER SANDUSKY
21845|UPPER TRACT
21846|UPSALA
21847|UPSON
21848|UPTON
21849|URANIA
21850|URAVAN
21851|URBAN
21852|URBANA
21853|URBANCREST
21854|URBANDALE
21855|URBANETTE
21856|URBANK
21857|URBANNA
21858|URIAH
21859|URICH
21860|URIE
21861|URSA
21862|URSINA
21863|URSINE
21864|USHER
21865|USK
21866|UTE
21867|UTE PARK
21868|UTICA
21869|UTLEYVILLE
21870|UTOPIA
21871|UTQIAĠVIK
21872|UTTING
21873|UTUADO
21874|UTUADO ZONA URBANA
21875|UVALDA
21876|UVALDE
21877|UVALDE ESTATES
21878|UYAK
21879|VACAVILLE
21880|VACHERIE
21881|VADER
21882|VADITO
21883|VADNAIS HEIGHTS
21884|VADO
21885|VAIDEN
21886|VAIL
21887|VAILS GATE
21888|VAIR
21889|VAIVA VO
21890|VAL VERDA
21891|VAL VERDE
21892|VAL VERDE PARK
21893|VALATIE
21894|VALDERS
21895|VALDESE
21896|VALDEZ
21897|VALDOSTA
21898|VALE
21899|VALE SUMMIT
21900|VALEENE
21901|VALENCIA
21902|VALENTINE
21903|VALERA
21904|VALERIA
21905|VALHALLA
21906|VALIER
21907|VALINDA
21908|VALKARIA
21909|VALLE
21910|VALLE CRUCIS
21911|VALLE VISTA
21912|VALLECITO
21913|VALLEJO
21914|VALLES MINES
21915|VALLEY
21916|VALLEY ACRES
21917|VALLEY BEND
21918|VALLEY BROOK
21919|VALLEY CENTER
21920|VALLEY CITY
21921|VALLEY COTTAGE
21922|VALLEY CREEK
21923|VALLEY FALLS
21924|VALLEY FORD
21925|VALLEY FORGE
21926|VALLEY GRANDE
21927|VALLEY GREEN
21928|VALLEY GROVE
21929|VALLEY HEAD
21930|VALLEY HI
21931|VALLEY HILL
21932|VALLEY HOME
21933|VALLEY MILLS
21934|VALLEY PARK
21935|VALLEY RANCH
21936|VALLEY SPRING
21937|VALLEY SPRINGS
21938|VALLEY STREAM
21939|VALLEY VIEW
21940|VALLEY VIEW PARK
21941|VALLEY WELLS
21942|VALLEY-HI
21943|VALLIANT
21944|VALLONIA
21945|VALMEYER
21946|VALMONT
21947|VALMORA
21948|VALMY
21949|VALPARAISO
21950|VALRICO
21951|VALTON
21952|VALUE
21953|VAMO
21954|VAN
21955|VAN ALSTYNE
21956|VAN BIBBER LAKE
21957|VAN BUREN
21958|VAN BUSKIRK
21959|VAN CORTLANDTVILLE
21960|VAN DYNE
21961|VAN ETTEN
21962|VAN HISEVILLE
21963|VAN HORN
21964|VAN HORNE
21965|VAN LEAR
21966|VAN METER
21967|VAN METRE
21968|VAN TASSELL
21969|VAN VLECK
21970|VAN VOORHIS
21971|VAN WERT
21972|VAN WYCK
21973|VAN ZANDT
21974|VANANDA
21975|VANCE
21976|VANCEBORO
21977|VANCEBURG
21978|VANCLEAVE
21979|VANCLEVE
21980|VANCOURT
21981|VANCOUVER
21982|VANDALIA
21983|VANDEMERE
21984|VANDENBERG VILLAGE
21985|VANDER
21986|VANDERBILT
21987|VANDERCOOK LAKE
21988|VANDERGRIFT
21989|VANDERPOOL
21990|VANDERVOORT
21991|VANDIVER
21992|VANDLING
21993|VANDUSER
21994|VANDYKE
21995|VANLEER
21996|VANLUE
21997|VANN CROSSROADS
21998|VANNDALE
21999|VANOSS
22000|VANPORT
22001|VANSANT
22002|VANTAGE
22003|VANZANT
22004|VARDAMAN
22005|VARINA
22006|VARNA
22007|VARNADO
22008|VARNAMTOWN
22009|VARNELL
22010|VARNER
22011|VARNVILLE
22012|VASHON
22013|VASHON HEIGHTS
22014|VASS
22015|VASSAR
22016|VAUCLUSE
22017|VAUDREUIL
22018|VAUGHAN
22019|VAUGHN
22020|VAUGHNS MILL
22021|VAUGHNSVILLE
22022|VAYAS
22023|VAYAS COMUNIDAD
22024|VEAL
22025|VEBLEN
22026|VEEDERSBURG
22027|VEGA
22028|VEGA ALTA
22029|VEGA ALTA ZONA URBANA
22030|VEGA BAJA
22031|VEGA BAJA ZONA URBANA
22032|VEGUITA
22033|VELARDE
22034|VELDA VILLAGE
22035|VELDA VILLAGE HILLS
22036|VELMA
22037|VELVA
22038|VENANGO
22039|VENEDOCIA
22040|VENEDY
22041|VENERSBORG
22042|VENETA
22043|VENETIAN VILLAGE
22044|VENETIE
22045|VENICE
22046|VENICE GARDENS
22047|VENTANA
22048|VENTNOR CITY
22049|VENTRESS
22050|VENTURA
22051|VENTURIA
22052|VENUS
22053|VERA
22054|VERA CRUZ
22055|VERADALE
22056|VERBENA
22057|VERDA
22058|VERDE VILLAGE
22059|VERDEL
22060|VERDEMONT
22061|VERDEN
22062|VERDERY
22063|VERDI
22064|VERDIGRE
22065|VERDIGRIS
22066|VERDON
22067|VERDUNVILLE
22068|VERGAS
22069|VERGENNES
22070|VERHALEN
22071|VERLOT
22072|VERMILION
22073|VERMILLION
22074|VERMONT
22075|VERMONT HEIGHTS
22076|VERMONTVILLE
22077|VERNA
22078|VERNAL
22079|VERNDALE
22080|VERNE
22081|VERNON
22082|VERNON CENTER
22083|VERNON HILLS
22084|VERNON VALLEY
22085|VERNONBURG
22086|VERNONIA
22087|VERO BEACH
22088|VERONA
22089|VERPLANCK
22090|VERRET
22091|VERSAILLES
22092|VESPER
22093|VESTA
22094|VESTABURG
22095|VESTAL CENTER
22096|VESTAVIA HILLS
22097|VESUVIUS
22098|VETAL
22099|VETERAN
22100|VEVAY
22101|VEYO
22102|VIAN
22103|VIBBARD
22104|VIBORAS
22105|VIBORG
22106|VIBURNUM
22107|VICCO
22108|VICHY
22109|VICI
22110|VICK
22111|VICKERY
22112|VICKSBURG
22113|VICTOR
22114|VICTORIA
22115|VICTORVILLE
22116|VICTORY GARDENS
22117|VICTORY LAKES
22118|VICTORY MILLS
22119|VIDA
22120|VIDAL
22121|VIDAL JUNCTION
22122|VIDALIA
22123|VIDAURRI
22124|VIDETTE
22125|VIDOR
22126|VIDRINE
22127|VIENNA
22128|VIENNA BEND
22129|VIEQUES
22130|VIEQUES COMUNIDAD
22131|VIEQUES ZONA URBANA
22132|VIEW PARK
22133|VIEWFIELD
22134|VIGIL
22135|VIGO PARK
22136|VIGUS
22137|VIKING
22138|VILANO BEACH
22139|VILAS
22140|VILLA
22141|VILLA DEL SOL
22142|VILLA GROVE
22143|VILLA HEIGHTS
22144|VILLA HILLS
22145|VILLA PANCHO
22146|VILLA PARK
22147|VILLA RICA
22148|VILLA RIDGE
22149|VILLA VERDE
22150|VILLAGE GREEN
22151|VILLAGE MILLS
22152|VILLAGE OF THE BRANCH
22153|VILLAGE SAINT GEORGE
22154|VILLAGE SHIRES
22155|VILLAGE SPRINGS
22156|VILLALBA
22157|VILLALBA ZONA URBANA
22158|VILLANO BEACH
22159|VILLANOVA
22160|VILLANUEVA
22161|VILLARD
22162|VILLAS
22163|VILLE PLATTE
22164|VILLEGREEN
22165|VILLISCA
22166|VILONIA
22167|VIMY RIDGE
22168|VINA
22169|VINCENNES
22170|VINCENT
22171|VINCENTOWN
22172|VINCO
22173|VINE GROVE
22174|VINE HILL
22175|VINEGAR BEND
22176|VINELAND
22177|VINEYARD
22178|VINEYARD HAVEN
22179|VINEYARDS
22180|VINING
22181|VININGS
22182|VINITA
22183|VINITA PARK
22184|VINITA TERRACE
22185|VINLAND
22186|VINSON
22187|VINTON
22188|VINTONDALE
22189|VIOLA
22190|VIOLET
22191|VIOLET HILL
22192|VIPER
22193|VIRDEN
22194|VIRGELLE
22195|VIRGIE
22196|VIRGIL
22197|VIRGILINA
22198|VIRGIN
22199|VIRGINIA
22200|VIRGINIA BEACH
22201|VIRGINIA CITY
22202|VIRGINIA GARDENS
22203|VIRGINVILLE
22204|VIROQUA
22205|VISALIA
22206|VISTA
22207|VISTA CENTER
22208|VISTA SANTA ROSA
22209|VISTA WEST
22210|VIVIAN
22211|VOCA
22212|VOLANT
22213|VOLBORG
22214|VOLCANO
22215|VOLENS
22216|VOLENTE
22217|VOLGA
22218|VOLIN
22219|VOLLAND
22220|VOLLMAR
22221|VOLO
22222|VOLT
22223|VOLTA
22224|VOLTAIRE
22225|VON ORMY
22226|VONA
22227|VONORE
22228|VOORHEES
22229|VOORHEESVILLE
22230|VOORHIES
22231|VORTEX
22232|VOSS
22233|VOSSBURG
22234|VOTAW
22235|VOWINCKEL
22236|VREDENBURGH
22237|VULCAN
22238|VYA
22239|VÁZQUEZ
22240|VÁZQUEZ COMUNIDAD
22241|WABASH
22242|WABASHA
22243|WABASSO
22244|WABASSO BEACH
22245|WABAUNSEE
22246|WABBASEKA
22247|WABENO
22248|WABUSKA
22249|WACCABUC
22250|WACHAPREAGUE
22251|WACISSA
22252|WACO
22253|WACONIA
22254|WACOUSTA
22255|WACOUTA
22256|WADDINGTON
22257|WADDY
22258|WADE
22259|WADE HAMPTON
22260|WADENA
22261|WADESBORO
22262|WADESVILLE
22263|WADING RIVER
22264|WADLEY
22265|WADSWORTH
22266|WAELDER
22267|WAGARVILLE
22268|WAGENER
22269|WAGGAMAN
22270|WAGGONER
22271|WAGNER
22272|WAGON MOUND
22273|WAGONER
22274|WAGONTIRE
22275|WAGRAM
22276|WAGSTAFF
22277|WAH KEENEY PARK
22278|WAHAK HOTRONTK
22279|WAHIAWĀ
22280|WAHKON
22281|WAHNETA
22282|WAHOO
22283|WAHPETON
22284|WAHSATCH
22285|WAIAKOA
22286|WAIALUA
22287|WAIEHU
22288|WAIHEʻE
22289|WAIKAPŪ
22290|WAIKOLOA VILLAGE
22291|WAIKĀNE
22292|WAILEA
22293|WAILUA
22294|WAILUA HOMESTEADS
22295|WAILUKU
22296|WAIMALU
22297|WAIMEA
22298|WAIMĀNALO
22299|WAIMĀNALO BEACH
22300|WAINAKU
22301|WAINIHA
22302|WAINSCOTT
22303|WAINWRIGHT
22304|WAIPAHU
22305|WAIPIʻO
22306|WAIPIʻO ACRES
22307|WAITE HILL
22308|WAITE PARK
22309|WAITEVILLE
22310|WAITSBURG
22311|WAITSFIELD
22312|WAIʻANAE
22313|WAIʻŌHINU
22314|WAKA
22315|WAKARUSA
22316|WAKE FOREST
22317|WAKE VILLAGE
22318|WAKEENEY
22319|WAKEFIELD
22320|WAKEMAN
22321|WAKENDA
22322|WAKITA
22323|WAKONDA
22324|WAKPALA
22325|WAKULLA
22326|WAKULLA BEACH
22327|WALAPAI
22328|WALBRIDGE
22329|WALCOTT
22330|WALDEN
22331|WALDENBURG
22332|WALDO
22333|WALDOBORO
22334|WALDORF
22335|WALDPORT
22336|WALDRON
22337|WALDWICK
22338|WALES
22339|WALESKA
22340|WALFORD
22341|WALHALLA
22342|WALKER LAKE
22343|WALKER MILL
22344|WALKER VALLEY
22345|WALKERS MILL
22346|WALKERSVILLE
22347|WALKERTON
22348|WALKERTOWN
22349|WALKERVILLE
22350|WALL LAKE
22351|WALLA WALLA
22352|WALLACE
22353|WALLACE RIDGE
22354|WALLACETON
22355|WALLAND
22356|WALLBURG
22357|WALLED LAKE
22358|WALLENPAUPACK LAKE ESTATES
22359|WALLER
22360|WALLERVILLE
22361|WALLINGFORD
22362|WALLINGTON
22363|WALLINS CREEK
22364|WALLIS
22365|WALLKILL
22366|WALLOON LAKE
22367|WALLOWA
22368|WALLSBORO
22369|WALLSBURG
22370|WALLSTREET
22371|WALLULA
22372|WALNUT
22373|WALNUT BOTTOM
22374|WALNUT COVE
22375|WALNUT CREEK
22376|WALNUT GROVE
22377|WALNUT HEIGHTS
22378|WALNUT HILL
22379|WALNUT PARK
22380|WALNUT RIDGE
22381|WALNUT SHADE
22382|WALNUT SPRINGS
22383|WALNUTPORT
22384|WALNUTTOWN
22385|WALPOLE
22386|WALSENBURG
22387|WALSH
22388|WALSHVILLE
22389|WALSTONBURG
22390|WALTERBORO
22391|WALTERHILL
22392|WALTERS
22393|WALTERSVILLE
22394|WALTERVILLE
22395|WALTHALL
22396|WALTHAM
22397|WALTHILL
22398|WALTHOURVILLE
22399|WALTMAN
22400|WALTON
22401|WALTON HILLS
22402|WALTON PARK
22403|WALTONVILLE
22404|WALTREAK
22405|WALUM
22406|WALWORTH
22407|WAMAC
22408|WAMEGO
22409|WAMESIT
22410|WAMIC
22411|WAMPSVILLE
22412|WAMPUM
22413|WAMSUTTER
22414|WANAKAH
22415|WANAMASSA
22416|WANAMIE
22417|WANAMINGO
22418|WANAQUE
22419|WANATAH
22420|WANBLEE
22421|WANCHESE
22422|WANDA
22423|WANDEROOS
22424|WANDO
22425|WANETTE
22426|WANILLA
22427|WANN
22428|WANNASKA
22429|WANNEE
22430|WANSHIP
22431|WANTAGH
22432|WAPAKONETA
22433|WAPANUCKA
22434|WAPATO
22435|WAPELLA
22436|WAPELLO
22437|WAPINITIA
22438|WAPITI
22439|WAPLES
22440|WAPPINGERS FALLS
22441|WAR
22442|WAR EAGLE
22443|WARBA
22444|WARD COVE
22445|WARD RIDGE
22446|WARD SPRINGS
22447|WARDA
22448|WARDELL
22449|WARDEN
22450|WARDENSVILLE
22451|WARDNER
22452|WARDSVILLE
22453|WARDVILLE
22454|WARE
22455|WARE PLACE
22456|WARE SHOALS
22457|WAREHAM CENTER
22458|WARESBORO
22459|WARETOWN
22460|WARFIELD
22461|WARING
22462|WARM BEACH
22463|WARM MINERAL SPRINGS
22464|WARM RIVER
22465|WARM SPRINGS
22466|WARMAN
22467|WARMINSTER
22468|WARMINSTER HEIGHTS
22469|WARNER
22470|WARNER ROBINS
22471|WARNER SPRINGS
22472|WARNERTON
22473|WARR ACRES
22474|WARREN
22475|WARREN CITY
22476|WARREN PARK
22477|WARRENDALE
22478|WARRENS
22479|WARRENS CORNERS
22480|WARRENSBURG
22481|WARRENSVILLE
22482|WARRENSVILLE HEIGHTS
22483|WARRENTON
22484|WARRENVILLE
22485|WARRINGTON
22486|WARRIOR
22487|WARRIOR RUN
22488|WARRIORS MARK
22489|WARROAD
22490|WARSAW
22491|WARSON WOODS
22492|WARTBURG
22493|WARTHEN
22494|WARTRACE
22495|WARWICK
22496|WASCO
22497|WASECA
22498|WASHAM
22499|WASHBURN
22500|WASHINGTON
22501|WASHINGTON BORO
22502|WASHINGTON COURT HOUSE
22503|WASHINGTON GROVE
22504|WASHINGTON HEIGHTS
22505|WASHINGTON MILLS
22506|WASHINGTON PARK
22507|WASHINGTON TERRACE
22508|WASHINGTONVILLE
22509|WASHOE
22510|WASHOE CITY
22511|WASHOUGAL
22512|WASHTA
22513|WASHTUCNA
22514|WASILLA
22515|WASKISH
22516|WASKOM
22517|WASOLA
22518|WASSON
22519|WASTA
22520|WASTELLA
22521|WATAGA
22522|WATAUGA
22523|WATCH HILL
22524|WATCHTOWER
22525|WATCHUNG
22526|WATER MILL
22527|WATER VALLEY
22528|WATERBURY
22529|WATEREE
22530|WATERFALL
22531|WATERFLOW
22532|WATERFORD
22533|WATERFORD WORKS
22534|WATERLOO
22535|WATERMAN
22536|WATERPROOF
22537|WATERSMEET
22538|WATERTOWN
22539|WATERVIEW
22540|WATERVILLE
22541|WATERVLIET
22542|WATFORD CITY
22543|WATHA
22544|WATHENA
22545|WATKINS
22546|WATKINS GLEN
22547|WATKINSVILLE
22548|WATONGA
22549|WATOVA
22550|WATROUS
22551|WATSEKA
22552|WATSON
22553|WATSONTOWN
22554|WATSONVILLE
22555|WATTENBERG
22556|WATTERS
22557|WATTERSON PARK
22558|WATTIS
22559|WATTS
22560|WATTSBURG
22561|WATTSVILLE
22562|WAUBAY
22563|WAUBEKA
22564|WAUBUN
22565|WAUCHULA
22566|WAUCOMA
22567|WAUCONDA
22568|WAUCOUSTA
22569|WAUHILLAU
22570|WAUKAU
22571|WAUKEE
22572|WAUKEENAH
22573|WAUKEGAN
22574|WAUKENA
22575|WAUKESHA
22576|WAUKOMIS
22577|WAUKON
22578|WAUMANDEE
22579|WAUNA
22580|WAUNAKEE
22581|WAUNETA
22582|WAUPACA
22583|WAUPUN
22584|WAUREGAN
22585|WAURIKA
22586|WAUSA
22587|WAUSAU
22588|WAUSAUKEE
22589|WAUSEON
22590|WAUTAUGA BEACH
22591|WAUTOMA
22592|WAUWATOSA
22593|WAUZEKA
22594|WAVELAND
22595|WAVERLY
22596|WAVERLY HALL
22597|WAVES
22598|WAWINA
22599|WAWONA
22600|WAXAHACHIE
22601|WAXHAW
22602|WAYAN
22603|WAYCROSS
22604|WAYLAND
22605|WAYMART
22606|WAYNE
22607|WAYNE CITY
22608|WAYNE HEIGHTS
22609|WAYNE LAKES PARK
22610|WAYNESBORO
22611|WAYNESBURG
22612|WAYNESFIELD
22613|WAYNESVILLE
22614|WAYNETOWN
22615|WAYNOKA
22616|WAYSIDE
22617|WAYZATA
22618|WEATHERBY
22619|WEATHERBY LAKE
22620|WEATHERFORD
22621|WEATHERLY
22622|WEATHERS
22623|WEATHERSBY
22624|WEATOGUE
22625|WEAUBLEAU
22626|WEAVER
22627|WEAVERVILLE
22628|WEBB
22629|WEBB CITY
22630|WEBBER
22631|WEBBERS FALLS
22632|WEBBERVILLE
22633|WEBBVILLE
22634|WEBER
22635|WEBER CITY
22636|WEBSTER
22637|WEBSTER CITY
22638|WEBSTER GROVES
22639|WEBSTER SPRINGS
22640|WEBSTERS CORNERS
22641|WEBSTERS CROSSING
22642|WEBSTERVILLE
22643|WECHES
22644|WEDDINGTON
22645|WEDGEFIELD
22646|WEDGES CORNER
22647|WEDOWEE
22648|WEDRON
22649|WEED
22650|WEED HEIGHTS
22651|WEEDONVILLE
22652|WEEDPATCH
22653|WEEDSPORT
22654|WEEDVILLE
22655|WEEHAWKEN
22656|WEEKAPAUG
22657|WEEKI WACHEE
22658|WEEKI WACHEE GARDENS
22659|WEEKSVILLE
22660|WEEPING WATER
22661|WEESATCHE
22662|WEGDAHL
22663|WEIDMAN
22664|WEIGELSTOWN
22665|WEIMAR
22666|WEINER
22667|WEINERT
22668|WEINGARTEN
22669|WEIPPE
22670|WEIR
22671|WEIRSDALE
22672|WEIRTON
22673|WEISER
22674|WEISSERT
22675|WEISSPORT
22676|WEKIWA SPRINGS
22677|WELAKA
22678|WELBY
22679|WELCH
22680|WELDA
22681|WELDON
22682|WELDON SPRING
22683|WELDON SPRING HEIGHTS
22684|WELDONA
22685|WELEETKA
22686|WELLBORN
22687|WELLERSBURG
22688|WELLESLEY
22689|WELLFLEET
22690|WELLFORD
22691|WELLING
22692|WELLINGTON
22693|WELLMAN
22694|WELLPINIT
22695|WELLS
22696|WELLS BRANCH
22697|WELLS RIVER
22698|WELLSBORO
22699|WELLSBURG
22700|WELLSFORD
22701|WELLSTON
22702|WELLSVILLE
22703|WELLTON
22704|WELOKĀ
22705|WELSH
22706|WELSHFIELD
22707|WELTON
22708|WELTY
22709|WENASOGA
22710|WENATCHEE
22711|WENDEL
22712|WENDELL
22713|WENDELVILLE
22714|WENDEN
22715|WENDOVER
22716|WENDTE
22717|WENONA
22718|WENONAH
22719|WENTWORTH
22720|WENTZVILLE
22721|WEOGUFKA
22722|WEONA
22723|WEOTT
22724|WERLEY
22725|WERNERSVILLE
22726|WESCOSVILLE
22727|WESKAN
22728|WESLACO
22729|WESLEY
22730|WESLEY CHAPEL
22731|WESLEY HILLS
22732|WESLEYVILLE
22733|WESSINGTON
22734|WESSINGTON SPRINGS
22735|WESSON
22736|WEST
22737|WEST ACTON
22738|WEST ALEXANDER
22739|WEST ALEXANDRIA
22740|WEST ALLIS
22741|WEST ALTO BONITO COLONIA
22742|WEST ALTON
22743|WEST AMANA
22744|WEST ATHENS
22745|WEST BABYLON
22746|WEST BADEN SPRINGS
22747|WEST BARABOO
22748|WEST BARNSTABLE
22749|WEST BAY
22750|WEST BAY SHORE
22751|WEST BELMAR
22752|WEST BEND
22753|WEST BERLIN
22754|WEST BISHOP
22755|WEST BLOCTON
22756|WEST BLOOMFIELD
22757|WEST BOUNTIFUL
22758|WEST BOXFORD
22759|WEST BRADENTON
22760|WEST BRANCH
22761|WEST BRATTLEBORO
22762|WEST BRISTOL
22763|WEST BROOKFIELD
22764|WEST BROOKLYN
22765|WEST BROWNSVILLE
22766|WEST BUECHEL
22767|WEST BURKE
22768|WEST BURLINGTON
22769|WEST CANTON
22770|WEST CAPE MAY
22771|WEST CARROLLTON
22772|WEST CARSON
22773|WEST CARTHAGE
22774|WEST CHATHAM
22775|WEST CHAZY
22776|WEST CHESTER
22777|WEST CHICAGO
22778|WEST CITY
22779|WEST COLLEGE CORNER
22780|WEST COLUMBIA
22781|WEST CONCORD
22782|WEST CONSHOHOCKEN
22783|WEST COVINA
22784|WEST CREEK
22785|WEST CROSSETT
22786|WEST DECATUR
22787|WEST DELAND
22788|WEST DENNIS
22789|WEST DENTON
22790|WEST DEPTFORD
22791|WEST DES MOINES
22792|WEST DOVER
22793|WEST DUNDEE
22794|WEST EASTON
22795|WEST ELIZABETH
22796|WEST ELKTON
22797|WEST ELMIRA
22798|WEST END
22799|WEST FAIRVIEW
22800|WEST FALLS
22801|WEST FALLS CHURCH
22802|WEST FALMOUTH
22803|WEST FARGO
22804|WEST FARMINGTON
22805|WEST FORK
22806|WEST FORKS
22807|WEST FRANKFORT
22808|WEST FREEHOLD
22809|WEST FROSTPROOF
22810|WEST GILGO BEACH
22811|WEST GLACIER
22812|WEST GLENDIVE
22813|WEST GLENS FALLS
22814|WEST GREEN
22815|WEST GROVE
22816|WEST HAMBURG
22817|WEST HAMLIN
22818|WEST HAMPTON DUNES
22819|WEST HANOVER
22820|WEST HARRISON
22821|WEST HARTFORD
22822|WEST HATTIESBURG
22823|WEST HAVEN
22824|WEST HAVERSTRAW
22825|WEST HAVRE
22826|WEST HAZLETON
22827|WEST HELENA
22828|WEST HEMPSTEAD
22829|WEST HICKORY
22830|WEST HILL
22831|WEST HILLS
22832|WEST HOLLYWOOD
22833|WEST HOMESTEAD
22834|WEST HURLEY
22835|WEST ISHPEMING
22836|WEST ISLIP
22837|WEST JEFFERSON
22838|WEST JERSEY
22839|WEST JORDAN
22840|WEST KENNEBUNK
22841|WEST KINGSTON
22842|WEST KITTANNING
22843|WEST LAFAYETTE
22844|WEST LAKE HILLS
22845|WEST LAKE SAMMAMISH
22846|WEST LAKE WALES
22847|WEST LAUREL
22848|WEST LAWN
22849|WEST LEBANON
22850|WEST LEECHBURG
22851|WEST LEIPSIC
22852|WEST LIBERTY
22853|WEST LINCOLN
22854|WEST LINE
22855|WEST LINN
22856|WEST LITTLE RIVER
22857|WEST LIVINGSTON
22858|WEST LOGAN
22859|WEST LONG BRANCH
22860|WEST LOUISVILLE
22861|WEST MANCHESTER
22862|WEST MANSFIELD
22863|WEST MARION
22864|WEST MAYFIELD
22865|WEST MEDWAY
22866|WEST MELBOURNE
22867|WEST MEMPHIS
22868|WEST MENLO PARK
22869|WEST MIAMI
22870|WEST MIDDLESEX
22871|WEST MIDDLETOWN
22872|WEST MIFFLIN
22873|WEST MILFORD
22874|WEST MILLGROVE
22875|WEST MILTON
22876|WEST MILWAUKEE
22877|WEST MINERAL
22878|WEST MONROE
22879|WEST MOUNTAIN
22880|WEST MYSTIC
22881|WEST NANTICOKE
22882|WEST NEW YORK
22883|WEST NEWTON
22884|WEST NYACK
22885|WEST OCEAN CITY
22886|WEST ODESSA
22887|WEST OKOBOJI
22888|WEST ORANGE
22889|WEST PALM BEACH
22890|WEST PARK
22891|WEST PASCO
22892|WEST PAWLET
22893|WEST PEAVINE
22894|WEST PELZER
22895|WEST PENSACOLA
22896|WEST PEORIA
22897|WEST PERRINE
22898|WEST PIKE
22899|WEST PITTSBURG
22900|WEST PITTSTON
22901|WEST PLAINS
22902|WEST POCOMOKE
22903|WEST POINT
22904|WEST PORTSMOUTH
22905|WEST PUENTE VALLEY
22906|WEST RANCHO DOMINGUEZ
22907|WEST READING
22908|WEST RICHFIELD
22909|WEST RICHLAND
22910|WEST RIVERSIDE
22911|WEST ROXBURY
22912|WEST RUSHVILLE
22913|WEST RUTLAND
22914|WEST SACRAMENTO
22915|WEST SAINT PAUL
22916|WEST SALEM
22917|WEST SAMOSET
22918|WEST SAND LAKE
22919|WEST SAYVILLE
22920|WEST SCIO
22921|WEST SEBOEIS
22922|WEST SELMONT
22923|WEST SENECA
22924|WEST SHARYLAND
22925|WEST SHILOH
22926|WEST SILOAM SPRINGS
22927|WEST SIMSBURY
22928|WEST SLOPE
22929|WEST SMITHFIELD
22930|WEST SPRINGFIELD
22931|WEST STEWARTSTOWN
22932|WEST SULLIVAN
22933|WEST SUNBURY
22934|WEST SWANZEY
22935|WEST TAWAKONI
22936|WEST TERRE HAUTE
22937|WEST THUMB
22938|WEST TOPSHAM
22939|WEST UNION
22940|WEST UNITY
22941|WEST UNIVERSITY PLACE
22942|WEST UPTON
22943|WEST VALLEY
22944|WEST VALLEY CITY
22945|WEST VANDERGRIFT
22946|WEST VIEW
22947|WEST WAREHAM
22948|WEST WARWICK
22949|WEST WAYNESBURG
22950|WEST WENDOVER
22951|WEST WHITTIER
22952|WEST WILDWOOD
22953|WEST WINFIELD
22954|WEST WYOMING
22955|WEST WYOMISSING
22956|WEST YARMOUTH
22957|WEST YELLOWSTONE
22958|WEST YORK
22959|WESTACRES
22960|WESTBEND
22961|WESTBORO
22962|WESTBOROUGH
22963|WESTBROOK
22964|WESTBURY
22965|WESTBY
22966|WESTCHASE
22967|WESTCHESTER
22968|WESTCLIFFE
22969|WESTCREEK
22970|WESTDALE
22971|WESTEL
22972|WESTEND
22973|WESTERLY
22974|WESTERN
22975|WESTERN GROVE
22976|WESTERN HILLS
22977|WESTERN LAKE
22978|WESTERN SPRINGS
22979|WESTERNPORT
22980|WESTERVELT
22981|WESTERVILLE
22982|WESTFALL
22983|WESTFIELD
22984|WESTFIELD CENTER
22985|WESTFIR
22986|WESTGATE
22987|WESTHAMPTON
22988|WESTHAMPTON BEACH
22989|WESTHAVEN
22990|WESTHOFF
22991|WESTHOPE
22992|WESTLAKE
22993|WESTLAKE CORNER
22994|WESTLAKE VILLAGE
22995|WESTLAND
22996|WESTLEY
22997|WESTLINE
22998|WESTMERE
22999|WESTMINSTER
23000|WESTMONT
23001|WESTMORELAND
23002|WESTMORELAND CITY
23003|WESTMORLAND
23004|WESTOAK
23005|WESTON
23006|WESTON LAKES
23007|WESTON MILLS
23008|WESTOVER
23009|WESTOVER HILLS
23010|WESTPHALIA
23011|WESTPOINT
23012|WESTPORT
23013|WESTSIDE
23014|WESTTOWN
23015|WESTVALE
23016|WESTVIEW
23017|WESTVIEW CIRCLE
23018|WESTVILLE
23019|WESTWATER
23020|WESTWAY
23021|WESTWEGO
23022|WESTWOOD
23023|WESTWOOD HILLS
23024|WESTWOOD LAKE
23025|WETHERINGTON
23026|WETHERSFIELD
23027|WETMORE
23028|WETONKA
23029|WETUMKA
23030|WETUMPKA
23031|WEVER
23032|WEWAHITCHKA
23033|WEWEANTIC
23034|WEWELA
23035|WEWOKA
23036|WEXFORD
23037|WEYAUWEGA
23038|WEYERHAEUSER
23039|WEYERS CAVE
23040|WHALAN
23041|WHALE PASS
23042|WHALEYVILLE
23043|WHARNCLIFFE
23044|WHARTON
23045|WHAT CHEER
23046|WHATLEY
23047|WHEAT RIDGE
23048|WHEATCROFT
23049|WHEATFIELD
23050|WHEATLAND
23051|WHEATLEY
23052|WHEATLEY HEIGHTS
23053|WHEATON
23054|WHEELER
23055|WHEELER RIDGE
23056|WHEELER SPRINGS
23057|WHEELERSBURG
23058|WHEELESS
23059|WHEELING
23060|WHEELOCK
23061|WHEELWRIGHT
23062|WHELEN SPRINGS
23063|WHETSTONE
23064|WHIGHAM
23065|WHIPHOLT
23066|WHIPPANY
23067|WHIPPLE
23068|WHISKEY CREEK
23069|WHISPERING PINES
23070|WHITAKER
23071|WHITAKERS
23072|WHITE APPLE
23073|WHITE ASH
23074|WHITE BEAD
23075|WHITE BEAR BEACH
23076|WHITE BEAR LAKE
23077|WHITE BIRD
23078|WHITE BLUFF
23079|WHITE BUTTE
23080|WHITE CASTLE
23081|WHITE CENTER
23082|WHITE CHURCH
23083|WHITE CITY
23084|WHITE CLOUD
23085|WHITE CONE
23086|WHITE CREEK
23087|WHITE CRYSTAL BEACH
23088|WHITE DEER
23089|WHITE EARTH
23090|WHITE HALL
23091|WHITE HAVEN
23092|WHITE HEATH
23093|WHITE HILLS
23094|WHITE HORSE
23095|WHITE HORSE BEACH
23096|WHITE HOUSE
23097|WHITE ISLAND SHORES
23098|WHITE LAKE
23099|WHITE MARSH
23100|WHITE MEADOW LAKE
23101|WHITE MESA
23102|WHITE MILLS
23103|WHITE MOUNTAIN
23104|WHITE MOUNTAIN LAKE
23105|WHITE OAK
23106|WHITE OWL
23107|WHITE PIGEON
23108|WHITE PINE
23109|WHITE PINES
23110|WHITE PLAINS
23111|WHITE RIVER
23112|WHITE RIVER JUNCTION
23113|WHITE ROCK
23114|WHITE SALMON
23115|WHITE SANDS
23116|WHITE SETTLEMENT
23117|WHITE SHIELD
23118|WHITE SIGNAL
23119|WHITE SPRINGS
23120|WHITE STONE
23121|WHITE SULPHUR SPRINGS
23122|WHITE SWAN
23123|WHITE TOWER
23124|WHITE WATER
23125|WHITECLAY
23126|WHITEFACE
23127|WHITEFIELD
23128|WHITEFISH
23129|WHITEFISH BAY
23130|WHITEFLAT
23131|WHITEFORD
23132|WHITEHALL
23133|WHITEHAVEN
23134|WHITEHAWK
23135|WHITEHORSE
23136|WHITEHOUSE
23137|WHITEHOUSE STATION
23138|WHITELAND
23139|WHITELAW
23140|WHITEMARSH ISLAND
23141|WHITERIVER
23142|WHITEROCKS
23143|WHITES CITY
23144|WHITES LANDING
23145|WHITESBORO
23146|WHITESBURG
23147|WHITESIDE
23148|WHITESON
23149|WHITESTONE
23150|WHITESTONE LOGGING CAMP
23151|WHITESTOWN
23152|WHITESVILLE
23153|WHITETAIL
23154|WHITETHORN
23155|WHITETOP
23156|WHITEVILLE
23157|WHITEWATER
23158|WHITEWOOD
23159|WHITEWRIGHT
23160|WHITFIELD
23161|WHITHARRAL
23162|WHITING
23163|WHITINSVILLE
23164|WHITLASH
23165|WHITLEY CITY
23166|WHITLEY GARDENS
23167|WHITMAN
23168|WHITMAN SQUARE
23169|WHITMER
23170|WHITMIRE
23171|WHITMORE LAKE
23172|WHITMORE VILLAGE
23173|WHITNEL
23174|WHITNEY
23175|WHITNEY POINT
23176|WHITSETT
23177|WHITTAKER
23178|WHITTEMORE
23179|WHITTEN
23180|WHITTIER
23181|WHITTINGTON
23182|WHITTLESEY
23183|WHITWELL
23184|WHY
23185|WHYTE
23186|WIBAUX
23187|WICHITA
23188|WICHITA FALLS
23189|WICK
23190|WICKATUNK
23191|WICKENBURG
23192|WICKERHAM MANOR
23193|WICKERSHAM
23194|WICKES
23195|WICKETT
23196|WICKLIFFE
23197|WICKSVILLE
23198|WICOMICO CHURCH
23199|WICONISCO
23200|WIDE RUINS
23201|WIDEMAN
23202|WIDENER
23203|WIEDERKEHR VILLAGE
23204|WIGGINS
23205|WIGHTMANS GROVE
23206|WIGWAM
23207|WIKIEUP
23208|WILBER
23209|WILBERFORCE
23210|WILBRAHAM
23211|WILBUR
23212|WILBUR PARK
23213|WILBURTON
23214|WILBURTON NUMBER ONE
23215|WILBURTON NUMBER TWO
23216|WILCOX
23217|WILD CHERRY
23218|WILD HORSE
23219|WILD PEACH VILLAGE
23220|WILD ROSE
23221|WILDELL
23222|WILDER
23223|WILDERNESS
23224|WILDERSVILLE
23225|WILDERVILLE
23226|WILDOMAR
23227|WILDORADO
23228|WILDROSE
23229|WILDWOOD
23230|WILDWOOD CREST
23231|WILDWOOD LAKE
23232|WILEY
23233|WILEY FORD
23234|WILHOIT
23235|WILKES BARRE
23236|WILKES-BARRE
23237|WILKESBORO
23238|WILKESON
23239|WILKESVILLE
23240|WILKINSBURG
23241|WILKINSON
23242|WILKINSON HEIGHTS
23243|WILLACOOCHEE
23244|WILLAHA
23245|WILLAMINA
23246|WILLAPA
23247|WILLARD
23248|WILLARDS
23249|WILLCOX
23250|WILLERNIE
23251|WILLETTE
23252|WILLEY
23253|WILLHOIT
23254|WILLIAMS
23255|WILLIAMS BAY
23256|WILLIAMS CREEK
23257|WILLIAMS PARK
23258|WILLIAMSBURG
23259|WILLIAMSDALE
23260|WILLIAMSFIELD
23261|WILLIAMSON
23262|WILLIAMSPORT
23263|WILLIAMSTON
23264|WILLIAMSTOWN
23265|WILLIAMSVILLE
23266|WILLIFORD
23267|WILLIMANTIC
23268|WILLINGBORO
23269|WILLINGTON
23270|WILLIS
23271|WILLISBURG
23272|WILLISTON
23273|WILLISTON HIGHLANDS
23274|WILLISTON PARK
23275|WILLISVILLE
23276|WILLITS
23277|WILLMAR
23278|WILLOUGHBY
23279|WILLOUGHBY HILLS
23280|WILLOW
23281|WILLOW CANYON
23282|WILLOW CITY
23283|WILLOW CREEK
23284|WILLOW GLEN
23285|WILLOW GROVE
23286|WILLOW HILL
23287|WILLOW ISLAND
23288|WILLOW LAKE
23289|WILLOW OAK
23290|WILLOW PARK
23291|WILLOW RANCH
23292|WILLOW RIVER
23293|WILLOW RUN
23294|WILLOW SPRINGS
23295|WILLOW STREET
23296|WILLOW VALLEY
23297|WILLOWBROOK
23298|WILLOWDALE
23299|WILLOWICK
23300|WILLOWS
23301|WILLOWVILLE
23302|WILLS POINT
23303|WILLSBORO
23304|WILLSBORO POINT
23305|WILLSHIRE
23306|WILMA
23307|WILMAR
23308|WILMER
23309|WILMERDING
23310|WILMETTE
23311|WILMINGTON
23312|WILMINGTON ISLAND
23313|WILMINGTON MANOR
23314|WILMONT
23315|WILMORE
23316|WILMOT
23317|WILNA
23318|WILNO
23319|WILROADS GARDENS
23320|WILSALL
23321|WILSEY
23322|WILSEYVILLE
23323|WILSON
23324|WILSON CITY
23325|WILSON CREEK
23326|WILSONIA
23327|WILSONS
23328|WILSONS MILLS
23329|WILSONVILLE
23330|WILTON
23331|WILTON CENTER
23332|WILTON MANORS
23333|WIMAUMA
23334|WIMBERLEY
23335|WIMBLEDON
23336|WIMER
23337|WINAMAC
23338|WINBORN
23339|WINCHELL
23340|WINCHENDON
23341|WINCHESTER
23342|WINCHESTER BAY
23343|WIND GAP
23344|WIND LAKE
23345|WIND POINT
23346|WIND RIDGE
23347|WINDBER
23348|WINDCREST
23349|WINDEMERE
23350|WINDER
23351|WINDERMERE
23352|WINDFALL
23353|WINDHAM
23354|WINDHORST
23355|WINDMILL
23356|WINDOM
23357|WINDOW ROCK
23358|WINDSOR
23359|WINDSOR FOREST
23360|WINDSOR HEIGHTS
23361|WINDSOR HILLS
23362|WINDSOR LOCKS
23363|WINDSOR MILL
23364|WINDSOR PLACE
23365|WINDTHORST
23366|WINDY HILLS
23367|WINDYVILLE
23368|WINESBURG
23369|WINFALL
23370|WINFIELD
23371|WINFRED
23372|WING
23373|WINGATE
23374|WINGER
23375|WINGO
23376|WINIFRED
23377|WINIGAN
23378|WINK
23379|WINKELMAN
23380|WINLOCK
23381|WINN
23382|WINNABOW
23383|WINNEBAGO
23384|WINNECONNE
23385|WINNEMUCCA
23386|WINNER
23387|WINNETKA
23388|WINNETOON
23389|WINNETT
23390|WINNFIELD
23391|WINNIE
23392|WINNSBORO
23393|WINNSBORO MILLS
23394|WINOKUR
23395|WINONA
23396|WINONA LAKE
23397|WINOOSKI
23398|WINSIDE
23399|WINSLOW
23400|WINSLOW WEST
23401|WINSTED
23402|WINSTON
23403|WINSTON SALEM
23404|WINSTON-SALEM
23405|WINSTONVILLE
23406|WINTER
23407|WINTER BEACH
23408|WINTER GARDEN
23409|WINTER GARDENS
23410|WINTER HARBOR
23411|WINTER HAVEN
23412|WINTER PARK
23413|WINTER SPRINGS
23414|WINTERBORO
23415|WINTERGREEN
23416|WINTERHAVEN
23417|WINTERPOCK
23418|WINTERPORT
23419|WINTERS
23420|WINTERSBURG
23421|WINTERSET
23422|WINTERSTOWN
23423|WINTERSVILLE
23424|WINTERVILLE
23425|WINTHROP
23426|WINTHROP HARBOR
23427|WINTON
23428|WIOTA
23429|WIRT
23430|WISACKY
23431|WISCASSET
23432|WISCON
23433|WISCONSIN DELLS
23434|WISCONSIN RAPIDS
23435|WISDOM
23436|WISE
23437|WISE RIVER
23438|WISEMAN
23439|WISHEK
23440|WISHRAM
23441|WISNER
23442|WISTER
23443|WITCO
23444|WITHAMSVILLE
23445|WITHEE
23446|WITHERBEE
23447|WITHERS
23448|WITHROW
23449|WITMER
23450|WITOKA
23451|WITT
23452|WITTEN
23453|WITTENBERG
23454|WITTER
23455|WITTMAN
23456|WITTMANN
23457|WITTS SPRINGS
23458|WIXOM
23459|WIXON VALLEY
23460|WOBURN
23461|WODEN
23462|WOFFORD HEIGHTS
23463|WOLBACH
23464|WOLCOTT
23465|WOLCOTTVILLE
23466|WOLF
23467|WOLF BAYOU
23468|WOLF CREEK
23469|WOLF LAKE
23470|WOLF POINT
23471|WOLF SUMMIT
23472|WOLF TRAP
23473|WOLFDALE
23474|WOLFE CITY
23475|WOLFEBORO
23476|WOLFFORTH
23477|WOLFHURST
23478|WOLFLAKE
23479|WOLFORD
23480|WOLLOCHET
23481|WOLSEY
23482|WOLVERINE
23483|WOLVERINE LAKE
23484|WOLVERTON
23485|WOMELSDORF
23486|WOMENS BAY
23487|WONDER LAKE
23488|WONDERVU
23489|WONEWOC
23490|WONNIE
23491|WOOD
23492|WOOD DALE
23493|WOOD HEIGHTS
23494|WOOD LAKE
23495|WOOD RIVER
23496|WOOD VILLAGE
23497|WOOD-LYNNE
23498|WOOD-RIDGE
23499|WOODACRE
23500|WOODALL
23501|WOODARDVILLE
23502|WOODBERRY
23503|WOODBINE
23504|WOODBOURNE
23505|WOODBRANCH
23506|WOODBRIDGE
23507|WOODBURN
23508|WOODBURY
23509|WOODBURY HEIGHTS
23510|WOODCLIFF LAKE
23511|WOODCOCK
23512|WOODCREEK
23513|WOODCREST
23514|WOODFIELD
23515|WOODFIN
23516|WOODFORD
23517|WOODFORDS
23518|WOODHAVEN
23519|WOODHULL
23520|WOODINVILLE
23521|WOODLAKE
23522|WOODLAND
23523|WOODLAND BEACH
23524|WOODLAND HEIGHTS
23525|WOODLAND HILLS
23526|WOODLAND MILLS
23527|WOODLAND PARK
23528|WOODLAWN
23529|WOODLAWN BEACH
23530|WOODLAWN HEIGHTS
23531|WOODLAWN PARK
23532|WOODLEAF
23533|WOODLOCH
23534|WOODLYN
23535|WOODMAN
23536|WOODMERE
23537|WOODMONT
23538|WOODMONT BEACH
23539|WOODMOOR
23540|WOODMORE
23541|WOODPORT
23542|WOODRIDGE
23543|WOODROW
23544|WOODRUFF
23545|WOODS BAY
23546|WOODS CREEK
23547|WOODS CROSS
23548|WOODS HOLE
23549|WOODS LANDING
23550|WOODS TAVERN
23551|WOODSBORO
23552|WOODSBURGH
23553|WOODSDALE
23554|WOODSFIELD
23555|WOODSIDE
23556|WOODSON TERRACE
23557|WOODSTOCK
23558|WOODSTON
23559|WOODSTOWN
23560|WOODSVILLE
23561|WOODVILLE
23562|WOODWARD
23563|WOODWAY
23564|WOODWORTH
23565|WOODY CREEK
23566|WOOL MARKET
23567|WOOLDRIDGE
23568|WOOLSEY
23569|WOOLSTOCK
23570|WOOLWINE
23571|WOONSOCKET
23572|WOOSTER
23573|WOOSUNG
23574|WORCESTER
23575|WORDEN
23576|WORLAND
23577|WORLEY
23578|WORMLEYSBURG
23579|WORTH
23580|WORTHAM
23581|WORTHING
23582|WORTHINGTON
23583|WORTHINGTON HILLS
23584|WORTHINGTON SPRINGS
23585|WORTHVILLE
23586|WORTON
23587|WOUNDED KNEE
23588|WOXALL
23589|WRANGELL
23590|WRAY
23591|WREN
23592|WRENS
23593|WRENSHALL
23594|WRIGHT
23595|WRIGHT CITY
23596|WRIGHTS CORNERS
23597|WRIGHTSBORO
23598|WRIGHTSTOWN
23599|WRIGHTSVILLE
23600|WRIGHTSVILLE BEACH
23601|WRIGHTWOOD
23602|WRIGLEY
23603|WURTLAND
23604|WURTSBORO
23605|WYACONDA
23606|WYALUSING
23607|WYANDANCH
23608|WYANDOTTE
23609|WYANET
23610|WYANO
23611|WYARNO
23612|WYATT
23613|WYATTE
23614|WYATTVILLE
23615|WYE
23616|WYE MILLS
23617|WYEVILLE
23618|WYKOFF
23619|WYLANDVILLE
23620|WYLDWOOD
23621|WYLIE
23622|WYLLIESBURG
23623|WYMAN
23624|WYMER
23625|WYMORE
23626|WYNANTSKILL
23627|WYNCOTE
23628|WYNDHAM
23629|WYNDMERE
23630|WYNDMOOR
23631|WYNNBURG
23632|WYNNE
23633|WYNNEDALE
23634|WYNNEWOOD
23635|WYNONA
23636|WYNOT
23637|WYOCENA
23638|WYODAK
23639|WYOLA
23640|WYOMING
23641|WYOMISSING
23642|WYOMISSING HILLS
23643|WYTHEVILLE
23644|WYTOPITLOCK
23645|XENIA
23646|Y CITY
23647|Y-O RANCH
23648|YAAK
23649|YABUCOA
23650|YABUCOA ZONA URBANA
23651|YACHATS
23652|YACOLT
23653|YADKIN VALLEY
23654|YADKINVILLE
23655|YAH-TA-HEY
23656|YAKIMA
23657|YAKUTAT
23658|YALAHA
23659|YALE
23660|YAMHILL
23661|YAMPA
23662|YAMPAI
23663|YANCEY
23664|YANCEYVILLE
23665|YANCOPIN
23666|YANKEE HILL
23667|YANKEE LAKE
23668|YANKEETOWN
23669|YANKTON
23670|YANTIS
23671|YANUSH
23672|YAPHANK
23673|YARBO
23674|YARBOROUGH LANDING
23675|YARDLEY
23676|YARDVILLE
23677|YARMOUTH
23678|YARMOUTH PORT
23679|YARNELL
23680|YARROW POINT
23681|YARROWSBURG
23682|YATES
23683|YATES CENTER
23684|YATES CITY
23685|YATESBORO
23686|YATESVILLE
23687|YAUCO
23688|YAUCO ZONA URBANA
23689|YAUREL
23690|YAUREL COMUNIDAD
23691|YAZOO CITY
23692|YEADON
23693|YEAGER
23694|YEAGERTOWN
23695|YEDDO
23696|YEEHAW JUNCTION
23697|YELLOW BLUFF
23698|YELLOW JACKET
23699|YELLOW LAKE
23700|YELLOW PINE
23701|YELLOW SPRINGS
23702|YELLVILLE
23703|YELM
23704|YEMASSEE
23705|YEOMAN
23706|YERINGTON
23707|YERKES
23708|YERMO
23709|YESO
23710|YETTEM
23711|YETTER
23712|YEWED
23713|YOAKUM
23714|YOCEMENTO
23715|YODER
23716|YOE
23717|YOGAVILLE
23718|YOLO
23719|YOMAN
23720|YONAH
23721|YONCALLA
23722|YONKERS
23723|YORBA LINDA
23724|YORK
23725|YORK CENTER
23726|YORK HARBOR
23727|YORK HAVEN
23728|YORK HAVEN ANCHORAGE
23729|YORK SPRINGS
23730|YORKANA
23731|YORKETOWN
23732|YORKFIELD
23733|YORKLYN
23734|YORKSHIRE
23735|YORKTOWN
23736|YORKTOWN HEIGHTS
23737|YORKVILLE
23738|YOSEMITE
23739|YOSEMITE LAKES
23740|YOUNG
23741|YOUNG AMERICA
23742|YOUNG HARRIS
23743|YOUNGSTOWN
23744|YOUNGSVILLE
23745|YOUNGTOWN
23746|YOUNGWOOD
23747|YOUNTVILLE
23748|YPSILANTI
23749|YREKA
23750|YSCLOSKEY
23751|YUBA
23752|YUBA CITY
23753|YUCAIPA
23754|YUCCA
23755|YUCCA VALLEY
23756|YUKON
23757|YULEE
23758|YUMA
23759|YUTAN
23760|YZNAGA
23761|ZACHARY
23762|ZAFRA
23763|ZAG
23764|ZAHL
23765|ZALESKI
23766|ZALMA
23767|ZAMA
23768|ZANE
23769|ZANESFIELD
23770|ZANESVILLE
23771|ZAP
23772|ZAPATA
23773|ZAPATA RANCH
23774|ZAREPHATH
23775|ZAVALLA
23776|ZAYANTE
23777|ZEARING
23778|ZEB
23779|ZEBA
23780|ZEBINA
23781|ZEBULON
23782|ZEELAND
23783|ZEIGLER
23784|ZELA
23785|ZELIENOPLE
23786|ZELL
23787|ZELLWOOD
23788|ZEMPLE
23789|ZENA
23790|ZENDA
23791|ZENITH
23792|ZEPHYR
23793|ZEPHYR COVE
23794|ZEPHYRHILLS
23795|ZIA PUEBLO
23796|ZIHLMAN
23797|ZILLAH
23798|ZILWAUKEE
23799|ZIM
23800|ZIMMERMAN
23801|ZINC
23802|ZION
23803|ZIONSVILLE
23804|ZITA
23805|ZOAR
23806|ZOLFO SPRINGS
23807|ZONA
23808|ZORTMAN
23809|ZUEHL
23810|ZUMBRO FALLS
23811|ZUMBROTA
23812|ZUNI
23813|ZUNI PUEBLO
23814|ZURICH
23815|ZWINGLE
23816|ZWOLLE
23817|ĀHUIMANU
23818|ĀINALOA
23819|ŌMAʻO
23820|ŌʻŌKALA
