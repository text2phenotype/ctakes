C0364968|T201|LN|2823-3|LNC2HPO|Hyperkalemia|Hyperkalemia
C0364968|T201|MTH_LN|2823-3|LNC2HPO|Hyperkalemia|Hyperkalemia
C0364968|T201|DN|2823-3|LNC2HPO|Hyperkalemia|Hyperkalemia
C0364968|T201|OSN|2823-3|LNC2HPO|Hyperkalemia|Hyperkalemia
C0364968|T201|LC|2823-3|LNC2HPO|Hyperkalemia|Hyperkalemia
C0364968|T201|LN|2823-3|LNC2HPO|Hypokalemia|Hypokalemia
C0364968|T201|MTH_LN|2823-3|LNC2HPO|Hypokalemia|Hypokalemia
C0364968|T201|DN|2823-3|LNC2HPO|Hypokalemia|Hypokalemia
C0364968|T201|OSN|2823-3|LNC2HPO|Hypokalemia|Hypokalemia
C0364968|T201|LC|2823-3|LNC2HPO|Hypokalemia|Hypokalemia
C0364207|T201|LN|2075-0|LNC2HPO|Hyperchloremia|Hyperchloremia
C0364207|T201|MTH_LN|2075-0|LNC2HPO|Hyperchloremia|Hyperchloremia
C0364207|T201|DN|2075-0|LNC2HPO|Hyperchloremia|Hyperchloremia
C0364207|T201|OSN|2075-0|LNC2HPO|Hyperchloremia|Hyperchloremia
C0364207|T201|LC|2075-0|LNC2HPO|Hyperchloremia|Hyperchloremia
C0364207|T201|LN|2075-0|LNC2HPO|Hypochloremia|Hypochloremia
C0364207|T201|MTH_LN|2075-0|LNC2HPO|Hypochloremia|Hypochloremia
C0364207|T201|DN|2075-0|LNC2HPO|Hypochloremia|Hypochloremia
C0364207|T201|OSN|2075-0|LNC2HPO|Hypochloremia|Hypochloremia
C0364207|T201|LC|2075-0|LNC2HPO|Hypochloremia|Hypochloremia
C0362994|T201|OSN|777-3|LNC2HPO|Thrombocytosis|Thrombocytosis
C0362994|T201|LN|777-3|LNC2HPO|Thrombocytosis|Thrombocytosis
C0362994|T201|DN|777-3|LNC2HPO|Thrombocytosis|Thrombocytosis
C0362994|T201|MTH_LN|777-3|LNC2HPO|Thrombocytosis|Thrombocytosis
C0362994|T201|LC|777-3|LNC2HPO|Thrombocytosis|Thrombocytosis
C0362994|T201|OSN|777-3|LNC2HPO|Thrombocythemia|Thrombocythemia
C0362994|T201|LN|777-3|LNC2HPO|Thrombocythemia|Thrombocythemia
C0362994|T201|DN|777-3|LNC2HPO|Thrombocythemia|Thrombocythemia
C0362994|T201|MTH_LN|777-3|LNC2HPO|Thrombocythemia|Thrombocythemia
C0362994|T201|LC|777-3|LNC2HPO|Thrombocythemia|Thrombocythemia
C0362994|T201|OSN|777-3|LNC2HPO|Thrombocythaemia|Thrombocythaemia
C0362994|T201|LN|777-3|LNC2HPO|Thrombocythaemia|Thrombocythaemia
C0362994|T201|DN|777-3|LNC2HPO|Thrombocythaemia|Thrombocythaemia
C0362994|T201|MTH_LN|777-3|LNC2HPO|Thrombocythaemia|Thrombocythaemia
C0362994|T201|LC|777-3|LNC2HPO|Thrombocythaemia|Thrombocythaemia
C0362994|T201|OSN|777-3|LNC2HPO|Thrombocytopenia|Thrombocytopenia
C0362994|T201|LN|777-3|LNC2HPO|Thrombocytopenia|Thrombocytopenia
C0362994|T201|DN|777-3|LNC2HPO|Thrombocytopenia|Thrombocytopenia
C0362994|T201|MTH_LN|777-3|LNC2HPO|Thrombocytopenia|Thrombocytopenia
C0362994|T201|LC|777-3|LNC2HPO|Thrombocytopenia|Thrombocytopenia
C0362908|T201|LN|787-2|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C0362908|T201|MTH_LN|787-2|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C0362908|T201|LC|787-2|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C0362908|T201|DN|787-2|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C0362908|T201|OSN|787-2|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C0362908|T201|LN|787-2|LNC2HPO|Microcytosis|Microcytosis
C0362908|T201|MTH_LN|787-2|LNC2HPO|Microcytosis|Microcytosis
C0362908|T201|LC|787-2|LNC2HPO|Microcytosis|Microcytosis
C0362908|T201|DN|787-2|LNC2HPO|Microcytosis|Microcytosis
C0362908|T201|OSN|787-2|LNC2HPO|Microcytosis|Microcytosis
C0365095|T201|LN|2951-2|LNC2HPO|Hypernatremia|Hypernatremia
C0365095|T201|MTH_LN|2951-2|LNC2HPO|Hypernatremia|Hypernatremia
C0365095|T201|DN|2951-2|LNC2HPO|Hypernatremia|Hypernatremia
C0365095|T201|OSN|2951-2|LNC2HPO|Hypernatremia|Hypernatremia
C0365095|T201|LC|2951-2|LNC2HPO|Hypernatremia|Hypernatremia
C0365095|T201|LN|2951-2|LNC2HPO|Hyponatremia|Hyponatremia
C0365095|T201|MTH_LN|2951-2|LNC2HPO|Hyponatremia|Hyponatremia
C0365095|T201|DN|2951-2|LNC2HPO|Hyponatremia|Hyponatremia
C0365095|T201|OSN|2951-2|LNC2HPO|Hyponatremia|Hyponatremia
C0365095|T201|LC|2951-2|LNC2HPO|Hyponatremia|Hyponatremia
C0484731|T201|MTH_LN|2345-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0484731|T201|LN|2345-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0484731|T201|DN|2345-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0484731|T201|OSN|2345-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0484731|T201|LC|2345-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0484731|T201|MTH_LN|2345-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0484731|T201|LN|2345-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0484731|T201|DN|2345-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0484731|T201|OSN|2345-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0484731|T201|LC|2345-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0484731|T201|MTH_LN|2345-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0484731|T201|LN|2345-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0484731|T201|DN|2345-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0484731|T201|OSN|2345-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0484731|T201|LC|2345-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0800968|T201|LC|17861-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0800968|T201|MTH_LN|17861-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0800968|T201|LN|17861-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0800968|T201|DN|17861-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0800968|T201|OSN|17861-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0800968|T201|LC|17861-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0800968|T201|MTH_LN|17861-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0800968|T201|LN|17861-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0800968|T201|DN|17861-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0800968|T201|OSN|17861-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0800968|T201|LC|17861-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0800968|T201|MTH_LN|17861-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0800968|T201|LN|17861-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0800968|T201|DN|17861-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0800968|T201|OSN|17861-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0800968|T201|LC|17861-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0800968|T201|MTH_LN|17861-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0800968|T201|LN|17861-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0800968|T201|DN|17861-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0800968|T201|OSN|17861-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364160|T201|LN|2028-9|LNC2HPO|Hypercapnia|Hypercapnia
C0364160|T201|MTH_LN|2028-9|LNC2HPO|Hypercapnia|Hypercapnia
C0364160|T201|DN|2028-9|LNC2HPO|Hypercapnia|Hypercapnia
C0364160|T201|OSN|2028-9|LNC2HPO|Hypercapnia|Hypercapnia
C0364160|T201|LC|2028-9|LNC2HPO|Hypercapnia|Hypercapnia
C0364160|T201|LN|2028-9|LNC2HPO|Hypercarbia|Hypercarbia
C0364160|T201|MTH_LN|2028-9|LNC2HPO|Hypercarbia|Hypercarbia
C0364160|T201|DN|2028-9|LNC2HPO|Hypercarbia|Hypercarbia
C0364160|T201|OSN|2028-9|LNC2HPO|Hypercarbia|Hypercarbia
C0364160|T201|LC|2028-9|LNC2HPO|Hypercarbia|Hypercarbia
C0364160|T201|LN|2028-9|LNC2HPO|Hypocapnia|Hypocapnia
C0364160|T201|MTH_LN|2028-9|LNC2HPO|Hypocapnia|Hypocapnia
C0364160|T201|DN|2028-9|LNC2HPO|Hypocapnia|Hypocapnia
C0364160|T201|OSN|2028-9|LNC2HPO|Hypocapnia|Hypocapnia
C0364160|T201|LC|2028-9|LNC2HPO|Hypocapnia|Hypocapnia
C0364160|T201|LN|2028-9|LNC2HPO|Hypocarbia|Hypocarbia
C0364160|T201|MTH_LN|2028-9|LNC2HPO|Hypocarbia|Hypocarbia
C0364160|T201|DN|2028-9|LNC2HPO|Hypocarbia|Hypocarbia
C0364160|T201|OSN|2028-9|LNC2HPO|Hypocarbia|Hypocarbia
C0364160|T201|LC|2028-9|LNC2HPO|Hypocarbia|Hypocarbia
C1315182|T201|MTH_LN|32623-1|LNC2HPO|Large platelets|Large platelets
C1315182|T201|DN|32623-1|LNC2HPO|Large platelets|Large platelets
C1315182|T201|LN|32623-1|LNC2HPO|Large platelets|Large platelets
C1315182|T201|LC|32623-1|LNC2HPO|Large platelets|Large platelets
C1315182|T201|OSN|32623-1|LNC2HPO|Large platelets|Large platelets
C1315182|T201|MTH_LN|32623-1|LNC2HPO|Small platelet size|Small platelet size
C1315182|T201|DN|32623-1|LNC2HPO|Small platelet size|Small platelet size
C1315182|T201|LN|32623-1|LNC2HPO|Small platelet size|Small platelet size
C1315182|T201|LC|32623-1|LNC2HPO|Small platelet size|Small platelet size
C1315182|T201|OSN|32623-1|LNC2HPO|Small platelet size|Small platelet size
C1315182|T201|MTH_LN|32623-1|LNC2HPO|Small platelets size|Small platelets size
C1315182|T201|DN|32623-1|LNC2HPO|Small platelets size|Small platelets size
C1315182|T201|LN|32623-1|LNC2HPO|Small platelets size|Small platelets size
C1315182|T201|LC|32623-1|LNC2HPO|Small platelets size|Small platelets size
C1315182|T201|OSN|32623-1|LNC2HPO|Small platelets size|Small platelets size
C1315182|T201|MTH_LN|32623-1|LNC2HPO|Small platelets|Small platelets
C1315182|T201|DN|32623-1|LNC2HPO|Small platelets|Small platelets
C1315182|T201|LN|32623-1|LNC2HPO|Small platelets|Small platelets
C1315182|T201|LC|32623-1|LNC2HPO|Small platelets|Small platelets
C1315182|T201|OSN|32623-1|LNC2HPO|Small platelets|Small platelets
C0802053|T201|LC|19123-9|LNC2HPO|Hypermagnesemia|Hypermagnesemia
C0802053|T201|MTH_LN|19123-9|LNC2HPO|Hypermagnesemia|Hypermagnesemia
C0802053|T201|LN|19123-9|LNC2HPO|Hypermagnesemia|Hypermagnesemia
C0802053|T201|DN|19123-9|LNC2HPO|Hypermagnesemia|Hypermagnesemia
C0802053|T201|OSN|19123-9|LNC2HPO|Hypermagnesemia|Hypermagnesemia
C0802053|T201|LC|19123-9|LNC2HPO|Hypomagnesemia|Hypomagnesemia
C0802053|T201|MTH_LN|19123-9|LNC2HPO|Hypomagnesemia|Hypomagnesemia
C0802053|T201|LN|19123-9|LNC2HPO|Hypomagnesemia|Hypomagnesemia
C0802053|T201|DN|19123-9|LNC2HPO|Hypomagnesemia|Hypomagnesemia
C0802053|T201|OSN|19123-9|LNC2HPO|Hypomagnesemia|Hypomagnesemia
C0484430|T201|LN|6690-2|LNC2HPO|Leukocytosis|Leukocytosis
C0484430|T201|DN|6690-2|LNC2HPO|Leukocytosis|Leukocytosis
C0484430|T201|OSN|6690-2|LNC2HPO|Leukocytosis|Leukocytosis
C0484430|T201|MTH_LN|6690-2|LNC2HPO|Leukocytosis|Leukocytosis
C0484430|T201|LC|6690-2|LNC2HPO|Leukocytosis|Leukocytosis
C0484430|T201|LN|6690-2|LNC2HPO|Leukopenia|Leukopenia
C0484430|T201|DN|6690-2|LNC2HPO|Leukopenia|Leukopenia
C0484430|T201|OSN|6690-2|LNC2HPO|Leukopenia|Leukopenia
C0484430|T201|MTH_LN|6690-2|LNC2HPO|Leukopenia|Leukopenia
C0484430|T201|LC|6690-2|LNC2HPO|Leukopenia|Leukopenia
C1370010|T201|MTH_LN|2777-1|LNC2HPO|Hyperphosphatemia|Hyperphosphatemia
C1370010|T201|LN|2777-1|LNC2HPO|Hyperphosphatemia|Hyperphosphatemia
C1370010|T201|DN|2777-1|LNC2HPO|Hyperphosphatemia|Hyperphosphatemia
C1370010|T201|OSN|2777-1|LNC2HPO|Hyperphosphatemia|Hyperphosphatemia
C1370010|T201|LC|2777-1|LNC2HPO|Hyperphosphatemia|Hyperphosphatemia
C1370010|T201|MTH_LN|2777-1|LNC2HPO|Hypophosphatemia|Hypophosphatemia
C1370010|T201|LN|2777-1|LNC2HPO|Hypophosphatemia|Hypophosphatemia
C1370010|T201|DN|2777-1|LNC2HPO|Hypophosphatemia|Hypophosphatemia
C1370010|T201|OSN|2777-1|LNC2HPO|Hypophosphatemia|Hypophosphatemia
C1370010|T201|LC|2777-1|LNC2HPO|Hypophosphatemia|Hypophosphatemia
C1370010|T201|MTH_LN|2777-1|LNC2HPO|Hypophosphataemia|Hypophosphataemia
C1370010|T201|LN|2777-1|LNC2HPO|Hypophosphataemia|Hypophosphataemia
C1370010|T201|DN|2777-1|LNC2HPO|Hypophosphataemia|Hypophosphataemia
C1370010|T201|OSN|2777-1|LNC2HPO|Hypophosphataemia|Hypophosphataemia
C1370010|T201|LC|2777-1|LNC2HPO|Hypophosphataemia|Hypophosphataemia
C0550846|T201|LN|12227-5|LNC2HPO|Leukocytosis|Leukocytosis
C0550846|T201|DN|12227-5|LNC2HPO|Leukocytosis|Leukocytosis
C0550846|T201|OSN|12227-5|LNC2HPO|Leukocytosis|Leukocytosis
C0550846|T201|MTH_LN|12227-5|LNC2HPO|Leukocytosis|Leukocytosis
C0550846|T201|LC|12227-5|LNC2HPO|Leukocytosis|Leukocytosis
C0550846|T201|LN|12227-5|LNC2HPO|Leukopenia|Leukopenia
C0550846|T201|DN|12227-5|LNC2HPO|Leukopenia|Leukopenia
C0550846|T201|OSN|12227-5|LNC2HPO|Leukopenia|Leukopenia
C0550846|T201|MTH_LN|12227-5|LNC2HPO|Leukopenia|Leukopenia
C0550846|T201|LC|12227-5|LNC2HPO|Leukopenia|Leukopenia
C0362958|T201|LN|742-7|LNC2HPO|Monocytosis|Monocytosis
C0362958|T201|DN|742-7|LNC2HPO|Monocytosis|Monocytosis
C0362958|T201|OSN|742-7|LNC2HPO|Monocytosis|Monocytosis
C0362958|T201|MTH_LN|742-7|LNC2HPO|Monocytosis|Monocytosis
C0362958|T201|LC|742-7|LNC2HPO|Monocytosis|Monocytosis
C0362958|T201|LN|742-7|LNC2HPO|Monocytopenia|Monocytopenia
C0362958|T201|DN|742-7|LNC2HPO|Monocytopenia|Monocytopenia
C0362958|T201|OSN|742-7|LNC2HPO|Monocytopenia|Monocytopenia
C0362958|T201|MTH_LN|742-7|LNC2HPO|Monocytopenia|Monocytopenia
C0362958|T201|LC|742-7|LNC2HPO|Monocytopenia|Monocytopenia
C0362947|T201|LN|731-0|LNC2HPO|Lymphocytosis|Lymphocytosis
C0362947|T201|DN|731-0|LNC2HPO|Lymphocytosis|Lymphocytosis
C0362947|T201|OSN|731-0|LNC2HPO|Lymphocytosis|Lymphocytosis
C0362947|T201|MTH_LN|731-0|LNC2HPO|Lymphocytosis|Lymphocytosis
C0362947|T201|LC|731-0|LNC2HPO|Lymphocytosis|Lymphocytosis
C0362947|T201|LN|731-0|LNC2HPO|Lymphopenia|Lymphopenia
C0362947|T201|DN|731-0|LNC2HPO|Lymphopenia|Lymphopenia
C0362947|T201|OSN|731-0|LNC2HPO|Lymphopenia|Lymphopenia
C0362947|T201|MTH_LN|731-0|LNC2HPO|Lymphopenia|Lymphopenia
C0362947|T201|LC|731-0|LNC2HPO|Lymphopenia|Lymphopenia
C0362947|T201|LN|731-0|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0362947|T201|DN|731-0|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0362947|T201|OSN|731-0|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0362947|T201|MTH_LN|731-0|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0362947|T201|LC|731-0|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0362947|T201|LN|731-0|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0362947|T201|DN|731-0|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0362947|T201|OSN|731-0|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0362947|T201|MTH_LN|731-0|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0362947|T201|LC|731-0|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0798246|T201|LN|15074-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0798246|T201|MTH_LN|15074-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0798246|T201|DN|15074-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0798246|T201|OSN|15074-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0798246|T201|LC|15074-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0798246|T201|LN|15074-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0798246|T201|MTH_LN|15074-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0798246|T201|DN|15074-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0798246|T201|OSN|15074-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0798246|T201|LC|15074-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0798246|T201|LN|15074-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0798246|T201|MTH_LN|15074-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0798246|T201|DN|15074-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0798246|T201|OSN|15074-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0798246|T201|LC|15074-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1954230|T201|LN|48643-1|LNC2HPO|Impaired renal creatinine clearance|Impaired renal creatinine clearance
C1954230|T201|MTH_LN|48643-1|LNC2HPO|Impaired renal creatinine clearance|Impaired renal creatinine clearance
C1954230|T201|LC|48643-1|LNC2HPO|Impaired renal creatinine clearance|Impaired renal creatinine clearance
C1954230|T201|OSN|48643-1|LNC2HPO|Impaired renal creatinine clearance|Impaired renal creatinine clearance
C1954230|T201|DN|48643-1|LNC2HPO|Impaired renal creatinine clearance|Impaired renal creatinine clearance
C1954228|T201|LN|48642-3|LNC2HPO|Impaired renal creatinine clearance|Impaired renal creatinine clearance
C1954228|T201|LC|48642-3|LNC2HPO|Impaired renal creatinine clearance|Impaired renal creatinine clearance
C1954228|T201|OSN|48642-3|LNC2HPO|Impaired renal creatinine clearance|Impaired renal creatinine clearance
C1954228|T201|MTH_LN|48642-3|LNC2HPO|Impaired renal creatinine clearance|Impaired renal creatinine clearance
C1954228|T201|DN|48642-3|LNC2HPO|Impaired renal creatinine clearance|Impaired renal creatinine clearance
C0364480|T201|LN|2340-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0364480|T201|OSN|2340-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0364480|T201|LC|2340-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0364480|T201|MTH_LN|2340-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0364480|T201|DN|2340-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0364480|T201|LN|2340-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0364480|T201|OSN|2340-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0364480|T201|LC|2340-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0364480|T201|MTH_LN|2340-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0364480|T201|DN|2340-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0364480|T201|LN|2340-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0364480|T201|OSN|2340-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0364480|T201|LC|2340-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0364480|T201|MTH_LN|2340-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0364480|T201|DN|2340-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942437|T201|LN|26474-7|LNC2HPO|Lymphocytosis|Lymphocytosis
C0942437|T201|DN|26474-7|LNC2HPO|Lymphocytosis|Lymphocytosis
C0942437|T201|OSN|26474-7|LNC2HPO|Lymphocytosis|Lymphocytosis
C0942437|T201|MTH_LN|26474-7|LNC2HPO|Lymphocytosis|Lymphocytosis
C0942437|T201|LC|26474-7|LNC2HPO|Lymphocytosis|Lymphocytosis
C0942437|T201|LN|26474-7|LNC2HPO|Lymphopenia|Lymphopenia
C0942437|T201|DN|26474-7|LNC2HPO|Lymphopenia|Lymphopenia
C0942437|T201|OSN|26474-7|LNC2HPO|Lymphopenia|Lymphopenia
C0942437|T201|MTH_LN|26474-7|LNC2HPO|Lymphopenia|Lymphopenia
C0942437|T201|LC|26474-7|LNC2HPO|Lymphopenia|Lymphopenia
C0942437|T201|LN|26474-7|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0942437|T201|DN|26474-7|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0942437|T201|OSN|26474-7|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0942437|T201|MTH_LN|26474-7|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0942437|T201|LC|26474-7|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0942437|T201|LN|26474-7|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0942437|T201|DN|26474-7|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0942437|T201|OSN|26474-7|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0942437|T201|MTH_LN|26474-7|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0942437|T201|LC|26474-7|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0364479|T201|LN|2339-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0364479|T201|MTH_LN|2339-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0364479|T201|DN|2339-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0364479|T201|OSN|2339-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0364479|T201|LC|2339-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0364479|T201|LN|2339-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0364479|T201|MTH_LN|2339-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0364479|T201|DN|2339-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0364479|T201|OSN|2339-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0364479|T201|LC|2339-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0364479|T201|LN|2339-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0364479|T201|MTH_LN|2339-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0364479|T201|DN|2339-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0364479|T201|OSN|2339-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0364479|T201|LC|2339-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942446|T201|LN|26484-6|LNC2HPO|Monocytosis|Monocytosis
C0942446|T201|DN|26484-6|LNC2HPO|Monocytosis|Monocytosis
C0942446|T201|OSN|26484-6|LNC2HPO|Monocytosis|Monocytosis
C0942446|T201|MTH_LN|26484-6|LNC2HPO|Monocytosis|Monocytosis
C0942446|T201|LC|26484-6|LNC2HPO|Monocytosis|Monocytosis
C0942446|T201|LN|26484-6|LNC2HPO|Monocytopenia|Monocytopenia
C0942446|T201|DN|26484-6|LNC2HPO|Monocytopenia|Monocytopenia
C0942446|T201|OSN|26484-6|LNC2HPO|Monocytopenia|Monocytopenia
C0942446|T201|MTH_LN|26484-6|LNC2HPO|Monocytopenia|Monocytopenia
C0942446|T201|LC|26484-6|LNC2HPO|Monocytopenia|Monocytopenia
C0942447|T201|LN|26485-3|LNC2HPO|Monocytosis|Monocytosis
C0942447|T201|OSN|26485-3|LNC2HPO|Monocytosis|Monocytosis
C0942447|T201|DN|26485-3|LNC2HPO|Monocytosis|Monocytosis
C0942447|T201|MTH_LN|26485-3|LNC2HPO|Monocytosis|Monocytosis
C0942447|T201|LC|26485-3|LNC2HPO|Monocytosis|Monocytosis
C0942447|T201|LN|26485-3|LNC2HPO|Monocytopenia|Monocytopenia
C0942447|T201|OSN|26485-3|LNC2HPO|Monocytopenia|Monocytopenia
C0942447|T201|DN|26485-3|LNC2HPO|Monocytopenia|Monocytopenia
C0942447|T201|MTH_LN|26485-3|LNC2HPO|Monocytopenia|Monocytopenia
C0942447|T201|LC|26485-3|LNC2HPO|Monocytopenia|Monocytopenia
C0942461|T201|LN|26499-4|LNC2HPO|Neutrophilia|Neutrophilia
C0942461|T201|DN|26499-4|LNC2HPO|Neutrophilia|Neutrophilia
C0942461|T201|OSN|26499-4|LNC2HPO|Neutrophilia|Neutrophilia
C0942461|T201|MTH_LN|26499-4|LNC2HPO|Neutrophilia|Neutrophilia
C0942461|T201|LC|26499-4|LNC2HPO|Neutrophilia|Neutrophilia
C0942461|T201|LN|26499-4|LNC2HPO|Neutropenia|Neutropenia
C0942461|T201|DN|26499-4|LNC2HPO|Neutropenia|Neutropenia
C0942461|T201|OSN|26499-4|LNC2HPO|Neutropenia|Neutropenia
C0942461|T201|MTH_LN|26499-4|LNC2HPO|Neutropenia|Neutropenia
C0942461|T201|LC|26499-4|LNC2HPO|Neutropenia|Neutropenia
C0942461|T201|LN|26499-4|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0942461|T201|DN|26499-4|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0942461|T201|OSN|26499-4|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0942461|T201|MTH_LN|26499-4|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0942461|T201|LC|26499-4|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0362900|T201|LN|711-2|LNC2HPO|Eosinophilia|Eosinophilia
C0362900|T201|DN|711-2|LNC2HPO|Eosinophilia|Eosinophilia
C0362900|T201|OSN|711-2|LNC2HPO|Eosinophilia|Eosinophilia
C0362900|T201|MTH_LN|711-2|LNC2HPO|Eosinophilia|Eosinophilia
C0362900|T201|LC|711-2|LNC2HPO|Eosinophilia|Eosinophilia
C0362901|T201|LN|712-0|LNC2HPO|Eosinophilia|Eosinophilia
C0362901|T201|DN|712-0|LNC2HPO|Eosinophilia|Eosinophilia
C0362901|T201|OSN|712-0|LNC2HPO|Eosinophilia|Eosinophilia
C0362901|T201|MTH_LN|712-0|LNC2HPO|Eosinophilia|Eosinophilia
C0362901|T201|LC|712-0|LNC2HPO|Eosinophilia|Eosinophilia
C0362968|T201|OSN|751-8|LNC2HPO|Neutrophilia|Neutrophilia
C0362968|T201|LN|751-8|LNC2HPO|Neutrophilia|Neutrophilia
C0362968|T201|DN|751-8|LNC2HPO|Neutrophilia|Neutrophilia
C0362968|T201|MTH_LN|751-8|LNC2HPO|Neutrophilia|Neutrophilia
C0362968|T201|LC|751-8|LNC2HPO|Neutrophilia|Neutrophilia
C0362968|T201|OSN|751-8|LNC2HPO|Neutropenia|Neutropenia
C0362968|T201|LN|751-8|LNC2HPO|Neutropenia|Neutropenia
C0362968|T201|DN|751-8|LNC2HPO|Neutropenia|Neutropenia
C0362968|T201|MTH_LN|751-8|LNC2HPO|Neutropenia|Neutropenia
C0362968|T201|LC|751-8|LNC2HPO|Neutropenia|Neutropenia
C0362968|T201|OSN|751-8|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0362968|T201|LN|751-8|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0362968|T201|DN|751-8|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0362968|T201|MTH_LN|751-8|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0362968|T201|LC|751-8|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0364489|T201|LN|2349-9|LNC2HPO|Glycosuria|Glycosuria
C0364489|T201|MTH_LN|2349-9|LNC2HPO|Glycosuria|Glycosuria
C0364489|T201|DN|2349-9|LNC2HPO|Glycosuria|Glycosuria
C0364489|T201|OSN|2349-9|LNC2HPO|Glycosuria|Glycosuria
C0364489|T201|LC|2349-9|LNC2HPO|Glycosuria|Glycosuria
C0364489|T201|LN|2349-9|LNC2HPO|Glucosuria|Glucosuria
C0364489|T201|MTH_LN|2349-9|LNC2HPO|Glucosuria|Glucosuria
C0364489|T201|DN|2349-9|LNC2HPO|Glucosuria|Glucosuria
C0364489|T201|OSN|2349-9|LNC2HPO|Glucosuria|Glucosuria
C0364489|T201|LC|2349-9|LNC2HPO|Glucosuria|Glucosuria
C0363885|T201|LN|1751-7|LNC2HPO|Hyperalbuminemia|Hyperalbuminemia
C0363885|T201|DN|1751-7|LNC2HPO|Hyperalbuminemia|Hyperalbuminemia
C0363885|T201|MTH_LN|1751-7|LNC2HPO|Hyperalbuminemia|Hyperalbuminemia
C0363885|T201|OSN|1751-7|LNC2HPO|Hyperalbuminemia|Hyperalbuminemia
C0363885|T201|LC|1751-7|LNC2HPO|Hyperalbuminemia|Hyperalbuminemia
C0363885|T201|LN|1751-7|LNC2HPO|Hyperalbuminaemia|Hyperalbuminaemia
C0363885|T201|DN|1751-7|LNC2HPO|Hyperalbuminaemia|Hyperalbuminaemia
C0363885|T201|MTH_LN|1751-7|LNC2HPO|Hyperalbuminaemia|Hyperalbuminaemia
C0363885|T201|OSN|1751-7|LNC2HPO|Hyperalbuminaemia|Hyperalbuminaemia
C0363885|T201|LC|1751-7|LNC2HPO|Hyperalbuminaemia|Hyperalbuminaemia
C0363885|T201|LN|1751-7|LNC2HPO|Hypoalbuminemia|Hypoalbuminemia
C0363885|T201|DN|1751-7|LNC2HPO|Hypoalbuminemia|Hypoalbuminemia
C0363885|T201|MTH_LN|1751-7|LNC2HPO|Hypoalbuminemia|Hypoalbuminemia
C0363885|T201|OSN|1751-7|LNC2HPO|Hypoalbuminemia|Hypoalbuminemia
C0363885|T201|LC|1751-7|LNC2HPO|Hypoalbuminemia|Hypoalbuminemia
C0363885|T201|LN|1751-7|LNC2HPO|Hypoalbuminaemia|Hypoalbuminaemia
C0363885|T201|DN|1751-7|LNC2HPO|Hypoalbuminaemia|Hypoalbuminaemia
C0363885|T201|MTH_LN|1751-7|LNC2HPO|Hypoalbuminaemia|Hypoalbuminaemia
C0363885|T201|OSN|1751-7|LNC2HPO|Hypoalbuminaemia|Hypoalbuminaemia
C0363885|T201|LC|1751-7|LNC2HPO|Hypoalbuminaemia|Hypoalbuminaemia
C0364708|T201|MTH_LN|2093-3|LNC2HPO|Hypercholesterolemia|Hypercholesterolemia
C0364708|T201|LN|2093-3|LNC2HPO|Hypercholesterolemia|Hypercholesterolemia
C0364708|T201|DN|2093-3|LNC2HPO|Hypercholesterolemia|Hypercholesterolemia
C0364708|T201|OSN|2093-3|LNC2HPO|Hypercholesterolemia|Hypercholesterolemia
C0364708|T201|LC|2093-3|LNC2HPO|Hypercholesterolemia|Hypercholesterolemia
C0364708|T201|MTH_LN|2093-3|LNC2HPO|Hypocholesterolemia|Hypocholesterolemia
C0364708|T201|LN|2093-3|LNC2HPO|Hypocholesterolemia|Hypocholesterolemia
C0364708|T201|DN|2093-3|LNC2HPO|Hypocholesterolemia|Hypocholesterolemia
C0364708|T201|OSN|2093-3|LNC2HPO|Hypocholesterolemia|Hypocholesterolemia
C0364708|T201|LC|2093-3|LNC2HPO|Hypocholesterolemia|Hypocholesterolemia
C0484638|T201|MTH_LN|6768-6|LNC2HPO|Hyperphosphatasia|Hyperphosphatasia
C0484638|T201|LN|6768-6|LNC2HPO|Hyperphosphatasia|Hyperphosphatasia
C0484638|T201|DN|6768-6|LNC2HPO|Hyperphosphatasia|Hyperphosphatasia
C0484638|T201|OSN|6768-6|LNC2HPO|Hyperphosphatasia|Hyperphosphatasia
C0484638|T201|LC|6768-6|LNC2HPO|Hyperphosphatasia|Hyperphosphatasia
C0484638|T201|MTH_LN|6768-6|LNC2HPO|Hyperphosphatasemia|Hyperphosphatasemia
C0484638|T201|LN|6768-6|LNC2HPO|Hyperphosphatasemia|Hyperphosphatasemia
C0484638|T201|DN|6768-6|LNC2HPO|Hyperphosphatasemia|Hyperphosphatasemia
C0484638|T201|OSN|6768-6|LNC2HPO|Hyperphosphatasemia|Hyperphosphatasemia
C0484638|T201|LC|6768-6|LNC2HPO|Hyperphosphatasemia|Hyperphosphatasemia
C1316377|T201|LN|33914-3|LNC2HPO|Impaired renal creatinine clearance|Impaired renal creatinine clearance
C1316377|T201|MTH_LN|33914-3|LNC2HPO|Impaired renal creatinine clearance|Impaired renal creatinine clearance
C1316377|T201|LC|33914-3|LNC2HPO|Impaired renal creatinine clearance|Impaired renal creatinine clearance
C1316377|T201|DN|33914-3|LNC2HPO|Impaired renal creatinine clearance|Impaired renal creatinine clearance
C1316377|T201|OSN|33914-3|LNC2HPO|Impaired renal creatinine clearance|Impaired renal creatinine clearance
C0365029|T201|LN|2885-2|LNC2HPO|Hyperproteinemia|Hyperproteinemia
C0365029|T201|DN|2885-2|LNC2HPO|Hyperproteinemia|Hyperproteinemia
C0365029|T201|MTH_LN|2885-2|LNC2HPO|Hyperproteinemia|Hyperproteinemia
C0365029|T201|OSN|2885-2|LNC2HPO|Hyperproteinemia|Hyperproteinemia
C0365029|T201|LC|2885-2|LNC2HPO|Hyperproteinemia|Hyperproteinemia
C0365029|T201|LN|2885-2|LNC2HPO|Hypoproteinemia|Hypoproteinemia
C0365029|T201|DN|2885-2|LNC2HPO|Hypoproteinemia|Hypoproteinemia
C0365029|T201|MTH_LN|2885-2|LNC2HPO|Hypoproteinemia|Hypoproteinemia
C0365029|T201|OSN|2885-2|LNC2HPO|Hypoproteinemia|Hypoproteinemia
C0365029|T201|LC|2885-2|LNC2HPO|Hypoproteinemia|Hypoproteinemia
C0482694|T201|LN|5902-2|LNC2HPO|Prolonged prothrombin time|Prolonged prothrombin time
C0482694|T201|OSN|5902-2|LNC2HPO|Prolonged prothrombin time|Prolonged prothrombin time
C0482694|T201|LC|5902-2|LNC2HPO|Prolonged prothrombin time|Prolonged prothrombin time
C0482694|T201|DN|5902-2|LNC2HPO|Prolonged prothrombin time|Prolonged prothrombin time
C0482694|T201|MTH_LN|5902-2|LNC2HPO|Prolonged prothrombin time|Prolonged prothrombin time
C0482694|T201|LN|5902-2|LNC2HPO|Prolonged PT|Prolonged PT
C0482694|T201|OSN|5902-2|LNC2HPO|Prolonged PT|Prolonged PT
C0482694|T201|LC|5902-2|LNC2HPO|Prolonged PT|Prolonged PT
C0482694|T201|DN|5902-2|LNC2HPO|Prolonged PT|Prolonged PT
C0482694|T201|MTH_LN|5902-2|LNC2HPO|Prolonged PT|Prolonged PT
C0482694|T201|LN|5902-2|LNC2HPO|increased international normalised ratio|increased international normalised ratio
C0482694|T201|OSN|5902-2|LNC2HPO|increased international normalised ratio|increased international normalised ratio
C0482694|T201|LC|5902-2|LNC2HPO|increased international normalised ratio|increased international normalised ratio
C0482694|T201|DN|5902-2|LNC2HPO|increased international normalised ratio|increased international normalised ratio
C0482694|T201|MTH_LN|5902-2|LNC2HPO|increased international normalised ratio|increased international normalised ratio
C0362890|T201|LN|702-1|LNC2HPO|Anisocytosis|Anisocytosis
C0362890|T201|MTH_LN|702-1|LNC2HPO|Anisocytosis|Anisocytosis
C0362890|T201|DN|702-1|LNC2HPO|Anisocytosis|Anisocytosis
C0362890|T201|OSN|702-1|LNC2HPO|Anisocytosis|Anisocytosis
C0362890|T201|LC|702-1|LNC2HPO|Anisocytosis|Anisocytosis
C0881213|T201|LN|23860-0|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C0881213|T201|DN|23860-0|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C0881213|T201|OSN|23860-0|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C0881213|T201|MTH_LN|23860-0|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C0881213|T201|LC|23860-0|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C0881213|T201|LN|23860-0|LNC2HPO|Microcytosis|Microcytosis
C0881213|T201|DN|23860-0|LNC2HPO|Microcytosis|Microcytosis
C0881213|T201|OSN|23860-0|LNC2HPO|Microcytosis|Microcytosis
C0881213|T201|MTH_LN|23860-0|LNC2HPO|Microcytosis|Microcytosis
C0881213|T201|LC|23860-0|LNC2HPO|Microcytosis|Microcytosis
C0803268|T201|LN|20454-5|LNC2HPO|Proteinuria|Proteinuria
C0803268|T201|MTH_LN|20454-5|LNC2HPO|Proteinuria|Proteinuria
C0803268|T201|DN|20454-5|LNC2HPO|Proteinuria|Proteinuria
C0803268|T201|OSN|20454-5|LNC2HPO|Proteinuria|Proteinuria
C0803268|T201|LC|20454-5|LNC2HPO|Proteinuria|Proteinuria
C0362954|T201|LN|738-5|LNC2HPO|Macrocytic anemia|Macrocytic anemia
C0362954|T201|MTH_LN|738-5|LNC2HPO|Macrocytic anemia|Macrocytic anemia
C0362954|T201|DN|738-5|LNC2HPO|Macrocytic anemia|Macrocytic anemia
C0362954|T201|OSN|738-5|LNC2HPO|Macrocytic anemia|Macrocytic anemia
C0362954|T201|LC|738-5|LNC2HPO|Macrocytic anemia|Macrocytic anemia
C0362957|T201|LN|741-9|LNC2HPO|Microcytic anemia|Microcytic anemia
C0362957|T201|MTH_LN|741-9|LNC2HPO|Microcytic anemia|Microcytic anemia
C0362957|T201|DN|741-9|LNC2HPO|Microcytic anemia|Microcytic anemia
C0362957|T201|OSN|741-9|LNC2HPO|Microcytic anemia|Microcytic anemia
C0362957|T201|LC|741-9|LNC2HPO|Microcytic anemia|Microcytic anemia
C2736146|T201|LN|57735-3|LNC2HPO|Proteinuria|Proteinuria
C2736146|T201|MTH_LN|57735-3|LNC2HPO|Proteinuria|Proteinuria
C2736146|T201|DN|57735-3|LNC2HPO|Proteinuria|Proteinuria
C2736146|T201|OSN|57735-3|LNC2HPO|Proteinuria|Proteinuria
C2736146|T201|LC|57735-3|LNC2HPO|Proteinuria|Proteinuria
C0364714|T201|LC|2571-8|LNC2HPO|Dyslipidemia|Dyslipidemia
C0364714|T201|DN|2571-8|LNC2HPO|Dyslipidemia|Dyslipidemia
C0364714|T201|MTH_LN|2571-8|LNC2HPO|Dyslipidemia|Dyslipidemia
C0364714|T201|LN|2571-8|LNC2HPO|Dyslipidemia|Dyslipidemia
C0364714|T201|OSN|2571-8|LNC2HPO|Dyslipidemia|Dyslipidemia
C0364714|T201|LC|2571-8|LNC2HPO|Hypertriglyceridemia|Hypertriglyceridemia
C0364714|T201|DN|2571-8|LNC2HPO|Hypertriglyceridemia|Hypertriglyceridemia
C0364714|T201|MTH_LN|2571-8|LNC2HPO|Hypertriglyceridemia|Hypertriglyceridemia
C0364714|T201|LN|2571-8|LNC2HPO|Hypertriglyceridemia|Hypertriglyceridemia
C0364714|T201|OSN|2571-8|LNC2HPO|Hypertriglyceridemia|Hypertriglyceridemia
C0364714|T201|LC|2571-8|LNC2HPO|Hypotriglyceridemia|Hypotriglyceridemia
C0364714|T201|DN|2571-8|LNC2HPO|Hypotriglyceridemia|Hypotriglyceridemia
C0364714|T201|MTH_LN|2571-8|LNC2HPO|Hypotriglyceridemia|Hypotriglyceridemia
C0364714|T201|LN|2571-8|LNC2HPO|Hypotriglyceridemia|Hypotriglyceridemia
C0364714|T201|OSN|2571-8|LNC2HPO|Hypotriglyceridemia|Hypotriglyceridemia
C0364151|T201|LN|2019-8|LNC2HPO|Hypercapnia|Hypercapnia
C0364151|T201|MTH_LN|2019-8|LNC2HPO|Hypercapnia|Hypercapnia
C0364151|T201|DN|2019-8|LNC2HPO|Hypercapnia|Hypercapnia
C0364151|T201|LC|2019-8|LNC2HPO|Hypercapnia|Hypercapnia
C0364151|T201|OSN|2019-8|LNC2HPO|Hypercapnia|Hypercapnia
C0364151|T201|LN|2019-8|LNC2HPO|Hypercarbia|Hypercarbia
C0364151|T201|MTH_LN|2019-8|LNC2HPO|Hypercarbia|Hypercarbia
C0364151|T201|DN|2019-8|LNC2HPO|Hypercarbia|Hypercarbia
C0364151|T201|LC|2019-8|LNC2HPO|Hypercarbia|Hypercarbia
C0364151|T201|OSN|2019-8|LNC2HPO|Hypercarbia|Hypercarbia
C0364151|T201|LN|2019-8|LNC2HPO|Hypocapnia|Hypocapnia
C0364151|T201|MTH_LN|2019-8|LNC2HPO|Hypocapnia|Hypocapnia
C0364151|T201|DN|2019-8|LNC2HPO|Hypocapnia|Hypocapnia
C0364151|T201|LC|2019-8|LNC2HPO|Hypocapnia|Hypocapnia
C0364151|T201|OSN|2019-8|LNC2HPO|Hypocapnia|Hypocapnia
C0364151|T201|LN|2019-8|LNC2HPO|Hypocarbia|Hypocarbia
C0364151|T201|MTH_LN|2019-8|LNC2HPO|Hypocarbia|Hypocarbia
C0364151|T201|DN|2019-8|LNC2HPO|Hypocarbia|Hypocarbia
C0364151|T201|LC|2019-8|LNC2HPO|Hypocarbia|Hypocarbia
C0364151|T201|OSN|2019-8|LNC2HPO|Hypocarbia|Hypocarbia
C0365091|T201|LN|2947-0|LNC2HPO|Hypernatremia|Hypernatremia
C0365091|T201|MTH_LN|2947-0|LNC2HPO|Hypernatremia|Hypernatremia
C0365091|T201|DN|2947-0|LNC2HPO|Hypernatremia|Hypernatremia
C0365091|T201|OSN|2947-0|LNC2HPO|Hypernatremia|Hypernatremia
C0365091|T201|LC|2947-0|LNC2HPO|Hypernatremia|Hypernatremia
C0365091|T201|LN|2947-0|LNC2HPO|Hyponatremia|Hyponatremia
C0365091|T201|MTH_LN|2947-0|LNC2HPO|Hyponatremia|Hyponatremia
C0365091|T201|DN|2947-0|LNC2HPO|Hyponatremia|Hyponatremia
C0365091|T201|OSN|2947-0|LNC2HPO|Hyponatremia|Hyponatremia
C0365091|T201|LC|2947-0|LNC2HPO|Hyponatremia|Hyponatremia
C0364411|T201|LC|2276-4|LNC2HPO|Hyperferritinaemia|Hyperferritinaemia
C0364411|T201|DN|2276-4|LNC2HPO|Hyperferritinaemia|Hyperferritinaemia
C0364411|T201|MTH_LN|2276-4|LNC2HPO|Hyperferritinaemia|Hyperferritinaemia
C0364411|T201|LN|2276-4|LNC2HPO|Hyperferritinaemia|Hyperferritinaemia
C0364411|T201|OSN|2276-4|LNC2HPO|Hyperferritinaemia|Hyperferritinaemia
C0364411|T201|LC|2276-4|LNC2HPO|Hyperferritinemia|Hyperferritinemia
C0364411|T201|DN|2276-4|LNC2HPO|Hyperferritinemia|Hyperferritinemia
C0364411|T201|MTH_LN|2276-4|LNC2HPO|Hyperferritinemia|Hyperferritinemia
C0364411|T201|LN|2276-4|LNC2HPO|Hyperferritinemia|Hyperferritinemia
C0364411|T201|OSN|2276-4|LNC2HPO|Hyperferritinemia|Hyperferritinemia
C0368042|T201|LN|5803-2|LNC2HPO|Acid base imbalance|Acid base imbalance
C0368042|T201|DN|5803-2|LNC2HPO|Acid base imbalance|Acid base imbalance
C0368042|T201|MTH_LN|5803-2|LNC2HPO|Acid base imbalance|Acid base imbalance
C0368042|T201|OSN|5803-2|LNC2HPO|Acid base imbalance|Acid base imbalance
C0368042|T201|LC|5803-2|LNC2HPO|Acid base imbalance|Acid base imbalance
C0368042|T201|LN|5803-2|LNC2HPO|Alkalemia|Alkalemia
C0368042|T201|DN|5803-2|LNC2HPO|Alkalemia|Alkalemia
C0368042|T201|MTH_LN|5803-2|LNC2HPO|Alkalemia|Alkalemia
C0368042|T201|OSN|5803-2|LNC2HPO|Alkalemia|Alkalemia
C0368042|T201|LC|5803-2|LNC2HPO|Alkalemia|Alkalemia
C0368042|T201|LN|5803-2|LNC2HPO|Acidemia|Acidemia
C0368042|T201|DN|5803-2|LNC2HPO|Acidemia|Acidemia
C0368042|T201|MTH_LN|5803-2|LNC2HPO|Acidemia|Acidemia
C0368042|T201|OSN|5803-2|LNC2HPO|Acidemia|Acidemia
C0368042|T201|LC|5803-2|LNC2HPO|Acidemia|Acidemia
C0364961|T201|LN|6298-4|LNC2HPO|Hyperkalemia|Hyperkalemia
C0364961|T201|MTH_LN|6298-4|LNC2HPO|Hyperkalemia|Hyperkalemia
C0364961|T201|DN|6298-4|LNC2HPO|Hyperkalemia|Hyperkalemia
C0364961|T201|OSN|6298-4|LNC2HPO|Hyperkalemia|Hyperkalemia
C0364961|T201|LC|6298-4|LNC2HPO|Hyperkalemia|Hyperkalemia
C0364961|T201|LN|6298-4|LNC2HPO|Hypokalemia|Hypokalemia
C0364961|T201|MTH_LN|6298-4|LNC2HPO|Hypokalemia|Hypokalemia
C0364961|T201|DN|6298-4|LNC2HPO|Hypokalemia|Hypokalemia
C0364961|T201|OSN|6298-4|LNC2HPO|Hypokalemia|Hypokalemia
C0364961|T201|LC|6298-4|LNC2HPO|Hypokalemia|Hypokalemia
C0550239|T201|LN|12180-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0550239|T201|DN|12180-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0550239|T201|MTH_LN|12180-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0550239|T201|OSN|12180-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0550239|T201|LC|12180-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0550239|T201|LN|12180-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0550239|T201|DN|12180-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0550239|T201|MTH_LN|12180-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0550239|T201|OSN|12180-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0550239|T201|LC|12180-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0550239|T201|LN|12180-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0550239|T201|DN|12180-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0550239|T201|MTH_LN|12180-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0550239|T201|OSN|12180-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0550239|T201|LC|12180-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0550239|T201|LN|12180-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0550239|T201|DN|12180-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0550239|T201|MTH_LN|12180-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0550239|T201|OSN|12180-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0550239|T201|LC|12180-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0550242|T201|LN|13444-5|LNC2HPO|Hypercalcemia|Hypercalcemia
C0550242|T201|OSN|13444-5|LNC2HPO|Hypercalcemia|Hypercalcemia
C0550242|T201|MTH_LN|13444-5|LNC2HPO|Hypercalcemia|Hypercalcemia
C0550242|T201|DN|13444-5|LNC2HPO|Hypercalcemia|Hypercalcemia
C0550242|T201|LC|13444-5|LNC2HPO|Hypercalcemia|Hypercalcemia
C0550242|T201|LN|13444-5|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0550242|T201|OSN|13444-5|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0550242|T201|MTH_LN|13444-5|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0550242|T201|DN|13444-5|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0550242|T201|LC|13444-5|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0550242|T201|LN|13444-5|LNC2HPO|Hypocalcemia|Hypocalcemia
C0550242|T201|OSN|13444-5|LNC2HPO|Hypocalcemia|Hypocalcemia
C0550242|T201|MTH_LN|13444-5|LNC2HPO|Hypocalcemia|Hypocalcemia
C0550242|T201|DN|13444-5|LNC2HPO|Hypocalcemia|Hypocalcemia
C0550242|T201|LC|13444-5|LNC2HPO|Hypocalcemia|Hypocalcemia
C0550242|T201|LN|13444-5|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0550242|T201|OSN|13444-5|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0550242|T201|MTH_LN|13444-5|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0550242|T201|DN|13444-5|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0550242|T201|LC|13444-5|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0797147|T201|LN|13959-2|LNC2HPO|Hypercalcemia|Hypercalcemia
C0797147|T201|DN|13959-2|LNC2HPO|Hypercalcemia|Hypercalcemia
C0797147|T201|MTH_LN|13959-2|LNC2HPO|Hypercalcemia|Hypercalcemia
C0797147|T201|OSN|13959-2|LNC2HPO|Hypercalcemia|Hypercalcemia
C0797147|T201|LC|13959-2|LNC2HPO|Hypercalcemia|Hypercalcemia
C0797147|T201|LN|13959-2|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0797147|T201|DN|13959-2|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0797147|T201|MTH_LN|13959-2|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0797147|T201|OSN|13959-2|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0797147|T201|LC|13959-2|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0797147|T201|LN|13959-2|LNC2HPO|Hypocalcemia|Hypocalcemia
C0797147|T201|DN|13959-2|LNC2HPO|Hypocalcemia|Hypocalcemia
C0797147|T201|MTH_LN|13959-2|LNC2HPO|Hypocalcemia|Hypocalcemia
C0797147|T201|OSN|13959-2|LNC2HPO|Hypocalcemia|Hypocalcemia
C0797147|T201|LC|13959-2|LNC2HPO|Hypocalcemia|Hypocalcemia
C0797147|T201|LN|13959-2|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0797147|T201|DN|13959-2|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0797147|T201|MTH_LN|13959-2|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0797147|T201|OSN|13959-2|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0797147|T201|LC|13959-2|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0799677|T201|LN|16526-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0799677|T201|MTH_LN|16526-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0799677|T201|OSN|16526-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0799677|T201|DN|16526-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0799677|T201|LC|16526-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0799677|T201|LN|16526-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0799677|T201|MTH_LN|16526-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0799677|T201|OSN|16526-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0799677|T201|DN|16526-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0799677|T201|LC|16526-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0799677|T201|LN|16526-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0799677|T201|MTH_LN|16526-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0799677|T201|OSN|16526-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0799677|T201|DN|16526-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0799677|T201|LC|16526-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0799677|T201|LN|16526-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0799677|T201|MTH_LN|16526-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0799677|T201|OSN|16526-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0799677|T201|DN|16526-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0799677|T201|LC|16526-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0800970|T201|LC|17863-2|LNC2HPO|Hypercalcemia|Hypercalcemia
C0800970|T201|DN|17863-2|LNC2HPO|Hypercalcemia|Hypercalcemia
C0800970|T201|MTH_LN|17863-2|LNC2HPO|Hypercalcemia|Hypercalcemia
C0800970|T201|LN|17863-2|LNC2HPO|Hypercalcemia|Hypercalcemia
C0800970|T201|OSN|17863-2|LNC2HPO|Hypercalcemia|Hypercalcemia
C0800970|T201|LC|17863-2|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0800970|T201|DN|17863-2|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0800970|T201|MTH_LN|17863-2|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0800970|T201|LN|17863-2|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0800970|T201|OSN|17863-2|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0800970|T201|LC|17863-2|LNC2HPO|Hypocalcemia|Hypocalcemia
C0800970|T201|DN|17863-2|LNC2HPO|Hypocalcemia|Hypocalcemia
C0800970|T201|MTH_LN|17863-2|LNC2HPO|Hypocalcemia|Hypocalcemia
C0800970|T201|LN|17863-2|LNC2HPO|Hypocalcemia|Hypocalcemia
C0800970|T201|OSN|17863-2|LNC2HPO|Hypocalcemia|Hypocalcemia
C0800970|T201|LC|17863-2|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0800970|T201|DN|17863-2|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0800970|T201|MTH_LN|17863-2|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0800970|T201|LN|17863-2|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0800970|T201|OSN|17863-2|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0801327|T201|LN|18281-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0801327|T201|DN|18281-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0801327|T201|MTH_LN|18281-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0801327|T201|OSN|18281-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0801327|T201|LC|18281-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0801327|T201|LN|18281-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0801327|T201|DN|18281-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0801327|T201|MTH_LN|18281-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0801327|T201|OSN|18281-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0801327|T201|LC|18281-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0801327|T201|LN|18281-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0801327|T201|DN|18281-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0801327|T201|MTH_LN|18281-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0801327|T201|OSN|18281-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0801327|T201|LC|18281-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0801327|T201|LN|18281-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0801327|T201|DN|18281-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0801327|T201|MTH_LN|18281-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0801327|T201|OSN|18281-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0801327|T201|LC|18281-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0812462|T201|LN|19072-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C0812462|T201|DN|19072-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C0812462|T201|MTH_LN|19072-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C0812462|T201|OSN|19072-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C0812462|T201|LC|19072-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C0812462|T201|LN|19072-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0812462|T201|DN|19072-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0812462|T201|MTH_LN|19072-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0812462|T201|OSN|19072-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0812462|T201|LC|19072-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0812462|T201|LN|19072-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C0812462|T201|DN|19072-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C0812462|T201|MTH_LN|19072-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C0812462|T201|OSN|19072-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C0812462|T201|LC|19072-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C0812462|T201|LN|19072-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0812462|T201|DN|19072-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0812462|T201|MTH_LN|19072-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0812462|T201|OSN|19072-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0812462|T201|LC|19072-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364129|T201|LN|1996-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C0364129|T201|MTH_LN|1996-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C0364129|T201|DN|1996-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C0364129|T201|OSN|1996-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C0364129|T201|LC|1996-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C0364129|T201|LN|1996-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0364129|T201|MTH_LN|1996-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0364129|T201|DN|1996-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0364129|T201|OSN|1996-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0364129|T201|LC|1996-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0364129|T201|LN|1996-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C0364129|T201|MTH_LN|1996-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C0364129|T201|DN|1996-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C0364129|T201|OSN|1996-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C0364129|T201|LC|1996-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C0364129|T201|LN|1996-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364129|T201|MTH_LN|1996-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364129|T201|DN|1996-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364129|T201|OSN|1996-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364129|T201|LC|1996-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1507674|T201|LN|38230-9|LNC2HPO|Hypercalcemia|Hypercalcemia
C1507674|T201|DN|38230-9|LNC2HPO|Hypercalcemia|Hypercalcemia
C1507674|T201|OSN|38230-9|LNC2HPO|Hypercalcemia|Hypercalcemia
C1507674|T201|MTH_LN|38230-9|LNC2HPO|Hypercalcemia|Hypercalcemia
C1507674|T201|LC|38230-9|LNC2HPO|Hypercalcemia|Hypercalcemia
C1507674|T201|LN|38230-9|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1507674|T201|DN|38230-9|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1507674|T201|OSN|38230-9|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1507674|T201|MTH_LN|38230-9|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1507674|T201|LC|38230-9|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1507674|T201|LN|38230-9|LNC2HPO|Hypocalcemia|Hypocalcemia
C1507674|T201|DN|38230-9|LNC2HPO|Hypocalcemia|Hypocalcemia
C1507674|T201|OSN|38230-9|LNC2HPO|Hypocalcemia|Hypocalcemia
C1507674|T201|MTH_LN|38230-9|LNC2HPO|Hypocalcemia|Hypocalcemia
C1507674|T201|LC|38230-9|LNC2HPO|Hypocalcemia|Hypocalcemia
C1507674|T201|LN|38230-9|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1507674|T201|DN|38230-9|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1507674|T201|OSN|38230-9|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1507674|T201|MTH_LN|38230-9|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1507674|T201|LC|38230-9|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1642581|T201|LN|41644-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C1642581|T201|DN|41644-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C1642581|T201|OSN|41644-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C1642581|T201|MTH_LN|41644-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C1642581|T201|LC|41644-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C1642581|T201|LN|41644-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1642581|T201|DN|41644-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1642581|T201|OSN|41644-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1642581|T201|MTH_LN|41644-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1642581|T201|LC|41644-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1642581|T201|LN|41644-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C1642581|T201|DN|41644-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C1642581|T201|OSN|41644-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C1642581|T201|MTH_LN|41644-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C1642581|T201|LC|41644-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C1642581|T201|LN|41644-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1642581|T201|DN|41644-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1642581|T201|OSN|41644-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1642581|T201|MTH_LN|41644-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1642581|T201|LC|41644-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1651491|T201|LN|41645-3|LNC2HPO|Hypercalcemia|Hypercalcemia
C1651491|T201|DN|41645-3|LNC2HPO|Hypercalcemia|Hypercalcemia
C1651491|T201|OSN|41645-3|LNC2HPO|Hypercalcemia|Hypercalcemia
C1651491|T201|MTH_LN|41645-3|LNC2HPO|Hypercalcemia|Hypercalcemia
C1651491|T201|LC|41645-3|LNC2HPO|Hypercalcemia|Hypercalcemia
C1651491|T201|LN|41645-3|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1651491|T201|DN|41645-3|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1651491|T201|OSN|41645-3|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1651491|T201|MTH_LN|41645-3|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1651491|T201|LC|41645-3|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1651491|T201|LN|41645-3|LNC2HPO|Hypocalcemia|Hypocalcemia
C1651491|T201|DN|41645-3|LNC2HPO|Hypocalcemia|Hypocalcemia
C1651491|T201|OSN|41645-3|LNC2HPO|Hypocalcemia|Hypocalcemia
C1651491|T201|MTH_LN|41645-3|LNC2HPO|Hypocalcemia|Hypocalcemia
C1651491|T201|LC|41645-3|LNC2HPO|Hypocalcemia|Hypocalcemia
C1651491|T201|LN|41645-3|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1651491|T201|DN|41645-3|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1651491|T201|OSN|41645-3|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1651491|T201|MTH_LN|41645-3|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1651491|T201|LC|41645-3|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1641514|T201|LN|41646-1|LNC2HPO|Hypercalcemia|Hypercalcemia
C1641514|T201|DN|41646-1|LNC2HPO|Hypercalcemia|Hypercalcemia
C1641514|T201|OSN|41646-1|LNC2HPO|Hypercalcemia|Hypercalcemia
C1641514|T201|MTH_LN|41646-1|LNC2HPO|Hypercalcemia|Hypercalcemia
C1641514|T201|LC|41646-1|LNC2HPO|Hypercalcemia|Hypercalcemia
C1641514|T201|LN|41646-1|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1641514|T201|DN|41646-1|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1641514|T201|OSN|41646-1|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1641514|T201|MTH_LN|41646-1|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1641514|T201|LC|41646-1|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1641514|T201|LN|41646-1|LNC2HPO|Hypocalcemia|Hypocalcemia
C1641514|T201|DN|41646-1|LNC2HPO|Hypocalcemia|Hypocalcemia
C1641514|T201|OSN|41646-1|LNC2HPO|Hypocalcemia|Hypocalcemia
C1641514|T201|MTH_LN|41646-1|LNC2HPO|Hypocalcemia|Hypocalcemia
C1641514|T201|LC|41646-1|LNC2HPO|Hypocalcemia|Hypocalcemia
C1641514|T201|LN|41646-1|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1641514|T201|DN|41646-1|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1641514|T201|OSN|41646-1|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1641514|T201|MTH_LN|41646-1|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1641514|T201|LC|41646-1|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C5201128|T201|LC|42567-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C5201128|T201|DN|42567-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C5201128|T201|MTH_LN|42567-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C5201128|T201|OSN|42567-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C5201128|T201|LN|42567-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C5201128|T201|LC|42567-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C5201128|T201|DN|42567-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C5201128|T201|MTH_LN|42567-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C5201128|T201|OSN|42567-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C5201128|T201|LN|42567-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C5201128|T201|LC|42567-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C5201128|T201|DN|42567-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C5201128|T201|MTH_LN|42567-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C5201128|T201|OSN|42567-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C5201128|T201|LN|42567-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C5201128|T201|LC|42567-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C5201128|T201|DN|42567-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C5201128|T201|MTH_LN|42567-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C5201128|T201|OSN|42567-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C5201128|T201|LN|42567-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1639938|T201|LN|42593-4|LNC2HPO|Hypercalcemia|Hypercalcemia
C1639938|T201|DN|42593-4|LNC2HPO|Hypercalcemia|Hypercalcemia
C1639938|T201|OSN|42593-4|LNC2HPO|Hypercalcemia|Hypercalcemia
C1639938|T201|MTH_LN|42593-4|LNC2HPO|Hypercalcemia|Hypercalcemia
C1639938|T201|LC|42593-4|LNC2HPO|Hypercalcemia|Hypercalcemia
C1639938|T201|LN|42593-4|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1639938|T201|DN|42593-4|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1639938|T201|OSN|42593-4|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1639938|T201|MTH_LN|42593-4|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1639938|T201|LC|42593-4|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1639938|T201|LN|42593-4|LNC2HPO|Hypocalcemia|Hypocalcemia
C1639938|T201|DN|42593-4|LNC2HPO|Hypocalcemia|Hypocalcemia
C1639938|T201|OSN|42593-4|LNC2HPO|Hypocalcemia|Hypocalcemia
C1639938|T201|MTH_LN|42593-4|LNC2HPO|Hypocalcemia|Hypocalcemia
C1639938|T201|LC|42593-4|LNC2HPO|Hypocalcemia|Hypocalcemia
C1639938|T201|LN|42593-4|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1639938|T201|DN|42593-4|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1639938|T201|OSN|42593-4|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1639938|T201|MTH_LN|42593-4|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1639938|T201|LC|42593-4|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1633476|T201|LN|42857-3|LNC2HPO|Hypercalcemia|Hypercalcemia
C1633476|T201|DN|42857-3|LNC2HPO|Hypercalcemia|Hypercalcemia
C1633476|T201|OSN|42857-3|LNC2HPO|Hypercalcemia|Hypercalcemia
C1633476|T201|MTH_LN|42857-3|LNC2HPO|Hypercalcemia|Hypercalcemia
C1633476|T201|LC|42857-3|LNC2HPO|Hypercalcemia|Hypercalcemia
C1633476|T201|LN|42857-3|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1633476|T201|DN|42857-3|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1633476|T201|OSN|42857-3|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1633476|T201|MTH_LN|42857-3|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1633476|T201|LC|42857-3|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1633476|T201|LN|42857-3|LNC2HPO|Hypocalcemia|Hypocalcemia
C1633476|T201|DN|42857-3|LNC2HPO|Hypocalcemia|Hypocalcemia
C1633476|T201|OSN|42857-3|LNC2HPO|Hypocalcemia|Hypocalcemia
C1633476|T201|MTH_LN|42857-3|LNC2HPO|Hypocalcemia|Hypocalcemia
C1633476|T201|LC|42857-3|LNC2HPO|Hypocalcemia|Hypocalcemia
C1633476|T201|LN|42857-3|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1633476|T201|DN|42857-3|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1633476|T201|OSN|42857-3|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1633476|T201|MTH_LN|42857-3|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1633476|T201|LC|42857-3|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1717133|T201|LN|46099-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C1717133|T201|DN|46099-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C1717133|T201|OSN|46099-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C1717133|T201|MTH_LN|46099-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C1717133|T201|LC|46099-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C1717133|T201|LN|46099-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1717133|T201|DN|46099-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1717133|T201|OSN|46099-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1717133|T201|MTH_LN|46099-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1717133|T201|LC|46099-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1717133|T201|LN|46099-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C1717133|T201|DN|46099-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C1717133|T201|OSN|46099-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C1717133|T201|MTH_LN|46099-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C1717133|T201|LC|46099-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C1717133|T201|LN|46099-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1717133|T201|DN|46099-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1717133|T201|OSN|46099-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1717133|T201|MTH_LN|46099-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1717133|T201|LC|46099-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1952827|T201|LN|47596-2|LNC2HPO|Hypercalcemia|Hypercalcemia
C1952827|T201|DN|47596-2|LNC2HPO|Hypercalcemia|Hypercalcemia
C1952827|T201|OSN|47596-2|LNC2HPO|Hypercalcemia|Hypercalcemia
C1952827|T201|MTH_LN|47596-2|LNC2HPO|Hypercalcemia|Hypercalcemia
C1952827|T201|LC|47596-2|LNC2HPO|Hypercalcemia|Hypercalcemia
C1952827|T201|LN|47596-2|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1952827|T201|DN|47596-2|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1952827|T201|OSN|47596-2|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1952827|T201|MTH_LN|47596-2|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1952827|T201|LC|47596-2|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1952827|T201|LN|47596-2|LNC2HPO|Hypocalcemia|Hypocalcemia
C1952827|T201|DN|47596-2|LNC2HPO|Hypocalcemia|Hypocalcemia
C1952827|T201|OSN|47596-2|LNC2HPO|Hypocalcemia|Hypocalcemia
C1952827|T201|MTH_LN|47596-2|LNC2HPO|Hypocalcemia|Hypocalcemia
C1952827|T201|LC|47596-2|LNC2HPO|Hypocalcemia|Hypocalcemia
C1952827|T201|LN|47596-2|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1952827|T201|DN|47596-2|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1952827|T201|OSN|47596-2|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1952827|T201|MTH_LN|47596-2|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1952827|T201|LC|47596-2|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1952828|T201|LN|47597-0|LNC2HPO|Hypercalcemia|Hypercalcemia
C1952828|T201|DN|47597-0|LNC2HPO|Hypercalcemia|Hypercalcemia
C1952828|T201|OSN|47597-0|LNC2HPO|Hypercalcemia|Hypercalcemia
C1952828|T201|MTH_LN|47597-0|LNC2HPO|Hypercalcemia|Hypercalcemia
C1952828|T201|LC|47597-0|LNC2HPO|Hypercalcemia|Hypercalcemia
C1952828|T201|LN|47597-0|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1952828|T201|DN|47597-0|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1952828|T201|OSN|47597-0|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1952828|T201|MTH_LN|47597-0|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1952828|T201|LC|47597-0|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1952828|T201|LN|47597-0|LNC2HPO|Hypocalcemia|Hypocalcemia
C1952828|T201|DN|47597-0|LNC2HPO|Hypocalcemia|Hypocalcemia
C1952828|T201|OSN|47597-0|LNC2HPO|Hypocalcemia|Hypocalcemia
C1952828|T201|MTH_LN|47597-0|LNC2HPO|Hypocalcemia|Hypocalcemia
C1952828|T201|LC|47597-0|LNC2HPO|Hypocalcemia|Hypocalcemia
C1952828|T201|LN|47597-0|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1952828|T201|DN|47597-0|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1952828|T201|OSN|47597-0|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1952828|T201|MTH_LN|47597-0|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1952828|T201|LC|47597-0|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1952829|T201|LN|47598-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C1952829|T201|DN|47598-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C1952829|T201|OSN|47598-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C1952829|T201|MTH_LN|47598-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C1952829|T201|LC|47598-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C1952829|T201|LN|47598-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1952829|T201|DN|47598-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1952829|T201|OSN|47598-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1952829|T201|MTH_LN|47598-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1952829|T201|LC|47598-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1952829|T201|LN|47598-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C1952829|T201|DN|47598-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C1952829|T201|OSN|47598-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C1952829|T201|MTH_LN|47598-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C1952829|T201|LC|47598-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C1952829|T201|LN|47598-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1952829|T201|DN|47598-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1952829|T201|OSN|47598-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1952829|T201|MTH_LN|47598-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1952829|T201|LC|47598-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1977516|T201|LN|49765-1|LNC2HPO|Hypercalcemia|Hypercalcemia
C1977516|T201|DN|49765-1|LNC2HPO|Hypercalcemia|Hypercalcemia
C1977516|T201|MTH_LN|49765-1|LNC2HPO|Hypercalcemia|Hypercalcemia
C1977516|T201|OSN|49765-1|LNC2HPO|Hypercalcemia|Hypercalcemia
C1977516|T201|LC|49765-1|LNC2HPO|Hypercalcemia|Hypercalcemia
C1977516|T201|LN|49765-1|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1977516|T201|DN|49765-1|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1977516|T201|MTH_LN|49765-1|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1977516|T201|OSN|49765-1|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1977516|T201|LC|49765-1|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C1977516|T201|LN|49765-1|LNC2HPO|Hypocalcemia|Hypocalcemia
C1977516|T201|DN|49765-1|LNC2HPO|Hypocalcemia|Hypocalcemia
C1977516|T201|MTH_LN|49765-1|LNC2HPO|Hypocalcemia|Hypocalcemia
C1977516|T201|OSN|49765-1|LNC2HPO|Hypocalcemia|Hypocalcemia
C1977516|T201|LC|49765-1|LNC2HPO|Hypocalcemia|Hypocalcemia
C1977516|T201|LN|49765-1|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1977516|T201|DN|49765-1|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1977516|T201|MTH_LN|49765-1|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1977516|T201|OSN|49765-1|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C1977516|T201|LC|49765-1|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364264|T201|LC|2132-9|LNC2HPO|Vitamin B12 deficiency|Vitamin B12 deficiency
C0364264|T201|MTH_LN|2132-9|LNC2HPO|Vitamin B12 deficiency|Vitamin B12 deficiency
C0364264|T201|OSN|2132-9|LNC2HPO|Vitamin B12 deficiency|Vitamin B12 deficiency
C0364264|T201|LN|2132-9|LNC2HPO|Vitamin B12 deficiency|Vitamin B12 deficiency
C0364264|T201|DN|2132-9|LNC2HPO|Vitamin B12 deficiency|Vitamin B12 deficiency
C0803222|T201|LN|20407-3|LNC2HPO|Nitrituria|Nitrituria
C0803222|T201|MTH_LN|20407-3|LNC2HPO|Nitrituria|Nitrituria
C0803222|T201|DN|20407-3|LNC2HPO|Nitrituria|Nitrituria
C0803222|T201|OSN|20407-3|LNC2HPO|Nitrituria|Nitrituria
C0803222|T201|LC|20407-3|LNC2HPO|Nitrituria|Nitrituria
C1315181|T201|LN|32710-6|LNC2HPO|Nitrituria|Nitrituria
C1315181|T201|MTH_LN|32710-6|LNC2HPO|Nitrituria|Nitrituria
C1315181|T201|DN|32710-6|LNC2HPO|Nitrituria|Nitrituria
C1315181|T201|OSN|32710-6|LNC2HPO|Nitrituria|Nitrituria
C1315181|T201|LC|32710-6|LNC2HPO|Nitrituria|Nitrituria
C0364802|T201|LN|2657-5|LNC2HPO|Nitrituria|Nitrituria
C0364802|T201|MTH_LN|2657-5|LNC2HPO|Nitrituria|Nitrituria
C0364802|T201|DN|2657-5|LNC2HPO|Nitrituria|Nitrituria
C0364802|T201|OSN|2657-5|LNC2HPO|Nitrituria|Nitrituria
C0364802|T201|LC|2657-5|LNC2HPO|Nitrituria|Nitrituria
C1978485|T201|LN|50558-6|LNC2HPO|Nitrituria|Nitrituria
C1978485|T201|MTH_LN|50558-6|LNC2HPO|Nitrituria|Nitrituria
C1978485|T201|DN|50558-6|LNC2HPO|Nitrituria|Nitrituria
C1978485|T201|OSN|50558-6|LNC2HPO|Nitrituria|Nitrituria
C1978485|T201|LC|50558-6|LNC2HPO|Nitrituria|Nitrituria
C0368040|T201|LN|5802-4|LNC2HPO|Nitrituria|Nitrituria
C0368040|T201|MTH_LN|5802-4|LNC2HPO|Nitrituria|Nitrituria
C0368040|T201|DN|5802-4|LNC2HPO|Nitrituria|Nitrituria
C0368040|T201|OSN|5802-4|LNC2HPO|Nitrituria|Nitrituria
C0368040|T201|LC|5802-4|LNC2HPO|Nitrituria|Nitrituria
C1114065|T201|LN|30180-4|LNC2HPO|Basophilia|Basophilia
C1114065|T201|OSN|30180-4|LNC2HPO|Basophilia|Basophilia
C1114065|T201|DN|30180-4|LNC2HPO|Basophilia|Basophilia
C1114065|T201|MTH_LN|30180-4|LNC2HPO|Basophilia|Basophilia
C1114065|T201|LC|30180-4|LNC2HPO|Basophilia|Basophilia
C0798323|T201|LN|15152-2|LNC2HPO|Conjugated hyperbilirubinemia|Conjugated hyperbilirubinemia
C0798323|T201|DN|15152-2|LNC2HPO|Conjugated hyperbilirubinemia|Conjugated hyperbilirubinemia
C0798323|T201|MTH_LN|15152-2|LNC2HPO|Conjugated hyperbilirubinemia|Conjugated hyperbilirubinemia
C0798323|T201|OSN|15152-2|LNC2HPO|Conjugated hyperbilirubinemia|Conjugated hyperbilirubinemia
C0798323|T201|LC|15152-2|LNC2HPO|Conjugated hyperbilirubinemia|Conjugated hyperbilirubinemia
C0798323|T201|LN|15152-2|LNC2HPO|Direct hyperbilirubinemia|Direct hyperbilirubinemia
C0798323|T201|DN|15152-2|LNC2HPO|Direct hyperbilirubinemia|Direct hyperbilirubinemia
C0798323|T201|MTH_LN|15152-2|LNC2HPO|Direct hyperbilirubinemia|Direct hyperbilirubinemia
C0798323|T201|OSN|15152-2|LNC2HPO|Direct hyperbilirubinemia|Direct hyperbilirubinemia
C0798323|T201|LC|15152-2|LNC2HPO|Direct hyperbilirubinemia|Direct hyperbilirubinemia
C0942414|T201|LN|26444-0|LNC2HPO|Basophilia|Basophilia
C0942414|T201|DN|26444-0|LNC2HPO|Basophilia|Basophilia
C0942414|T201|OSN|26444-0|LNC2HPO|Basophilia|Basophilia
C0942414|T201|MTH_LN|26444-0|LNC2HPO|Basophilia|Basophilia
C0942414|T201|LC|26444-0|LNC2HPO|Basophilia|Basophilia
C0367985|T201|LN|5770-3|LNC2HPO|Bilirubinuria|Bilirubinuria
C0367985|T201|LC|5770-3|LNC2HPO|Bilirubinuria|Bilirubinuria
C0367985|T201|MTH_LN|5770-3|LNC2HPO|Bilirubinuria|Bilirubinuria
C0367985|T201|DN|5770-3|LNC2HPO|Bilirubinuria|Bilirubinuria
C0367985|T201|OSN|5770-3|LNC2HPO|Bilirubinuria|Bilirubinuria
C2607829|T201|LC|35209-6|LNC2HPO|Hyperferritinaemia|Hyperferritinaemia
C2607829|T201|DN|35209-6|LNC2HPO|Hyperferritinaemia|Hyperferritinaemia
C2607829|T201|MTH_LN|35209-6|LNC2HPO|Hyperferritinaemia|Hyperferritinaemia
C2607829|T201|LN|35209-6|LNC2HPO|Hyperferritinaemia|Hyperferritinaemia
C2607829|T201|OSN|35209-6|LNC2HPO|Hyperferritinaemia|Hyperferritinaemia
C2607829|T201|LC|35209-6|LNC2HPO|Hyperferritinemia|Hyperferritinemia
C2607829|T201|DN|35209-6|LNC2HPO|Hyperferritinemia|Hyperferritinemia
C2607829|T201|MTH_LN|35209-6|LNC2HPO|Hyperferritinemia|Hyperferritinemia
C2607829|T201|LN|35209-6|LNC2HPO|Hyperferritinemia|Hyperferritinemia
C2607829|T201|OSN|35209-6|LNC2HPO|Hyperferritinemia|Hyperferritinemia
C0803376|T201|LN|20567-4|LNC2HPO|Hyperferritinaemia|Hyperferritinaemia
C0803376|T201|OSN|20567-4|LNC2HPO|Hyperferritinaemia|Hyperferritinaemia
C0803376|T201|DN|20567-4|LNC2HPO|Hyperferritinaemia|Hyperferritinaemia
C0803376|T201|MTH_LN|20567-4|LNC2HPO|Hyperferritinaemia|Hyperferritinaemia
C0803376|T201|LC|20567-4|LNC2HPO|Hyperferritinaemia|Hyperferritinaemia
C0803376|T201|LN|20567-4|LNC2HPO|Hyperferritinemia|Hyperferritinemia
C0803376|T201|OSN|20567-4|LNC2HPO|Hyperferritinemia|Hyperferritinemia
C0803376|T201|DN|20567-4|LNC2HPO|Hyperferritinemia|Hyperferritinemia
C0803376|T201|MTH_LN|20567-4|LNC2HPO|Hyperferritinemia|Hyperferritinemia
C0803376|T201|LC|20567-4|LNC2HPO|Hyperferritinemia|Hyperferritinemia
C1978478|T201|LN|50551-1|LNC2HPO|Bilirubinuria|Bilirubinuria
C1978478|T201|LC|50551-1|LNC2HPO|Bilirubinuria|Bilirubinuria
C1978478|T201|MTH_LN|50551-1|LNC2HPO|Bilirubinuria|Bilirubinuria
C1978478|T201|DN|50551-1|LNC2HPO|Bilirubinuria|Bilirubinuria
C1978478|T201|OSN|50551-1|LNC2HPO|Bilirubinuria|Bilirubinuria
C0364110|T201|LN|1977-8|LNC2HPO|Bilirubinuria|Bilirubinuria
C0364110|T201|LC|1977-8|LNC2HPO|Bilirubinuria|Bilirubinuria
C0364110|T201|MTH_LN|1977-8|LNC2HPO|Bilirubinuria|Bilirubinuria
C0364110|T201|DN|1977-8|LNC2HPO|Bilirubinuria|Bilirubinuria
C0364110|T201|OSN|1977-8|LNC2HPO|Bilirubinuria|Bilirubinuria
C1715313|T201|LN|44033-9|LNC2HPO|Bilirubinuria|Bilirubinuria
C1715313|T201|LC|44033-9|LNC2HPO|Bilirubinuria|Bilirubinuria
C1715313|T201|MTH_LN|44033-9|LNC2HPO|Bilirubinuria|Bilirubinuria
C1715313|T201|DN|44033-9|LNC2HPO|Bilirubinuria|Bilirubinuria
C1715313|T201|OSN|44033-9|LNC2HPO|Bilirubinuria|Bilirubinuria
C0365032|T201|LN|2888-6|LNC2HPO|Proteinuria|Proteinuria
C0365032|T201|MTH_LN|2888-6|LNC2HPO|Proteinuria|Proteinuria
C0365032|T201|DN|2888-6|LNC2HPO|Proteinuria|Proteinuria
C0365032|T201|OSN|2888-6|LNC2HPO|Proteinuria|Proteinuria
C0365032|T201|LC|2888-6|LNC2HPO|Proteinuria|Proteinuria
C0550834|T201|LN|11151-8|LNC2HPO|Reticulocytosis|Reticulocytosis
C0550834|T201|DN|11151-8|LNC2HPO|Reticulocytosis|Reticulocytosis
C0550834|T201|MTH_LN|11151-8|LNC2HPO|Reticulocytosis|Reticulocytosis
C0550834|T201|LC|11151-8|LNC2HPO|Reticulocytosis|Reticulocytosis
C0550834|T201|OSN|11151-8|LNC2HPO|Reticulocytosis|Reticulocytosis
C0550834|T201|LN|11151-8|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0550834|T201|DN|11151-8|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0550834|T201|MTH_LN|11151-8|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0550834|T201|LC|11151-8|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0550834|T201|OSN|11151-8|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0550836|T201|LN|11153-4|LNC2HPO|Reticulocytosis|Reticulocytosis
C0550836|T201|DN|11153-4|LNC2HPO|Reticulocytosis|Reticulocytosis
C0550836|T201|MTH_LN|11153-4|LNC2HPO|Reticulocytosis|Reticulocytosis
C0550836|T201|LC|11153-4|LNC2HPO|Reticulocytosis|Reticulocytosis
C0550836|T201|OSN|11153-4|LNC2HPO|Reticulocytosis|Reticulocytosis
C0550836|T201|LN|11153-4|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0550836|T201|DN|11153-4|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0550836|T201|MTH_LN|11153-4|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0550836|T201|LC|11153-4|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0550836|T201|OSN|11153-4|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0550835|T201|LN|11271-4|LNC2HPO|Reticulocytosis|Reticulocytosis
C0550835|T201|DN|11271-4|LNC2HPO|Reticulocytosis|Reticulocytosis
C0550835|T201|MTH_LN|11271-4|LNC2HPO|Reticulocytosis|Reticulocytosis
C0550835|T201|LC|11271-4|LNC2HPO|Reticulocytosis|Reticulocytosis
C0550835|T201|OSN|11271-4|LNC2HPO|Reticulocytosis|Reticulocytosis
C0550835|T201|LN|11271-4|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0550835|T201|DN|11271-4|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0550835|T201|MTH_LN|11271-4|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0550835|T201|LC|11271-4|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0550835|T201|OSN|11271-4|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0549854|T201|LN|12250-7|LNC2HPO|Reticulocytosis|Reticulocytosis
C0549854|T201|DN|12250-7|LNC2HPO|Reticulocytosis|Reticulocytosis
C0549854|T201|OSN|12250-7|LNC2HPO|Reticulocytosis|Reticulocytosis
C0549854|T201|LC|12250-7|LNC2HPO|Reticulocytosis|Reticulocytosis
C0549854|T201|MTH_LN|12250-7|LNC2HPO|Reticulocytosis|Reticulocytosis
C0549854|T201|LN|12250-7|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0549854|T201|DN|12250-7|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0549854|T201|OSN|12250-7|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0549854|T201|LC|12250-7|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0549854|T201|MTH_LN|12250-7|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0796702|T201|LN|13508-7|LNC2HPO|Reticulocytosis|Reticulocytosis
C0796702|T201|DN|13508-7|LNC2HPO|Reticulocytosis|Reticulocytosis
C0796702|T201|MTH_LN|13508-7|LNC2HPO|Reticulocytosis|Reticulocytosis
C0796702|T201|LC|13508-7|LNC2HPO|Reticulocytosis|Reticulocytosis
C0796702|T201|OSN|13508-7|LNC2HPO|Reticulocytosis|Reticulocytosis
C0796702|T201|LN|13508-7|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0796702|T201|DN|13508-7|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0796702|T201|MTH_LN|13508-7|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0796702|T201|LC|13508-7|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0796702|T201|OSN|13508-7|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0797381|T201|LN|14196-0|LNC2HPO|Reticulocytosis|Reticulocytosis
C0797381|T201|DN|14196-0|LNC2HPO|Reticulocytosis|Reticulocytosis
C0797381|T201|OSN|14196-0|LNC2HPO|Reticulocytosis|Reticulocytosis
C0797381|T201|MTH_LN|14196-0|LNC2HPO|Reticulocytosis|Reticulocytosis
C0797381|T201|LC|14196-0|LNC2HPO|Reticulocytosis|Reticulocytosis
C0797381|T201|LN|14196-0|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0797381|T201|DN|14196-0|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0797381|T201|OSN|14196-0|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0797381|T201|MTH_LN|14196-0|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0797381|T201|LC|14196-0|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0800955|T201|LN|17848-3|LNC2HPO|Reticulocytosis|Reticulocytosis
C0800955|T201|DN|17848-3|LNC2HPO|Reticulocytosis|Reticulocytosis
C0800955|T201|OSN|17848-3|LNC2HPO|Reticulocytosis|Reticulocytosis
C0800955|T201|LC|17848-3|LNC2HPO|Reticulocytosis|Reticulocytosis
C0800955|T201|MTH_LN|17848-3|LNC2HPO|Reticulocytosis|Reticulocytosis
C0800955|T201|LN|17848-3|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0800955|T201|DN|17848-3|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0800955|T201|OSN|17848-3|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0800955|T201|LC|17848-3|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0800955|T201|MTH_LN|17848-3|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0800956|T201|LN|17849-1|LNC2HPO|Reticulocytosis|Reticulocytosis
C0800956|T201|DN|17849-1|LNC2HPO|Reticulocytosis|Reticulocytosis
C0800956|T201|MTH_LN|17849-1|LNC2HPO|Reticulocytosis|Reticulocytosis
C0800956|T201|OSN|17849-1|LNC2HPO|Reticulocytosis|Reticulocytosis
C0800956|T201|LC|17849-1|LNC2HPO|Reticulocytosis|Reticulocytosis
C0800956|T201|LN|17849-1|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0800956|T201|DN|17849-1|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0800956|T201|MTH_LN|17849-1|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0800956|T201|OSN|17849-1|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0800956|T201|LC|17849-1|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C1146797|T201|LN|31112-6|LNC2HPO|Reticulocytosis|Reticulocytosis
C1146797|T201|DN|31112-6|LNC2HPO|Reticulocytosis|Reticulocytosis
C1146797|T201|MTH_LN|31112-6|LNC2HPO|Reticulocytosis|Reticulocytosis
C1146797|T201|OSN|31112-6|LNC2HPO|Reticulocytosis|Reticulocytosis
C1146797|T201|LC|31112-6|LNC2HPO|Reticulocytosis|Reticulocytosis
C1146797|T201|LN|31112-6|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C1146797|T201|DN|31112-6|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C1146797|T201|MTH_LN|31112-6|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C1146797|T201|OSN|31112-6|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C1146797|T201|LC|31112-6|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C1624714|T201|LN|42758-3|LNC2HPO|Reticulocytosis|Reticulocytosis
C1624714|T201|DN|42758-3|LNC2HPO|Reticulocytosis|Reticulocytosis
C1624714|T201|OSN|42758-3|LNC2HPO|Reticulocytosis|Reticulocytosis
C1624714|T201|MTH_LN|42758-3|LNC2HPO|Reticulocytosis|Reticulocytosis
C1624714|T201|LC|42758-3|LNC2HPO|Reticulocytosis|Reticulocytosis
C1624714|T201|LN|42758-3|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C1624714|T201|DN|42758-3|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C1624714|T201|OSN|42758-3|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C1624714|T201|MTH_LN|42758-3|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C1624714|T201|LC|42758-3|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0366908|T201|LN|4679-7|LNC2HPO|Reticulocytosis|Reticulocytosis
C0366908|T201|DN|4679-7|LNC2HPO|Reticulocytosis|Reticulocytosis
C0366908|T201|OSN|4679-7|LNC2HPO|Reticulocytosis|Reticulocytosis
C0366908|T201|LC|4679-7|LNC2HPO|Reticulocytosis|Reticulocytosis
C0366908|T201|MTH_LN|4679-7|LNC2HPO|Reticulocytosis|Reticulocytosis
C0366908|T201|LN|4679-7|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0366908|T201|DN|4679-7|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0366908|T201|OSN|4679-7|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0366908|T201|LC|4679-7|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0366908|T201|MTH_LN|4679-7|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C2970267|T201|LN|60474-4|LNC2HPO|Reticulocytosis|Reticulocytosis
C2970267|T201|DN|60474-4|LNC2HPO|Reticulocytosis|Reticulocytosis
C2970267|T201|LC|60474-4|LNC2HPO|Reticulocytosis|Reticulocytosis
C2970267|T201|MTH_LN|60474-4|LNC2HPO|Reticulocytosis|Reticulocytosis
C2970267|T201|OSN|60474-4|LNC2HPO|Reticulocytosis|Reticulocytosis
C2970267|T201|LN|60474-4|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C2970267|T201|DN|60474-4|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C2970267|T201|LC|60474-4|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C2970267|T201|MTH_LN|60474-4|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C2970267|T201|OSN|60474-4|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0802054|T201|LC|19124-7|LNC2HPO|Hypermagnesiuria|Hypermagnesiuria
C0802054|T201|MTH_LN|19124-7|LNC2HPO|Hypermagnesiuria|Hypermagnesiuria
C0802054|T201|DN|19124-7|LNC2HPO|Hypermagnesiuria|Hypermagnesiuria
C0802054|T201|OSN|19124-7|LNC2HPO|Hypermagnesiuria|Hypermagnesiuria
C0802054|T201|LN|19124-7|LNC2HPO|Hypermagnesiuria|Hypermagnesiuria
C0802054|T201|LC|19124-7|LNC2HPO|Hypomagnesiuria|Hypomagnesiuria
C0802054|T201|MTH_LN|19124-7|LNC2HPO|Hypomagnesiuria|Hypomagnesiuria
C0802054|T201|DN|19124-7|LNC2HPO|Hypomagnesiuria|Hypomagnesiuria
C0802054|T201|OSN|19124-7|LNC2HPO|Hypomagnesiuria|Hypomagnesiuria
C0802054|T201|LN|19124-7|LNC2HPO|Hypomagnesiuria|Hypomagnesiuria
C0364612|T201|LN|2472-9|LNC2HPO|IgM deficiency|IgM deficiency
C0364612|T201|OSN|2472-9|LNC2HPO|IgM deficiency|IgM deficiency
C0364612|T201|MTH_LN|2472-9|LNC2HPO|IgM deficiency|IgM deficiency
C0364612|T201|LC|2472-9|LNC2HPO|IgM deficiency|IgM deficiency
C0364612|T201|DN|2472-9|LNC2HPO|IgM deficiency|IgM deficiency
C0945354|T201|LN|26450-7|LNC2HPO|Eosinophilia|Eosinophilia
C0945354|T201|OSN|26450-7|LNC2HPO|Eosinophilia|Eosinophilia
C0945354|T201|DN|26450-7|LNC2HPO|Eosinophilia|Eosinophilia
C0945354|T201|MTH_LN|26450-7|LNC2HPO|Eosinophilia|Eosinophilia
C0945354|T201|LC|26450-7|LNC2HPO|Eosinophilia|Eosinophilia
C0364538|T201|LN|2398-6|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C0364538|T201|MTH_LN|2398-6|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C0364538|T201|DN|2398-6|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C0364538|T201|OSN|2398-6|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C0364538|T201|LC|2398-6|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C3847305|T201|LN|74632-1|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C3847305|T201|OSN|74632-1|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C3847305|T201|LC|74632-1|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C3847305|T201|MTH_LN|74632-1|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C3847305|T201|DN|74632-1|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C0364539|T201|LN|2399-4|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C0364539|T201|MTH_LN|2399-4|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C0364539|T201|DN|2399-4|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C0364539|T201|OSN|2399-4|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C0364539|T201|LC|2399-4|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C2736145|T201|LN|57734-6|LNC2HPO|Ketonuria|Ketonuria
C2736145|T201|MTH_LN|57734-6|LNC2HPO|Ketonuria|Ketonuria
C2736145|T201|DN|57734-6|LNC2HPO|Ketonuria|Ketonuria
C2736145|T201|OSN|57734-6|LNC2HPO|Ketonuria|Ketonuria
C2736145|T201|LC|57734-6|LNC2HPO|Ketonuria|Ketonuria
C2736145|T201|LN|57734-6|LNC2HPO|Acetonuria|Acetonuria
C2736145|T201|MTH_LN|57734-6|LNC2HPO|Acetonuria|Acetonuria
C2736145|T201|DN|57734-6|LNC2HPO|Acetonuria|Acetonuria
C2736145|T201|OSN|57734-6|LNC2HPO|Acetonuria|Acetonuria
C2736145|T201|LC|57734-6|LNC2HPO|Acetonuria|Acetonuria
C2736145|T201|LN|57734-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C2736145|T201|MTH_LN|57734-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C2736145|T201|DN|57734-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C2736145|T201|OSN|57734-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C2736145|T201|LC|57734-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C2736145|T201|LN|57734-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C2736145|T201|MTH_LN|57734-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C2736145|T201|DN|57734-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C2736145|T201|OSN|57734-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C2736145|T201|LC|57734-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C0798130|T201|LN|14957-5|LNC2HPO|Microalbuminuria|Microalbuminuria
C0798130|T201|MTH_LN|14957-5|LNC2HPO|Microalbuminuria|Microalbuminuria
C0798130|T201|DN|14957-5|LNC2HPO|Microalbuminuria|Microalbuminuria
C0798130|T201|OSN|14957-5|LNC2HPO|Microalbuminuria|Microalbuminuria
C0798130|T201|LC|14957-5|LNC2HPO|Microalbuminuria|Microalbuminuria
C2926219|T201|LN|58448-2|LNC2HPO|Microalbuminuria|Microalbuminuria
C2926219|T201|DN|58448-2|LNC2HPO|Microalbuminuria|Microalbuminuria
C2926219|T201|MTH_LN|58448-2|LNC2HPO|Microalbuminuria|Microalbuminuria
C2926219|T201|LC|58448-2|LNC2HPO|Microalbuminuria|Microalbuminuria
C2926219|T201|OSN|58448-2|LNC2HPO|Microalbuminuria|Microalbuminuria
C0365099|T201|LN|2955-3|LNC2HPO|Hypernatriuria|Hypernatriuria
C0365099|T201|MTH_LN|2955-3|LNC2HPO|Hypernatriuria|Hypernatriuria
C0365099|T201|DN|2955-3|LNC2HPO|Hypernatriuria|Hypernatriuria
C0365099|T201|OSN|2955-3|LNC2HPO|Hypernatriuria|Hypernatriuria
C0365099|T201|LC|2955-3|LNC2HPO|Hypernatriuria|Hypernatriuria
C0365099|T201|LN|2955-3|LNC2HPO|Hyponatriuria|Hyponatriuria
C0365099|T201|MTH_LN|2955-3|LNC2HPO|Hyponatriuria|Hyponatriuria
C0365099|T201|DN|2955-3|LNC2HPO|Hyponatriuria|Hyponatriuria
C0365099|T201|OSN|2955-3|LNC2HPO|Hyponatriuria|Hyponatriuria
C0365099|T201|LC|2955-3|LNC2HPO|Hyponatriuria|Hyponatriuria
C0363974|T201|LN|1839-0|LNC2HPO|Hyperammonemia|Hyperammonemia
C0363974|T201|MTH_LN|1839-0|LNC2HPO|Hyperammonemia|Hyperammonemia
C0363974|T201|DN|1839-0|LNC2HPO|Hyperammonemia|Hyperammonemia
C0363974|T201|OSN|1839-0|LNC2HPO|Hyperammonemia|Hyperammonemia
C0363974|T201|LC|1839-0|LNC2HPO|Hyperammonemia|Hyperammonemia
C0363974|T201|LN|1839-0|LNC2HPO|Hypoammonemia|Hypoammonemia
C0363974|T201|MTH_LN|1839-0|LNC2HPO|Hypoammonemia|Hypoammonemia
C0363974|T201|DN|1839-0|LNC2HPO|Hypoammonemia|Hypoammonemia
C0363974|T201|OSN|1839-0|LNC2HPO|Hypoammonemia|Hypoammonemia
C0363974|T201|LC|1839-0|LNC2HPO|Hypoammonemia|Hypoammonemia
C0368530|T201|LN|600-7|LNC2HPO|Bacteremia|Bacteremia
C0368530|T201|DN|600-7|LNC2HPO|Bacteremia|Bacteremia
C0368530|T201|OSN|600-7|LNC2HPO|Bacteremia|Bacteremia
C0368530|T201|MTH_LN|600-7|LNC2HPO|Bacteremia|Bacteremia
C0368530|T201|LC|600-7|LNC2HPO|Bacteremia|Bacteremia
C0550261|T201|LN|12773-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0550261|T201|MTH_LN|12773-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0550261|T201|DN|12773-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0550261|T201|OSN|12773-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0550261|T201|LC|12773-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0550261|T201|LN|12773-8|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0550261|T201|MTH_LN|12773-8|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0550261|T201|DN|12773-8|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0550261|T201|OSN|12773-8|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0550261|T201|LC|12773-8|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0550264|T201|LN|13457-7|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0550264|T201|MTH_LN|13457-7|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0550264|T201|DN|13457-7|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0550264|T201|OSN|13457-7|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0550264|T201|LC|13457-7|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0550264|T201|LN|13457-7|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0550264|T201|MTH_LN|13457-7|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0550264|T201|DN|13457-7|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0550264|T201|OSN|13457-7|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0550264|T201|LC|13457-7|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0801307|T201|LN|18261-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0801307|T201|MTH_LN|18261-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0801307|T201|DN|18261-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0801307|T201|OSN|18261-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0801307|T201|LC|18261-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0801307|T201|LN|18261-8|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0801307|T201|MTH_LN|18261-8|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0801307|T201|DN|18261-8|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0801307|T201|OSN|18261-8|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0801307|T201|LC|18261-8|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0801308|T201|LN|18262-6|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0801308|T201|MTH_LN|18262-6|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0801308|T201|DN|18262-6|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0801308|T201|OSN|18262-6|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0801308|T201|LC|18262-6|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0801308|T201|LN|18262-6|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0801308|T201|MTH_LN|18262-6|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0801308|T201|DN|18262-6|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0801308|T201|OSN|18262-6|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0801308|T201|LC|18262-6|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0364225|T201|MTH_LN|2089-1|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0364225|T201|DN|2089-1|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0364225|T201|LN|2089-1|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0364225|T201|OSN|2089-1|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0364225|T201|LC|2089-1|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0364225|T201|MTH_LN|2089-1|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0364225|T201|DN|2089-1|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0364225|T201|LN|2089-1|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0364225|T201|OSN|2089-1|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0364225|T201|LC|2089-1|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0880253|T201|LN|22748-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0880253|T201|DN|22748-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0880253|T201|MTH_LN|22748-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0880253|T201|OSN|22748-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0880253|T201|LC|22748-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0880253|T201|LN|22748-8|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0880253|T201|DN|22748-8|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0880253|T201|MTH_LN|22748-8|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0880253|T201|OSN|22748-8|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0880253|T201|LC|22748-8|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C2603388|T201|DN|35198-1|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2603388|T201|MTH_LN|35198-1|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2603388|T201|LN|35198-1|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2603388|T201|OSN|35198-1|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2603388|T201|LC|35198-1|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2603388|T201|DN|35198-1|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C2603388|T201|MTH_LN|35198-1|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C2603388|T201|LN|35198-1|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C2603388|T201|OSN|35198-1|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C2603388|T201|LC|35198-1|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C1543545|T201|LN|39469-2|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1543545|T201|DN|39469-2|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1543545|T201|OSN|39469-2|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1543545|T201|MTH_LN|39469-2|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1543545|T201|LC|39469-2|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1543545|T201|LN|39469-2|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C1543545|T201|DN|39469-2|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C1543545|T201|OSN|39469-2|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C1543545|T201|MTH_LN|39469-2|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C1543545|T201|LC|39469-2|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C1954896|T201|LN|49132-4|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1954896|T201|DN|49132-4|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1954896|T201|MTH_LN|49132-4|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1954896|T201|OSN|49132-4|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1954896|T201|LC|49132-4|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1954896|T201|LN|49132-4|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C1954896|T201|DN|49132-4|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C1954896|T201|MTH_LN|49132-4|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C1954896|T201|OSN|49132-4|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C1954896|T201|LC|49132-4|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C2708273|T201|LN|55440-2|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2708273|T201|DN|55440-2|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2708273|T201|LC|55440-2|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2708273|T201|OSN|55440-2|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2708273|T201|MTH_LN|55440-2|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2708273|T201|LN|55440-2|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C2708273|T201|DN|55440-2|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C2708273|T201|LC|55440-2|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C2708273|T201|OSN|55440-2|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C2708273|T201|MTH_LN|55440-2|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C3481704|T201|LN|69419-0|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C3481704|T201|MTH_LN|69419-0|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C3481704|T201|OSN|69419-0|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C3481704|T201|LC|69419-0|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C3481704|T201|DN|69419-0|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C3481704|T201|LN|69419-0|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C3481704|T201|MTH_LN|69419-0|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C3481704|T201|OSN|69419-0|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C3481704|T201|LC|69419-0|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C3481704|T201|DN|69419-0|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C4531914|T201|LN|86911-5|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C4531914|T201|OSN|86911-5|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C4531914|T201|LC|86911-5|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C4531914|T201|MTH_LN|86911-5|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C4531914|T201|LN|86911-5|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C4531914|T201|OSN|86911-5|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C4531914|T201|LC|86911-5|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C4531914|T201|MTH_LN|86911-5|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0365023|T201|LN|2880-3|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C0365023|T201|MTH_LN|2880-3|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C0365023|T201|DN|2880-3|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C0365023|T201|OSN|2880-3|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C0365023|T201|LC|2880-3|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C0365023|T201|LN|2880-3|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C0365023|T201|MTH_LN|2880-3|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C0365023|T201|DN|2880-3|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C0365023|T201|OSN|2880-3|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C0365023|T201|LC|2880-3|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C4037678|T201|LN|76665-9|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C4037678|T201|OSN|76665-9|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C4037678|T201|MTH_LN|76665-9|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C4037678|T201|LC|76665-9|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C4037678|T201|DN|76665-9|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C4037678|T201|LN|76665-9|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C4037678|T201|OSN|76665-9|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C4037678|T201|MTH_LN|76665-9|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C4037678|T201|LC|76665-9|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C4037678|T201|DN|76665-9|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C4037677|T201|LN|76666-7|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C4037677|T201|OSN|76666-7|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C4037677|T201|MTH_LN|76666-7|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C4037677|T201|LC|76666-7|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C4037677|T201|DN|76666-7|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C4037677|T201|LN|76666-7|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C4037677|T201|OSN|76666-7|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C4037677|T201|MTH_LN|76666-7|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C4037677|T201|LC|76666-7|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C4037677|T201|DN|76666-7|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C4037676|T201|LN|76667-5|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C4037676|T201|OSN|76667-5|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C4037676|T201|LC|76667-5|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C4037676|T201|MTH_LN|76667-5|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C4037676|T201|DN|76667-5|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C4037676|T201|LN|76667-5|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C4037676|T201|OSN|76667-5|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C4037676|T201|LC|76667-5|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C4037676|T201|MTH_LN|76667-5|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C4037676|T201|DN|76667-5|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C4037570|T201|LN|76668-3|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C4037570|T201|LC|76668-3|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C4037570|T201|MTH_LN|76668-3|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C4037570|T201|OSN|76668-3|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C4037570|T201|DN|76668-3|LNC2HPO|Hyperproteinorrhachia|Hyperproteinorrhachia
C4037570|T201|LN|76668-3|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C4037570|T201|LC|76668-3|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C4037570|T201|MTH_LN|76668-3|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C4037570|T201|OSN|76668-3|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C4037570|T201|DN|76668-3|LNC2HPO|Hypoproteinorrhachia|Hypoproteinorrhachia
C0364482|T201|LN|2342-4|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C0364482|T201|MTH_LN|2342-4|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C0364482|T201|DN|2342-4|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C0364482|T201|OSN|2342-4|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C0364482|T201|LC|2342-4|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C0364482|T201|LN|2342-4|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C0364482|T201|MTH_LN|2342-4|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C0364482|T201|DN|2342-4|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C0364482|T201|OSN|2342-4|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C0364482|T201|LC|2342-4|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C0797918|T201|LN|14744-7|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C0797918|T201|MTH_LN|14744-7|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C0797918|T201|DN|14744-7|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C0797918|T201|OSN|14744-7|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C0797918|T201|LC|14744-7|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C0797918|T201|LN|14744-7|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C0797918|T201|MTH_LN|14744-7|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C0797918|T201|DN|14744-7|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C0797918|T201|OSN|14744-7|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C0797918|T201|LC|14744-7|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C4037569|T201|LN|76669-1|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C4037569|T201|OSN|76669-1|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C4037569|T201|LC|76669-1|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C4037569|T201|MTH_LN|76669-1|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C4037569|T201|DN|76669-1|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C4037569|T201|LN|76669-1|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C4037569|T201|OSN|76669-1|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C4037569|T201|LC|76669-1|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C4037569|T201|MTH_LN|76669-1|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C4037569|T201|DN|76669-1|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C4037568|T201|LN|76670-9|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C4037568|T201|MTH_LN|76670-9|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C4037568|T201|OSN|76670-9|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C4037568|T201|LC|76670-9|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C4037568|T201|DN|76670-9|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C4037568|T201|LN|76670-9|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C4037568|T201|MTH_LN|76670-9|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C4037568|T201|OSN|76670-9|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C4037568|T201|LC|76670-9|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C4037568|T201|DN|76670-9|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C4037567|T201|LN|76671-7|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C4037567|T201|MTH_LN|76671-7|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C4037567|T201|LC|76671-7|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C4037567|T201|OSN|76671-7|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C4037567|T201|DN|76671-7|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C4037567|T201|LN|76671-7|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C4037567|T201|MTH_LN|76671-7|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C4037567|T201|LC|76671-7|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C4037567|T201|OSN|76671-7|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C4037567|T201|DN|76671-7|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C4037566|T201|LN|76672-5|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C4037566|T201|LC|76672-5|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C4037566|T201|MTH_LN|76672-5|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C4037566|T201|OSN|76672-5|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C4037566|T201|DN|76672-5|LNC2HPO|Hyperglycorrhachia|Hyperglycorrhachia
C4037566|T201|LN|76672-5|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C4037566|T201|LC|76672-5|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C4037566|T201|MTH_LN|76672-5|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C4037566|T201|OSN|76672-5|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C4037566|T201|DN|76672-5|LNC2HPO|Hypoglycorrhachia|Hypoglycorrhachia
C0484581|T201|LN|10449-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0484581|T201|MTH_LN|10449-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0484581|T201|DN|10449-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0484581|T201|OSN|10449-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0484581|T201|LC|10449-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0484581|T201|LN|10449-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0484581|T201|MTH_LN|10449-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0484581|T201|DN|10449-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0484581|T201|OSN|10449-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0484581|T201|LC|10449-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0484581|T201|LN|10449-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0484581|T201|MTH_LN|10449-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0484581|T201|DN|10449-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0484581|T201|OSN|10449-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0484581|T201|LC|10449-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0484599|T201|LN|10450-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0484599|T201|MTH_LN|10450-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0484599|T201|DN|10450-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0484599|T201|OSN|10450-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0484599|T201|LC|10450-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0484599|T201|LN|10450-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0484599|T201|MTH_LN|10450-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0484599|T201|DN|10450-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0484599|T201|OSN|10450-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0484599|T201|LC|10450-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0484599|T201|LN|10450-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0484599|T201|MTH_LN|10450-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0484599|T201|DN|10450-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0484599|T201|OSN|10450-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0484599|T201|LC|10450-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549973|T201|LN|10832-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549973|T201|MTH_LN|10832-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549973|T201|DN|10832-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549973|T201|OSN|10832-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549973|T201|LC|10832-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549973|T201|LN|10832-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549973|T201|MTH_LN|10832-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549973|T201|DN|10832-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549973|T201|OSN|10832-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549973|T201|LC|10832-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549973|T201|LN|10832-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549973|T201|MTH_LN|10832-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549973|T201|DN|10832-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549973|T201|OSN|10832-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549973|T201|LC|10832-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549989|T201|LN|11032-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549989|T201|MTH_LN|11032-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549989|T201|DN|11032-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549989|T201|OSN|11032-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549989|T201|LC|11032-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549989|T201|LN|11032-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549989|T201|MTH_LN|11032-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549989|T201|DN|11032-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549989|T201|OSN|11032-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549989|T201|LC|11032-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549989|T201|LN|11032-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549989|T201|MTH_LN|11032-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549989|T201|DN|11032-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549989|T201|OSN|11032-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549989|T201|LC|11032-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550357|T201|LN|11142-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550357|T201|MTH_LN|11142-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550357|T201|DN|11142-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550357|T201|OSN|11142-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550357|T201|LC|11142-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550357|T201|LN|11142-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550357|T201|MTH_LN|11142-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550357|T201|DN|11142-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550357|T201|OSN|11142-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550357|T201|LC|11142-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550357|T201|LN|11142-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550357|T201|MTH_LN|11142-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550357|T201|DN|11142-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550357|T201|OSN|11142-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550357|T201|LC|11142-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550363|T201|LN|11143-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550363|T201|DN|11143-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550363|T201|MTH_LN|11143-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550363|T201|OSN|11143-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550363|T201|LC|11143-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550363|T201|LN|11143-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550363|T201|DN|11143-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550363|T201|MTH_LN|11143-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550363|T201|OSN|11143-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550363|T201|LC|11143-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550363|T201|LN|11143-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550363|T201|DN|11143-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550363|T201|MTH_LN|11143-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550363|T201|OSN|11143-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550363|T201|LC|11143-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549981|T201|LN|12610-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549981|T201|MTH_LN|12610-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549981|T201|DN|12610-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549981|T201|OSN|12610-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549981|T201|LC|12610-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549981|T201|LN|12610-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549981|T201|MTH_LN|12610-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549981|T201|DN|12610-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549981|T201|OSN|12610-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549981|T201|LC|12610-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549981|T201|LN|12610-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549981|T201|MTH_LN|12610-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549981|T201|DN|12610-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549981|T201|OSN|12610-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549981|T201|LC|12610-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550366|T201|LN|12611-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550366|T201|MTH_LN|12611-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550366|T201|DN|12611-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550366|T201|OSN|12611-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550366|T201|LC|12611-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550366|T201|LN|12611-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550366|T201|MTH_LN|12611-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550366|T201|DN|12611-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550366|T201|OSN|12611-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550366|T201|LC|12611-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550366|T201|LN|12611-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550366|T201|MTH_LN|12611-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550366|T201|DN|12611-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550366|T201|OSN|12611-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550366|T201|LC|12611-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550000|T201|LN|12614-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550000|T201|MTH_LN|12614-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550000|T201|DN|12614-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550000|T201|OSN|12614-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550000|T201|LC|12614-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550000|T201|LN|12614-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550000|T201|MTH_LN|12614-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550000|T201|DN|12614-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550000|T201|OSN|12614-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550000|T201|LC|12614-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550000|T201|LN|12614-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550000|T201|MTH_LN|12614-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550000|T201|DN|12614-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550000|T201|OSN|12614-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550000|T201|LC|12614-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549978|T201|LN|12615-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549978|T201|MTH_LN|12615-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549978|T201|DN|12615-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549978|T201|OSN|12615-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549978|T201|LC|12615-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549978|T201|LN|12615-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549978|T201|MTH_LN|12615-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549978|T201|DN|12615-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549978|T201|OSN|12615-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549978|T201|LC|12615-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549978|T201|LN|12615-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549978|T201|MTH_LN|12615-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549978|T201|DN|12615-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549978|T201|OSN|12615-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549978|T201|LC|12615-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549983|T201|LN|12616-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549983|T201|MTH_LN|12616-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549983|T201|DN|12616-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549983|T201|OSN|12616-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549983|T201|LC|12616-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549983|T201|LN|12616-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549983|T201|MTH_LN|12616-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549983|T201|DN|12616-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549983|T201|OSN|12616-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549983|T201|LC|12616-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549983|T201|LN|12616-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549983|T201|MTH_LN|12616-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549983|T201|DN|12616-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549983|T201|OSN|12616-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549983|T201|LC|12616-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549986|T201|LN|12617-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549986|T201|MTH_LN|12617-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549986|T201|DN|12617-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549986|T201|OSN|12617-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549986|T201|LC|12617-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549986|T201|LN|12617-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549986|T201|MTH_LN|12617-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549986|T201|DN|12617-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549986|T201|OSN|12617-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549986|T201|LC|12617-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549986|T201|LN|12617-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549986|T201|MTH_LN|12617-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549986|T201|DN|12617-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549986|T201|OSN|12617-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549986|T201|LC|12617-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549991|T201|LN|12618-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549991|T201|MTH_LN|12618-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549991|T201|DN|12618-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549991|T201|OSN|12618-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549991|T201|LC|12618-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549991|T201|LN|12618-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549991|T201|MTH_LN|12618-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549991|T201|DN|12618-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549991|T201|OSN|12618-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549991|T201|LC|12618-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549991|T201|LN|12618-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549991|T201|MTH_LN|12618-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549991|T201|DN|12618-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549991|T201|OSN|12618-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549991|T201|LC|12618-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549993|T201|LN|12619-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549993|T201|MTH_LN|12619-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549993|T201|DN|12619-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549993|T201|OSN|12619-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549993|T201|LC|12619-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549993|T201|LN|12619-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549993|T201|MTH_LN|12619-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549993|T201|DN|12619-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549993|T201|OSN|12619-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549993|T201|LC|12619-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549993|T201|LN|12619-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549993|T201|MTH_LN|12619-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549993|T201|DN|12619-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549993|T201|OSN|12619-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549993|T201|LC|12619-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549995|T201|LN|12620-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549995|T201|MTH_LN|12620-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549995|T201|DN|12620-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549995|T201|OSN|12620-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549995|T201|LC|12620-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549995|T201|LN|12620-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549995|T201|MTH_LN|12620-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549995|T201|DN|12620-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549995|T201|OSN|12620-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549995|T201|LC|12620-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549995|T201|LN|12620-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549995|T201|MTH_LN|12620-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549995|T201|DN|12620-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549995|T201|OSN|12620-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549995|T201|LC|12620-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550005|T201|LN|12621-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550005|T201|MTH_LN|12621-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550005|T201|DN|12621-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550005|T201|OSN|12621-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550005|T201|LC|12621-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550005|T201|LN|12621-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550005|T201|MTH_LN|12621-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550005|T201|DN|12621-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550005|T201|OSN|12621-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550005|T201|LC|12621-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550005|T201|LN|12621-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550005|T201|MTH_LN|12621-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550005|T201|DN|12621-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550005|T201|OSN|12621-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550005|T201|LC|12621-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549967|T201|LN|12622-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549967|T201|MTH_LN|12622-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549967|T201|DN|12622-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549967|T201|OSN|12622-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549967|T201|LC|12622-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549967|T201|LN|12622-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549967|T201|MTH_LN|12622-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549967|T201|DN|12622-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549967|T201|OSN|12622-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549967|T201|LC|12622-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549967|T201|LN|12622-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549967|T201|MTH_LN|12622-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549967|T201|DN|12622-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549967|T201|OSN|12622-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549967|T201|LC|12622-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549968|T201|LN|12623-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549968|T201|MTH_LN|12623-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549968|T201|DN|12623-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549968|T201|OSN|12623-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549968|T201|LC|12623-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549968|T201|LN|12623-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549968|T201|MTH_LN|12623-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549968|T201|DN|12623-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549968|T201|OSN|12623-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549968|T201|LC|12623-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549968|T201|LN|12623-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549968|T201|MTH_LN|12623-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549968|T201|DN|12623-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549968|T201|OSN|12623-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549968|T201|LC|12623-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549970|T201|LN|12624-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549970|T201|MTH_LN|12624-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549970|T201|DN|12624-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549970|T201|OSN|12624-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549970|T201|LC|12624-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549970|T201|LN|12624-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549970|T201|MTH_LN|12624-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549970|T201|DN|12624-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549970|T201|OSN|12624-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549970|T201|LC|12624-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549970|T201|LN|12624-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549970|T201|MTH_LN|12624-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549970|T201|DN|12624-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549970|T201|OSN|12624-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549970|T201|LC|12624-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549971|T201|LN|12625-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549971|T201|MTH_LN|12625-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549971|T201|DN|12625-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549971|T201|OSN|12625-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549971|T201|LC|12625-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549971|T201|LN|12625-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549971|T201|MTH_LN|12625-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549971|T201|DN|12625-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549971|T201|OSN|12625-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549971|T201|LC|12625-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549971|T201|LN|12625-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549971|T201|MTH_LN|12625-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549971|T201|DN|12625-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549971|T201|OSN|12625-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549971|T201|LC|12625-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549972|T201|LN|12626-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549972|T201|MTH_LN|12626-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549972|T201|DN|12626-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549972|T201|OSN|12626-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549972|T201|LC|12626-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549972|T201|LN|12626-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549972|T201|MTH_LN|12626-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549972|T201|DN|12626-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549972|T201|OSN|12626-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549972|T201|LC|12626-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549972|T201|LN|12626-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549972|T201|MTH_LN|12626-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549972|T201|DN|12626-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549972|T201|OSN|12626-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549972|T201|LC|12626-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549976|T201|LN|12627-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549976|T201|MTH_LN|12627-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549976|T201|DN|12627-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549976|T201|OSN|12627-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549976|T201|LC|12627-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549976|T201|LN|12627-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549976|T201|MTH_LN|12627-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549976|T201|DN|12627-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549976|T201|OSN|12627-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549976|T201|LC|12627-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549976|T201|LN|12627-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549976|T201|MTH_LN|12627-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549976|T201|DN|12627-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549976|T201|OSN|12627-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549976|T201|LC|12627-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550006|T201|LN|12638-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550006|T201|DN|12638-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550006|T201|MTH_LN|12638-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550006|T201|OSN|12638-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550006|T201|LC|12638-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550006|T201|LN|12638-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550006|T201|DN|12638-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550006|T201|MTH_LN|12638-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550006|T201|OSN|12638-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550006|T201|LC|12638-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550006|T201|LN|12638-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550006|T201|DN|12638-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550006|T201|MTH_LN|12638-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550006|T201|OSN|12638-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550006|T201|LC|12638-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549974|T201|LN|12639-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549974|T201|MTH_LN|12639-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549974|T201|DN|12639-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549974|T201|OSN|12639-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549974|T201|LC|12639-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549974|T201|LN|12639-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549974|T201|MTH_LN|12639-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549974|T201|DN|12639-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549974|T201|OSN|12639-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549974|T201|LC|12639-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549974|T201|LN|12639-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549974|T201|MTH_LN|12639-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549974|T201|DN|12639-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549974|T201|OSN|12639-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549974|T201|LC|12639-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549994|T201|LN|12640-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549994|T201|MTH_LN|12640-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549994|T201|DN|12640-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549994|T201|OSN|12640-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549994|T201|LC|12640-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549994|T201|LN|12640-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549994|T201|MTH_LN|12640-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549994|T201|DN|12640-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549994|T201|OSN|12640-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549994|T201|LC|12640-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549994|T201|LN|12640-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549994|T201|MTH_LN|12640-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549994|T201|DN|12640-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549994|T201|OSN|12640-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549994|T201|LC|12640-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549999|T201|LN|12641-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549999|T201|MTH_LN|12641-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549999|T201|DN|12641-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549999|T201|OSN|12641-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549999|T201|LC|12641-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549999|T201|LN|12641-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549999|T201|MTH_LN|12641-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549999|T201|DN|12641-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549999|T201|OSN|12641-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549999|T201|LC|12641-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549999|T201|LN|12641-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549999|T201|MTH_LN|12641-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549999|T201|DN|12641-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549999|T201|OSN|12641-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549999|T201|LC|12641-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549997|T201|LN|12642-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549997|T201|MTH_LN|12642-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549997|T201|DN|12642-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549997|T201|OSN|12642-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549997|T201|LC|12642-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549997|T201|LN|12642-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549997|T201|MTH_LN|12642-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549997|T201|DN|12642-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549997|T201|OSN|12642-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549997|T201|LC|12642-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549997|T201|LN|12642-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549997|T201|MTH_LN|12642-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549997|T201|DN|12642-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549997|T201|OSN|12642-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549997|T201|LC|12642-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550001|T201|LN|12643-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550001|T201|MTH_LN|12643-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550001|T201|DN|12643-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550001|T201|OSN|12643-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550001|T201|LC|12643-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550001|T201|LN|12643-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550001|T201|MTH_LN|12643-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550001|T201|DN|12643-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550001|T201|OSN|12643-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550001|T201|LC|12643-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550001|T201|LN|12643-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550001|T201|MTH_LN|12643-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550001|T201|DN|12643-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550001|T201|OSN|12643-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550001|T201|LC|12643-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550004|T201|LN|12644-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550004|T201|MTH_LN|12644-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550004|T201|DN|12644-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550004|T201|OSN|12644-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550004|T201|LC|12644-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550004|T201|LN|12644-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550004|T201|MTH_LN|12644-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550004|T201|DN|12644-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550004|T201|OSN|12644-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550004|T201|LC|12644-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550004|T201|LN|12644-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550004|T201|MTH_LN|12644-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550004|T201|DN|12644-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550004|T201|OSN|12644-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550004|T201|LC|12644-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549964|T201|LN|12645-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549964|T201|MTH_LN|12645-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549964|T201|DN|12645-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549964|T201|OSN|12645-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549964|T201|LC|12645-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549964|T201|LN|12645-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549964|T201|MTH_LN|12645-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549964|T201|DN|12645-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549964|T201|OSN|12645-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549964|T201|LC|12645-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549964|T201|LN|12645-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549964|T201|MTH_LN|12645-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549964|T201|DN|12645-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549964|T201|OSN|12645-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549964|T201|LC|12645-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549977|T201|LN|12646-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549977|T201|MTH_LN|12646-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549977|T201|DN|12646-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549977|T201|OSN|12646-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549977|T201|LC|12646-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549977|T201|LN|12646-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549977|T201|MTH_LN|12646-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549977|T201|DN|12646-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549977|T201|OSN|12646-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549977|T201|LC|12646-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549977|T201|LN|12646-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549977|T201|MTH_LN|12646-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549977|T201|DN|12646-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549977|T201|OSN|12646-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549977|T201|LC|12646-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549969|T201|LN|12647-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549969|T201|MTH_LN|12647-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549969|T201|DN|12647-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549969|T201|OSN|12647-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549969|T201|LC|12647-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549969|T201|LN|12647-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549969|T201|MTH_LN|12647-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549969|T201|DN|12647-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549969|T201|OSN|12647-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549969|T201|LC|12647-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549969|T201|LN|12647-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549969|T201|MTH_LN|12647-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549969|T201|DN|12647-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549969|T201|OSN|12647-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549969|T201|LC|12647-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549975|T201|LN|12648-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549975|T201|DN|12648-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549975|T201|MTH_LN|12648-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549975|T201|OSN|12648-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549975|T201|LC|12648-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549975|T201|LN|12648-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549975|T201|DN|12648-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549975|T201|MTH_LN|12648-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549975|T201|OSN|12648-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549975|T201|LC|12648-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549975|T201|LN|12648-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549975|T201|DN|12648-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549975|T201|MTH_LN|12648-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549975|T201|OSN|12648-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549975|T201|LC|12648-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549996|T201|LN|12649-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549996|T201|DN|12649-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549996|T201|MTH_LN|12649-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549996|T201|OSN|12649-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549996|T201|LC|12649-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549996|T201|LN|12649-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549996|T201|DN|12649-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549996|T201|MTH_LN|12649-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549996|T201|OSN|12649-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549996|T201|LC|12649-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549996|T201|LN|12649-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549996|T201|DN|12649-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549996|T201|MTH_LN|12649-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549996|T201|OSN|12649-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549996|T201|LC|12649-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549985|T201|LN|12650-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549985|T201|DN|12650-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549985|T201|MTH_LN|12650-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549985|T201|OSN|12650-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549985|T201|LC|12650-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549985|T201|LN|12650-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549985|T201|DN|12650-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549985|T201|MTH_LN|12650-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549985|T201|OSN|12650-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549985|T201|LC|12650-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549985|T201|LN|12650-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549985|T201|DN|12650-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549985|T201|MTH_LN|12650-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549985|T201|OSN|12650-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549985|T201|LC|12650-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549966|T201|LN|12651-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549966|T201|MTH_LN|12651-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549966|T201|DN|12651-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549966|T201|OSN|12651-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549966|T201|LC|12651-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549966|T201|LN|12651-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549966|T201|MTH_LN|12651-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549966|T201|DN|12651-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549966|T201|OSN|12651-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549966|T201|LC|12651-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549966|T201|LN|12651-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549966|T201|MTH_LN|12651-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549966|T201|DN|12651-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549966|T201|OSN|12651-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549966|T201|LC|12651-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549982|T201|LN|12652-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549982|T201|MTH_LN|12652-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549982|T201|DN|12652-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549982|T201|OSN|12652-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549982|T201|LC|12652-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549982|T201|LN|12652-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549982|T201|MTH_LN|12652-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549982|T201|DN|12652-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549982|T201|OSN|12652-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549982|T201|LC|12652-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549982|T201|LN|12652-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549982|T201|MTH_LN|12652-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549982|T201|DN|12652-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549982|T201|OSN|12652-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549982|T201|LC|12652-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550002|T201|LN|12653-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550002|T201|MTH_LN|12653-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550002|T201|DN|12653-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550002|T201|OSN|12653-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550002|T201|LC|12653-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0550002|T201|LN|12653-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550002|T201|MTH_LN|12653-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550002|T201|DN|12653-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550002|T201|OSN|12653-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550002|T201|LC|12653-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0550002|T201|LN|12653-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550002|T201|MTH_LN|12653-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550002|T201|DN|12653-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550002|T201|OSN|12653-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0550002|T201|LC|12653-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549965|T201|LN|12654-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549965|T201|MTH_LN|12654-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549965|T201|DN|12654-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549965|T201|OSN|12654-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549965|T201|LC|12654-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549965|T201|LN|12654-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549965|T201|MTH_LN|12654-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549965|T201|DN|12654-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549965|T201|OSN|12654-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549965|T201|LC|12654-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549965|T201|LN|12654-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549965|T201|MTH_LN|12654-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549965|T201|DN|12654-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549965|T201|OSN|12654-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549965|T201|LC|12654-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549980|T201|LN|12655-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549980|T201|MTH_LN|12655-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549980|T201|DN|12655-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549980|T201|OSN|12655-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549980|T201|LC|12655-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549980|T201|LN|12655-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549980|T201|MTH_LN|12655-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549980|T201|DN|12655-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549980|T201|OSN|12655-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549980|T201|LC|12655-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549980|T201|LN|12655-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549980|T201|MTH_LN|12655-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549980|T201|DN|12655-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549980|T201|OSN|12655-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549980|T201|LC|12655-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549990|T201|LN|12656-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549990|T201|MTH_LN|12656-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549990|T201|DN|12656-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549990|T201|OSN|12656-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549990|T201|LC|12656-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549990|T201|LN|12656-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549990|T201|MTH_LN|12656-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549990|T201|DN|12656-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549990|T201|OSN|12656-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549990|T201|LC|12656-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549990|T201|LN|12656-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549990|T201|MTH_LN|12656-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549990|T201|DN|12656-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549990|T201|OSN|12656-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549990|T201|LC|12656-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549988|T201|LN|12657-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549988|T201|MTH_LN|12657-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549988|T201|DN|12657-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549988|T201|OSN|12657-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549988|T201|LC|12657-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549988|T201|LN|12657-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549988|T201|MTH_LN|12657-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549988|T201|DN|12657-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549988|T201|OSN|12657-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549988|T201|LC|12657-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549988|T201|LN|12657-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549988|T201|MTH_LN|12657-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549988|T201|DN|12657-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549988|T201|OSN|12657-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549988|T201|LC|12657-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549992|T201|LN|12658-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549992|T201|MTH_LN|12658-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549992|T201|DN|12658-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549992|T201|OSN|12658-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549992|T201|LC|12658-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549992|T201|LN|12658-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549992|T201|MTH_LN|12658-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549992|T201|DN|12658-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549992|T201|OSN|12658-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549992|T201|LC|12658-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549992|T201|LN|12658-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549992|T201|MTH_LN|12658-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549992|T201|DN|12658-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549992|T201|OSN|12658-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549992|T201|LC|12658-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549998|T201|LN|12659-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549998|T201|MTH_LN|12659-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549998|T201|DN|12659-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549998|T201|OSN|12659-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549998|T201|LC|12659-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0549998|T201|LN|12659-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549998|T201|MTH_LN|12659-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549998|T201|DN|12659-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549998|T201|OSN|12659-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549998|T201|LC|12659-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0549998|T201|LN|12659-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549998|T201|MTH_LN|12659-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549998|T201|DN|12659-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549998|T201|OSN|12659-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0549998|T201|LC|12659-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0796797|T201|LN|13606-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0796797|T201|MTH_LN|13606-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0796797|T201|DN|13606-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0796797|T201|OSN|13606-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0796797|T201|LC|13606-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0796797|T201|LN|13606-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0796797|T201|MTH_LN|13606-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0796797|T201|DN|13606-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0796797|T201|OSN|13606-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0796797|T201|LC|13606-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0796797|T201|LN|13606-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0796797|T201|MTH_LN|13606-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0796797|T201|DN|13606-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0796797|T201|OSN|13606-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0796797|T201|LC|13606-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0796798|T201|LN|13607-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0796798|T201|MTH_LN|13607-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0796798|T201|DN|13607-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0796798|T201|OSN|13607-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0796798|T201|LC|13607-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0796798|T201|LN|13607-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0796798|T201|MTH_LN|13607-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0796798|T201|DN|13607-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0796798|T201|OSN|13607-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0796798|T201|LC|13607-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0796798|T201|LN|13607-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0796798|T201|MTH_LN|13607-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0796798|T201|DN|13607-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0796798|T201|OSN|13607-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0796798|T201|LC|13607-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797054|T201|LN|13865-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797054|T201|DN|13865-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797054|T201|OSN|13865-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797054|T201|MTH_LN|13865-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797054|T201|LC|13865-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797054|T201|LN|13865-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797054|T201|DN|13865-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797054|T201|OSN|13865-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797054|T201|MTH_LN|13865-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797054|T201|LC|13865-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797054|T201|LN|13865-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797054|T201|DN|13865-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797054|T201|OSN|13865-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797054|T201|MTH_LN|13865-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797054|T201|LC|13865-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797055|T201|LN|13866-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797055|T201|MTH_LN|13866-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797055|T201|DN|13866-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797055|T201|OSN|13866-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797055|T201|LC|13866-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797055|T201|LN|13866-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797055|T201|MTH_LN|13866-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797055|T201|DN|13866-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797055|T201|OSN|13866-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797055|T201|LC|13866-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797055|T201|LN|13866-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797055|T201|MTH_LN|13866-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797055|T201|DN|13866-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797055|T201|OSN|13866-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797055|T201|LC|13866-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797323|T201|LN|14137-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797323|T201|MTH_LN|14137-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797323|T201|DN|14137-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797323|T201|OSN|14137-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797323|T201|LC|14137-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797323|T201|LN|14137-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797323|T201|MTH_LN|14137-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797323|T201|DN|14137-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797323|T201|OSN|14137-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797323|T201|LC|14137-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797323|T201|LN|14137-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797323|T201|MTH_LN|14137-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797323|T201|DN|14137-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797323|T201|OSN|14137-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797323|T201|LC|14137-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797917|T201|LN|14743-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797917|T201|MTH_LN|14743-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797917|T201|DN|14743-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797917|T201|OSN|14743-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797917|T201|LC|14743-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797917|T201|LN|14743-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797917|T201|MTH_LN|14743-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797917|T201|DN|14743-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797917|T201|OSN|14743-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797917|T201|LC|14743-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797917|T201|LN|14743-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797917|T201|MTH_LN|14743-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797917|T201|DN|14743-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797917|T201|OSN|14743-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797917|T201|LC|14743-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797923|T201|LN|14749-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797923|T201|MTH_LN|14749-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797923|T201|DN|14749-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797923|T201|OSN|14749-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797923|T201|LC|14749-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797923|T201|LN|14749-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797923|T201|MTH_LN|14749-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797923|T201|DN|14749-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797923|T201|OSN|14749-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797923|T201|LC|14749-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797923|T201|LN|14749-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797923|T201|MTH_LN|14749-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797923|T201|DN|14749-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797923|T201|OSN|14749-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797923|T201|LC|14749-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797925|T201|LN|14751-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797925|T201|DN|14751-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797925|T201|OSN|14751-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797925|T201|MTH_LN|14751-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797925|T201|LC|14751-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797925|T201|LN|14751-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797925|T201|DN|14751-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797925|T201|OSN|14751-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797925|T201|MTH_LN|14751-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797925|T201|LC|14751-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797925|T201|LN|14751-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797925|T201|DN|14751-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797925|T201|OSN|14751-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797925|T201|MTH_LN|14751-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797925|T201|LC|14751-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797926|T201|LN|14752-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797926|T201|DN|14752-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797926|T201|OSN|14752-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797926|T201|MTH_LN|14752-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797926|T201|LC|14752-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797926|T201|LN|14752-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797926|T201|DN|14752-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797926|T201|OSN|14752-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797926|T201|MTH_LN|14752-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797926|T201|LC|14752-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797926|T201|LN|14752-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797926|T201|DN|14752-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797926|T201|OSN|14752-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797926|T201|MTH_LN|14752-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797926|T201|LC|14752-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797927|T201|LN|14753-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797927|T201|MTH_LN|14753-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797927|T201|DN|14753-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797927|T201|OSN|14753-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797927|T201|LC|14753-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797927|T201|LN|14753-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797927|T201|MTH_LN|14753-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797927|T201|DN|14753-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797927|T201|OSN|14753-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797927|T201|LC|14753-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797927|T201|LN|14753-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797927|T201|MTH_LN|14753-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797927|T201|DN|14753-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797927|T201|OSN|14753-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797927|T201|LC|14753-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797928|T201|LN|14754-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797928|T201|MTH_LN|14754-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797928|T201|DN|14754-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797928|T201|OSN|14754-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797928|T201|LC|14754-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797928|T201|LN|14754-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797928|T201|MTH_LN|14754-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797928|T201|DN|14754-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797928|T201|OSN|14754-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797928|T201|LC|14754-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797928|T201|LN|14754-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797928|T201|MTH_LN|14754-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797928|T201|DN|14754-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797928|T201|OSN|14754-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797928|T201|LC|14754-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797929|T201|LN|14755-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797929|T201|MTH_LN|14755-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797929|T201|DN|14755-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797929|T201|OSN|14755-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797929|T201|LC|14755-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797929|T201|LN|14755-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797929|T201|MTH_LN|14755-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797929|T201|DN|14755-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797929|T201|OSN|14755-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797929|T201|LC|14755-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797929|T201|LN|14755-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797929|T201|MTH_LN|14755-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797929|T201|DN|14755-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797929|T201|OSN|14755-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797929|T201|LC|14755-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797930|T201|LN|14756-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797930|T201|DN|14756-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797930|T201|MTH_LN|14756-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797930|T201|OSN|14756-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797930|T201|LC|14756-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797930|T201|LN|14756-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797930|T201|DN|14756-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797930|T201|MTH_LN|14756-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797930|T201|OSN|14756-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797930|T201|LC|14756-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797930|T201|LN|14756-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797930|T201|DN|14756-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797930|T201|MTH_LN|14756-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797930|T201|OSN|14756-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797930|T201|LC|14756-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797931|T201|LN|14757-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797931|T201|MTH_LN|14757-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797931|T201|DN|14757-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797931|T201|OSN|14757-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797931|T201|LC|14757-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797931|T201|LN|14757-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797931|T201|MTH_LN|14757-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797931|T201|DN|14757-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797931|T201|OSN|14757-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797931|T201|LC|14757-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797931|T201|LN|14757-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797931|T201|MTH_LN|14757-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797931|T201|DN|14757-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797931|T201|OSN|14757-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797931|T201|LC|14757-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797932|T201|LN|14758-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797932|T201|MTH_LN|14758-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797932|T201|DN|14758-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797932|T201|OSN|14758-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797932|T201|LC|14758-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797932|T201|LN|14758-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797932|T201|MTH_LN|14758-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797932|T201|DN|14758-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797932|T201|OSN|14758-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797932|T201|LC|14758-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797932|T201|LN|14758-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797932|T201|MTH_LN|14758-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797932|T201|DN|14758-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797932|T201|OSN|14758-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797932|T201|LC|14758-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797933|T201|LN|14759-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797933|T201|DN|14759-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797933|T201|MTH_LN|14759-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797933|T201|OSN|14759-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797933|T201|LC|14759-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797933|T201|LN|14759-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797933|T201|DN|14759-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797933|T201|MTH_LN|14759-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797933|T201|OSN|14759-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797933|T201|LC|14759-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797933|T201|LN|14759-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797933|T201|DN|14759-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797933|T201|MTH_LN|14759-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797933|T201|OSN|14759-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797933|T201|LC|14759-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797934|T201|LN|14760-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797934|T201|MTH_LN|14760-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797934|T201|DN|14760-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797934|T201|OSN|14760-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797934|T201|LC|14760-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797934|T201|LN|14760-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797934|T201|MTH_LN|14760-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797934|T201|DN|14760-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797934|T201|OSN|14760-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797934|T201|LC|14760-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797934|T201|LN|14760-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797934|T201|MTH_LN|14760-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797934|T201|DN|14760-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797934|T201|OSN|14760-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797934|T201|LC|14760-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797935|T201|LN|14761-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797935|T201|MTH_LN|14761-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797935|T201|DN|14761-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797935|T201|OSN|14761-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797935|T201|LC|14761-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797935|T201|LN|14761-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797935|T201|MTH_LN|14761-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797935|T201|DN|14761-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797935|T201|OSN|14761-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797935|T201|LC|14761-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797935|T201|LN|14761-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797935|T201|MTH_LN|14761-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797935|T201|DN|14761-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797935|T201|OSN|14761-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797935|T201|LC|14761-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797936|T201|LN|14762-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797936|T201|MTH_LN|14762-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797936|T201|DN|14762-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797936|T201|OSN|14762-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797936|T201|LC|14762-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797936|T201|LN|14762-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797936|T201|MTH_LN|14762-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797936|T201|DN|14762-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797936|T201|OSN|14762-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797936|T201|LC|14762-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797936|T201|LN|14762-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797936|T201|MTH_LN|14762-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797936|T201|DN|14762-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797936|T201|OSN|14762-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797936|T201|LC|14762-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797937|T201|LN|14763-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797937|T201|DN|14763-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797937|T201|MTH_LN|14763-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797937|T201|OSN|14763-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797937|T201|LC|14763-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797937|T201|LN|14763-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797937|T201|DN|14763-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797937|T201|MTH_LN|14763-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797937|T201|OSN|14763-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797937|T201|LC|14763-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797937|T201|LN|14763-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797937|T201|DN|14763-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797937|T201|MTH_LN|14763-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797937|T201|OSN|14763-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797937|T201|LC|14763-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797938|T201|LN|14764-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797938|T201|MTH_LN|14764-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797938|T201|DN|14764-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797938|T201|OSN|14764-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797938|T201|LC|14764-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797938|T201|LN|14764-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797938|T201|MTH_LN|14764-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797938|T201|DN|14764-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797938|T201|OSN|14764-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797938|T201|LC|14764-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797938|T201|LN|14764-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797938|T201|MTH_LN|14764-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797938|T201|DN|14764-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797938|T201|OSN|14764-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797938|T201|LC|14764-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797939|T201|LN|14765-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797939|T201|DN|14765-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797939|T201|MTH_LN|14765-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797939|T201|OSN|14765-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797939|T201|LC|14765-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797939|T201|LN|14765-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797939|T201|DN|14765-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797939|T201|MTH_LN|14765-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797939|T201|OSN|14765-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797939|T201|LC|14765-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797939|T201|LN|14765-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797939|T201|DN|14765-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797939|T201|MTH_LN|14765-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797939|T201|OSN|14765-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797939|T201|LC|14765-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797940|T201|LN|14766-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797940|T201|DN|14766-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797940|T201|MTH_LN|14766-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797940|T201|OSN|14766-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797940|T201|LC|14766-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797940|T201|LN|14766-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797940|T201|DN|14766-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797940|T201|MTH_LN|14766-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797940|T201|OSN|14766-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797940|T201|LC|14766-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797940|T201|LN|14766-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797940|T201|DN|14766-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797940|T201|MTH_LN|14766-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797940|T201|OSN|14766-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797940|T201|LC|14766-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797941|T201|LN|14767-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797941|T201|DN|14767-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797941|T201|MTH_LN|14767-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797941|T201|OSN|14767-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797941|T201|LC|14767-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797941|T201|LN|14767-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797941|T201|DN|14767-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797941|T201|MTH_LN|14767-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797941|T201|OSN|14767-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797941|T201|LC|14767-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797941|T201|LN|14767-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797941|T201|DN|14767-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797941|T201|MTH_LN|14767-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797941|T201|OSN|14767-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797941|T201|LC|14767-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797942|T201|LN|14768-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797942|T201|MTH_LN|14768-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797942|T201|DN|14768-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797942|T201|OSN|14768-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797942|T201|LC|14768-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797942|T201|LN|14768-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797942|T201|MTH_LN|14768-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797942|T201|DN|14768-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797942|T201|OSN|14768-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797942|T201|LC|14768-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797942|T201|LN|14768-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797942|T201|MTH_LN|14768-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797942|T201|DN|14768-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797942|T201|OSN|14768-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797942|T201|LC|14768-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797943|T201|LN|14769-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797943|T201|DN|14769-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797943|T201|MTH_LN|14769-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797943|T201|OSN|14769-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797943|T201|LC|14769-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797943|T201|LN|14769-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797943|T201|DN|14769-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797943|T201|MTH_LN|14769-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797943|T201|OSN|14769-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797943|T201|LC|14769-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797943|T201|LN|14769-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797943|T201|DN|14769-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797943|T201|MTH_LN|14769-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797943|T201|OSN|14769-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797943|T201|LC|14769-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797945|T201|LN|14771-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797945|T201|MTH_LN|14771-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797945|T201|DN|14771-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797945|T201|OSN|14771-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797945|T201|LC|14771-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797945|T201|LN|14771-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797945|T201|MTH_LN|14771-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797945|T201|DN|14771-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797945|T201|OSN|14771-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797945|T201|LC|14771-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797945|T201|LN|14771-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797945|T201|MTH_LN|14771-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797945|T201|DN|14771-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797945|T201|OSN|14771-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797945|T201|LC|14771-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363626|T201|LN|1492-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363626|T201|DN|1492-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363626|T201|OSN|1492-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363626|T201|MTH_LN|1492-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363626|T201|LC|1492-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363626|T201|LN|1492-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363626|T201|DN|1492-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363626|T201|OSN|1492-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363626|T201|MTH_LN|1492-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363626|T201|LC|1492-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363626|T201|LN|1492-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363626|T201|DN|1492-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363626|T201|OSN|1492-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363626|T201|MTH_LN|1492-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363626|T201|LC|1492-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363627|T201|LN|1493-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363627|T201|DN|1493-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363627|T201|OSN|1493-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363627|T201|MTH_LN|1493-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363627|T201|LC|1493-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363627|T201|LN|1493-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363627|T201|DN|1493-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363627|T201|OSN|1493-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363627|T201|MTH_LN|1493-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363627|T201|LC|1493-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363627|T201|LN|1493-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363627|T201|DN|1493-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363627|T201|OSN|1493-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363627|T201|MTH_LN|1493-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363627|T201|LC|1493-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363628|T201|LN|1494-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363628|T201|DN|1494-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363628|T201|OSN|1494-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363628|T201|MTH_LN|1494-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363628|T201|LC|1494-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363628|T201|LN|1494-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363628|T201|DN|1494-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363628|T201|OSN|1494-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363628|T201|MTH_LN|1494-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363628|T201|LC|1494-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363628|T201|LN|1494-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363628|T201|DN|1494-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363628|T201|OSN|1494-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363628|T201|MTH_LN|1494-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363628|T201|LC|1494-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482534|T201|LN|1496-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482534|T201|DN|1496-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482534|T201|OSN|1496-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482534|T201|MTH_LN|1496-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482534|T201|LC|1496-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482534|T201|LN|1496-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482534|T201|DN|1496-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482534|T201|OSN|1496-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482534|T201|MTH_LN|1496-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482534|T201|LC|1496-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482534|T201|LN|1496-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482534|T201|DN|1496-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482534|T201|OSN|1496-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482534|T201|MTH_LN|1496-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482534|T201|LC|1496-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363631|T201|LN|1497-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363631|T201|DN|1497-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363631|T201|OSN|1497-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363631|T201|MTH_LN|1497-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363631|T201|LC|1497-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363631|T201|LN|1497-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363631|T201|DN|1497-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363631|T201|OSN|1497-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363631|T201|MTH_LN|1497-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363631|T201|LC|1497-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363631|T201|LN|1497-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363631|T201|DN|1497-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363631|T201|OSN|1497-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363631|T201|MTH_LN|1497-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363631|T201|LC|1497-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363632|T201|LN|1498-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363632|T201|DN|1498-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363632|T201|MTH_LN|1498-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363632|T201|OSN|1498-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363632|T201|LC|1498-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363632|T201|LN|1498-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363632|T201|DN|1498-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363632|T201|MTH_LN|1498-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363632|T201|OSN|1498-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363632|T201|LC|1498-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363632|T201|LN|1498-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363632|T201|DN|1498-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363632|T201|MTH_LN|1498-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363632|T201|OSN|1498-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363632|T201|LC|1498-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363633|T201|LN|1499-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363633|T201|DN|1499-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363633|T201|MTH_LN|1499-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363633|T201|OSN|1499-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363633|T201|LC|1499-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363633|T201|LN|1499-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363633|T201|DN|1499-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363633|T201|MTH_LN|1499-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363633|T201|OSN|1499-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363633|T201|LC|1499-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363633|T201|LN|1499-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363633|T201|DN|1499-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363633|T201|MTH_LN|1499-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363633|T201|OSN|1499-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363633|T201|LC|1499-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0798168|T201|LN|14995-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0798168|T201|MTH_LN|14995-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0798168|T201|DN|14995-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0798168|T201|OSN|14995-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0798168|T201|LC|14995-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0798168|T201|LN|14995-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0798168|T201|MTH_LN|14995-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0798168|T201|DN|14995-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0798168|T201|OSN|14995-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0798168|T201|LC|14995-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0798168|T201|LN|14995-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0798168|T201|MTH_LN|14995-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0798168|T201|DN|14995-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0798168|T201|OSN|14995-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0798168|T201|LC|14995-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0798169|T201|LN|14996-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0798169|T201|DN|14996-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0798169|T201|MTH_LN|14996-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0798169|T201|OSN|14996-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0798169|T201|LC|14996-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0798169|T201|LN|14996-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0798169|T201|DN|14996-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0798169|T201|MTH_LN|14996-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0798169|T201|OSN|14996-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0798169|T201|LC|14996-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0798169|T201|LN|14996-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0798169|T201|DN|14996-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0798169|T201|MTH_LN|14996-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0798169|T201|OSN|14996-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0798169|T201|LC|14996-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363634|T201|LN|1500-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363634|T201|DN|1500-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363634|T201|MTH_LN|1500-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363634|T201|OSN|1500-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363634|T201|LC|1500-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363634|T201|LN|1500-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363634|T201|DN|1500-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363634|T201|MTH_LN|1500-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363634|T201|OSN|1500-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363634|T201|LC|1500-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363634|T201|LN|1500-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363634|T201|DN|1500-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363634|T201|MTH_LN|1500-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363634|T201|OSN|1500-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363634|T201|LC|1500-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363635|T201|LN|1501-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363635|T201|MTH_LN|1501-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363635|T201|DN|1501-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363635|T201|OSN|1501-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363635|T201|LC|1501-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363635|T201|LN|1501-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363635|T201|MTH_LN|1501-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363635|T201|DN|1501-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363635|T201|OSN|1501-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363635|T201|LC|1501-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363635|T201|LN|1501-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363635|T201|MTH_LN|1501-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363635|T201|DN|1501-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363635|T201|OSN|1501-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363635|T201|LC|1501-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363637|T201|LN|1503-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363637|T201|MTH_LN|1503-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363637|T201|DN|1503-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363637|T201|OSN|1503-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363637|T201|LC|1503-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363637|T201|LN|1503-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363637|T201|MTH_LN|1503-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363637|T201|DN|1503-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363637|T201|OSN|1503-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363637|T201|LC|1503-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363637|T201|LN|1503-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363637|T201|MTH_LN|1503-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363637|T201|DN|1503-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363637|T201|OSN|1503-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363637|T201|LC|1503-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363638|T201|LN|1504-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363638|T201|MTH_LN|1504-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363638|T201|DN|1504-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363638|T201|OSN|1504-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363638|T201|LC|1504-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363638|T201|LN|1504-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363638|T201|MTH_LN|1504-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363638|T201|DN|1504-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363638|T201|OSN|1504-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363638|T201|LC|1504-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363638|T201|LN|1504-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363638|T201|MTH_LN|1504-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363638|T201|DN|1504-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363638|T201|OSN|1504-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363638|T201|LC|1504-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363640|T201|LN|1506-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363640|T201|DN|1506-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363640|T201|MTH_LN|1506-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363640|T201|OSN|1506-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363640|T201|LC|1506-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363640|T201|LN|1506-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363640|T201|DN|1506-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363640|T201|MTH_LN|1506-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363640|T201|OSN|1506-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363640|T201|LC|1506-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363640|T201|LN|1506-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363640|T201|DN|1506-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363640|T201|MTH_LN|1506-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363640|T201|OSN|1506-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363640|T201|LC|1506-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363641|T201|LN|1507-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363641|T201|MTH_LN|1507-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363641|T201|DN|1507-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363641|T201|OSN|1507-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363641|T201|LC|1507-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363641|T201|LN|1507-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363641|T201|MTH_LN|1507-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363641|T201|DN|1507-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363641|T201|OSN|1507-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363641|T201|LC|1507-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363641|T201|LN|1507-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363641|T201|MTH_LN|1507-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363641|T201|DN|1507-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363641|T201|OSN|1507-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363641|T201|LC|1507-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363644|T201|MTH_LN|1510-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363644|T201|DN|1510-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363644|T201|LN|1510-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363644|T201|OSN|1510-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363644|T201|LC|1510-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363644|T201|MTH_LN|1510-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363644|T201|DN|1510-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363644|T201|LN|1510-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363644|T201|OSN|1510-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363644|T201|LC|1510-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363644|T201|MTH_LN|1510-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363644|T201|DN|1510-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363644|T201|LN|1510-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363644|T201|OSN|1510-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363644|T201|LC|1510-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363645|T201|LN|1512-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363645|T201|DN|1512-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363645|T201|MTH_LN|1512-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363645|T201|OSN|1512-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363645|T201|LC|1512-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363645|T201|LN|1512-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363645|T201|DN|1512-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363645|T201|MTH_LN|1512-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363645|T201|OSN|1512-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363645|T201|LC|1512-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363645|T201|LN|1512-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363645|T201|DN|1512-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363645|T201|MTH_LN|1512-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363645|T201|OSN|1512-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363645|T201|LC|1512-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363646|T201|LN|1513-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363646|T201|DN|1513-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363646|T201|MTH_LN|1513-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363646|T201|OSN|1513-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363646|T201|LC|1513-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363646|T201|LN|1513-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363646|T201|DN|1513-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363646|T201|MTH_LN|1513-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363646|T201|OSN|1513-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363646|T201|LC|1513-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363646|T201|LN|1513-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363646|T201|DN|1513-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363646|T201|MTH_LN|1513-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363646|T201|OSN|1513-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363646|T201|LC|1513-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363647|T201|LN|1514-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363647|T201|MTH_LN|1514-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363647|T201|DN|1514-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363647|T201|OSN|1514-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363647|T201|LC|1514-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363647|T201|LN|1514-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363647|T201|MTH_LN|1514-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363647|T201|DN|1514-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363647|T201|OSN|1514-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363647|T201|LC|1514-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363647|T201|LN|1514-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363647|T201|MTH_LN|1514-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363647|T201|DN|1514-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363647|T201|OSN|1514-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363647|T201|LC|1514-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363649|T201|LN|1516-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363649|T201|MTH_LN|1516-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363649|T201|DN|1516-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363649|T201|OSN|1516-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363649|T201|LC|1516-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363649|T201|LN|1516-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363649|T201|MTH_LN|1516-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363649|T201|DN|1516-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363649|T201|OSN|1516-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363649|T201|LC|1516-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363649|T201|LN|1516-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363649|T201|MTH_LN|1516-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363649|T201|DN|1516-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363649|T201|OSN|1516-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363649|T201|LC|1516-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363650|T201|LN|1517-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363650|T201|DN|1517-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363650|T201|MTH_LN|1517-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363650|T201|OSN|1517-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363650|T201|LC|1517-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363650|T201|LN|1517-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363650|T201|DN|1517-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363650|T201|MTH_LN|1517-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363650|T201|OSN|1517-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363650|T201|LC|1517-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363650|T201|LN|1517-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363650|T201|DN|1517-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363650|T201|MTH_LN|1517-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363650|T201|OSN|1517-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363650|T201|LC|1517-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363651|T201|LN|1518-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363651|T201|MTH_LN|1518-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363651|T201|DN|1518-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363651|T201|OSN|1518-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363651|T201|LC|1518-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363651|T201|LN|1518-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363651|T201|MTH_LN|1518-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363651|T201|DN|1518-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363651|T201|OSN|1518-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363651|T201|LC|1518-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363651|T201|LN|1518-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363651|T201|MTH_LN|1518-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363651|T201|DN|1518-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363651|T201|OSN|1518-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363651|T201|LC|1518-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363653|T201|LN|1520-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363653|T201|MTH_LN|1520-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363653|T201|DN|1520-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363653|T201|OSN|1520-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363653|T201|LC|1520-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363653|T201|LN|1520-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363653|T201|MTH_LN|1520-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363653|T201|DN|1520-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363653|T201|OSN|1520-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363653|T201|LC|1520-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363653|T201|LN|1520-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363653|T201|MTH_LN|1520-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363653|T201|DN|1520-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363653|T201|OSN|1520-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363653|T201|LC|1520-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482535|T201|LN|1521-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482535|T201|MTH_LN|1521-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482535|T201|DN|1521-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482535|T201|OSN|1521-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482535|T201|LC|1521-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482535|T201|LN|1521-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482535|T201|MTH_LN|1521-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482535|T201|DN|1521-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482535|T201|OSN|1521-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482535|T201|LC|1521-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482535|T201|LN|1521-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482535|T201|MTH_LN|1521-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482535|T201|DN|1521-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482535|T201|OSN|1521-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482535|T201|LC|1521-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363655|T201|LN|1522-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363655|T201|DN|1522-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363655|T201|MTH_LN|1522-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363655|T201|OSN|1522-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363655|T201|LC|1522-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363655|T201|LN|1522-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363655|T201|DN|1522-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363655|T201|MTH_LN|1522-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363655|T201|OSN|1522-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363655|T201|LC|1522-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363655|T201|LN|1522-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363655|T201|DN|1522-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363655|T201|MTH_LN|1522-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363655|T201|OSN|1522-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363655|T201|LC|1522-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363656|T201|LN|1523-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363656|T201|DN|1523-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363656|T201|MTH_LN|1523-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363656|T201|OSN|1523-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363656|T201|LC|1523-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363656|T201|LN|1523-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363656|T201|DN|1523-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363656|T201|MTH_LN|1523-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363656|T201|OSN|1523-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363656|T201|LC|1523-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363656|T201|LN|1523-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363656|T201|DN|1523-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363656|T201|MTH_LN|1523-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363656|T201|OSN|1523-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363656|T201|LC|1523-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482536|T201|LN|1524-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482536|T201|DN|1524-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482536|T201|MTH_LN|1524-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482536|T201|OSN|1524-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482536|T201|LC|1524-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482536|T201|LN|1524-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482536|T201|DN|1524-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482536|T201|MTH_LN|1524-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482536|T201|OSN|1524-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482536|T201|LC|1524-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482536|T201|LN|1524-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482536|T201|DN|1524-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482536|T201|MTH_LN|1524-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482536|T201|OSN|1524-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482536|T201|LC|1524-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363658|T201|LN|1525-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363658|T201|MTH_LN|1525-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363658|T201|DN|1525-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363658|T201|OSN|1525-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363658|T201|LC|1525-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363658|T201|LN|1525-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363658|T201|MTH_LN|1525-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363658|T201|DN|1525-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363658|T201|OSN|1525-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363658|T201|LC|1525-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363658|T201|LN|1525-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363658|T201|MTH_LN|1525-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363658|T201|DN|1525-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363658|T201|OSN|1525-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363658|T201|LC|1525-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363659|T201|LN|1526-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363659|T201|DN|1526-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363659|T201|MTH_LN|1526-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363659|T201|OSN|1526-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363659|T201|LC|1526-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363659|T201|LN|1526-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363659|T201|DN|1526-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363659|T201|MTH_LN|1526-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363659|T201|OSN|1526-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363659|T201|LC|1526-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363659|T201|LN|1526-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363659|T201|DN|1526-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363659|T201|MTH_LN|1526-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363659|T201|OSN|1526-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363659|T201|LC|1526-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482537|T201|LN|1527-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482537|T201|MTH_LN|1527-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482537|T201|DN|1527-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482537|T201|OSN|1527-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482537|T201|LC|1527-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482537|T201|LN|1527-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482537|T201|MTH_LN|1527-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482537|T201|DN|1527-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482537|T201|OSN|1527-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482537|T201|LC|1527-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482537|T201|LN|1527-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482537|T201|MTH_LN|1527-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482537|T201|DN|1527-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482537|T201|OSN|1527-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482537|T201|LC|1527-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363661|T201|MTH_LN|1528-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363661|T201|DN|1528-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363661|T201|LN|1528-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363661|T201|OSN|1528-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363661|T201|LC|1528-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363661|T201|MTH_LN|1528-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363661|T201|DN|1528-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363661|T201|LN|1528-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363661|T201|OSN|1528-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363661|T201|LC|1528-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363661|T201|MTH_LN|1528-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363661|T201|DN|1528-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363661|T201|LN|1528-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363661|T201|OSN|1528-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363661|T201|LC|1528-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363662|T201|LN|1530-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363662|T201|MTH_LN|1530-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363662|T201|DN|1530-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363662|T201|OSN|1530-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363662|T201|LC|1530-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363662|T201|LN|1530-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363662|T201|MTH_LN|1530-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363662|T201|DN|1530-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363662|T201|OSN|1530-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363662|T201|LC|1530-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363662|T201|LN|1530-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363662|T201|MTH_LN|1530-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363662|T201|DN|1530-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363662|T201|OSN|1530-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363662|T201|LC|1530-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363665|T201|LN|1533-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363665|T201|DN|1533-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363665|T201|MTH_LN|1533-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363665|T201|OSN|1533-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363665|T201|LC|1533-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363665|T201|LN|1533-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363665|T201|DN|1533-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363665|T201|MTH_LN|1533-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363665|T201|OSN|1533-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363665|T201|LC|1533-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363665|T201|LN|1533-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363665|T201|DN|1533-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363665|T201|MTH_LN|1533-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363665|T201|OSN|1533-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363665|T201|LC|1533-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363666|T201|LN|1534-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363666|T201|DN|1534-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363666|T201|MTH_LN|1534-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363666|T201|OSN|1534-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363666|T201|LC|1534-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363666|T201|LN|1534-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363666|T201|DN|1534-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363666|T201|MTH_LN|1534-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363666|T201|OSN|1534-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363666|T201|LC|1534-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363666|T201|LN|1534-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363666|T201|DN|1534-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363666|T201|MTH_LN|1534-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363666|T201|OSN|1534-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363666|T201|LC|1534-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363667|T201|LN|1535-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363667|T201|DN|1535-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363667|T201|MTH_LN|1535-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363667|T201|OSN|1535-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363667|T201|LC|1535-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363667|T201|LN|1535-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363667|T201|DN|1535-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363667|T201|MTH_LN|1535-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363667|T201|OSN|1535-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363667|T201|LC|1535-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363667|T201|LN|1535-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363667|T201|DN|1535-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363667|T201|MTH_LN|1535-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363667|T201|OSN|1535-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363667|T201|LC|1535-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363668|T201|LN|1536-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363668|T201|DN|1536-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363668|T201|MTH_LN|1536-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363668|T201|OSN|1536-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363668|T201|LC|1536-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363668|T201|LN|1536-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363668|T201|DN|1536-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363668|T201|MTH_LN|1536-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363668|T201|OSN|1536-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363668|T201|LC|1536-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363668|T201|LN|1536-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363668|T201|DN|1536-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363668|T201|MTH_LN|1536-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363668|T201|OSN|1536-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363668|T201|LC|1536-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363669|T201|LN|1537-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363669|T201|DN|1537-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363669|T201|MTH_LN|1537-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363669|T201|OSN|1537-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363669|T201|LC|1537-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363669|T201|LN|1537-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363669|T201|DN|1537-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363669|T201|MTH_LN|1537-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363669|T201|OSN|1537-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363669|T201|LC|1537-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363669|T201|LN|1537-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363669|T201|DN|1537-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363669|T201|MTH_LN|1537-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363669|T201|OSN|1537-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363669|T201|LC|1537-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363671|T201|LN|1539-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363671|T201|DN|1539-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363671|T201|MTH_LN|1539-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363671|T201|OSN|1539-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363671|T201|LC|1539-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363671|T201|LN|1539-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363671|T201|DN|1539-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363671|T201|MTH_LN|1539-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363671|T201|OSN|1539-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363671|T201|LC|1539-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363671|T201|LN|1539-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363671|T201|DN|1539-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363671|T201|MTH_LN|1539-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363671|T201|OSN|1539-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363671|T201|LC|1539-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363672|T201|LN|1540-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363672|T201|MTH_LN|1540-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363672|T201|DN|1540-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363672|T201|OSN|1540-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363672|T201|LC|1540-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363672|T201|LN|1540-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363672|T201|MTH_LN|1540-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363672|T201|DN|1540-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363672|T201|OSN|1540-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363672|T201|LC|1540-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363672|T201|LN|1540-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363672|T201|MTH_LN|1540-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363672|T201|DN|1540-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363672|T201|OSN|1540-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363672|T201|LC|1540-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363674|T201|LN|1542-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363674|T201|MTH_LN|1542-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363674|T201|DN|1542-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363674|T201|OSN|1542-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363674|T201|LC|1542-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363674|T201|LN|1542-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363674|T201|MTH_LN|1542-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363674|T201|DN|1542-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363674|T201|OSN|1542-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363674|T201|LC|1542-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363674|T201|LN|1542-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363674|T201|MTH_LN|1542-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363674|T201|DN|1542-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363674|T201|OSN|1542-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363674|T201|LC|1542-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363675|T201|LN|1543-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363675|T201|DN|1543-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363675|T201|MTH_LN|1543-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363675|T201|OSN|1543-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363675|T201|LC|1543-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363675|T201|LN|1543-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363675|T201|DN|1543-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363675|T201|MTH_LN|1543-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363675|T201|OSN|1543-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363675|T201|LC|1543-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363675|T201|LN|1543-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363675|T201|DN|1543-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363675|T201|MTH_LN|1543-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363675|T201|OSN|1543-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363675|T201|LC|1543-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0700436|T201|LN|1544-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0700436|T201|MTH_LN|1544-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0700436|T201|DN|1544-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0700436|T201|OSN|1544-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0700436|T201|LC|1544-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0700436|T201|LN|1544-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0700436|T201|MTH_LN|1544-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0700436|T201|DN|1544-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0700436|T201|OSN|1544-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0700436|T201|LC|1544-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0700436|T201|LN|1544-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0700436|T201|MTH_LN|1544-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0700436|T201|DN|1544-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0700436|T201|OSN|1544-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0700436|T201|LC|1544-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363678|T201|LN|1547-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363678|T201|DN|1547-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363678|T201|MTH_LN|1547-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363678|T201|OSN|1547-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363678|T201|LC|1547-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363678|T201|LN|1547-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363678|T201|DN|1547-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363678|T201|MTH_LN|1547-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363678|T201|OSN|1547-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363678|T201|LC|1547-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363678|T201|LN|1547-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363678|T201|DN|1547-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363678|T201|MTH_LN|1547-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363678|T201|OSN|1547-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363678|T201|LC|1547-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482538|T201|LN|1548-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482538|T201|DN|1548-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482538|T201|MTH_LN|1548-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482538|T201|OSN|1548-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482538|T201|LC|1548-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482538|T201|LN|1548-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482538|T201|DN|1548-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482538|T201|MTH_LN|1548-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482538|T201|OSN|1548-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482538|T201|LC|1548-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482538|T201|LN|1548-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482538|T201|DN|1548-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482538|T201|MTH_LN|1548-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482538|T201|OSN|1548-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482538|T201|LC|1548-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482539|T201|LN|1549-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482539|T201|DN|1549-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482539|T201|MTH_LN|1549-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482539|T201|OSN|1549-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482539|T201|LC|1549-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482539|T201|LN|1549-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482539|T201|DN|1549-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482539|T201|MTH_LN|1549-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482539|T201|OSN|1549-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482539|T201|LC|1549-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482539|T201|LN|1549-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482539|T201|DN|1549-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482539|T201|MTH_LN|1549-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482539|T201|OSN|1549-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482539|T201|LC|1549-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482540|T201|LN|1550-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482540|T201|DN|1550-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482540|T201|MTH_LN|1550-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482540|T201|OSN|1550-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482540|T201|LC|1550-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482540|T201|LN|1550-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482540|T201|DN|1550-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482540|T201|MTH_LN|1550-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482540|T201|OSN|1550-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482540|T201|LC|1550-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482540|T201|LN|1550-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482540|T201|DN|1550-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482540|T201|MTH_LN|1550-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482540|T201|OSN|1550-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482540|T201|LC|1550-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482541|T201|LN|1551-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482541|T201|DN|1551-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482541|T201|MTH_LN|1551-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482541|T201|OSN|1551-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482541|T201|LC|1551-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482541|T201|LN|1551-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482541|T201|DN|1551-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482541|T201|MTH_LN|1551-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482541|T201|OSN|1551-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482541|T201|LC|1551-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482541|T201|LN|1551-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482541|T201|DN|1551-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482541|T201|MTH_LN|1551-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482541|T201|OSN|1551-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482541|T201|LC|1551-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482542|T201|LN|1552-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482542|T201|DN|1552-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482542|T201|MTH_LN|1552-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482542|T201|OSN|1552-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482542|T201|LC|1552-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482542|T201|LN|1552-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482542|T201|DN|1552-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482542|T201|MTH_LN|1552-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482542|T201|OSN|1552-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482542|T201|LC|1552-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482542|T201|LN|1552-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482542|T201|DN|1552-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482542|T201|MTH_LN|1552-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482542|T201|OSN|1552-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482542|T201|LC|1552-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482543|T201|LN|1553-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482543|T201|DN|1553-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482543|T201|MTH_LN|1553-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482543|T201|OSN|1553-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482543|T201|LC|1553-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482543|T201|LN|1553-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482543|T201|DN|1553-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482543|T201|MTH_LN|1553-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482543|T201|OSN|1553-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482543|T201|LC|1553-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482543|T201|LN|1553-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482543|T201|DN|1553-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482543|T201|MTH_LN|1553-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482543|T201|OSN|1553-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482543|T201|LC|1553-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363685|T201|LN|1554-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363685|T201|DN|1554-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363685|T201|MTH_LN|1554-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363685|T201|OSN|1554-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363685|T201|LC|1554-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363685|T201|LN|1554-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363685|T201|DN|1554-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363685|T201|MTH_LN|1554-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363685|T201|OSN|1554-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363685|T201|LC|1554-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0363685|T201|LN|1554-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363685|T201|DN|1554-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363685|T201|MTH_LN|1554-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363685|T201|OSN|1554-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0363685|T201|LC|1554-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799330|T201|LN|16165-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799330|T201|DN|16165-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799330|T201|MTH_LN|16165-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799330|T201|OSN|16165-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799330|T201|LC|16165-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799330|T201|LN|16165-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799330|T201|DN|16165-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799330|T201|MTH_LN|16165-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799330|T201|OSN|16165-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799330|T201|LC|16165-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799330|T201|LN|16165-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799330|T201|DN|16165-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799330|T201|MTH_LN|16165-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799330|T201|OSN|16165-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799330|T201|LC|16165-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799331|T201|LN|16166-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799331|T201|DN|16166-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799331|T201|MTH_LN|16166-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799331|T201|OSN|16166-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799331|T201|LC|16166-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799331|T201|LN|16166-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799331|T201|DN|16166-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799331|T201|MTH_LN|16166-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799331|T201|OSN|16166-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799331|T201|LC|16166-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799331|T201|LN|16166-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799331|T201|DN|16166-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799331|T201|MTH_LN|16166-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799331|T201|OSN|16166-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799331|T201|LC|16166-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799332|T201|LN|16167-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799332|T201|DN|16167-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799332|T201|MTH_LN|16167-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799332|T201|OSN|16167-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799332|T201|LC|16167-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799332|T201|LN|16167-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799332|T201|DN|16167-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799332|T201|MTH_LN|16167-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799332|T201|OSN|16167-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799332|T201|LC|16167-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799332|T201|LN|16167-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799332|T201|DN|16167-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799332|T201|MTH_LN|16167-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799332|T201|OSN|16167-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799332|T201|LC|16167-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799333|T201|LN|16168-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799333|T201|DN|16168-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799333|T201|MTH_LN|16168-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799333|T201|OSN|16168-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799333|T201|LC|16168-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799333|T201|LN|16168-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799333|T201|DN|16168-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799333|T201|MTH_LN|16168-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799333|T201|OSN|16168-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799333|T201|LC|16168-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799333|T201|LN|16168-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799333|T201|DN|16168-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799333|T201|MTH_LN|16168-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799333|T201|OSN|16168-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799333|T201|LC|16168-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799334|T201|LN|16169-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799334|T201|DN|16169-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799334|T201|MTH_LN|16169-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799334|T201|OSN|16169-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799334|T201|LC|16169-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799334|T201|LN|16169-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799334|T201|DN|16169-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799334|T201|MTH_LN|16169-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799334|T201|OSN|16169-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799334|T201|LC|16169-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799334|T201|LN|16169-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799334|T201|DN|16169-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799334|T201|MTH_LN|16169-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799334|T201|OSN|16169-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799334|T201|LC|16169-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799335|T201|LN|16170-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799335|T201|DN|16170-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799335|T201|MTH_LN|16170-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799335|T201|OSN|16170-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799335|T201|LC|16170-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0799335|T201|LN|16170-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799335|T201|DN|16170-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799335|T201|MTH_LN|16170-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799335|T201|OSN|16170-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799335|T201|LC|16170-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0799335|T201|LN|16170-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799335|T201|DN|16170-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799335|T201|MTH_LN|16170-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799335|T201|OSN|16170-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0799335|T201|LC|16170-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0800048|T201|LN|16914-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0800048|T201|DN|16914-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0800048|T201|MTH_LN|16914-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0800048|T201|OSN|16914-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0800048|T201|LC|16914-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0800048|T201|LN|16914-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0800048|T201|DN|16914-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0800048|T201|MTH_LN|16914-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0800048|T201|OSN|16914-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0800048|T201|LC|16914-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0800048|T201|LN|16914-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0800048|T201|DN|16914-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0800048|T201|MTH_LN|16914-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0800048|T201|OSN|16914-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0800048|T201|LC|16914-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0800049|T201|LN|16915-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0800049|T201|DN|16915-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0800049|T201|MTH_LN|16915-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0800049|T201|OSN|16915-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0800049|T201|LC|16915-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0800049|T201|LN|16915-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0800049|T201|DN|16915-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0800049|T201|MTH_LN|16915-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0800049|T201|OSN|16915-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0800049|T201|LC|16915-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0800049|T201|LN|16915-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0800049|T201|DN|16915-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0800049|T201|MTH_LN|16915-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0800049|T201|OSN|16915-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0800049|T201|LC|16915-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0800972|T201|LN|17865-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0800972|T201|MTH_LN|17865-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0800972|T201|DN|17865-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0800972|T201|OSN|17865-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0800972|T201|LC|17865-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0800972|T201|LN|17865-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0800972|T201|MTH_LN|17865-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0800972|T201|DN|17865-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0800972|T201|OSN|17865-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0800972|T201|LC|17865-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0800972|T201|LN|17865-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0800972|T201|MTH_LN|17865-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0800972|T201|DN|17865-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0800972|T201|OSN|17865-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0800972|T201|LC|17865-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0801384|T201|LN|18342-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0801384|T201|MTH_LN|18342-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0801384|T201|DN|18342-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0801384|T201|OSN|18342-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0801384|T201|LC|18342-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0801384|T201|LN|18342-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0801384|T201|MTH_LN|18342-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0801384|T201|DN|18342-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0801384|T201|OSN|18342-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0801384|T201|LC|18342-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0801384|T201|LN|18342-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0801384|T201|MTH_LN|18342-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0801384|T201|DN|18342-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0801384|T201|OSN|18342-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0801384|T201|LC|18342-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0801395|T201|LN|18353-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0801395|T201|MTH_LN|18353-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0801395|T201|DN|18353-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0801395|T201|OSN|18353-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0801395|T201|LC|18353-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0801395|T201|LN|18353-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0801395|T201|MTH_LN|18353-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0801395|T201|DN|18353-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0801395|T201|OSN|18353-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0801395|T201|LC|18353-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0801395|T201|LN|18353-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0801395|T201|MTH_LN|18353-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0801395|T201|DN|18353-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0801395|T201|OSN|18353-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0801395|T201|LC|18353-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0801396|T201|LN|18354-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0801396|T201|MTH_LN|18354-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0801396|T201|DN|18354-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0801396|T201|OSN|18354-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0801396|T201|LC|18354-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0801396|T201|LN|18354-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0801396|T201|MTH_LN|18354-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0801396|T201|DN|18354-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0801396|T201|OSN|18354-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0801396|T201|LC|18354-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0801396|T201|LN|18354-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0801396|T201|MTH_LN|18354-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0801396|T201|DN|18354-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0801396|T201|OSN|18354-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0801396|T201|LC|18354-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803251|T201|LN|20436-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803251|T201|MTH_LN|20436-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803251|T201|DN|20436-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803251|T201|OSN|20436-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803251|T201|LC|20436-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803251|T201|LN|20436-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803251|T201|MTH_LN|20436-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803251|T201|DN|20436-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803251|T201|OSN|20436-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803251|T201|LC|20436-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803251|T201|LN|20436-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803251|T201|MTH_LN|20436-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803251|T201|DN|20436-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803251|T201|OSN|20436-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803251|T201|LC|20436-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803252|T201|LN|20437-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803252|T201|MTH_LN|20437-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803252|T201|DN|20437-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803252|T201|OSN|20437-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803252|T201|LC|20437-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803252|T201|LN|20437-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803252|T201|MTH_LN|20437-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803252|T201|DN|20437-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803252|T201|OSN|20437-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803252|T201|LC|20437-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803252|T201|LN|20437-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803252|T201|MTH_LN|20437-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803252|T201|DN|20437-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803252|T201|OSN|20437-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803252|T201|LC|20437-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803253|T201|LN|20438-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803253|T201|MTH_LN|20438-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803253|T201|DN|20438-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803253|T201|OSN|20438-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803253|T201|LC|20438-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803253|T201|LN|20438-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803253|T201|MTH_LN|20438-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803253|T201|DN|20438-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803253|T201|OSN|20438-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803253|T201|LC|20438-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803253|T201|LN|20438-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803253|T201|MTH_LN|20438-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803253|T201|DN|20438-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803253|T201|OSN|20438-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803253|T201|LC|20438-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803254|T201|LN|20439-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803254|T201|MTH_LN|20439-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803254|T201|DN|20439-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803254|T201|OSN|20439-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803254|T201|LC|20439-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803254|T201|LN|20439-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803254|T201|MTH_LN|20439-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803254|T201|DN|20439-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803254|T201|OSN|20439-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803254|T201|LC|20439-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803254|T201|LN|20439-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803254|T201|MTH_LN|20439-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803254|T201|DN|20439-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803254|T201|OSN|20439-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803254|T201|LC|20439-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803255|T201|LN|20440-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803255|T201|DN|20440-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803255|T201|OSN|20440-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803255|T201|MTH_LN|20440-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803255|T201|LC|20440-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803255|T201|LN|20440-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803255|T201|DN|20440-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803255|T201|OSN|20440-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803255|T201|MTH_LN|20440-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803255|T201|LC|20440-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803255|T201|LN|20440-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803255|T201|DN|20440-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803255|T201|OSN|20440-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803255|T201|MTH_LN|20440-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803255|T201|LC|20440-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803256|T201|LN|20441-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803256|T201|DN|20441-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803256|T201|MTH_LN|20441-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803256|T201|OSN|20441-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803256|T201|LC|20441-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0803256|T201|LN|20441-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803256|T201|DN|20441-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803256|T201|MTH_LN|20441-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803256|T201|OSN|20441-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803256|T201|LC|20441-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0803256|T201|LN|20441-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803256|T201|DN|20441-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803256|T201|MTH_LN|20441-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803256|T201|OSN|20441-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0803256|T201|LC|20441-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0804102|T201|LN|21308-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0804102|T201|MTH_LN|21308-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0804102|T201|DN|21308-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0804102|T201|OSN|21308-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0804102|T201|LC|21308-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0804102|T201|LN|21308-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0804102|T201|MTH_LN|21308-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0804102|T201|DN|21308-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0804102|T201|OSN|21308-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0804102|T201|LC|21308-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0804102|T201|LN|21308-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0804102|T201|MTH_LN|21308-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0804102|T201|DN|21308-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0804102|T201|OSN|21308-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0804102|T201|LC|21308-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0804103|T201|LN|21309-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0804103|T201|MTH_LN|21309-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0804103|T201|DN|21309-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0804103|T201|OSN|21309-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0804103|T201|LC|21309-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0804103|T201|LN|21309-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0804103|T201|MTH_LN|21309-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0804103|T201|DN|21309-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0804103|T201|OSN|21309-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0804103|T201|LC|21309-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0804103|T201|LN|21309-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0804103|T201|MTH_LN|21309-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0804103|T201|DN|21309-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0804103|T201|OSN|21309-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0804103|T201|LC|21309-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0804104|T201|LN|21310-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0804104|T201|MTH_LN|21310-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0804104|T201|DN|21310-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0804104|T201|OSN|21310-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0804104|T201|LC|21310-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0804104|T201|LN|21310-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0804104|T201|MTH_LN|21310-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0804104|T201|DN|21310-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0804104|T201|OSN|21310-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0804104|T201|LC|21310-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0804104|T201|LN|21310-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0804104|T201|MTH_LN|21310-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0804104|T201|DN|21310-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0804104|T201|OSN|21310-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0804104|T201|LC|21310-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941756|T201|LN|25663-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941756|T201|DN|25663-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941756|T201|MTH_LN|25663-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941756|T201|OSN|25663-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941756|T201|LC|25663-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941756|T201|LN|25663-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941756|T201|DN|25663-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941756|T201|MTH_LN|25663-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941756|T201|OSN|25663-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941756|T201|LC|25663-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941756|T201|LN|25663-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941756|T201|DN|25663-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941756|T201|MTH_LN|25663-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941756|T201|OSN|25663-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941756|T201|LC|25663-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941758|T201|LN|25665-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941758|T201|DN|25665-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941758|T201|MTH_LN|25665-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941758|T201|OSN|25665-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941758|T201|LC|25665-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941758|T201|LN|25665-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941758|T201|DN|25665-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941758|T201|MTH_LN|25665-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941758|T201|OSN|25665-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941758|T201|LC|25665-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941758|T201|LN|25665-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941758|T201|DN|25665-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941758|T201|MTH_LN|25665-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941758|T201|OSN|25665-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941758|T201|LC|25665-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945252|T201|LN|25666-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945252|T201|DN|25666-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945252|T201|OSN|25666-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945252|T201|MTH_LN|25666-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945252|T201|LC|25666-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945252|T201|LN|25666-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945252|T201|DN|25666-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945252|T201|OSN|25666-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945252|T201|MTH_LN|25666-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945252|T201|LC|25666-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945252|T201|LN|25666-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945252|T201|DN|25666-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945252|T201|OSN|25666-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945252|T201|MTH_LN|25666-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945252|T201|LC|25666-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941760|T201|LN|25668-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941760|T201|DN|25668-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941760|T201|MTH_LN|25668-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941760|T201|OSN|25668-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941760|T201|LC|25668-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941760|T201|LN|25668-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941760|T201|DN|25668-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941760|T201|MTH_LN|25668-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941760|T201|OSN|25668-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941760|T201|LC|25668-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941760|T201|LN|25668-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941760|T201|DN|25668-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941760|T201|MTH_LN|25668-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941760|T201|OSN|25668-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941760|T201|LC|25668-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941761|T201|LN|25669-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941761|T201|DN|25669-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941761|T201|MTH_LN|25669-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941761|T201|OSN|25669-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941761|T201|LC|25669-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941761|T201|LN|25669-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941761|T201|DN|25669-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941761|T201|MTH_LN|25669-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941761|T201|OSN|25669-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941761|T201|LC|25669-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941761|T201|LN|25669-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941761|T201|DN|25669-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941761|T201|MTH_LN|25669-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941761|T201|OSN|25669-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941761|T201|LC|25669-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941763|T201|LN|25671-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941763|T201|DN|25671-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941763|T201|MTH_LN|25671-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941763|T201|OSN|25671-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941763|T201|LC|25671-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941763|T201|LN|25671-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941763|T201|DN|25671-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941763|T201|MTH_LN|25671-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941763|T201|OSN|25671-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941763|T201|LC|25671-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941763|T201|LN|25671-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941763|T201|DN|25671-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941763|T201|MTH_LN|25671-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941763|T201|OSN|25671-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941763|T201|LC|25671-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941764|T201|LN|25672-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941764|T201|DN|25672-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941764|T201|MTH_LN|25672-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941764|T201|OSN|25672-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941764|T201|LC|25672-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941764|T201|LN|25672-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941764|T201|DN|25672-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941764|T201|MTH_LN|25672-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941764|T201|OSN|25672-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941764|T201|LC|25672-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941764|T201|LN|25672-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941764|T201|DN|25672-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941764|T201|MTH_LN|25672-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941764|T201|OSN|25672-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941764|T201|LC|25672-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941765|T201|LN|25673-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941765|T201|DN|25673-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941765|T201|MTH_LN|25673-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941765|T201|OSN|25673-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941765|T201|LC|25673-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941765|T201|LN|25673-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941765|T201|DN|25673-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941765|T201|MTH_LN|25673-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941765|T201|OSN|25673-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941765|T201|LC|25673-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941765|T201|LN|25673-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941765|T201|DN|25673-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941765|T201|MTH_LN|25673-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941765|T201|OSN|25673-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941765|T201|LC|25673-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941766|T201|LN|25674-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941766|T201|DN|25674-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941766|T201|MTH_LN|25674-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941766|T201|OSN|25674-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941766|T201|LC|25674-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941766|T201|LN|25674-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941766|T201|DN|25674-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941766|T201|MTH_LN|25674-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941766|T201|OSN|25674-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941766|T201|LC|25674-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941766|T201|LN|25674-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941766|T201|DN|25674-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941766|T201|MTH_LN|25674-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941766|T201|OSN|25674-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941766|T201|LC|25674-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941768|T201|LN|25676-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941768|T201|DN|25676-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941768|T201|MTH_LN|25676-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941768|T201|OSN|25676-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941768|T201|LC|25676-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941768|T201|LN|25676-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941768|T201|DN|25676-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941768|T201|MTH_LN|25676-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941768|T201|OSN|25676-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941768|T201|LC|25676-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941768|T201|LN|25676-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941768|T201|DN|25676-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941768|T201|MTH_LN|25676-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941768|T201|OSN|25676-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941768|T201|LC|25676-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941769|T201|LN|25677-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941769|T201|DN|25677-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941769|T201|MTH_LN|25677-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941769|T201|OSN|25677-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941769|T201|LC|25677-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941769|T201|LN|25677-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941769|T201|DN|25677-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941769|T201|MTH_LN|25677-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941769|T201|OSN|25677-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941769|T201|LC|25677-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941769|T201|LN|25677-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941769|T201|DN|25677-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941769|T201|MTH_LN|25677-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941769|T201|OSN|25677-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941769|T201|LC|25677-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941770|T201|LN|25679-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941770|T201|DN|25679-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941770|T201|OSN|25679-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941770|T201|MTH_LN|25679-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941770|T201|LC|25679-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941770|T201|LN|25679-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941770|T201|DN|25679-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941770|T201|OSN|25679-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941770|T201|MTH_LN|25679-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941770|T201|LC|25679-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941770|T201|LN|25679-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941770|T201|DN|25679-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941770|T201|OSN|25679-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941770|T201|MTH_LN|25679-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941770|T201|LC|25679-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941771|T201|LN|25680-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941771|T201|DN|25680-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941771|T201|MTH_LN|25680-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941771|T201|OSN|25680-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941771|T201|LC|25680-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0941771|T201|LN|25680-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941771|T201|DN|25680-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941771|T201|MTH_LN|25680-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941771|T201|OSN|25680-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941771|T201|LC|25680-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0941771|T201|LN|25680-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941771|T201|DN|25680-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941771|T201|MTH_LN|25680-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941771|T201|OSN|25680-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0941771|T201|LC|25680-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942492|T201|LN|26539-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942492|T201|DN|26539-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942492|T201|MTH_LN|26539-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942492|T201|OSN|26539-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942492|T201|LC|26539-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942492|T201|LN|26539-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942492|T201|DN|26539-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942492|T201|MTH_LN|26539-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942492|T201|OSN|26539-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942492|T201|LC|26539-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942492|T201|LN|26539-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942492|T201|DN|26539-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942492|T201|MTH_LN|26539-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942492|T201|OSN|26539-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942492|T201|LC|26539-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942494|T201|LN|26541-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942494|T201|DN|26541-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942494|T201|MTH_LN|26541-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942494|T201|OSN|26541-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942494|T201|LC|26541-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942494|T201|LN|26541-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942494|T201|DN|26541-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942494|T201|MTH_LN|26541-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942494|T201|OSN|26541-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942494|T201|LC|26541-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942494|T201|LN|26541-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942494|T201|DN|26541-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942494|T201|MTH_LN|26541-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942494|T201|OSN|26541-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942494|T201|LC|26541-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942496|T201|LN|26543-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942496|T201|DN|26543-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942496|T201|MTH_LN|26543-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942496|T201|OSN|26543-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942496|T201|LC|26543-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942496|T201|LN|26543-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942496|T201|DN|26543-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942496|T201|MTH_LN|26543-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942496|T201|OSN|26543-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942496|T201|LC|26543-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942496|T201|LN|26543-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942496|T201|DN|26543-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942496|T201|MTH_LN|26543-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942496|T201|OSN|26543-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942496|T201|LC|26543-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942497|T201|LN|26544-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942497|T201|DN|26544-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942497|T201|MTH_LN|26544-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942497|T201|OSN|26544-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942497|T201|LC|26544-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942497|T201|LN|26544-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942497|T201|DN|26544-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942497|T201|MTH_LN|26544-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942497|T201|OSN|26544-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942497|T201|LC|26544-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942497|T201|LN|26544-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942497|T201|DN|26544-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942497|T201|MTH_LN|26544-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942497|T201|OSN|26544-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942497|T201|LC|26544-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942506|T201|LN|26554-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942506|T201|DN|26554-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942506|T201|OSN|26554-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942506|T201|MTH_LN|26554-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942506|T201|LC|26554-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942506|T201|LN|26554-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942506|T201|DN|26554-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942506|T201|OSN|26554-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942506|T201|MTH_LN|26554-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942506|T201|LC|26554-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942506|T201|LN|26554-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942506|T201|DN|26554-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942506|T201|OSN|26554-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942506|T201|MTH_LN|26554-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942506|T201|LC|26554-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942507|T201|LN|26555-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942507|T201|DN|26555-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942507|T201|MTH_LN|26555-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942507|T201|OSN|26555-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942507|T201|LC|26555-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942507|T201|LN|26555-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942507|T201|DN|26555-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942507|T201|MTH_LN|26555-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942507|T201|OSN|26555-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942507|T201|LC|26555-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942507|T201|LN|26555-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942507|T201|DN|26555-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942507|T201|MTH_LN|26555-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942507|T201|OSN|26555-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942507|T201|LC|26555-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942624|T201|LN|26695-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942624|T201|DN|26695-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942624|T201|MTH_LN|26695-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942624|T201|OSN|26695-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942624|T201|LC|26695-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942624|T201|LN|26695-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942624|T201|DN|26695-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942624|T201|MTH_LN|26695-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942624|T201|OSN|26695-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942624|T201|LC|26695-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942624|T201|LN|26695-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942624|T201|DN|26695-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942624|T201|MTH_LN|26695-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942624|T201|OSN|26695-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942624|T201|LC|26695-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0947224|T201|LN|26777-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0947224|T201|DN|26777-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0947224|T201|MTH_LN|26777-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0947224|T201|OSN|26777-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0947224|T201|LC|26777-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0947224|T201|LN|26777-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0947224|T201|DN|26777-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0947224|T201|MTH_LN|26777-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0947224|T201|OSN|26777-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0947224|T201|LC|26777-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0947224|T201|LN|26777-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0947224|T201|DN|26777-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0947224|T201|MTH_LN|26777-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0947224|T201|OSN|26777-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0947224|T201|LC|26777-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942692|T201|LN|26778-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942692|T201|DN|26778-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942692|T201|MTH_LN|26778-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942692|T201|OSN|26778-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942692|T201|LC|26778-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942692|T201|LN|26778-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942692|T201|DN|26778-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942692|T201|MTH_LN|26778-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942692|T201|OSN|26778-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942692|T201|LC|26778-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942692|T201|LN|26778-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942692|T201|DN|26778-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942692|T201|MTH_LN|26778-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942692|T201|OSN|26778-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942692|T201|LC|26778-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945403|T201|LN|26779-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945403|T201|DN|26779-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945403|T201|OSN|26779-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945403|T201|MTH_LN|26779-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945403|T201|LC|26779-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945403|T201|LN|26779-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945403|T201|DN|26779-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945403|T201|OSN|26779-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945403|T201|MTH_LN|26779-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945403|T201|LC|26779-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945403|T201|LN|26779-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945403|T201|DN|26779-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945403|T201|OSN|26779-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945403|T201|MTH_LN|26779-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945403|T201|LC|26779-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942693|T201|LN|26780-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942693|T201|DN|26780-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942693|T201|MTH_LN|26780-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942693|T201|OSN|26780-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942693|T201|LC|26780-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942693|T201|LN|26780-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942693|T201|DN|26780-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942693|T201|MTH_LN|26780-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942693|T201|OSN|26780-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942693|T201|LC|26780-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942693|T201|LN|26780-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942693|T201|DN|26780-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942693|T201|MTH_LN|26780-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942693|T201|OSN|26780-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942693|T201|LC|26780-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0947225|T201|LN|26781-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0947225|T201|DN|26781-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0947225|T201|MTH_LN|26781-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0947225|T201|OSN|26781-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0947225|T201|LC|26781-5|LNC2HPO|Hyperglycemia|Hyperglycemia
C0947225|T201|LN|26781-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0947225|T201|DN|26781-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0947225|T201|MTH_LN|26781-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0947225|T201|OSN|26781-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0947225|T201|LC|26781-5|LNC2HPO|Hypoglycemia|Hypoglycemia
C0947225|T201|LN|26781-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0947225|T201|DN|26781-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0947225|T201|MTH_LN|26781-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0947225|T201|OSN|26781-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0947225|T201|LC|26781-5|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945404|T201|LN|26782-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945404|T201|DN|26782-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945404|T201|MTH_LN|26782-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945404|T201|OSN|26782-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945404|T201|LC|26782-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945404|T201|LN|26782-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945404|T201|DN|26782-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945404|T201|MTH_LN|26782-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945404|T201|OSN|26782-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945404|T201|LC|26782-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945404|T201|LN|26782-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945404|T201|DN|26782-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945404|T201|MTH_LN|26782-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945404|T201|OSN|26782-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945404|T201|LC|26782-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942694|T201|LN|26783-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942694|T201|DN|26783-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942694|T201|MTH_LN|26783-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942694|T201|OSN|26783-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942694|T201|LC|26783-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942694|T201|LN|26783-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942694|T201|DN|26783-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942694|T201|MTH_LN|26783-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942694|T201|OSN|26783-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942694|T201|LC|26783-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942694|T201|LN|26783-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942694|T201|DN|26783-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942694|T201|MTH_LN|26783-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942694|T201|OSN|26783-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942694|T201|LC|26783-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942723|T201|LN|26817-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942723|T201|DN|26817-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942723|T201|MTH_LN|26817-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942723|T201|OSN|26817-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942723|T201|LC|26817-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942723|T201|LN|26817-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942723|T201|DN|26817-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942723|T201|MTH_LN|26817-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942723|T201|OSN|26817-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942723|T201|LC|26817-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942723|T201|LN|26817-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942723|T201|DN|26817-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942723|T201|MTH_LN|26817-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942723|T201|OSN|26817-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942723|T201|LC|26817-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942751|T201|LN|26853-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942751|T201|DN|26853-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942751|T201|MTH_LN|26853-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942751|T201|OSN|26853-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942751|T201|LC|26853-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942751|T201|LN|26853-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942751|T201|DN|26853-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942751|T201|MTH_LN|26853-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942751|T201|OSN|26853-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942751|T201|LC|26853-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942751|T201|LN|26853-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942751|T201|DN|26853-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942751|T201|MTH_LN|26853-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942751|T201|OSN|26853-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942751|T201|LC|26853-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942752|T201|LN|26854-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942752|T201|DN|26854-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942752|T201|MTH_LN|26854-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942752|T201|OSN|26854-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942752|T201|LC|26854-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0942752|T201|LN|26854-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942752|T201|DN|26854-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942752|T201|MTH_LN|26854-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942752|T201|OSN|26854-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942752|T201|LC|26854-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0942752|T201|LN|26854-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942752|T201|DN|26854-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942752|T201|MTH_LN|26854-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942752|T201|OSN|26854-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0942752|T201|LC|26854-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945506|T201|LN|27432-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945506|T201|DN|27432-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945506|T201|MTH_LN|27432-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945506|T201|OSN|27432-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945506|T201|LC|27432-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945506|T201|LN|27432-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945506|T201|DN|27432-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945506|T201|MTH_LN|27432-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945506|T201|OSN|27432-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945506|T201|LC|27432-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945506|T201|LN|27432-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945506|T201|DN|27432-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945506|T201|MTH_LN|27432-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945506|T201|OSN|27432-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945506|T201|LC|27432-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0947266|T201|LN|29329-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0947266|T201|DN|29329-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0947266|T201|MTH_LN|29329-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0947266|T201|OSN|29329-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0947266|T201|LC|29329-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C0947266|T201|LN|29329-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0947266|T201|DN|29329-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0947266|T201|MTH_LN|29329-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0947266|T201|OSN|29329-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0947266|T201|LC|29329-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C0947266|T201|LN|29329-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0947266|T201|DN|29329-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0947266|T201|MTH_LN|29329-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0947266|T201|OSN|29329-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0947266|T201|LC|29329-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0944796|T201|LN|29330-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0944796|T201|DN|29330-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0944796|T201|MTH_LN|29330-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0944796|T201|OSN|29330-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0944796|T201|LC|29330-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0944796|T201|LN|29330-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0944796|T201|DN|29330-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0944796|T201|MTH_LN|29330-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0944796|T201|OSN|29330-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0944796|T201|LC|29330-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C0944796|T201|LN|29330-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0944796|T201|DN|29330-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0944796|T201|MTH_LN|29330-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0944796|T201|OSN|29330-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0944796|T201|LC|29330-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0944797|T201|LN|29331-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0944797|T201|DN|29331-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0944797|T201|MTH_LN|29331-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0944797|T201|OSN|29331-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0944797|T201|LC|29331-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0944797|T201|LN|29331-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0944797|T201|DN|29331-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0944797|T201|MTH_LN|29331-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0944797|T201|OSN|29331-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0944797|T201|LC|29331-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0944797|T201|LN|29331-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0944797|T201|DN|29331-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0944797|T201|MTH_LN|29331-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0944797|T201|OSN|29331-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0944797|T201|LC|29331-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0944798|T201|LN|29332-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0944798|T201|DN|29332-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0944798|T201|OSN|29332-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0944798|T201|MTH_LN|29332-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0944798|T201|LC|29332-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0944798|T201|LN|29332-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0944798|T201|DN|29332-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0944798|T201|OSN|29332-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0944798|T201|MTH_LN|29332-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0944798|T201|LC|29332-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0944798|T201|LN|29332-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0944798|T201|DN|29332-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0944798|T201|OSN|29332-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0944798|T201|MTH_LN|29332-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0944798|T201|LC|29332-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945746|T201|LN|29412-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945746|T201|DN|29412-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945746|T201|MTH_LN|29412-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945746|T201|OSN|29412-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945746|T201|LC|29412-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C0945746|T201|LN|29412-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945746|T201|DN|29412-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945746|T201|MTH_LN|29412-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945746|T201|OSN|29412-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945746|T201|LC|29412-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C0945746|T201|LN|29412-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945746|T201|DN|29412-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945746|T201|MTH_LN|29412-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945746|T201|OSN|29412-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0945746|T201|LC|29412-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114129|T201|LN|30251-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114129|T201|DN|30251-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114129|T201|MTH_LN|30251-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114129|T201|OSN|30251-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114129|T201|LC|30251-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114129|T201|LN|30251-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114129|T201|DN|30251-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114129|T201|MTH_LN|30251-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114129|T201|OSN|30251-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114129|T201|LC|30251-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114129|T201|LN|30251-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114129|T201|DN|30251-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114129|T201|MTH_LN|30251-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114129|T201|OSN|30251-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114129|T201|LC|30251-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114130|T201|LN|30252-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114130|T201|DN|30252-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114130|T201|MTH_LN|30252-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114130|T201|OSN|30252-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114130|T201|LC|30252-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114130|T201|LN|30252-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114130|T201|DN|30252-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114130|T201|MTH_LN|30252-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114130|T201|OSN|30252-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114130|T201|LC|30252-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114130|T201|LN|30252-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114130|T201|DN|30252-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114130|T201|MTH_LN|30252-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114130|T201|OSN|30252-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114130|T201|LC|30252-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114131|T201|LN|30253-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114131|T201|DN|30253-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114131|T201|MTH_LN|30253-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114131|T201|OSN|30253-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114131|T201|LC|30253-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114131|T201|LN|30253-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114131|T201|DN|30253-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114131|T201|MTH_LN|30253-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114131|T201|OSN|30253-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114131|T201|LC|30253-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114131|T201|LN|30253-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114131|T201|DN|30253-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114131|T201|MTH_LN|30253-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114131|T201|OSN|30253-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114131|T201|LC|30253-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114140|T201|LN|30263-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114140|T201|DN|30263-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114140|T201|MTH_LN|30263-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114140|T201|OSN|30263-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114140|T201|LC|30263-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114140|T201|LN|30263-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114140|T201|DN|30263-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114140|T201|MTH_LN|30263-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114140|T201|OSN|30263-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114140|T201|LC|30263-8|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114140|T201|LN|30263-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114140|T201|DN|30263-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114140|T201|MTH_LN|30263-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114140|T201|OSN|30263-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114140|T201|LC|30263-8|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114881|T201|LN|30264-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114881|T201|DN|30264-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114881|T201|MTH_LN|30264-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114881|T201|OSN|30264-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114881|T201|LC|30264-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114881|T201|LN|30264-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114881|T201|DN|30264-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114881|T201|MTH_LN|30264-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114881|T201|OSN|30264-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114881|T201|LC|30264-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114881|T201|LN|30264-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114881|T201|DN|30264-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114881|T201|MTH_LN|30264-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114881|T201|OSN|30264-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114881|T201|LC|30264-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114141|T201|LN|30265-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114141|T201|DN|30265-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114141|T201|MTH_LN|30265-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114141|T201|OSN|30265-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114141|T201|LC|30265-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114141|T201|LN|30265-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114141|T201|DN|30265-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114141|T201|MTH_LN|30265-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114141|T201|OSN|30265-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114141|T201|LC|30265-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114141|T201|LN|30265-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114141|T201|DN|30265-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114141|T201|MTH_LN|30265-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114141|T201|OSN|30265-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114141|T201|LC|30265-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114882|T201|LN|30266-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114882|T201|DN|30266-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114882|T201|MTH_LN|30266-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114882|T201|OSN|30266-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114882|T201|LC|30266-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114882|T201|LN|30266-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114882|T201|DN|30266-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114882|T201|MTH_LN|30266-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114882|T201|OSN|30266-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114882|T201|LC|30266-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114882|T201|LN|30266-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114882|T201|DN|30266-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114882|T201|MTH_LN|30266-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114882|T201|OSN|30266-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114882|T201|LC|30266-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114142|T201|LN|30267-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114142|T201|DN|30267-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114142|T201|MTH_LN|30267-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114142|T201|OSN|30267-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114142|T201|LC|30267-9|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114142|T201|LN|30267-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114142|T201|DN|30267-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114142|T201|MTH_LN|30267-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114142|T201|OSN|30267-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114142|T201|LC|30267-9|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114142|T201|LN|30267-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114142|T201|DN|30267-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114142|T201|MTH_LN|30267-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114142|T201|OSN|30267-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114142|T201|LC|30267-9|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114209|T201|LN|30344-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114209|T201|DN|30344-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114209|T201|MTH_LN|30344-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114209|T201|OSN|30344-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114209|T201|LC|30344-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114209|T201|LN|30344-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114209|T201|DN|30344-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114209|T201|MTH_LN|30344-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114209|T201|OSN|30344-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114209|T201|LC|30344-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114209|T201|LN|30344-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114209|T201|DN|30344-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114209|T201|MTH_LN|30344-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114209|T201|OSN|30344-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114209|T201|LC|30344-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114210|T201|LN|30345-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114210|T201|DN|30345-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114210|T201|MTH_LN|30345-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114210|T201|OSN|30345-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114210|T201|LC|30345-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114210|T201|LN|30345-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114210|T201|DN|30345-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114210|T201|MTH_LN|30345-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114210|T201|OSN|30345-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114210|T201|LC|30345-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114210|T201|LN|30345-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114210|T201|DN|30345-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114210|T201|MTH_LN|30345-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114210|T201|OSN|30345-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114210|T201|LC|30345-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114892|T201|LN|30346-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114892|T201|DN|30346-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114892|T201|MTH_LN|30346-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114892|T201|OSN|30346-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114892|T201|LC|30346-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C1114892|T201|LN|30346-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114892|T201|DN|30346-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114892|T201|MTH_LN|30346-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114892|T201|OSN|30346-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114892|T201|LC|30346-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C1114892|T201|LN|30346-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114892|T201|DN|30346-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114892|T201|MTH_LN|30346-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114892|T201|OSN|30346-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1114892|T201|LC|30346-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148003|T201|LN|32319-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148003|T201|DN|32319-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148003|T201|MTH_LN|32319-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148003|T201|OSN|32319-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148003|T201|LC|32319-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148003|T201|LN|32319-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148003|T201|DN|32319-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148003|T201|MTH_LN|32319-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148003|T201|OSN|32319-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148003|T201|LC|32319-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148003|T201|LN|32319-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148003|T201|DN|32319-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148003|T201|MTH_LN|32319-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148003|T201|OSN|32319-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148003|T201|LC|32319-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148004|T201|LN|32320-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148004|T201|DN|32320-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148004|T201|MTH_LN|32320-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148004|T201|OSN|32320-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148004|T201|LC|32320-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148004|T201|LN|32320-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148004|T201|DN|32320-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148004|T201|MTH_LN|32320-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148004|T201|OSN|32320-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148004|T201|LC|32320-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148004|T201|LN|32320-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148004|T201|DN|32320-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148004|T201|MTH_LN|32320-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148004|T201|OSN|32320-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148004|T201|LC|32320-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148005|T201|LN|32321-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148005|T201|DN|32321-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148005|T201|MTH_LN|32321-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148005|T201|OSN|32321-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148005|T201|LC|32321-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148005|T201|LN|32321-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148005|T201|DN|32321-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148005|T201|MTH_LN|32321-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148005|T201|OSN|32321-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148005|T201|LC|32321-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148005|T201|LN|32321-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148005|T201|DN|32321-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148005|T201|MTH_LN|32321-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148005|T201|OSN|32321-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148005|T201|LC|32321-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148006|T201|LN|32322-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148006|T201|DN|32322-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148006|T201|MTH_LN|32322-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148006|T201|OSN|32322-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148006|T201|LC|32322-0|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148006|T201|LN|32322-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148006|T201|DN|32322-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148006|T201|MTH_LN|32322-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148006|T201|OSN|32322-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148006|T201|LC|32322-0|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148006|T201|LN|32322-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148006|T201|DN|32322-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148006|T201|MTH_LN|32322-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148006|T201|OSN|32322-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148006|T201|LC|32322-0|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148043|T201|LN|32359-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148043|T201|DN|32359-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148043|T201|MTH_LN|32359-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148043|T201|OSN|32359-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148043|T201|LC|32359-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C1148043|T201|LN|32359-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148043|T201|DN|32359-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148043|T201|MTH_LN|32359-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148043|T201|OSN|32359-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148043|T201|LC|32359-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C1148043|T201|LN|32359-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148043|T201|DN|32359-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148043|T201|MTH_LN|32359-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148043|T201|OSN|32359-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1148043|T201|LC|32359-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1315291|T201|LN|32820-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C1315291|T201|DN|32820-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C1315291|T201|MTH_LN|32820-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C1315291|T201|OSN|32820-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C1315291|T201|LC|32820-3|LNC2HPO|Hyperglycemia|Hyperglycemia
C1315291|T201|LN|32820-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C1315291|T201|DN|32820-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C1315291|T201|MTH_LN|32820-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C1315291|T201|OSN|32820-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C1315291|T201|LC|32820-3|LNC2HPO|Hypoglycemia|Hypoglycemia
C1315291|T201|LN|32820-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1315291|T201|DN|32820-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1315291|T201|MTH_LN|32820-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1315291|T201|OSN|32820-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1315291|T201|LC|32820-3|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1315495|T201|LN|33024-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C1315495|T201|DN|33024-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C1315495|T201|MTH_LN|33024-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C1315495|T201|OSN|33024-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C1315495|T201|LC|33024-1|LNC2HPO|Hyperglycemia|Hyperglycemia
C1315495|T201|LN|33024-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C1315495|T201|DN|33024-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C1315495|T201|MTH_LN|33024-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C1315495|T201|OSN|33024-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C1315495|T201|LC|33024-1|LNC2HPO|Hypoglycemia|Hypoglycemia
C1315495|T201|LN|33024-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1315495|T201|DN|33024-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1315495|T201|MTH_LN|33024-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1315495|T201|OSN|33024-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1315495|T201|LC|33024-1|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C2607836|T201|MTH_LN|35211-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C2607836|T201|DN|35211-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C2607836|T201|LN|35211-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C2607836|T201|OSN|35211-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C2607836|T201|LC|35211-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C2607836|T201|MTH_LN|35211-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C2607836|T201|DN|35211-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C2607836|T201|LN|35211-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C2607836|T201|OSN|35211-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C2607836|T201|LC|35211-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C2607836|T201|MTH_LN|35211-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C2607836|T201|DN|35211-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C2607836|T201|LN|35211-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C2607836|T201|OSN|35211-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C2607836|T201|LC|35211-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1543636|T201|LN|39561-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C1543636|T201|DN|39561-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C1543636|T201|MTH_LN|39561-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C1543636|T201|OSN|39561-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C1543636|T201|LC|39561-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C1543636|T201|LN|39561-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C1543636|T201|DN|39561-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C1543636|T201|MTH_LN|39561-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C1543636|T201|OSN|39561-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C1543636|T201|LC|39561-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C1543636|T201|LN|39561-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1543636|T201|DN|39561-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1543636|T201|MTH_LN|39561-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1543636|T201|OSN|39561-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1543636|T201|LC|39561-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1543637|T201|LN|39562-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C1543637|T201|DN|39562-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C1543637|T201|MTH_LN|39562-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C1543637|T201|OSN|39562-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C1543637|T201|LC|39562-4|LNC2HPO|Hyperglycemia|Hyperglycemia
C1543637|T201|LN|39562-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C1543637|T201|DN|39562-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C1543637|T201|MTH_LN|39562-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C1543637|T201|OSN|39562-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C1543637|T201|LC|39562-4|LNC2HPO|Hypoglycemia|Hypoglycemia
C1543637|T201|LN|39562-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1543637|T201|DN|39562-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1543637|T201|MTH_LN|39562-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1543637|T201|OSN|39562-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1543637|T201|LC|39562-4|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1543638|T201|LN|39563-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C1543638|T201|DN|39563-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C1543638|T201|MTH_LN|39563-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C1543638|T201|OSN|39563-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C1543638|T201|LC|39563-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C1543638|T201|LN|39563-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C1543638|T201|DN|39563-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C1543638|T201|MTH_LN|39563-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C1543638|T201|OSN|39563-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C1543638|T201|LC|39563-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C1543638|T201|LN|39563-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1543638|T201|DN|39563-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1543638|T201|MTH_LN|39563-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1543638|T201|OSN|39563-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1543638|T201|LC|39563-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0484416|T201|LN|7789-1|LNC2HPO|Acanthocytosis|Acanthocytosis
C0484416|T201|MTH_LN|7789-1|LNC2HPO|Acanthocytosis|Acanthocytosis
C0484416|T201|DN|7789-1|LNC2HPO|Acanthocytosis|Acanthocytosis
C0484416|T201|OSN|7789-1|LNC2HPO|Acanthocytosis|Acanthocytosis
C0484416|T201|LC|7789-1|LNC2HPO|Acanthocytosis|Acanthocytosis
C0484416|T201|LN|7789-1|LNC2HPO|Acanthocytes|Acanthocytes
C0484416|T201|MTH_LN|7789-1|LNC2HPO|Acanthocytes|Acanthocytes
C0484416|T201|DN|7789-1|LNC2HPO|Acanthocytes|Acanthocytes
C0484416|T201|OSN|7789-1|LNC2HPO|Acanthocytes|Acanthocytes
C0484416|T201|LC|7789-1|LNC2HPO|Acanthocytes|Acanthocytes
C0484416|T201|LN|7789-1|LNC2HPO|Red cell acanthocytosis|Red cell acanthocytosis
C0484416|T201|MTH_LN|7789-1|LNC2HPO|Red cell acanthocytosis|Red cell acanthocytosis
C0484416|T201|DN|7789-1|LNC2HPO|Red cell acanthocytosis|Red cell acanthocytosis
C0484416|T201|OSN|7789-1|LNC2HPO|Red cell acanthocytosis|Red cell acanthocytosis
C0484416|T201|LC|7789-1|LNC2HPO|Red cell acanthocytosis|Red cell acanthocytosis
C0801529|T201|LC|18488-7|LNC2HPO|Hypercalciuria|Hypercalciuria
C0801529|T201|MTH_LN|18488-7|LNC2HPO|Hypercalciuria|Hypercalciuria
C0801529|T201|DN|18488-7|LNC2HPO|Hypercalciuria|Hypercalciuria
C0801529|T201|OSN|18488-7|LNC2HPO|Hypercalciuria|Hypercalciuria
C0801529|T201|LN|18488-7|LNC2HPO|Hypercalciuria|Hypercalciuria
C0801529|T201|LC|18488-7|LNC2HPO|Hypercalcinuria|Hypercalcinuria
C0801529|T201|MTH_LN|18488-7|LNC2HPO|Hypercalcinuria|Hypercalcinuria
C0801529|T201|DN|18488-7|LNC2HPO|Hypercalcinuria|Hypercalcinuria
C0801529|T201|OSN|18488-7|LNC2HPO|Hypercalcinuria|Hypercalcinuria
C0801529|T201|LN|18488-7|LNC2HPO|Hypercalcinuria|Hypercalcinuria
C0801529|T201|LC|18488-7|LNC2HPO|Hypocalciuria|Hypocalciuria
C0801529|T201|MTH_LN|18488-7|LNC2HPO|Hypocalciuria|Hypocalciuria
C0801529|T201|DN|18488-7|LNC2HPO|Hypocalciuria|Hypocalciuria
C0801529|T201|OSN|18488-7|LNC2HPO|Hypocalciuria|Hypocalciuria
C0801529|T201|LN|18488-7|LNC2HPO|Hypocalciuria|Hypocalciuria
C0550042|T201|LN|12448-7|LNC2HPO|Ketonuria|Ketonuria
C0550042|T201|MTH_LN|12448-7|LNC2HPO|Ketonuria|Ketonuria
C0550042|T201|DN|12448-7|LNC2HPO|Ketonuria|Ketonuria
C0550042|T201|OSN|12448-7|LNC2HPO|Ketonuria|Ketonuria
C0550042|T201|LC|12448-7|LNC2HPO|Ketonuria|Ketonuria
C0550042|T201|LN|12448-7|LNC2HPO|Acetonuria|Acetonuria
C0550042|T201|MTH_LN|12448-7|LNC2HPO|Acetonuria|Acetonuria
C0550042|T201|DN|12448-7|LNC2HPO|Acetonuria|Acetonuria
C0550042|T201|OSN|12448-7|LNC2HPO|Acetonuria|Acetonuria
C0550042|T201|LC|12448-7|LNC2HPO|Acetonuria|Acetonuria
C0550042|T201|LN|12448-7|LNC2HPO|Ketoaciduria|Ketoaciduria
C0550042|T201|MTH_LN|12448-7|LNC2HPO|Ketoaciduria|Ketoaciduria
C0550042|T201|DN|12448-7|LNC2HPO|Ketoaciduria|Ketoaciduria
C0550042|T201|OSN|12448-7|LNC2HPO|Ketoaciduria|Ketoaciduria
C0550042|T201|LC|12448-7|LNC2HPO|Ketoaciduria|Ketoaciduria
C0550042|T201|LN|12448-7|LNC2HPO|Ketonaciduria|Ketonaciduria
C0550042|T201|MTH_LN|12448-7|LNC2HPO|Ketonaciduria|Ketonaciduria
C0550042|T201|DN|12448-7|LNC2HPO|Ketonaciduria|Ketonaciduria
C0550042|T201|OSN|12448-7|LNC2HPO|Ketonaciduria|Ketonaciduria
C0550042|T201|LC|12448-7|LNC2HPO|Ketonaciduria|Ketonaciduria
C0550043|T201|LN|12449-5|LNC2HPO|Ketonuria|Ketonuria
C0550043|T201|MTH_LN|12449-5|LNC2HPO|Ketonuria|Ketonuria
C0550043|T201|DN|12449-5|LNC2HPO|Ketonuria|Ketonuria
C0550043|T201|OSN|12449-5|LNC2HPO|Ketonuria|Ketonuria
C0550043|T201|LC|12449-5|LNC2HPO|Ketonuria|Ketonuria
C0550043|T201|LN|12449-5|LNC2HPO|Acetonuria|Acetonuria
C0550043|T201|MTH_LN|12449-5|LNC2HPO|Acetonuria|Acetonuria
C0550043|T201|DN|12449-5|LNC2HPO|Acetonuria|Acetonuria
C0550043|T201|OSN|12449-5|LNC2HPO|Acetonuria|Acetonuria
C0550043|T201|LC|12449-5|LNC2HPO|Acetonuria|Acetonuria
C0550043|T201|LN|12449-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C0550043|T201|MTH_LN|12449-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C0550043|T201|DN|12449-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C0550043|T201|OSN|12449-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C0550043|T201|LC|12449-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C0550043|T201|LN|12449-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C0550043|T201|MTH_LN|12449-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C0550043|T201|DN|12449-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C0550043|T201|OSN|12449-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C0550043|T201|LC|12449-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C0550044|T201|LN|12450-3|LNC2HPO|Ketonuria|Ketonuria
C0550044|T201|MTH_LN|12450-3|LNC2HPO|Ketonuria|Ketonuria
C0550044|T201|DN|12450-3|LNC2HPO|Ketonuria|Ketonuria
C0550044|T201|OSN|12450-3|LNC2HPO|Ketonuria|Ketonuria
C0550044|T201|LC|12450-3|LNC2HPO|Ketonuria|Ketonuria
C0550044|T201|LN|12450-3|LNC2HPO|Acetonuria|Acetonuria
C0550044|T201|MTH_LN|12450-3|LNC2HPO|Acetonuria|Acetonuria
C0550044|T201|DN|12450-3|LNC2HPO|Acetonuria|Acetonuria
C0550044|T201|OSN|12450-3|LNC2HPO|Acetonuria|Acetonuria
C0550044|T201|LC|12450-3|LNC2HPO|Acetonuria|Acetonuria
C0550044|T201|LN|12450-3|LNC2HPO|Ketoaciduria|Ketoaciduria
C0550044|T201|MTH_LN|12450-3|LNC2HPO|Ketoaciduria|Ketoaciduria
C0550044|T201|DN|12450-3|LNC2HPO|Ketoaciduria|Ketoaciduria
C0550044|T201|OSN|12450-3|LNC2HPO|Ketoaciduria|Ketoaciduria
C0550044|T201|LC|12450-3|LNC2HPO|Ketoaciduria|Ketoaciduria
C0550044|T201|LN|12450-3|LNC2HPO|Ketonaciduria|Ketonaciduria
C0550044|T201|MTH_LN|12450-3|LNC2HPO|Ketonaciduria|Ketonaciduria
C0550044|T201|DN|12450-3|LNC2HPO|Ketonaciduria|Ketonaciduria
C0550044|T201|OSN|12450-3|LNC2HPO|Ketonaciduria|Ketonaciduria
C0550044|T201|LC|12450-3|LNC2HPO|Ketonaciduria|Ketonaciduria
C0550045|T201|LN|12451-1|LNC2HPO|Ketonuria|Ketonuria
C0550045|T201|MTH_LN|12451-1|LNC2HPO|Ketonuria|Ketonuria
C0550045|T201|DN|12451-1|LNC2HPO|Ketonuria|Ketonuria
C0550045|T201|OSN|12451-1|LNC2HPO|Ketonuria|Ketonuria
C0550045|T201|LC|12451-1|LNC2HPO|Ketonuria|Ketonuria
C0550045|T201|LN|12451-1|LNC2HPO|Acetonuria|Acetonuria
C0550045|T201|MTH_LN|12451-1|LNC2HPO|Acetonuria|Acetonuria
C0550045|T201|DN|12451-1|LNC2HPO|Acetonuria|Acetonuria
C0550045|T201|OSN|12451-1|LNC2HPO|Acetonuria|Acetonuria
C0550045|T201|LC|12451-1|LNC2HPO|Acetonuria|Acetonuria
C0550045|T201|LN|12451-1|LNC2HPO|Ketoaciduria|Ketoaciduria
C0550045|T201|MTH_LN|12451-1|LNC2HPO|Ketoaciduria|Ketoaciduria
C0550045|T201|DN|12451-1|LNC2HPO|Ketoaciduria|Ketoaciduria
C0550045|T201|OSN|12451-1|LNC2HPO|Ketoaciduria|Ketoaciduria
C0550045|T201|LC|12451-1|LNC2HPO|Ketoaciduria|Ketoaciduria
C0550045|T201|LN|12451-1|LNC2HPO|Ketonaciduria|Ketonaciduria
C0550045|T201|MTH_LN|12451-1|LNC2HPO|Ketonaciduria|Ketonaciduria
C0550045|T201|DN|12451-1|LNC2HPO|Ketonaciduria|Ketonaciduria
C0550045|T201|OSN|12451-1|LNC2HPO|Ketonaciduria|Ketonaciduria
C0550045|T201|LC|12451-1|LNC2HPO|Ketonaciduria|Ketonaciduria
C0797324|T201|LN|14138-2|LNC2HPO|Ketonuria|Ketonuria
C0797324|T201|MTH_LN|14138-2|LNC2HPO|Ketonuria|Ketonuria
C0797324|T201|DN|14138-2|LNC2HPO|Ketonuria|Ketonuria
C0797324|T201|OSN|14138-2|LNC2HPO|Ketonuria|Ketonuria
C0797324|T201|LC|14138-2|LNC2HPO|Ketonuria|Ketonuria
C0797324|T201|LN|14138-2|LNC2HPO|Acetonuria|Acetonuria
C0797324|T201|MTH_LN|14138-2|LNC2HPO|Acetonuria|Acetonuria
C0797324|T201|DN|14138-2|LNC2HPO|Acetonuria|Acetonuria
C0797324|T201|OSN|14138-2|LNC2HPO|Acetonuria|Acetonuria
C0797324|T201|LC|14138-2|LNC2HPO|Acetonuria|Acetonuria
C0797324|T201|LN|14138-2|LNC2HPO|Ketoaciduria|Ketoaciduria
C0797324|T201|MTH_LN|14138-2|LNC2HPO|Ketoaciduria|Ketoaciduria
C0797324|T201|DN|14138-2|LNC2HPO|Ketoaciduria|Ketoaciduria
C0797324|T201|OSN|14138-2|LNC2HPO|Ketoaciduria|Ketoaciduria
C0797324|T201|LC|14138-2|LNC2HPO|Ketoaciduria|Ketoaciduria
C0797324|T201|LN|14138-2|LNC2HPO|Ketonaciduria|Ketonaciduria
C0797324|T201|MTH_LN|14138-2|LNC2HPO|Ketonaciduria|Ketonaciduria
C0797324|T201|DN|14138-2|LNC2HPO|Ketonaciduria|Ketonaciduria
C0797324|T201|OSN|14138-2|LNC2HPO|Ketonaciduria|Ketonaciduria
C0797324|T201|LC|14138-2|LNC2HPO|Ketonaciduria|Ketonaciduria
C0797325|T201|LN|14139-0|LNC2HPO|Ketonuria|Ketonuria
C0797325|T201|MTH_LN|14139-0|LNC2HPO|Ketonuria|Ketonuria
C0797325|T201|DN|14139-0|LNC2HPO|Ketonuria|Ketonuria
C0797325|T201|OSN|14139-0|LNC2HPO|Ketonuria|Ketonuria
C0797325|T201|LC|14139-0|LNC2HPO|Ketonuria|Ketonuria
C0797325|T201|LN|14139-0|LNC2HPO|Acetonuria|Acetonuria
C0797325|T201|MTH_LN|14139-0|LNC2HPO|Acetonuria|Acetonuria
C0797325|T201|DN|14139-0|LNC2HPO|Acetonuria|Acetonuria
C0797325|T201|OSN|14139-0|LNC2HPO|Acetonuria|Acetonuria
C0797325|T201|LC|14139-0|LNC2HPO|Acetonuria|Acetonuria
C0797325|T201|LN|14139-0|LNC2HPO|Ketoaciduria|Ketoaciduria
C0797325|T201|MTH_LN|14139-0|LNC2HPO|Ketoaciduria|Ketoaciduria
C0797325|T201|DN|14139-0|LNC2HPO|Ketoaciduria|Ketoaciduria
C0797325|T201|OSN|14139-0|LNC2HPO|Ketoaciduria|Ketoaciduria
C0797325|T201|LC|14139-0|LNC2HPO|Ketoaciduria|Ketoaciduria
C0797325|T201|LN|14139-0|LNC2HPO|Ketonaciduria|Ketonaciduria
C0797325|T201|MTH_LN|14139-0|LNC2HPO|Ketonaciduria|Ketonaciduria
C0797325|T201|DN|14139-0|LNC2HPO|Ketonaciduria|Ketonaciduria
C0797325|T201|OSN|14139-0|LNC2HPO|Ketonaciduria|Ketonaciduria
C0797325|T201|LC|14139-0|LNC2HPO|Ketonaciduria|Ketonaciduria
C0797326|T201|LN|14140-8|LNC2HPO|Ketonuria|Ketonuria
C0797326|T201|MTH_LN|14140-8|LNC2HPO|Ketonuria|Ketonuria
C0797326|T201|DN|14140-8|LNC2HPO|Ketonuria|Ketonuria
C0797326|T201|OSN|14140-8|LNC2HPO|Ketonuria|Ketonuria
C0797326|T201|LC|14140-8|LNC2HPO|Ketonuria|Ketonuria
C0797326|T201|LN|14140-8|LNC2HPO|Acetonuria|Acetonuria
C0797326|T201|MTH_LN|14140-8|LNC2HPO|Acetonuria|Acetonuria
C0797326|T201|DN|14140-8|LNC2HPO|Acetonuria|Acetonuria
C0797326|T201|OSN|14140-8|LNC2HPO|Acetonuria|Acetonuria
C0797326|T201|LC|14140-8|LNC2HPO|Acetonuria|Acetonuria
C0797326|T201|LN|14140-8|LNC2HPO|Ketoaciduria|Ketoaciduria
C0797326|T201|MTH_LN|14140-8|LNC2HPO|Ketoaciduria|Ketoaciduria
C0797326|T201|DN|14140-8|LNC2HPO|Ketoaciduria|Ketoaciduria
C0797326|T201|OSN|14140-8|LNC2HPO|Ketoaciduria|Ketoaciduria
C0797326|T201|LC|14140-8|LNC2HPO|Ketoaciduria|Ketoaciduria
C0797326|T201|LN|14140-8|LNC2HPO|Ketonaciduria|Ketonaciduria
C0797326|T201|MTH_LN|14140-8|LNC2HPO|Ketonaciduria|Ketonaciduria
C0797326|T201|DN|14140-8|LNC2HPO|Ketonaciduria|Ketonaciduria
C0797326|T201|OSN|14140-8|LNC2HPO|Ketonaciduria|Ketonaciduria
C0797326|T201|LC|14140-8|LNC2HPO|Ketonaciduria|Ketonaciduria
C0797327|T201|LN|14141-6|LNC2HPO|Ketonuria|Ketonuria
C0797327|T201|MTH_LN|14141-6|LNC2HPO|Ketonuria|Ketonuria
C0797327|T201|DN|14141-6|LNC2HPO|Ketonuria|Ketonuria
C0797327|T201|OSN|14141-6|LNC2HPO|Ketonuria|Ketonuria
C0797327|T201|LC|14141-6|LNC2HPO|Ketonuria|Ketonuria
C0797327|T201|LN|14141-6|LNC2HPO|Acetonuria|Acetonuria
C0797327|T201|MTH_LN|14141-6|LNC2HPO|Acetonuria|Acetonuria
C0797327|T201|DN|14141-6|LNC2HPO|Acetonuria|Acetonuria
C0797327|T201|OSN|14141-6|LNC2HPO|Acetonuria|Acetonuria
C0797327|T201|LC|14141-6|LNC2HPO|Acetonuria|Acetonuria
C0797327|T201|LN|14141-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C0797327|T201|MTH_LN|14141-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C0797327|T201|DN|14141-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C0797327|T201|OSN|14141-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C0797327|T201|LC|14141-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C0797327|T201|LN|14141-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C0797327|T201|MTH_LN|14141-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C0797327|T201|DN|14141-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C0797327|T201|OSN|14141-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C0797327|T201|LC|14141-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C0804149|T201|LN|21355-3|LNC2HPO|Ketonuria|Ketonuria
C0804149|T201|MTH_LN|21355-3|LNC2HPO|Ketonuria|Ketonuria
C0804149|T201|DN|21355-3|LNC2HPO|Ketonuria|Ketonuria
C0804149|T201|OSN|21355-3|LNC2HPO|Ketonuria|Ketonuria
C0804149|T201|LC|21355-3|LNC2HPO|Ketonuria|Ketonuria
C0804149|T201|LN|21355-3|LNC2HPO|Acetonuria|Acetonuria
C0804149|T201|MTH_LN|21355-3|LNC2HPO|Acetonuria|Acetonuria
C0804149|T201|DN|21355-3|LNC2HPO|Acetonuria|Acetonuria
C0804149|T201|OSN|21355-3|LNC2HPO|Acetonuria|Acetonuria
C0804149|T201|LC|21355-3|LNC2HPO|Acetonuria|Acetonuria
C0804149|T201|LN|21355-3|LNC2HPO|Ketoaciduria|Ketoaciduria
C0804149|T201|MTH_LN|21355-3|LNC2HPO|Ketoaciduria|Ketoaciduria
C0804149|T201|DN|21355-3|LNC2HPO|Ketoaciduria|Ketoaciduria
C0804149|T201|OSN|21355-3|LNC2HPO|Ketoaciduria|Ketoaciduria
C0804149|T201|LC|21355-3|LNC2HPO|Ketoaciduria|Ketoaciduria
C0804149|T201|LN|21355-3|LNC2HPO|Ketonaciduria|Ketonaciduria
C0804149|T201|MTH_LN|21355-3|LNC2HPO|Ketonaciduria|Ketonaciduria
C0804149|T201|DN|21355-3|LNC2HPO|Ketonaciduria|Ketonaciduria
C0804149|T201|OSN|21355-3|LNC2HPO|Ketonaciduria|Ketonaciduria
C0804149|T201|LC|21355-3|LNC2HPO|Ketonaciduria|Ketonaciduria
C0804150|T201|LN|21356-1|LNC2HPO|Ketonuria|Ketonuria
C0804150|T201|MTH_LN|21356-1|LNC2HPO|Ketonuria|Ketonuria
C0804150|T201|DN|21356-1|LNC2HPO|Ketonuria|Ketonuria
C0804150|T201|OSN|21356-1|LNC2HPO|Ketonuria|Ketonuria
C0804150|T201|LC|21356-1|LNC2HPO|Ketonuria|Ketonuria
C0804150|T201|LN|21356-1|LNC2HPO|Acetonuria|Acetonuria
C0804150|T201|MTH_LN|21356-1|LNC2HPO|Acetonuria|Acetonuria
C0804150|T201|DN|21356-1|LNC2HPO|Acetonuria|Acetonuria
C0804150|T201|OSN|21356-1|LNC2HPO|Acetonuria|Acetonuria
C0804150|T201|LC|21356-1|LNC2HPO|Acetonuria|Acetonuria
C0804150|T201|LN|21356-1|LNC2HPO|Ketoaciduria|Ketoaciduria
C0804150|T201|MTH_LN|21356-1|LNC2HPO|Ketoaciduria|Ketoaciduria
C0804150|T201|DN|21356-1|LNC2HPO|Ketoaciduria|Ketoaciduria
C0804150|T201|OSN|21356-1|LNC2HPO|Ketoaciduria|Ketoaciduria
C0804150|T201|LC|21356-1|LNC2HPO|Ketoaciduria|Ketoaciduria
C0804150|T201|LN|21356-1|LNC2HPO|Ketonaciduria|Ketonaciduria
C0804150|T201|MTH_LN|21356-1|LNC2HPO|Ketonaciduria|Ketonaciduria
C0804150|T201|DN|21356-1|LNC2HPO|Ketonaciduria|Ketonaciduria
C0804150|T201|OSN|21356-1|LNC2HPO|Ketonaciduria|Ketonaciduria
C0804150|T201|LC|21356-1|LNC2HPO|Ketonaciduria|Ketonaciduria
C0804151|T201|LN|21357-9|LNC2HPO|Ketonuria|Ketonuria
C0804151|T201|MTH_LN|21357-9|LNC2HPO|Ketonuria|Ketonuria
C0804151|T201|DN|21357-9|LNC2HPO|Ketonuria|Ketonuria
C0804151|T201|OSN|21357-9|LNC2HPO|Ketonuria|Ketonuria
C0804151|T201|LC|21357-9|LNC2HPO|Ketonuria|Ketonuria
C0804151|T201|LN|21357-9|LNC2HPO|Acetonuria|Acetonuria
C0804151|T201|MTH_LN|21357-9|LNC2HPO|Acetonuria|Acetonuria
C0804151|T201|DN|21357-9|LNC2HPO|Acetonuria|Acetonuria
C0804151|T201|OSN|21357-9|LNC2HPO|Acetonuria|Acetonuria
C0804151|T201|LC|21357-9|LNC2HPO|Acetonuria|Acetonuria
C0804151|T201|LN|21357-9|LNC2HPO|Ketoaciduria|Ketoaciduria
C0804151|T201|MTH_LN|21357-9|LNC2HPO|Ketoaciduria|Ketoaciduria
C0804151|T201|DN|21357-9|LNC2HPO|Ketoaciduria|Ketoaciduria
C0804151|T201|OSN|21357-9|LNC2HPO|Ketoaciduria|Ketoaciduria
C0804151|T201|LC|21357-9|LNC2HPO|Ketoaciduria|Ketoaciduria
C0804151|T201|LN|21357-9|LNC2HPO|Ketonaciduria|Ketonaciduria
C0804151|T201|MTH_LN|21357-9|LNC2HPO|Ketonaciduria|Ketonaciduria
C0804151|T201|DN|21357-9|LNC2HPO|Ketonaciduria|Ketonaciduria
C0804151|T201|OSN|21357-9|LNC2HPO|Ketonaciduria|Ketonaciduria
C0804151|T201|LC|21357-9|LNC2HPO|Ketonaciduria|Ketonaciduria
C0880212|T201|LN|22702-5|LNC2HPO|Ketonuria|Ketonuria
C0880212|T201|DN|22702-5|LNC2HPO|Ketonuria|Ketonuria
C0880212|T201|MTH_LN|22702-5|LNC2HPO|Ketonuria|Ketonuria
C0880212|T201|OSN|22702-5|LNC2HPO|Ketonuria|Ketonuria
C0880212|T201|LC|22702-5|LNC2HPO|Ketonuria|Ketonuria
C0880212|T201|LN|22702-5|LNC2HPO|Acetonuria|Acetonuria
C0880212|T201|DN|22702-5|LNC2HPO|Acetonuria|Acetonuria
C0880212|T201|MTH_LN|22702-5|LNC2HPO|Acetonuria|Acetonuria
C0880212|T201|OSN|22702-5|LNC2HPO|Acetonuria|Acetonuria
C0880212|T201|LC|22702-5|LNC2HPO|Acetonuria|Acetonuria
C0880212|T201|LN|22702-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C0880212|T201|DN|22702-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C0880212|T201|MTH_LN|22702-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C0880212|T201|OSN|22702-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C0880212|T201|LC|22702-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C0880212|T201|LN|22702-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C0880212|T201|DN|22702-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C0880212|T201|MTH_LN|22702-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C0880212|T201|OSN|22702-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C0880212|T201|LC|22702-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C0364654|T201|LN|2513-0|LNC2HPO|Ketonemia|Ketonemia
C0364654|T201|MTH_LN|2513-0|LNC2HPO|Ketonemia|Ketonemia
C0364654|T201|DN|2513-0|LNC2HPO|Ketonemia|Ketonemia
C0364654|T201|OSN|2513-0|LNC2HPO|Ketonemia|Ketonemia
C0364654|T201|LC|2513-0|LNC2HPO|Ketonemia|Ketonemia
C0364654|T201|LN|2513-0|LNC2HPO|Hyperketonemia|Hyperketonemia
C0364654|T201|MTH_LN|2513-0|LNC2HPO|Hyperketonemia|Hyperketonemia
C0364654|T201|DN|2513-0|LNC2HPO|Hyperketonemia|Hyperketonemia
C0364654|T201|OSN|2513-0|LNC2HPO|Hyperketonemia|Hyperketonemia
C0364654|T201|LC|2513-0|LNC2HPO|Hyperketonemia|Hyperketonemia
C0941792|T201|LN|25705-5|LNC2HPO|Ketonuria|Ketonuria
C0941792|T201|MTH_LN|25705-5|LNC2HPO|Ketonuria|Ketonuria
C0941792|T201|DN|25705-5|LNC2HPO|Ketonuria|Ketonuria
C0941792|T201|OSN|25705-5|LNC2HPO|Ketonuria|Ketonuria
C0941792|T201|LC|25705-5|LNC2HPO|Ketonuria|Ketonuria
C0941792|T201|LN|25705-5|LNC2HPO|Acetonuria|Acetonuria
C0941792|T201|MTH_LN|25705-5|LNC2HPO|Acetonuria|Acetonuria
C0941792|T201|DN|25705-5|LNC2HPO|Acetonuria|Acetonuria
C0941792|T201|OSN|25705-5|LNC2HPO|Acetonuria|Acetonuria
C0941792|T201|LC|25705-5|LNC2HPO|Acetonuria|Acetonuria
C0941792|T201|LN|25705-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C0941792|T201|MTH_LN|25705-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C0941792|T201|DN|25705-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C0941792|T201|OSN|25705-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C0941792|T201|LC|25705-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C0941792|T201|LN|25705-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C0941792|T201|MTH_LN|25705-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C0941792|T201|DN|25705-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C0941792|T201|OSN|25705-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C0941792|T201|LC|25705-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C0941793|T201|LN|25706-3|LNC2HPO|Ketonuria|Ketonuria
C0941793|T201|DN|25706-3|LNC2HPO|Ketonuria|Ketonuria
C0941793|T201|MTH_LN|25706-3|LNC2HPO|Ketonuria|Ketonuria
C0941793|T201|OSN|25706-3|LNC2HPO|Ketonuria|Ketonuria
C0941793|T201|LC|25706-3|LNC2HPO|Ketonuria|Ketonuria
C0941793|T201|LN|25706-3|LNC2HPO|Acetonuria|Acetonuria
C0941793|T201|DN|25706-3|LNC2HPO|Acetonuria|Acetonuria
C0941793|T201|MTH_LN|25706-3|LNC2HPO|Acetonuria|Acetonuria
C0941793|T201|OSN|25706-3|LNC2HPO|Acetonuria|Acetonuria
C0941793|T201|LC|25706-3|LNC2HPO|Acetonuria|Acetonuria
C0941793|T201|LN|25706-3|LNC2HPO|Ketoaciduria|Ketoaciduria
C0941793|T201|DN|25706-3|LNC2HPO|Ketoaciduria|Ketoaciduria
C0941793|T201|MTH_LN|25706-3|LNC2HPO|Ketoaciduria|Ketoaciduria
C0941793|T201|OSN|25706-3|LNC2HPO|Ketoaciduria|Ketoaciduria
C0941793|T201|LC|25706-3|LNC2HPO|Ketoaciduria|Ketoaciduria
C0941793|T201|LN|25706-3|LNC2HPO|Ketonaciduria|Ketonaciduria
C0941793|T201|DN|25706-3|LNC2HPO|Ketonaciduria|Ketonaciduria
C0941793|T201|MTH_LN|25706-3|LNC2HPO|Ketonaciduria|Ketonaciduria
C0941793|T201|OSN|25706-3|LNC2HPO|Ketonaciduria|Ketonaciduria
C0941793|T201|LC|25706-3|LNC2HPO|Ketonaciduria|Ketonaciduria
C0941794|T201|LN|25707-1|LNC2HPO|Ketonuria|Ketonuria
C0941794|T201|DN|25707-1|LNC2HPO|Ketonuria|Ketonuria
C0941794|T201|MTH_LN|25707-1|LNC2HPO|Ketonuria|Ketonuria
C0941794|T201|OSN|25707-1|LNC2HPO|Ketonuria|Ketonuria
C0941794|T201|LC|25707-1|LNC2HPO|Ketonuria|Ketonuria
C0941794|T201|LN|25707-1|LNC2HPO|Acetonuria|Acetonuria
C0941794|T201|DN|25707-1|LNC2HPO|Acetonuria|Acetonuria
C0941794|T201|MTH_LN|25707-1|LNC2HPO|Acetonuria|Acetonuria
C0941794|T201|OSN|25707-1|LNC2HPO|Acetonuria|Acetonuria
C0941794|T201|LC|25707-1|LNC2HPO|Acetonuria|Acetonuria
C0941794|T201|LN|25707-1|LNC2HPO|Ketoaciduria|Ketoaciduria
C0941794|T201|DN|25707-1|LNC2HPO|Ketoaciduria|Ketoaciduria
C0941794|T201|MTH_LN|25707-1|LNC2HPO|Ketoaciduria|Ketoaciduria
C0941794|T201|OSN|25707-1|LNC2HPO|Ketoaciduria|Ketoaciduria
C0941794|T201|LC|25707-1|LNC2HPO|Ketoaciduria|Ketoaciduria
C0941794|T201|LN|25707-1|LNC2HPO|Ketonaciduria|Ketonaciduria
C0941794|T201|DN|25707-1|LNC2HPO|Ketonaciduria|Ketonaciduria
C0941794|T201|MTH_LN|25707-1|LNC2HPO|Ketonaciduria|Ketonaciduria
C0941794|T201|OSN|25707-1|LNC2HPO|Ketonaciduria|Ketonaciduria
C0941794|T201|LC|25707-1|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942779|T201|LN|26884-7|LNC2HPO|Ketonuria|Ketonuria
C0942779|T201|MTH_LN|26884-7|LNC2HPO|Ketonuria|Ketonuria
C0942779|T201|DN|26884-7|LNC2HPO|Ketonuria|Ketonuria
C0942779|T201|OSN|26884-7|LNC2HPO|Ketonuria|Ketonuria
C0942779|T201|LC|26884-7|LNC2HPO|Ketonuria|Ketonuria
C0942779|T201|LN|26884-7|LNC2HPO|Acetonuria|Acetonuria
C0942779|T201|MTH_LN|26884-7|LNC2HPO|Acetonuria|Acetonuria
C0942779|T201|DN|26884-7|LNC2HPO|Acetonuria|Acetonuria
C0942779|T201|OSN|26884-7|LNC2HPO|Acetonuria|Acetonuria
C0942779|T201|LC|26884-7|LNC2HPO|Acetonuria|Acetonuria
C0942779|T201|LN|26884-7|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942779|T201|MTH_LN|26884-7|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942779|T201|DN|26884-7|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942779|T201|OSN|26884-7|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942779|T201|LC|26884-7|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942779|T201|LN|26884-7|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942779|T201|MTH_LN|26884-7|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942779|T201|DN|26884-7|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942779|T201|OSN|26884-7|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942779|T201|LC|26884-7|LNC2HPO|Ketonaciduria|Ketonaciduria
C0945443|T201|LN|27028-0|LNC2HPO|Ketonuria|Ketonuria
C0945443|T201|MTH_LN|27028-0|LNC2HPO|Ketonuria|Ketonuria
C0945443|T201|DN|27028-0|LNC2HPO|Ketonuria|Ketonuria
C0945443|T201|OSN|27028-0|LNC2HPO|Ketonuria|Ketonuria
C0945443|T201|LC|27028-0|LNC2HPO|Ketonuria|Ketonuria
C0945443|T201|LN|27028-0|LNC2HPO|Acetonuria|Acetonuria
C0945443|T201|MTH_LN|27028-0|LNC2HPO|Acetonuria|Acetonuria
C0945443|T201|DN|27028-0|LNC2HPO|Acetonuria|Acetonuria
C0945443|T201|OSN|27028-0|LNC2HPO|Acetonuria|Acetonuria
C0945443|T201|LC|27028-0|LNC2HPO|Acetonuria|Acetonuria
C0945443|T201|LN|27028-0|LNC2HPO|Ketoaciduria|Ketoaciduria
C0945443|T201|MTH_LN|27028-0|LNC2HPO|Ketoaciduria|Ketoaciduria
C0945443|T201|DN|27028-0|LNC2HPO|Ketoaciduria|Ketoaciduria
C0945443|T201|OSN|27028-0|LNC2HPO|Ketoaciduria|Ketoaciduria
C0945443|T201|LC|27028-0|LNC2HPO|Ketoaciduria|Ketoaciduria
C0945443|T201|LN|27028-0|LNC2HPO|Ketonaciduria|Ketonaciduria
C0945443|T201|MTH_LN|27028-0|LNC2HPO|Ketonaciduria|Ketonaciduria
C0945443|T201|DN|27028-0|LNC2HPO|Ketonaciduria|Ketonaciduria
C0945443|T201|OSN|27028-0|LNC2HPO|Ketonaciduria|Ketonaciduria
C0945443|T201|LC|27028-0|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942905|T201|LN|27040-5|LNC2HPO|Ketonuria|Ketonuria
C0942905|T201|MTH_LN|27040-5|LNC2HPO|Ketonuria|Ketonuria
C0942905|T201|DN|27040-5|LNC2HPO|Ketonuria|Ketonuria
C0942905|T201|OSN|27040-5|LNC2HPO|Ketonuria|Ketonuria
C0942905|T201|LC|27040-5|LNC2HPO|Ketonuria|Ketonuria
C0942905|T201|LN|27040-5|LNC2HPO|Acetonuria|Acetonuria
C0942905|T201|MTH_LN|27040-5|LNC2HPO|Acetonuria|Acetonuria
C0942905|T201|DN|27040-5|LNC2HPO|Acetonuria|Acetonuria
C0942905|T201|OSN|27040-5|LNC2HPO|Acetonuria|Acetonuria
C0942905|T201|LC|27040-5|LNC2HPO|Acetonuria|Acetonuria
C0942905|T201|LN|27040-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942905|T201|MTH_LN|27040-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942905|T201|DN|27040-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942905|T201|OSN|27040-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942905|T201|LC|27040-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942905|T201|LN|27040-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942905|T201|MTH_LN|27040-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942905|T201|DN|27040-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942905|T201|OSN|27040-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942905|T201|LC|27040-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942922|T201|LN|27062-9|LNC2HPO|Ketonuria|Ketonuria
C0942922|T201|MTH_LN|27062-9|LNC2HPO|Ketonuria|Ketonuria
C0942922|T201|DN|27062-9|LNC2HPO|Ketonuria|Ketonuria
C0942922|T201|OSN|27062-9|LNC2HPO|Ketonuria|Ketonuria
C0942922|T201|LC|27062-9|LNC2HPO|Ketonuria|Ketonuria
C0942922|T201|LN|27062-9|LNC2HPO|Acetonuria|Acetonuria
C0942922|T201|MTH_LN|27062-9|LNC2HPO|Acetonuria|Acetonuria
C0942922|T201|DN|27062-9|LNC2HPO|Acetonuria|Acetonuria
C0942922|T201|OSN|27062-9|LNC2HPO|Acetonuria|Acetonuria
C0942922|T201|LC|27062-9|LNC2HPO|Acetonuria|Acetonuria
C0942922|T201|LN|27062-9|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942922|T201|MTH_LN|27062-9|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942922|T201|DN|27062-9|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942922|T201|OSN|27062-9|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942922|T201|LC|27062-9|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942922|T201|LN|27062-9|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942922|T201|MTH_LN|27062-9|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942922|T201|DN|27062-9|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942922|T201|OSN|27062-9|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942922|T201|LC|27062-9|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942925|T201|LN|27065-2|LNC2HPO|Ketonuria|Ketonuria
C0942925|T201|MTH_LN|27065-2|LNC2HPO|Ketonuria|Ketonuria
C0942925|T201|DN|27065-2|LNC2HPO|Ketonuria|Ketonuria
C0942925|T201|OSN|27065-2|LNC2HPO|Ketonuria|Ketonuria
C0942925|T201|LC|27065-2|LNC2HPO|Ketonuria|Ketonuria
C0942925|T201|LN|27065-2|LNC2HPO|Acetonuria|Acetonuria
C0942925|T201|MTH_LN|27065-2|LNC2HPO|Acetonuria|Acetonuria
C0942925|T201|DN|27065-2|LNC2HPO|Acetonuria|Acetonuria
C0942925|T201|OSN|27065-2|LNC2HPO|Acetonuria|Acetonuria
C0942925|T201|LC|27065-2|LNC2HPO|Acetonuria|Acetonuria
C0942925|T201|LN|27065-2|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942925|T201|MTH_LN|27065-2|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942925|T201|DN|27065-2|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942925|T201|OSN|27065-2|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942925|T201|LC|27065-2|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942925|T201|LN|27065-2|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942925|T201|MTH_LN|27065-2|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942925|T201|DN|27065-2|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942925|T201|OSN|27065-2|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942925|T201|LC|27065-2|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942926|T201|LN|27066-0|LNC2HPO|Ketonuria|Ketonuria
C0942926|T201|MTH_LN|27066-0|LNC2HPO|Ketonuria|Ketonuria
C0942926|T201|DN|27066-0|LNC2HPO|Ketonuria|Ketonuria
C0942926|T201|OSN|27066-0|LNC2HPO|Ketonuria|Ketonuria
C0942926|T201|LC|27066-0|LNC2HPO|Ketonuria|Ketonuria
C0942926|T201|LN|27066-0|LNC2HPO|Acetonuria|Acetonuria
C0942926|T201|MTH_LN|27066-0|LNC2HPO|Acetonuria|Acetonuria
C0942926|T201|DN|27066-0|LNC2HPO|Acetonuria|Acetonuria
C0942926|T201|OSN|27066-0|LNC2HPO|Acetonuria|Acetonuria
C0942926|T201|LC|27066-0|LNC2HPO|Acetonuria|Acetonuria
C0942926|T201|LN|27066-0|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942926|T201|MTH_LN|27066-0|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942926|T201|DN|27066-0|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942926|T201|OSN|27066-0|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942926|T201|LC|27066-0|LNC2HPO|Ketoaciduria|Ketoaciduria
C0942926|T201|LN|27066-0|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942926|T201|MTH_LN|27066-0|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942926|T201|DN|27066-0|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942926|T201|OSN|27066-0|LNC2HPO|Ketonaciduria|Ketonaciduria
C0942926|T201|LC|27066-0|LNC2HPO|Ketonaciduria|Ketonaciduria
C1148231|T201|LN|32547-2|LNC2HPO|Ketonemia|Ketonemia
C1148231|T201|DN|32547-2|LNC2HPO|Ketonemia|Ketonemia
C1148231|T201|MTH_LN|32547-2|LNC2HPO|Ketonemia|Ketonemia
C1148231|T201|OSN|32547-2|LNC2HPO|Ketonemia|Ketonemia
C1148231|T201|LC|32547-2|LNC2HPO|Ketonemia|Ketonemia
C1148231|T201|LN|32547-2|LNC2HPO|Hyperketonemia|Hyperketonemia
C1148231|T201|DN|32547-2|LNC2HPO|Hyperketonemia|Hyperketonemia
C1148231|T201|MTH_LN|32547-2|LNC2HPO|Hyperketonemia|Hyperketonemia
C1148231|T201|OSN|32547-2|LNC2HPO|Hyperketonemia|Hyperketonemia
C1148231|T201|LC|32547-2|LNC2HPO|Hyperketonemia|Hyperketonemia
C1315514|T201|LN|33043-1|LNC2HPO|Ketonuria|Ketonuria
C1315514|T201|MTH_LN|33043-1|LNC2HPO|Ketonuria|Ketonuria
C1315514|T201|DN|33043-1|LNC2HPO|Ketonuria|Ketonuria
C1315514|T201|OSN|33043-1|LNC2HPO|Ketonuria|Ketonuria
C1315514|T201|LC|33043-1|LNC2HPO|Ketonuria|Ketonuria
C1315514|T201|LN|33043-1|LNC2HPO|Acetonuria|Acetonuria
C1315514|T201|MTH_LN|33043-1|LNC2HPO|Acetonuria|Acetonuria
C1315514|T201|DN|33043-1|LNC2HPO|Acetonuria|Acetonuria
C1315514|T201|OSN|33043-1|LNC2HPO|Acetonuria|Acetonuria
C1315514|T201|LC|33043-1|LNC2HPO|Acetonuria|Acetonuria
C1315514|T201|LN|33043-1|LNC2HPO|Ketoaciduria|Ketoaciduria
C1315514|T201|MTH_LN|33043-1|LNC2HPO|Ketoaciduria|Ketoaciduria
C1315514|T201|DN|33043-1|LNC2HPO|Ketoaciduria|Ketoaciduria
C1315514|T201|OSN|33043-1|LNC2HPO|Ketoaciduria|Ketoaciduria
C1315514|T201|LC|33043-1|LNC2HPO|Ketoaciduria|Ketoaciduria
C1315514|T201|LN|33043-1|LNC2HPO|Ketonaciduria|Ketonaciduria
C1315514|T201|MTH_LN|33043-1|LNC2HPO|Ketonaciduria|Ketonaciduria
C1315514|T201|DN|33043-1|LNC2HPO|Ketonaciduria|Ketonaciduria
C1315514|T201|OSN|33043-1|LNC2HPO|Ketonaciduria|Ketonaciduria
C1315514|T201|LC|33043-1|LNC2HPO|Ketonaciduria|Ketonaciduria
C1315529|T201|LN|33058-9|LNC2HPO|Ketonemia|Ketonemia
C1315529|T201|DN|33058-9|LNC2HPO|Ketonemia|Ketonemia
C1315529|T201|MTH_LN|33058-9|LNC2HPO|Ketonemia|Ketonemia
C1315529|T201|OSN|33058-9|LNC2HPO|Ketonemia|Ketonemia
C1315529|T201|LC|33058-9|LNC2HPO|Ketonemia|Ketonemia
C1315529|T201|LN|33058-9|LNC2HPO|Hyperketonemia|Hyperketonemia
C1315529|T201|DN|33058-9|LNC2HPO|Hyperketonemia|Hyperketonemia
C1315529|T201|MTH_LN|33058-9|LNC2HPO|Hyperketonemia|Hyperketonemia
C1315529|T201|OSN|33058-9|LNC2HPO|Hyperketonemia|Hyperketonemia
C1315529|T201|LC|33058-9|LNC2HPO|Hyperketonemia|Hyperketonemia
C1316366|T201|LN|33903-6|LNC2HPO|Ketonuria|Ketonuria
C1316366|T201|MTH_LN|33903-6|LNC2HPO|Ketonuria|Ketonuria
C1316366|T201|DN|33903-6|LNC2HPO|Ketonuria|Ketonuria
C1316366|T201|OSN|33903-6|LNC2HPO|Ketonuria|Ketonuria
C1316366|T201|LC|33903-6|LNC2HPO|Ketonuria|Ketonuria
C1316366|T201|LN|33903-6|LNC2HPO|Acetonuria|Acetonuria
C1316366|T201|MTH_LN|33903-6|LNC2HPO|Acetonuria|Acetonuria
C1316366|T201|DN|33903-6|LNC2HPO|Acetonuria|Acetonuria
C1316366|T201|OSN|33903-6|LNC2HPO|Acetonuria|Acetonuria
C1316366|T201|LC|33903-6|LNC2HPO|Acetonuria|Acetonuria
C1316366|T201|LN|33903-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C1316366|T201|MTH_LN|33903-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C1316366|T201|DN|33903-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C1316366|T201|OSN|33903-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C1316366|T201|LC|33903-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C1316366|T201|LN|33903-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C1316366|T201|MTH_LN|33903-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C1316366|T201|DN|33903-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C1316366|T201|OSN|33903-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C1316366|T201|LC|33903-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C1526494|T201|LN|38493-3|LNC2HPO|Ketonemia|Ketonemia
C1526494|T201|DN|38493-3|LNC2HPO|Ketonemia|Ketonemia
C1526494|T201|MTH_LN|38493-3|LNC2HPO|Ketonemia|Ketonemia
C1526494|T201|OSN|38493-3|LNC2HPO|Ketonemia|Ketonemia
C1526494|T201|LC|38493-3|LNC2HPO|Ketonemia|Ketonemia
C1526494|T201|LN|38493-3|LNC2HPO|Hyperketonemia|Hyperketonemia
C1526494|T201|DN|38493-3|LNC2HPO|Hyperketonemia|Hyperketonemia
C1526494|T201|MTH_LN|38493-3|LNC2HPO|Hyperketonemia|Hyperketonemia
C1526494|T201|OSN|38493-3|LNC2HPO|Hyperketonemia|Hyperketonemia
C1526494|T201|LC|38493-3|LNC2HPO|Hyperketonemia|Hyperketonemia
C1977522|T201|LN|49779-2|LNC2HPO|Ketonuria|Ketonuria
C1977522|T201|DN|49779-2|LNC2HPO|Ketonuria|Ketonuria
C1977522|T201|MTH_LN|49779-2|LNC2HPO|Ketonuria|Ketonuria
C1977522|T201|OSN|49779-2|LNC2HPO|Ketonuria|Ketonuria
C1977522|T201|LC|49779-2|LNC2HPO|Ketonuria|Ketonuria
C1977522|T201|LN|49779-2|LNC2HPO|Acetonuria|Acetonuria
C1977522|T201|DN|49779-2|LNC2HPO|Acetonuria|Acetonuria
C1977522|T201|MTH_LN|49779-2|LNC2HPO|Acetonuria|Acetonuria
C1977522|T201|OSN|49779-2|LNC2HPO|Acetonuria|Acetonuria
C1977522|T201|LC|49779-2|LNC2HPO|Acetonuria|Acetonuria
C1977522|T201|LN|49779-2|LNC2HPO|Ketoaciduria|Ketoaciduria
C1977522|T201|DN|49779-2|LNC2HPO|Ketoaciduria|Ketoaciduria
C1977522|T201|MTH_LN|49779-2|LNC2HPO|Ketoaciduria|Ketoaciduria
C1977522|T201|OSN|49779-2|LNC2HPO|Ketoaciduria|Ketoaciduria
C1977522|T201|LC|49779-2|LNC2HPO|Ketoaciduria|Ketoaciduria
C1977522|T201|LN|49779-2|LNC2HPO|Ketonaciduria|Ketonaciduria
C1977522|T201|DN|49779-2|LNC2HPO|Ketonaciduria|Ketonaciduria
C1977522|T201|MTH_LN|49779-2|LNC2HPO|Ketonaciduria|Ketonaciduria
C1977522|T201|OSN|49779-2|LNC2HPO|Ketonaciduria|Ketonaciduria
C1977522|T201|LC|49779-2|LNC2HPO|Ketonaciduria|Ketonaciduria
C1978484|T201|LN|50557-8|LNC2HPO|Ketonuria|Ketonuria
C1978484|T201|DN|50557-8|LNC2HPO|Ketonuria|Ketonuria
C1978484|T201|OSN|50557-8|LNC2HPO|Ketonuria|Ketonuria
C1978484|T201|MTH_LN|50557-8|LNC2HPO|Ketonuria|Ketonuria
C1978484|T201|LC|50557-8|LNC2HPO|Ketonuria|Ketonuria
C1978484|T201|LN|50557-8|LNC2HPO|Acetonuria|Acetonuria
C1978484|T201|DN|50557-8|LNC2HPO|Acetonuria|Acetonuria
C1978484|T201|OSN|50557-8|LNC2HPO|Acetonuria|Acetonuria
C1978484|T201|MTH_LN|50557-8|LNC2HPO|Acetonuria|Acetonuria
C1978484|T201|LC|50557-8|LNC2HPO|Acetonuria|Acetonuria
C1978484|T201|LN|50557-8|LNC2HPO|Ketoaciduria|Ketoaciduria
C1978484|T201|DN|50557-8|LNC2HPO|Ketoaciduria|Ketoaciduria
C1978484|T201|OSN|50557-8|LNC2HPO|Ketoaciduria|Ketoaciduria
C1978484|T201|MTH_LN|50557-8|LNC2HPO|Ketoaciduria|Ketoaciduria
C1978484|T201|LC|50557-8|LNC2HPO|Ketoaciduria|Ketoaciduria
C1978484|T201|LN|50557-8|LNC2HPO|Ketonaciduria|Ketonaciduria
C1978484|T201|DN|50557-8|LNC2HPO|Ketonaciduria|Ketonaciduria
C1978484|T201|OSN|50557-8|LNC2HPO|Ketonaciduria|Ketonaciduria
C1978484|T201|MTH_LN|50557-8|LNC2HPO|Ketonaciduria|Ketonaciduria
C1978484|T201|LC|50557-8|LNC2HPO|Ketonaciduria|Ketonaciduria
C2361549|T201|LN|53061-8|LNC2HPO|Ketonemia|Ketonemia
C2361549|T201|DN|53061-8|LNC2HPO|Ketonemia|Ketonemia
C2361549|T201|OSN|53061-8|LNC2HPO|Ketonemia|Ketonemia
C2361549|T201|MTH_LN|53061-8|LNC2HPO|Ketonemia|Ketonemia
C2361549|T201|LC|53061-8|LNC2HPO|Ketonemia|Ketonemia
C2361549|T201|LN|53061-8|LNC2HPO|Hyperketonemia|Hyperketonemia
C2361549|T201|DN|53061-8|LNC2HPO|Hyperketonemia|Hyperketonemia
C2361549|T201|OSN|53061-8|LNC2HPO|Hyperketonemia|Hyperketonemia
C2361549|T201|MTH_LN|53061-8|LNC2HPO|Hyperketonemia|Hyperketonemia
C2361549|T201|LC|53061-8|LNC2HPO|Hyperketonemia|Hyperketonemia
C0368032|T201|LN|5797-6|LNC2HPO|Ketonuria|Ketonuria
C0368032|T201|MTH_LN|5797-6|LNC2HPO|Ketonuria|Ketonuria
C0368032|T201|DN|5797-6|LNC2HPO|Ketonuria|Ketonuria
C0368032|T201|OSN|5797-6|LNC2HPO|Ketonuria|Ketonuria
C0368032|T201|LC|5797-6|LNC2HPO|Ketonuria|Ketonuria
C0368032|T201|LN|5797-6|LNC2HPO|Acetonuria|Acetonuria
C0368032|T201|MTH_LN|5797-6|LNC2HPO|Acetonuria|Acetonuria
C0368032|T201|DN|5797-6|LNC2HPO|Acetonuria|Acetonuria
C0368032|T201|OSN|5797-6|LNC2HPO|Acetonuria|Acetonuria
C0368032|T201|LC|5797-6|LNC2HPO|Acetonuria|Acetonuria
C0368032|T201|LN|5797-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C0368032|T201|MTH_LN|5797-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C0368032|T201|DN|5797-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C0368032|T201|OSN|5797-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C0368032|T201|LC|5797-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C0368032|T201|LN|5797-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C0368032|T201|MTH_LN|5797-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C0368032|T201|DN|5797-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C0368032|T201|OSN|5797-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C0368032|T201|LC|5797-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C2925731|T201|LN|59158-6|LNC2HPO|Ketonuria|Ketonuria
C2925731|T201|DN|59158-6|LNC2HPO|Ketonuria|Ketonuria
C2925731|T201|OSN|59158-6|LNC2HPO|Ketonuria|Ketonuria
C2925731|T201|LC|59158-6|LNC2HPO|Ketonuria|Ketonuria
C2925731|T201|MTH_LN|59158-6|LNC2HPO|Ketonuria|Ketonuria
C2925731|T201|LN|59158-6|LNC2HPO|Acetonuria|Acetonuria
C2925731|T201|DN|59158-6|LNC2HPO|Acetonuria|Acetonuria
C2925731|T201|OSN|59158-6|LNC2HPO|Acetonuria|Acetonuria
C2925731|T201|LC|59158-6|LNC2HPO|Acetonuria|Acetonuria
C2925731|T201|MTH_LN|59158-6|LNC2HPO|Acetonuria|Acetonuria
C2925731|T201|LN|59158-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C2925731|T201|DN|59158-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C2925731|T201|OSN|59158-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C2925731|T201|LC|59158-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C2925731|T201|MTH_LN|59158-6|LNC2HPO|Ketoaciduria|Ketoaciduria
C2925731|T201|LN|59158-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C2925731|T201|DN|59158-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C2925731|T201|OSN|59158-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C2925731|T201|LC|59158-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C2925731|T201|MTH_LN|59158-6|LNC2HPO|Ketonaciduria|Ketonaciduria
C3172442|T201|LN|63371-9|LNC2HPO|Ketonuria|Ketonuria
C3172442|T201|OSN|63371-9|LNC2HPO|Ketonuria|Ketonuria
C3172442|T201|LC|63371-9|LNC2HPO|Ketonuria|Ketonuria
C3172442|T201|MTH_LN|63371-9|LNC2HPO|Ketonuria|Ketonuria
C3172442|T201|DN|63371-9|LNC2HPO|Ketonuria|Ketonuria
C3172442|T201|LN|63371-9|LNC2HPO|Acetonuria|Acetonuria
C3172442|T201|OSN|63371-9|LNC2HPO|Acetonuria|Acetonuria
C3172442|T201|LC|63371-9|LNC2HPO|Acetonuria|Acetonuria
C3172442|T201|MTH_LN|63371-9|LNC2HPO|Acetonuria|Acetonuria
C3172442|T201|DN|63371-9|LNC2HPO|Acetonuria|Acetonuria
C3172442|T201|LN|63371-9|LNC2HPO|Ketoaciduria|Ketoaciduria
C3172442|T201|OSN|63371-9|LNC2HPO|Ketoaciduria|Ketoaciduria
C3172442|T201|LC|63371-9|LNC2HPO|Ketoaciduria|Ketoaciduria
C3172442|T201|MTH_LN|63371-9|LNC2HPO|Ketoaciduria|Ketoaciduria
C3172442|T201|DN|63371-9|LNC2HPO|Ketoaciduria|Ketoaciduria
C3172442|T201|LN|63371-9|LNC2HPO|Ketonaciduria|Ketonaciduria
C3172442|T201|OSN|63371-9|LNC2HPO|Ketonaciduria|Ketonaciduria
C3172442|T201|LC|63371-9|LNC2HPO|Ketonaciduria|Ketonaciduria
C3172442|T201|MTH_LN|63371-9|LNC2HPO|Ketonaciduria|Ketonaciduria
C3172442|T201|DN|63371-9|LNC2HPO|Ketonaciduria|Ketonaciduria
C3172443|T201|LN|63372-7|LNC2HPO|Ketonuria|Ketonuria
C3172443|T201|OSN|63372-7|LNC2HPO|Ketonuria|Ketonuria
C3172443|T201|LC|63372-7|LNC2HPO|Ketonuria|Ketonuria
C3172443|T201|MTH_LN|63372-7|LNC2HPO|Ketonuria|Ketonuria
C3172443|T201|DN|63372-7|LNC2HPO|Ketonuria|Ketonuria
C3172443|T201|LN|63372-7|LNC2HPO|Acetonuria|Acetonuria
C3172443|T201|OSN|63372-7|LNC2HPO|Acetonuria|Acetonuria
C3172443|T201|LC|63372-7|LNC2HPO|Acetonuria|Acetonuria
C3172443|T201|MTH_LN|63372-7|LNC2HPO|Acetonuria|Acetonuria
C3172443|T201|DN|63372-7|LNC2HPO|Acetonuria|Acetonuria
C3172443|T201|LN|63372-7|LNC2HPO|Ketoaciduria|Ketoaciduria
C3172443|T201|OSN|63372-7|LNC2HPO|Ketoaciduria|Ketoaciduria
C3172443|T201|LC|63372-7|LNC2HPO|Ketoaciduria|Ketoaciduria
C3172443|T201|MTH_LN|63372-7|LNC2HPO|Ketoaciduria|Ketoaciduria
C3172443|T201|DN|63372-7|LNC2HPO|Ketoaciduria|Ketoaciduria
C3172443|T201|LN|63372-7|LNC2HPO|Ketonaciduria|Ketonaciduria
C3172443|T201|OSN|63372-7|LNC2HPO|Ketonaciduria|Ketonaciduria
C3172443|T201|LC|63372-7|LNC2HPO|Ketonaciduria|Ketonaciduria
C3172443|T201|MTH_LN|63372-7|LNC2HPO|Ketonaciduria|Ketonaciduria
C3172443|T201|DN|63372-7|LNC2HPO|Ketonaciduria|Ketonaciduria
C3172444|T201|LN|63373-5|LNC2HPO|Ketonuria|Ketonuria
C3172444|T201|OSN|63373-5|LNC2HPO|Ketonuria|Ketonuria
C3172444|T201|LC|63373-5|LNC2HPO|Ketonuria|Ketonuria
C3172444|T201|MTH_LN|63373-5|LNC2HPO|Ketonuria|Ketonuria
C3172444|T201|DN|63373-5|LNC2HPO|Ketonuria|Ketonuria
C3172444|T201|LN|63373-5|LNC2HPO|Acetonuria|Acetonuria
C3172444|T201|OSN|63373-5|LNC2HPO|Acetonuria|Acetonuria
C3172444|T201|LC|63373-5|LNC2HPO|Acetonuria|Acetonuria
C3172444|T201|MTH_LN|63373-5|LNC2HPO|Acetonuria|Acetonuria
C3172444|T201|DN|63373-5|LNC2HPO|Acetonuria|Acetonuria
C3172444|T201|LN|63373-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C3172444|T201|OSN|63373-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C3172444|T201|LC|63373-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C3172444|T201|MTH_LN|63373-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C3172444|T201|DN|63373-5|LNC2HPO|Ketoaciduria|Ketoaciduria
C3172444|T201|LN|63373-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C3172444|T201|OSN|63373-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C3172444|T201|LC|63373-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C3172444|T201|MTH_LN|63373-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C3172444|T201|DN|63373-5|LNC2HPO|Ketonaciduria|Ketonaciduria
C3262796|T201|LN|68955-4|LNC2HPO|Ketonemia|Ketonemia
C3262796|T201|OSN|68955-4|LNC2HPO|Ketonemia|Ketonemia
C3262796|T201|DN|68955-4|LNC2HPO|Ketonemia|Ketonemia
C3262796|T201|LC|68955-4|LNC2HPO|Ketonemia|Ketonemia
C3262796|T201|MTH_LN|68955-4|LNC2HPO|Ketonemia|Ketonemia
C3262796|T201|LN|68955-4|LNC2HPO|Hyperketonemia|Hyperketonemia
C3262796|T201|OSN|68955-4|LNC2HPO|Hyperketonemia|Hyperketonemia
C3262796|T201|DN|68955-4|LNC2HPO|Hyperketonemia|Hyperketonemia
C3262796|T201|LC|68955-4|LNC2HPO|Hyperketonemia|Hyperketonemia
C3262796|T201|MTH_LN|68955-4|LNC2HPO|Hyperketonemia|Hyperketonemia
C0364210|T201|LN|2078-4|LNC2HPO|Hyperchloriduria|Hyperchloriduria
C0364210|T201|MTH_LN|2078-4|LNC2HPO|Hyperchloriduria|Hyperchloriduria
C0364210|T201|DN|2078-4|LNC2HPO|Hyperchloriduria|Hyperchloriduria
C0364210|T201|OSN|2078-4|LNC2HPO|Hyperchloriduria|Hyperchloriduria
C0364210|T201|LC|2078-4|LNC2HPO|Hyperchloriduria|Hyperchloriduria
C0364210|T201|LN|2078-4|LNC2HPO|Hypochloriduria|Hypochloriduria
C0364210|T201|MTH_LN|2078-4|LNC2HPO|Hypochloriduria|Hypochloriduria
C0364210|T201|DN|2078-4|LNC2HPO|Hypochloriduria|Hypochloriduria
C0364210|T201|OSN|2078-4|LNC2HPO|Hypochloriduria|Hypochloriduria
C0364210|T201|LC|2078-4|LNC2HPO|Hypochloriduria|Hypochloriduria
C0367401|T201|LN|5117-7|LNC2HPO|Cryoglobulinemia|Cryoglobulinemia
C0367401|T201|MTH_LN|5117-7|LNC2HPO|Cryoglobulinemia|Cryoglobulinemia
C0367401|T201|DN|5117-7|LNC2HPO|Cryoglobulinemia|Cryoglobulinemia
C0367401|T201|OSN|5117-7|LNC2HPO|Cryoglobulinemia|Cryoglobulinemia
C0367401|T201|LC|5117-7|LNC2HPO|Cryoglobulinemia|Cryoglobulinemia
C0367401|T201|LN|5117-7|LNC2HPO|Cryoprecipitable immune complexes|Cryoprecipitable immune complexes
C0367401|T201|MTH_LN|5117-7|LNC2HPO|Cryoprecipitable immune complexes|Cryoprecipitable immune complexes
C0367401|T201|DN|5117-7|LNC2HPO|Cryoprecipitable immune complexes|Cryoprecipitable immune complexes
C0367401|T201|OSN|5117-7|LNC2HPO|Cryoprecipitable immune complexes|Cryoprecipitable immune complexes
C0367401|T201|LC|5117-7|LNC2HPO|Cryoprecipitable immune complexes|Cryoprecipitable immune complexes
C0484575|T201|LN|10332-5|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484575|T201|DN|10332-5|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484575|T201|MTH_LN|10332-5|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484575|T201|OSN|10332-5|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484575|T201|LC|10332-5|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484575|T201|LN|10332-5|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484575|T201|DN|10332-5|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484575|T201|MTH_LN|10332-5|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484575|T201|OSN|10332-5|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484575|T201|LC|10332-5|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484575|T201|LN|10332-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484575|T201|DN|10332-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484575|T201|MTH_LN|10332-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484575|T201|OSN|10332-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484575|T201|LC|10332-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484575|T201|LN|10332-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484575|T201|DN|10332-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484575|T201|MTH_LN|10332-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484575|T201|OSN|10332-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484575|T201|LC|10332-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484575|T201|LN|10332-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484575|T201|DN|10332-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484575|T201|MTH_LN|10332-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484575|T201|OSN|10332-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484575|T201|LC|10332-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0797041|T201|LN|13852-9|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C0797041|T201|DN|13852-9|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C0797041|T201|MTH_LN|13852-9|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C0797041|T201|OSN|13852-9|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C0797041|T201|LC|13852-9|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C0797041|T201|LN|13852-9|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C0797041|T201|DN|13852-9|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C0797041|T201|MTH_LN|13852-9|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C0797041|T201|OSN|13852-9|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C0797041|T201|LC|13852-9|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C0797044|T201|LN|13855-2|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C0797044|T201|DN|13855-2|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C0797044|T201|MTH_LN|13855-2|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C0797044|T201|OSN|13855-2|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C0797044|T201|LC|13855-2|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C0797044|T201|LN|13855-2|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C0797044|T201|DN|13855-2|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C0797044|T201|MTH_LN|13855-2|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C0797044|T201|OSN|13855-2|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C0797044|T201|LC|13855-2|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C0482485|T201|LN|1401-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482485|T201|DN|1401-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482485|T201|MTH_LN|1401-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482485|T201|OSN|1401-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482485|T201|LC|1401-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482485|T201|LN|1401-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482485|T201|DN|1401-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482485|T201|MTH_LN|1401-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482485|T201|OSN|1401-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482485|T201|LC|1401-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482485|T201|LN|1401-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482485|T201|DN|1401-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482485|T201|MTH_LN|1401-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482485|T201|OSN|1401-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482485|T201|LC|1401-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482486|T201|LN|1402-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482486|T201|DN|1402-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482486|T201|MTH_LN|1402-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482486|T201|OSN|1402-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482486|T201|LC|1402-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482486|T201|LN|1402-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482486|T201|DN|1402-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482486|T201|MTH_LN|1402-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482486|T201|OSN|1402-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482486|T201|LC|1402-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482486|T201|LN|1402-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482486|T201|DN|1402-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482486|T201|MTH_LN|1402-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482486|T201|OSN|1402-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482486|T201|LC|1402-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482487|T201|LN|1403-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482487|T201|DN|1403-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482487|T201|MTH_LN|1403-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482487|T201|OSN|1403-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482487|T201|LC|1403-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482487|T201|LN|1403-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482487|T201|DN|1403-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482487|T201|MTH_LN|1403-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482487|T201|OSN|1403-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482487|T201|LC|1403-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482487|T201|LN|1403-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482487|T201|DN|1403-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482487|T201|MTH_LN|1403-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482487|T201|OSN|1403-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482487|T201|LC|1403-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482489|T201|LN|1408-4|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482489|T201|DN|1408-4|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482489|T201|MTH_LN|1408-4|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482489|T201|OSN|1408-4|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482489|T201|LC|1408-4|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482489|T201|LN|1408-4|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482489|T201|DN|1408-4|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482489|T201|MTH_LN|1408-4|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482489|T201|OSN|1408-4|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482489|T201|LC|1408-4|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482489|T201|LN|1408-4|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482489|T201|DN|1408-4|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482489|T201|MTH_LN|1408-4|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482489|T201|OSN|1408-4|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482489|T201|LC|1408-4|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482490|T201|LN|1409-2|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482490|T201|DN|1409-2|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482490|T201|MTH_LN|1409-2|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482490|T201|OSN|1409-2|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482490|T201|LC|1409-2|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482490|T201|LN|1409-2|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482490|T201|DN|1409-2|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482490|T201|MTH_LN|1409-2|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482490|T201|OSN|1409-2|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482490|T201|LC|1409-2|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482490|T201|LN|1409-2|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482490|T201|DN|1409-2|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482490|T201|MTH_LN|1409-2|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482490|T201|OSN|1409-2|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482490|T201|LC|1409-2|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482493|T201|LN|1413-4|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482493|T201|DN|1413-4|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482493|T201|MTH_LN|1413-4|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482493|T201|OSN|1413-4|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482493|T201|LC|1413-4|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482493|T201|LN|1413-4|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482493|T201|DN|1413-4|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482493|T201|MTH_LN|1413-4|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482493|T201|OSN|1413-4|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482493|T201|LC|1413-4|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482493|T201|LN|1413-4|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482493|T201|DN|1413-4|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482493|T201|MTH_LN|1413-4|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482493|T201|OSN|1413-4|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482493|T201|LC|1413-4|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482495|T201|LN|1416-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482495|T201|DN|1416-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482495|T201|MTH_LN|1416-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482495|T201|OSN|1416-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482495|T201|LC|1416-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482495|T201|LN|1416-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482495|T201|DN|1416-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482495|T201|MTH_LN|1416-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482495|T201|OSN|1416-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482495|T201|LC|1416-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482495|T201|LN|1416-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482495|T201|DN|1416-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482495|T201|MTH_LN|1416-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482495|T201|OSN|1416-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482495|T201|LC|1416-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482496|T201|LN|1417-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482496|T201|DN|1417-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482496|T201|MTH_LN|1417-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482496|T201|OSN|1417-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482496|T201|LC|1417-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482496|T201|LN|1417-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482496|T201|DN|1417-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482496|T201|MTH_LN|1417-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482496|T201|OSN|1417-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482496|T201|LC|1417-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482496|T201|LN|1417-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482496|T201|DN|1417-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482496|T201|MTH_LN|1417-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482496|T201|OSN|1417-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482496|T201|LC|1417-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482497|T201|LN|1418-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482497|T201|DN|1418-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482497|T201|MTH_LN|1418-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482497|T201|OSN|1418-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482497|T201|LC|1418-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482497|T201|LN|1418-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482497|T201|DN|1418-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482497|T201|MTH_LN|1418-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482497|T201|OSN|1418-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482497|T201|LC|1418-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482497|T201|LN|1418-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482497|T201|DN|1418-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482497|T201|MTH_LN|1418-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482497|T201|OSN|1418-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482497|T201|LC|1418-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482498|T201|LN|1421-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482498|T201|DN|1421-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482498|T201|MTH_LN|1421-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482498|T201|OSN|1421-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482498|T201|LC|1421-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482498|T201|LN|1421-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482498|T201|DN|1421-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482498|T201|MTH_LN|1421-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482498|T201|OSN|1421-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482498|T201|LC|1421-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482498|T201|LN|1421-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482498|T201|DN|1421-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482498|T201|MTH_LN|1421-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482498|T201|OSN|1421-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482498|T201|LC|1421-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482499|T201|LN|1422-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482499|T201|DN|1422-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482499|T201|MTH_LN|1422-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482499|T201|OSN|1422-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482499|T201|LC|1422-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482499|T201|LN|1422-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482499|T201|DN|1422-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482499|T201|MTH_LN|1422-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482499|T201|OSN|1422-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482499|T201|LC|1422-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482499|T201|LN|1422-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482499|T201|DN|1422-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482499|T201|MTH_LN|1422-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482499|T201|OSN|1422-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482499|T201|LC|1422-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482501|T201|LN|1426-6|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482501|T201|DN|1426-6|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482501|T201|MTH_LN|1426-6|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482501|T201|OSN|1426-6|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482501|T201|LC|1426-6|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482501|T201|LN|1426-6|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482501|T201|DN|1426-6|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482501|T201|MTH_LN|1426-6|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482501|T201|OSN|1426-6|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482501|T201|LC|1426-6|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482501|T201|LN|1426-6|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482501|T201|DN|1426-6|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482501|T201|MTH_LN|1426-6|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482501|T201|OSN|1426-6|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482501|T201|LC|1426-6|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482504|T201|LN|1430-8|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482504|T201|DN|1430-8|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482504|T201|MTH_LN|1430-8|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482504|T201|OSN|1430-8|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482504|T201|LC|1430-8|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482504|T201|LN|1430-8|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482504|T201|DN|1430-8|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482504|T201|MTH_LN|1430-8|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482504|T201|OSN|1430-8|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482504|T201|LC|1430-8|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482504|T201|LN|1430-8|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482504|T201|DN|1430-8|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482504|T201|MTH_LN|1430-8|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482504|T201|OSN|1430-8|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482504|T201|LC|1430-8|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482508|T201|LN|1438-1|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482508|T201|DN|1438-1|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482508|T201|MTH_LN|1438-1|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482508|T201|OSN|1438-1|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482508|T201|LC|1438-1|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482508|T201|LN|1438-1|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482508|T201|DN|1438-1|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482508|T201|MTH_LN|1438-1|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482508|T201|OSN|1438-1|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482508|T201|LC|1438-1|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482508|T201|LN|1438-1|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482508|T201|DN|1438-1|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482508|T201|MTH_LN|1438-1|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482508|T201|OSN|1438-1|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482508|T201|LC|1438-1|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482513|T201|LN|1447-2|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482513|T201|DN|1447-2|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482513|T201|MTH_LN|1447-2|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482513|T201|OSN|1447-2|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482513|T201|LC|1447-2|LNC2HPO|Hypocortisolism|Hypocortisolism
C0482513|T201|LN|1447-2|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482513|T201|DN|1447-2|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482513|T201|MTH_LN|1447-2|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482513|T201|OSN|1447-2|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482513|T201|LC|1447-2|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0482513|T201|LN|1447-2|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482513|T201|DN|1447-2|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482513|T201|MTH_LN|1447-2|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482513|T201|OSN|1447-2|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0482513|T201|LC|1447-2|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0881654|T201|LN|24389-9|LNC2HPO|Cushing syndrome|Cushing syndrome
C0881654|T201|DN|24389-9|LNC2HPO|Cushing syndrome|Cushing syndrome
C0881654|T201|MTH_LN|24389-9|LNC2HPO|Cushing syndrome|Cushing syndrome
C0881654|T201|OSN|24389-9|LNC2HPO|Cushing syndrome|Cushing syndrome
C0881654|T201|LC|24389-9|LNC2HPO|Cushing syndrome|Cushing syndrome
C0881654|T201|LN|24389-9|LNC2HPO|Hypercortisolism|Hypercortisolism
C0881654|T201|DN|24389-9|LNC2HPO|Hypercortisolism|Hypercortisolism
C0881654|T201|MTH_LN|24389-9|LNC2HPO|Hypercortisolism|Hypercortisolism
C0881654|T201|OSN|24389-9|LNC2HPO|Hypercortisolism|Hypercortisolism
C0881654|T201|LC|24389-9|LNC2HPO|Hypercortisolism|Hypercortisolism
C0881654|T201|LN|24389-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C0881654|T201|DN|24389-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C0881654|T201|MTH_LN|24389-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C0881654|T201|OSN|24389-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C0881654|T201|LC|24389-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C0881654|T201|LN|24389-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0881654|T201|DN|24389-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0881654|T201|MTH_LN|24389-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0881654|T201|OSN|24389-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0881654|T201|LC|24389-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0881654|T201|LN|24389-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0881654|T201|DN|24389-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0881654|T201|MTH_LN|24389-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0881654|T201|OSN|24389-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0881654|T201|LC|24389-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1978030|T201|LN|50171-8|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C1978030|T201|DN|50171-8|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C1978030|T201|OSN|50171-8|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C1978030|T201|MTH_LN|50171-8|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C1978030|T201|LC|50171-8|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C1978030|T201|LN|50171-8|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C1978030|T201|DN|50171-8|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C1978030|T201|OSN|50171-8|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C1978030|T201|MTH_LN|50171-8|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C1978030|T201|LC|50171-8|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C1978031|T201|LN|50172-6|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C1978031|T201|DN|50172-6|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C1978031|T201|OSN|50172-6|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C1978031|T201|MTH_LN|50172-6|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C1978031|T201|LC|50172-6|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C1978031|T201|LN|50172-6|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C1978031|T201|DN|50172-6|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C1978031|T201|OSN|50172-6|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C1978031|T201|MTH_LN|50172-6|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C1978031|T201|LC|50172-6|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C1978032|T201|LN|50173-4|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C1978032|T201|DN|50173-4|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C1978032|T201|MTH_LN|50173-4|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C1978032|T201|OSN|50173-4|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C1978032|T201|LC|50173-4|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C1978032|T201|LN|50173-4|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C1978032|T201|DN|50173-4|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C1978032|T201|MTH_LN|50173-4|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C1978032|T201|OSN|50173-4|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C1978032|T201|LC|50173-4|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C1369886|T201|MTH_LN|35094-2|LNC2HPO|Hypertension|Hypertension
C1369886|T201|LN|35094-2|LNC2HPO|Hypertension|Hypertension
C1369886|T201|LC|35094-2|LNC2HPO|Hypertension|Hypertension
C1369886|T201|OSN|35094-2|LNC2HPO|Hypertension|Hypertension
C1369886|T201|MTH_LN|35094-2|LNC2HPO|Systemic hypertension|Systemic hypertension
C1369886|T201|LN|35094-2|LNC2HPO|Systemic hypertension|Systemic hypertension
C1369886|T201|LC|35094-2|LNC2HPO|Systemic hypertension|Systemic hypertension
C1369886|T201|OSN|35094-2|LNC2HPO|Systemic hypertension|Systemic hypertension
C1369886|T201|MTH_LN|35094-2|LNC2HPO|Hypotension|Hypotension
C1369886|T201|LN|35094-2|LNC2HPO|Hypotension|Hypotension
C1369886|T201|LC|35094-2|LNC2HPO|Hypotension|Hypotension
C1369886|T201|OSN|35094-2|LNC2HPO|Hypotension|Hypotension
C1369886|T201|MTH_LN|35094-2|LNC2HPO|Arterial hypotension|Arterial hypotension
C1369886|T201|LN|35094-2|LNC2HPO|Arterial hypotension|Arterial hypotension
C1369886|T201|LC|35094-2|LNC2HPO|Arterial hypotension|Arterial hypotension
C1369886|T201|OSN|35094-2|LNC2HPO|Arterial hypotension|Arterial hypotension
C0362892|T201|LN|704-7|LNC2HPO|Basophilia|Basophilia
C0362892|T201|DN|704-7|LNC2HPO|Basophilia|Basophilia
C0362892|T201|OSN|704-7|LNC2HPO|Basophilia|Basophilia
C0362892|T201|MTH_LN|704-7|LNC2HPO|Basophilia|Basophilia
C0362892|T201|LC|704-7|LNC2HPO|Basophilia|Basophilia
C0362893|T201|LN|705-4|LNC2HPO|Basophilia|Basophilia
C0362893|T201|DN|705-4|LNC2HPO|Basophilia|Basophilia
C0362893|T201|OSN|705-4|LNC2HPO|Basophilia|Basophilia
C0362893|T201|MTH_LN|705-4|LNC2HPO|Basophilia|Basophilia
C0362893|T201|LC|705-4|LNC2HPO|Basophilia|Basophilia
C0367984|T201|LN|5769-5|LNC2HPO|Bacteriuria|Bacteriuria
C0367984|T201|DN|5769-5|LNC2HPO|Bacteriuria|Bacteriuria
C0367984|T201|MTH_LN|5769-5|LNC2HPO|Bacteriuria|Bacteriuria
C0367984|T201|OSN|5769-5|LNC2HPO|Bacteriuria|Bacteriuria
C0367984|T201|LC|5769-5|LNC2HPO|Bacteriuria|Bacteriuria
C0798106|T201|LN|14933-6|LNC2HPO|Hyperuricemia|Hyperuricemia
C0798106|T201|MTH_LN|14933-6|LNC2HPO|Hyperuricemia|Hyperuricemia
C0798106|T201|DN|14933-6|LNC2HPO|Hyperuricemia|Hyperuricemia
C0798106|T201|OSN|14933-6|LNC2HPO|Hyperuricemia|Hyperuricemia
C0798106|T201|LC|14933-6|LNC2HPO|Hyperuricemia|Hyperuricemia
C0798106|T201|LN|14933-6|LNC2HPO|Hyperuricaemia|Hyperuricaemia
C0798106|T201|MTH_LN|14933-6|LNC2HPO|Hyperuricaemia|Hyperuricaemia
C0798106|T201|DN|14933-6|LNC2HPO|Hyperuricaemia|Hyperuricaemia
C0798106|T201|OSN|14933-6|LNC2HPO|Hyperuricaemia|Hyperuricaemia
C0798106|T201|LC|14933-6|LNC2HPO|Hyperuricaemia|Hyperuricaemia
C0798106|T201|LN|14933-6|LNC2HPO|Hypouricemia|Hypouricemia
C0798106|T201|MTH_LN|14933-6|LNC2HPO|Hypouricemia|Hypouricemia
C0798106|T201|DN|14933-6|LNC2HPO|Hypouricemia|Hypouricemia
C0798106|T201|OSN|14933-6|LNC2HPO|Hypouricemia|Hypouricemia
C0798106|T201|LC|14933-6|LNC2HPO|Hypouricemia|Hypouricemia
C2363286|T201|MTH_LN|35232-8|LNC2HPO|Hyperuricemia|Hyperuricemia
C2363286|T201|DN|35232-8|LNC2HPO|Hyperuricemia|Hyperuricemia
C2363286|T201|LN|35232-8|LNC2HPO|Hyperuricemia|Hyperuricemia
C2363286|T201|OSN|35232-8|LNC2HPO|Hyperuricemia|Hyperuricemia
C2363286|T201|LC|35232-8|LNC2HPO|Hyperuricemia|Hyperuricemia
C2363286|T201|MTH_LN|35232-8|LNC2HPO|Hyperuricaemia|Hyperuricaemia
C2363286|T201|DN|35232-8|LNC2HPO|Hyperuricaemia|Hyperuricaemia
C2363286|T201|LN|35232-8|LNC2HPO|Hyperuricaemia|Hyperuricaemia
C2363286|T201|OSN|35232-8|LNC2HPO|Hyperuricaemia|Hyperuricaemia
C2363286|T201|LC|35232-8|LNC2HPO|Hyperuricaemia|Hyperuricaemia
C2363286|T201|MTH_LN|35232-8|LNC2HPO|Hypouricemia|Hypouricemia
C2363286|T201|DN|35232-8|LNC2HPO|Hypouricemia|Hypouricemia
C2363286|T201|LN|35232-8|LNC2HPO|Hypouricemia|Hypouricemia
C2363286|T201|OSN|35232-8|LNC2HPO|Hypouricemia|Hypouricemia
C2363286|T201|LC|35232-8|LNC2HPO|Hypouricemia|Hypouricemia
C1315270|T201|LN|32799-9|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C1315270|T201|OSN|32799-9|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C1315270|T201|MTH_LN|32799-9|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C1315270|T201|DN|32799-9|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C1315270|T201|LC|32799-9|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C1715600|T201|LN|44366-3|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C1715600|T201|OSN|44366-3|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C1715600|T201|MTH_LN|44366-3|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C1715600|T201|DN|44366-3|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C1715600|T201|LC|44366-3|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C1715601|T201|LN|44367-1|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C1715601|T201|DN|44367-1|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C1715601|T201|OSN|44367-1|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C1715601|T201|LC|44367-1|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C1715601|T201|MTH_LN|44367-1|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C1717153|T201|LN|46132-7|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C1717153|T201|DN|46132-7|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C1717153|T201|MTH_LN|46132-7|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C1717153|T201|OSN|46132-7|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C1717153|T201|LC|46132-7|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C3847306|T201|LN|74631-3|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C3847306|T201|OSN|74631-3|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C3847306|T201|MTH_LN|74631-3|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C3847306|T201|LC|74631-3|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C3847306|T201|DN|74631-3|LNC2HPO|Urinary glycosaminoglycan excretion|Urinary glycosaminoglycan excretion
C0881655|T201|LN|24390-7|LNC2HPO|Cushing syndrome|Cushing syndrome
C0881655|T201|DN|24390-7|LNC2HPO|Cushing syndrome|Cushing syndrome
C0881655|T201|MTH_LN|24390-7|LNC2HPO|Cushing syndrome|Cushing syndrome
C0881655|T201|OSN|24390-7|LNC2HPO|Cushing syndrome|Cushing syndrome
C0881655|T201|LC|24390-7|LNC2HPO|Cushing syndrome|Cushing syndrome
C0881655|T201|LN|24390-7|LNC2HPO|Hypercortisolism|Hypercortisolism
C0881655|T201|DN|24390-7|LNC2HPO|Hypercortisolism|Hypercortisolism
C0881655|T201|MTH_LN|24390-7|LNC2HPO|Hypercortisolism|Hypercortisolism
C0881655|T201|OSN|24390-7|LNC2HPO|Hypercortisolism|Hypercortisolism
C0881655|T201|LC|24390-7|LNC2HPO|Hypercortisolism|Hypercortisolism
C0881655|T201|LN|24390-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0881655|T201|DN|24390-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0881655|T201|MTH_LN|24390-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0881655|T201|OSN|24390-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0881655|T201|LC|24390-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0881655|T201|LN|24390-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0881655|T201|DN|24390-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0881655|T201|MTH_LN|24390-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0881655|T201|OSN|24390-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0881655|T201|LC|24390-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0881655|T201|LN|24390-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0881655|T201|DN|24390-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0881655|T201|MTH_LN|24390-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0881655|T201|OSN|24390-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0881655|T201|LC|24390-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0881656|T201|LN|24391-5|LNC2HPO|Cushing syndrome|Cushing syndrome
C0881656|T201|DN|24391-5|LNC2HPO|Cushing syndrome|Cushing syndrome
C0881656|T201|MTH_LN|24391-5|LNC2HPO|Cushing syndrome|Cushing syndrome
C0881656|T201|OSN|24391-5|LNC2HPO|Cushing syndrome|Cushing syndrome
C0881656|T201|LC|24391-5|LNC2HPO|Cushing syndrome|Cushing syndrome
C0881656|T201|LN|24391-5|LNC2HPO|Hypercortisolism|Hypercortisolism
C0881656|T201|DN|24391-5|LNC2HPO|Hypercortisolism|Hypercortisolism
C0881656|T201|MTH_LN|24391-5|LNC2HPO|Hypercortisolism|Hypercortisolism
C0881656|T201|OSN|24391-5|LNC2HPO|Hypercortisolism|Hypercortisolism
C0881656|T201|LC|24391-5|LNC2HPO|Hypercortisolism|Hypercortisolism
C0881656|T201|LN|24391-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0881656|T201|DN|24391-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0881656|T201|MTH_LN|24391-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0881656|T201|OSN|24391-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0881656|T201|LC|24391-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0881656|T201|LN|24391-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0881656|T201|DN|24391-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0881656|T201|MTH_LN|24391-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0881656|T201|OSN|24391-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0881656|T201|LC|24391-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0881656|T201|LN|24391-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0881656|T201|DN|24391-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0881656|T201|MTH_LN|24391-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0881656|T201|OSN|24391-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0881656|T201|LC|24391-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942484|T201|LN|26528-0|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942484|T201|DN|26528-0|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942484|T201|MTH_LN|26528-0|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942484|T201|OSN|26528-0|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942484|T201|LC|26528-0|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942484|T201|LN|26528-0|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942484|T201|DN|26528-0|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942484|T201|MTH_LN|26528-0|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942484|T201|OSN|26528-0|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942484|T201|LC|26528-0|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942484|T201|LN|26528-0|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942484|T201|DN|26528-0|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942484|T201|MTH_LN|26528-0|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942484|T201|OSN|26528-0|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942484|T201|LC|26528-0|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942484|T201|LN|26528-0|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942484|T201|DN|26528-0|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942484|T201|MTH_LN|26528-0|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942484|T201|OSN|26528-0|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942484|T201|LC|26528-0|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942484|T201|LN|26528-0|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942484|T201|DN|26528-0|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942484|T201|MTH_LN|26528-0|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942484|T201|OSN|26528-0|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942484|T201|LC|26528-0|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942485|T201|LN|26529-8|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942485|T201|DN|26529-8|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942485|T201|MTH_LN|26529-8|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942485|T201|OSN|26529-8|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942485|T201|LC|26529-8|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942485|T201|LN|26529-8|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942485|T201|DN|26529-8|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942485|T201|MTH_LN|26529-8|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942485|T201|OSN|26529-8|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942485|T201|LC|26529-8|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942485|T201|LN|26529-8|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942485|T201|DN|26529-8|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942485|T201|MTH_LN|26529-8|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942485|T201|OSN|26529-8|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942485|T201|LC|26529-8|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942485|T201|LN|26529-8|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942485|T201|DN|26529-8|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942485|T201|MTH_LN|26529-8|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942485|T201|OSN|26529-8|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942485|T201|LC|26529-8|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942485|T201|LN|26529-8|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942485|T201|DN|26529-8|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942485|T201|MTH_LN|26529-8|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942485|T201|OSN|26529-8|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942485|T201|LC|26529-8|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942486|T201|LN|26530-6|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942486|T201|DN|26530-6|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942486|T201|MTH_LN|26530-6|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942486|T201|OSN|26530-6|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942486|T201|LC|26530-6|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942486|T201|LN|26530-6|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942486|T201|DN|26530-6|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942486|T201|MTH_LN|26530-6|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942486|T201|OSN|26530-6|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942486|T201|LC|26530-6|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942486|T201|LN|26530-6|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942486|T201|DN|26530-6|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942486|T201|MTH_LN|26530-6|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942486|T201|OSN|26530-6|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942486|T201|LC|26530-6|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942486|T201|LN|26530-6|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942486|T201|DN|26530-6|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942486|T201|MTH_LN|26530-6|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942486|T201|OSN|26530-6|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942486|T201|LC|26530-6|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942486|T201|LN|26530-6|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942486|T201|DN|26530-6|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942486|T201|MTH_LN|26530-6|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942486|T201|OSN|26530-6|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942486|T201|LC|26530-6|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942487|T201|LN|26531-4|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942487|T201|DN|26531-4|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942487|T201|MTH_LN|26531-4|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942487|T201|OSN|26531-4|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942487|T201|LC|26531-4|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942487|T201|LN|26531-4|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942487|T201|DN|26531-4|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942487|T201|MTH_LN|26531-4|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942487|T201|OSN|26531-4|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942487|T201|LC|26531-4|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942487|T201|LN|26531-4|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942487|T201|DN|26531-4|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942487|T201|MTH_LN|26531-4|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942487|T201|OSN|26531-4|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942487|T201|LC|26531-4|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942487|T201|LN|26531-4|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942487|T201|DN|26531-4|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942487|T201|MTH_LN|26531-4|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942487|T201|OSN|26531-4|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942487|T201|LC|26531-4|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942487|T201|LN|26531-4|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942487|T201|DN|26531-4|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942487|T201|MTH_LN|26531-4|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942487|T201|OSN|26531-4|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942487|T201|LC|26531-4|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0947220|T201|LN|26532-2|LNC2HPO|Cushing syndrome|Cushing syndrome
C0947220|T201|DN|26532-2|LNC2HPO|Cushing syndrome|Cushing syndrome
C0947220|T201|MTH_LN|26532-2|LNC2HPO|Cushing syndrome|Cushing syndrome
C0947220|T201|OSN|26532-2|LNC2HPO|Cushing syndrome|Cushing syndrome
C0947220|T201|LC|26532-2|LNC2HPO|Cushing syndrome|Cushing syndrome
C0947220|T201|LN|26532-2|LNC2HPO|Hypercortisolism|Hypercortisolism
C0947220|T201|DN|26532-2|LNC2HPO|Hypercortisolism|Hypercortisolism
C0947220|T201|MTH_LN|26532-2|LNC2HPO|Hypercortisolism|Hypercortisolism
C0947220|T201|OSN|26532-2|LNC2HPO|Hypercortisolism|Hypercortisolism
C0947220|T201|LC|26532-2|LNC2HPO|Hypercortisolism|Hypercortisolism
C0947220|T201|LN|26532-2|LNC2HPO|Hypocortisolism|Hypocortisolism
C0947220|T201|DN|26532-2|LNC2HPO|Hypocortisolism|Hypocortisolism
C0947220|T201|MTH_LN|26532-2|LNC2HPO|Hypocortisolism|Hypocortisolism
C0947220|T201|OSN|26532-2|LNC2HPO|Hypocortisolism|Hypocortisolism
C0947220|T201|LC|26532-2|LNC2HPO|Hypocortisolism|Hypocortisolism
C0947220|T201|LN|26532-2|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0947220|T201|DN|26532-2|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0947220|T201|MTH_LN|26532-2|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0947220|T201|OSN|26532-2|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0947220|T201|LC|26532-2|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0947220|T201|LN|26532-2|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0947220|T201|DN|26532-2|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0947220|T201|MTH_LN|26532-2|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0947220|T201|OSN|26532-2|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0947220|T201|LC|26532-2|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0945367|T201|LN|26533-0|LNC2HPO|Cushing syndrome|Cushing syndrome
C0945367|T201|DN|26533-0|LNC2HPO|Cushing syndrome|Cushing syndrome
C0945367|T201|MTH_LN|26533-0|LNC2HPO|Cushing syndrome|Cushing syndrome
C0945367|T201|OSN|26533-0|LNC2HPO|Cushing syndrome|Cushing syndrome
C0945367|T201|LC|26533-0|LNC2HPO|Cushing syndrome|Cushing syndrome
C0945367|T201|LN|26533-0|LNC2HPO|Hypercortisolism|Hypercortisolism
C0945367|T201|DN|26533-0|LNC2HPO|Hypercortisolism|Hypercortisolism
C0945367|T201|MTH_LN|26533-0|LNC2HPO|Hypercortisolism|Hypercortisolism
C0945367|T201|OSN|26533-0|LNC2HPO|Hypercortisolism|Hypercortisolism
C0945367|T201|LC|26533-0|LNC2HPO|Hypercortisolism|Hypercortisolism
C0945367|T201|LN|26533-0|LNC2HPO|Hypocortisolism|Hypocortisolism
C0945367|T201|DN|26533-0|LNC2HPO|Hypocortisolism|Hypocortisolism
C0945367|T201|MTH_LN|26533-0|LNC2HPO|Hypocortisolism|Hypocortisolism
C0945367|T201|OSN|26533-0|LNC2HPO|Hypocortisolism|Hypocortisolism
C0945367|T201|LC|26533-0|LNC2HPO|Hypocortisolism|Hypocortisolism
C0945367|T201|LN|26533-0|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0945367|T201|DN|26533-0|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0945367|T201|MTH_LN|26533-0|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0945367|T201|OSN|26533-0|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0945367|T201|LC|26533-0|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0945367|T201|LN|26533-0|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0945367|T201|DN|26533-0|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0945367|T201|MTH_LN|26533-0|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0945367|T201|OSN|26533-0|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0945367|T201|LC|26533-0|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942488|T201|LN|26534-8|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942488|T201|DN|26534-8|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942488|T201|MTH_LN|26534-8|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942488|T201|OSN|26534-8|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942488|T201|LC|26534-8|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942488|T201|LN|26534-8|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942488|T201|DN|26534-8|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942488|T201|MTH_LN|26534-8|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942488|T201|OSN|26534-8|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942488|T201|LC|26534-8|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942488|T201|LN|26534-8|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942488|T201|DN|26534-8|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942488|T201|MTH_LN|26534-8|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942488|T201|OSN|26534-8|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942488|T201|LC|26534-8|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942488|T201|LN|26534-8|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942488|T201|DN|26534-8|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942488|T201|MTH_LN|26534-8|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942488|T201|OSN|26534-8|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942488|T201|LC|26534-8|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942488|T201|LN|26534-8|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942488|T201|DN|26534-8|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942488|T201|MTH_LN|26534-8|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942488|T201|OSN|26534-8|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942488|T201|LC|26534-8|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942489|T201|LN|26535-5|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942489|T201|DN|26535-5|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942489|T201|MTH_LN|26535-5|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942489|T201|OSN|26535-5|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942489|T201|LC|26535-5|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942489|T201|LN|26535-5|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942489|T201|DN|26535-5|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942489|T201|MTH_LN|26535-5|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942489|T201|OSN|26535-5|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942489|T201|LC|26535-5|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942489|T201|LN|26535-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942489|T201|DN|26535-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942489|T201|MTH_LN|26535-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942489|T201|OSN|26535-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942489|T201|LC|26535-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942489|T201|LN|26535-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942489|T201|DN|26535-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942489|T201|MTH_LN|26535-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942489|T201|OSN|26535-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942489|T201|LC|26535-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942489|T201|LN|26535-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942489|T201|DN|26535-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942489|T201|MTH_LN|26535-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942489|T201|OSN|26535-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942489|T201|LC|26535-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942490|T201|LN|26536-3|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942490|T201|DN|26536-3|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942490|T201|MTH_LN|26536-3|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942490|T201|OSN|26536-3|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942490|T201|LC|26536-3|LNC2HPO|Cushing syndrome|Cushing syndrome
C0942490|T201|LN|26536-3|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942490|T201|DN|26536-3|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942490|T201|MTH_LN|26536-3|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942490|T201|OSN|26536-3|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942490|T201|LC|26536-3|LNC2HPO|Hypercortisolism|Hypercortisolism
C0942490|T201|LN|26536-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942490|T201|DN|26536-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942490|T201|MTH_LN|26536-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942490|T201|OSN|26536-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942490|T201|LC|26536-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C0942490|T201|LN|26536-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942490|T201|DN|26536-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942490|T201|MTH_LN|26536-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942490|T201|OSN|26536-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942490|T201|LC|26536-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0942490|T201|LN|26536-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942490|T201|DN|26536-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942490|T201|MTH_LN|26536-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942490|T201|OSN|26536-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0942490|T201|LC|26536-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1316528|T201|LN|34065-3|LNC2HPO|Cushing syndrome|Cushing syndrome
C1316528|T201|MTH_LN|34065-3|LNC2HPO|Cushing syndrome|Cushing syndrome
C1316528|T201|LC|34065-3|LNC2HPO|Cushing syndrome|Cushing syndrome
C1316528|T201|DN|34065-3|LNC2HPO|Cushing syndrome|Cushing syndrome
C1316528|T201|OSN|34065-3|LNC2HPO|Cushing syndrome|Cushing syndrome
C1316528|T201|LN|34065-3|LNC2HPO|Hypercortisolism|Hypercortisolism
C1316528|T201|MTH_LN|34065-3|LNC2HPO|Hypercortisolism|Hypercortisolism
C1316528|T201|LC|34065-3|LNC2HPO|Hypercortisolism|Hypercortisolism
C1316528|T201|DN|34065-3|LNC2HPO|Hypercortisolism|Hypercortisolism
C1316528|T201|OSN|34065-3|LNC2HPO|Hypercortisolism|Hypercortisolism
C1316528|T201|LN|34065-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C1316528|T201|MTH_LN|34065-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C1316528|T201|LC|34065-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C1316528|T201|DN|34065-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C1316528|T201|OSN|34065-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C1316528|T201|LN|34065-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1316528|T201|MTH_LN|34065-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1316528|T201|LC|34065-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1316528|T201|DN|34065-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1316528|T201|OSN|34065-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1316528|T201|LN|34065-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1316528|T201|MTH_LN|34065-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1316528|T201|LC|34065-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1316528|T201|DN|34065-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1316528|T201|OSN|34065-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1316938|T201|LN|34476-2|LNC2HPO|Cushing syndrome|Cushing syndrome
C1316938|T201|DN|34476-2|LNC2HPO|Cushing syndrome|Cushing syndrome
C1316938|T201|MTH_LN|34476-2|LNC2HPO|Cushing syndrome|Cushing syndrome
C1316938|T201|OSN|34476-2|LNC2HPO|Cushing syndrome|Cushing syndrome
C1316938|T201|LC|34476-2|LNC2HPO|Cushing syndrome|Cushing syndrome
C1316938|T201|LN|34476-2|LNC2HPO|Hypercortisolism|Hypercortisolism
C1316938|T201|DN|34476-2|LNC2HPO|Hypercortisolism|Hypercortisolism
C1316938|T201|MTH_LN|34476-2|LNC2HPO|Hypercortisolism|Hypercortisolism
C1316938|T201|OSN|34476-2|LNC2HPO|Hypercortisolism|Hypercortisolism
C1316938|T201|LC|34476-2|LNC2HPO|Hypercortisolism|Hypercortisolism
C1316938|T201|LN|34476-2|LNC2HPO|Hypocortisolism|Hypocortisolism
C1316938|T201|DN|34476-2|LNC2HPO|Hypocortisolism|Hypocortisolism
C1316938|T201|MTH_LN|34476-2|LNC2HPO|Hypocortisolism|Hypocortisolism
C1316938|T201|OSN|34476-2|LNC2HPO|Hypocortisolism|Hypocortisolism
C1316938|T201|LC|34476-2|LNC2HPO|Hypocortisolism|Hypocortisolism
C1316938|T201|LN|34476-2|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1316938|T201|DN|34476-2|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1316938|T201|MTH_LN|34476-2|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1316938|T201|OSN|34476-2|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1316938|T201|LC|34476-2|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1316938|T201|LN|34476-2|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1316938|T201|DN|34476-2|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1316938|T201|MTH_LN|34476-2|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1316938|T201|OSN|34476-2|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1316938|T201|LC|34476-2|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1649478|T201|LN|41407-8|LNC2HPO|Cushing syndrome|Cushing syndrome
C1649478|T201|DN|41407-8|LNC2HPO|Cushing syndrome|Cushing syndrome
C1649478|T201|OSN|41407-8|LNC2HPO|Cushing syndrome|Cushing syndrome
C1649478|T201|MTH_LN|41407-8|LNC2HPO|Cushing syndrome|Cushing syndrome
C1649478|T201|LC|41407-8|LNC2HPO|Cushing syndrome|Cushing syndrome
C1649478|T201|LN|41407-8|LNC2HPO|Hypercortisolism|Hypercortisolism
C1649478|T201|DN|41407-8|LNC2HPO|Hypercortisolism|Hypercortisolism
C1649478|T201|OSN|41407-8|LNC2HPO|Hypercortisolism|Hypercortisolism
C1649478|T201|MTH_LN|41407-8|LNC2HPO|Hypercortisolism|Hypercortisolism
C1649478|T201|LC|41407-8|LNC2HPO|Hypercortisolism|Hypercortisolism
C1649478|T201|LN|41407-8|LNC2HPO|Hypocortisolism|Hypocortisolism
C1649478|T201|DN|41407-8|LNC2HPO|Hypocortisolism|Hypocortisolism
C1649478|T201|OSN|41407-8|LNC2HPO|Hypocortisolism|Hypocortisolism
C1649478|T201|MTH_LN|41407-8|LNC2HPO|Hypocortisolism|Hypocortisolism
C1649478|T201|LC|41407-8|LNC2HPO|Hypocortisolism|Hypocortisolism
C1649478|T201|LN|41407-8|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1649478|T201|DN|41407-8|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1649478|T201|OSN|41407-8|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1649478|T201|MTH_LN|41407-8|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1649478|T201|LC|41407-8|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1649478|T201|LN|41407-8|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1649478|T201|DN|41407-8|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1649478|T201|OSN|41407-8|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1649478|T201|MTH_LN|41407-8|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1649478|T201|LC|41407-8|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1952839|T201|LN|47608-5|LNC2HPO|Cushing syndrome|Cushing syndrome
C1952839|T201|DN|47608-5|LNC2HPO|Cushing syndrome|Cushing syndrome
C1952839|T201|OSN|47608-5|LNC2HPO|Cushing syndrome|Cushing syndrome
C1952839|T201|MTH_LN|47608-5|LNC2HPO|Cushing syndrome|Cushing syndrome
C1952839|T201|LC|47608-5|LNC2HPO|Cushing syndrome|Cushing syndrome
C1952839|T201|LN|47608-5|LNC2HPO|Hypercortisolism|Hypercortisolism
C1952839|T201|DN|47608-5|LNC2HPO|Hypercortisolism|Hypercortisolism
C1952839|T201|OSN|47608-5|LNC2HPO|Hypercortisolism|Hypercortisolism
C1952839|T201|MTH_LN|47608-5|LNC2HPO|Hypercortisolism|Hypercortisolism
C1952839|T201|LC|47608-5|LNC2HPO|Hypercortisolism|Hypercortisolism
C1952839|T201|LN|47608-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C1952839|T201|DN|47608-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C1952839|T201|OSN|47608-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C1952839|T201|MTH_LN|47608-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C1952839|T201|LC|47608-5|LNC2HPO|Hypocortisolism|Hypocortisolism
C1952839|T201|LN|47608-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1952839|T201|DN|47608-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1952839|T201|OSN|47608-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1952839|T201|MTH_LN|47608-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1952839|T201|LC|47608-5|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1952839|T201|LN|47608-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1952839|T201|DN|47608-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1952839|T201|OSN|47608-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1952839|T201|MTH_LN|47608-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1952839|T201|LC|47608-5|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1953170|T201|LN|47850-3|LNC2HPO|Cushing syndrome|Cushing syndrome
C1953170|T201|DN|47850-3|LNC2HPO|Cushing syndrome|Cushing syndrome
C1953170|T201|MTH_LN|47850-3|LNC2HPO|Cushing syndrome|Cushing syndrome
C1953170|T201|OSN|47850-3|LNC2HPO|Cushing syndrome|Cushing syndrome
C1953170|T201|LC|47850-3|LNC2HPO|Cushing syndrome|Cushing syndrome
C1953170|T201|LN|47850-3|LNC2HPO|Hypercortisolism|Hypercortisolism
C1953170|T201|DN|47850-3|LNC2HPO|Hypercortisolism|Hypercortisolism
C1953170|T201|MTH_LN|47850-3|LNC2HPO|Hypercortisolism|Hypercortisolism
C1953170|T201|OSN|47850-3|LNC2HPO|Hypercortisolism|Hypercortisolism
C1953170|T201|LC|47850-3|LNC2HPO|Hypercortisolism|Hypercortisolism
C1953170|T201|LN|47850-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C1953170|T201|DN|47850-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C1953170|T201|MTH_LN|47850-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C1953170|T201|OSN|47850-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C1953170|T201|LC|47850-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C1953170|T201|LN|47850-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1953170|T201|DN|47850-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1953170|T201|MTH_LN|47850-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1953170|T201|OSN|47850-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1953170|T201|LC|47850-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1953170|T201|LN|47850-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1953170|T201|DN|47850-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1953170|T201|MTH_LN|47850-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1953170|T201|OSN|47850-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1953170|T201|LC|47850-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1977844|T201|LN|49968-1|LNC2HPO|Cushing syndrome|Cushing syndrome
C1977844|T201|OSN|49968-1|LNC2HPO|Cushing syndrome|Cushing syndrome
C1977844|T201|DN|49968-1|LNC2HPO|Cushing syndrome|Cushing syndrome
C1977844|T201|MTH_LN|49968-1|LNC2HPO|Cushing syndrome|Cushing syndrome
C1977844|T201|LC|49968-1|LNC2HPO|Cushing syndrome|Cushing syndrome
C1977844|T201|LN|49968-1|LNC2HPO|Hypercortisolism|Hypercortisolism
C1977844|T201|OSN|49968-1|LNC2HPO|Hypercortisolism|Hypercortisolism
C1977844|T201|DN|49968-1|LNC2HPO|Hypercortisolism|Hypercortisolism
C1977844|T201|MTH_LN|49968-1|LNC2HPO|Hypercortisolism|Hypercortisolism
C1977844|T201|LC|49968-1|LNC2HPO|Hypercortisolism|Hypercortisolism
C1977844|T201|LN|49968-1|LNC2HPO|Hypocortisolism|Hypocortisolism
C1977844|T201|OSN|49968-1|LNC2HPO|Hypocortisolism|Hypocortisolism
C1977844|T201|DN|49968-1|LNC2HPO|Hypocortisolism|Hypocortisolism
C1977844|T201|MTH_LN|49968-1|LNC2HPO|Hypocortisolism|Hypocortisolism
C1977844|T201|LC|49968-1|LNC2HPO|Hypocortisolism|Hypocortisolism
C1977844|T201|LN|49968-1|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1977844|T201|OSN|49968-1|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1977844|T201|DN|49968-1|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1977844|T201|MTH_LN|49968-1|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1977844|T201|LC|49968-1|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1977844|T201|LN|49968-1|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1977844|T201|OSN|49968-1|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1977844|T201|DN|49968-1|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1977844|T201|MTH_LN|49968-1|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1977844|T201|LC|49968-1|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1977845|T201|LN|49969-9|LNC2HPO|Cushing syndrome|Cushing syndrome
C1977845|T201|OSN|49969-9|LNC2HPO|Cushing syndrome|Cushing syndrome
C1977845|T201|DN|49969-9|LNC2HPO|Cushing syndrome|Cushing syndrome
C1977845|T201|MTH_LN|49969-9|LNC2HPO|Cushing syndrome|Cushing syndrome
C1977845|T201|LC|49969-9|LNC2HPO|Cushing syndrome|Cushing syndrome
C1977845|T201|LN|49969-9|LNC2HPO|Hypercortisolism|Hypercortisolism
C1977845|T201|OSN|49969-9|LNC2HPO|Hypercortisolism|Hypercortisolism
C1977845|T201|DN|49969-9|LNC2HPO|Hypercortisolism|Hypercortisolism
C1977845|T201|MTH_LN|49969-9|LNC2HPO|Hypercortisolism|Hypercortisolism
C1977845|T201|LC|49969-9|LNC2HPO|Hypercortisolism|Hypercortisolism
C1977845|T201|LN|49969-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C1977845|T201|OSN|49969-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C1977845|T201|DN|49969-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C1977845|T201|MTH_LN|49969-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C1977845|T201|LC|49969-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C1977845|T201|LN|49969-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1977845|T201|OSN|49969-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1977845|T201|DN|49969-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1977845|T201|MTH_LN|49969-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1977845|T201|LC|49969-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C1977845|T201|LN|49969-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1977845|T201|OSN|49969-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1977845|T201|DN|49969-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1977845|T201|MTH_LN|49969-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C1977845|T201|LC|49969-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C2706775|T201|LN|54213-4|LNC2HPO|Cushing syndrome|Cushing syndrome
C2706775|T201|DN|54213-4|LNC2HPO|Cushing syndrome|Cushing syndrome
C2706775|T201|OSN|54213-4|LNC2HPO|Cushing syndrome|Cushing syndrome
C2706775|T201|MTH_LN|54213-4|LNC2HPO|Cushing syndrome|Cushing syndrome
C2706775|T201|LC|54213-4|LNC2HPO|Cushing syndrome|Cushing syndrome
C2706775|T201|LN|54213-4|LNC2HPO|Hypercortisolism|Hypercortisolism
C2706775|T201|DN|54213-4|LNC2HPO|Hypercortisolism|Hypercortisolism
C2706775|T201|OSN|54213-4|LNC2HPO|Hypercortisolism|Hypercortisolism
C2706775|T201|MTH_LN|54213-4|LNC2HPO|Hypercortisolism|Hypercortisolism
C2706775|T201|LC|54213-4|LNC2HPO|Hypercortisolism|Hypercortisolism
C2706775|T201|LN|54213-4|LNC2HPO|Hypocortisolism|Hypocortisolism
C2706775|T201|DN|54213-4|LNC2HPO|Hypocortisolism|Hypocortisolism
C2706775|T201|OSN|54213-4|LNC2HPO|Hypocortisolism|Hypocortisolism
C2706775|T201|MTH_LN|54213-4|LNC2HPO|Hypocortisolism|Hypocortisolism
C2706775|T201|LC|54213-4|LNC2HPO|Hypocortisolism|Hypocortisolism
C2706775|T201|LN|54213-4|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C2706775|T201|DN|54213-4|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C2706775|T201|OSN|54213-4|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C2706775|T201|MTH_LN|54213-4|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C2706775|T201|LC|54213-4|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C2706775|T201|LN|54213-4|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C2706775|T201|DN|54213-4|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C2706775|T201|OSN|54213-4|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C2706775|T201|MTH_LN|54213-4|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C2706775|T201|LC|54213-4|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C2706777|T201|LN|54215-9|LNC2HPO|Cushing syndrome|Cushing syndrome
C2706777|T201|DN|54215-9|LNC2HPO|Cushing syndrome|Cushing syndrome
C2706777|T201|OSN|54215-9|LNC2HPO|Cushing syndrome|Cushing syndrome
C2706777|T201|MTH_LN|54215-9|LNC2HPO|Cushing syndrome|Cushing syndrome
C2706777|T201|LC|54215-9|LNC2HPO|Cushing syndrome|Cushing syndrome
C2706777|T201|LN|54215-9|LNC2HPO|Hypercortisolism|Hypercortisolism
C2706777|T201|DN|54215-9|LNC2HPO|Hypercortisolism|Hypercortisolism
C2706777|T201|OSN|54215-9|LNC2HPO|Hypercortisolism|Hypercortisolism
C2706777|T201|MTH_LN|54215-9|LNC2HPO|Hypercortisolism|Hypercortisolism
C2706777|T201|LC|54215-9|LNC2HPO|Hypercortisolism|Hypercortisolism
C2706777|T201|LN|54215-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C2706777|T201|DN|54215-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C2706777|T201|OSN|54215-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C2706777|T201|MTH_LN|54215-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C2706777|T201|LC|54215-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C2706777|T201|LN|54215-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C2706777|T201|DN|54215-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C2706777|T201|OSN|54215-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C2706777|T201|MTH_LN|54215-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C2706777|T201|LC|54215-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C2706777|T201|LN|54215-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C2706777|T201|DN|54215-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C2706777|T201|OSN|54215-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C2706777|T201|MTH_LN|54215-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C2706777|T201|LC|54215-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484571|T201|LN|9612-3|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484571|T201|DN|9612-3|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484571|T201|MTH_LN|9612-3|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484571|T201|OSN|9612-3|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484571|T201|LC|9612-3|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484571|T201|LN|9612-3|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484571|T201|DN|9612-3|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484571|T201|MTH_LN|9612-3|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484571|T201|OSN|9612-3|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484571|T201|LC|9612-3|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484571|T201|LN|9612-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484571|T201|DN|9612-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484571|T201|MTH_LN|9612-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484571|T201|OSN|9612-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484571|T201|LC|9612-3|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484571|T201|LN|9612-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484571|T201|DN|9612-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484571|T201|MTH_LN|9612-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484571|T201|OSN|9612-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484571|T201|LC|9612-3|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484571|T201|LN|9612-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484571|T201|DN|9612-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484571|T201|MTH_LN|9612-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484571|T201|OSN|9612-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484571|T201|LC|9612-3|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484572|T201|LN|9613-1|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484572|T201|DN|9613-1|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484572|T201|MTH_LN|9613-1|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484572|T201|OSN|9613-1|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484572|T201|LC|9613-1|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484572|T201|LN|9613-1|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484572|T201|DN|9613-1|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484572|T201|MTH_LN|9613-1|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484572|T201|OSN|9613-1|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484572|T201|LC|9613-1|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484572|T201|LN|9613-1|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484572|T201|DN|9613-1|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484572|T201|MTH_LN|9613-1|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484572|T201|OSN|9613-1|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484572|T201|LC|9613-1|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484572|T201|LN|9613-1|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484572|T201|DN|9613-1|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484572|T201|MTH_LN|9613-1|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484572|T201|OSN|9613-1|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484572|T201|LC|9613-1|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484572|T201|LN|9613-1|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484572|T201|DN|9613-1|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484572|T201|MTH_LN|9613-1|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484572|T201|OSN|9613-1|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484572|T201|LC|9613-1|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484573|T201|LN|9614-9|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484573|T201|DN|9614-9|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484573|T201|MTH_LN|9614-9|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484573|T201|OSN|9614-9|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484573|T201|LC|9614-9|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484573|T201|LN|9614-9|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484573|T201|DN|9614-9|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484573|T201|MTH_LN|9614-9|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484573|T201|OSN|9614-9|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484573|T201|LC|9614-9|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484573|T201|LN|9614-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484573|T201|DN|9614-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484573|T201|MTH_LN|9614-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484573|T201|OSN|9614-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484573|T201|LC|9614-9|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484573|T201|LN|9614-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484573|T201|DN|9614-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484573|T201|MTH_LN|9614-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484573|T201|OSN|9614-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484573|T201|LC|9614-9|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484573|T201|LN|9614-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484573|T201|DN|9614-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484573|T201|MTH_LN|9614-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484573|T201|OSN|9614-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484573|T201|LC|9614-9|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484574|T201|LN|9615-6|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484574|T201|DN|9615-6|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484574|T201|OSN|9615-6|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484574|T201|MTH_LN|9615-6|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484574|T201|LC|9615-6|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484574|T201|LN|9615-6|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484574|T201|DN|9615-6|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484574|T201|OSN|9615-6|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484574|T201|MTH_LN|9615-6|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484574|T201|LC|9615-6|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484574|T201|LN|9615-6|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484574|T201|DN|9615-6|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484574|T201|OSN|9615-6|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484574|T201|MTH_LN|9615-6|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484574|T201|LC|9615-6|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484574|T201|LN|9615-6|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484574|T201|DN|9615-6|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484574|T201|OSN|9615-6|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484574|T201|MTH_LN|9615-6|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484574|T201|LC|9615-6|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484574|T201|LN|9615-6|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484574|T201|DN|9615-6|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484574|T201|OSN|9615-6|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484574|T201|MTH_LN|9615-6|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484574|T201|LC|9615-6|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0365228|T201|LC|3084-1|LNC2HPO|Hyperuricemia|Hyperuricemia
C0365228|T201|MTH_LN|3084-1|LNC2HPO|Hyperuricemia|Hyperuricemia
C0365228|T201|LN|3084-1|LNC2HPO|Hyperuricemia|Hyperuricemia
C0365228|T201|DN|3084-1|LNC2HPO|Hyperuricemia|Hyperuricemia
C0365228|T201|OSN|3084-1|LNC2HPO|Hyperuricemia|Hyperuricemia
C0365228|T201|LC|3084-1|LNC2HPO|Hyperuricaemia|Hyperuricaemia
C0365228|T201|MTH_LN|3084-1|LNC2HPO|Hyperuricaemia|Hyperuricaemia
C0365228|T201|LN|3084-1|LNC2HPO|Hyperuricaemia|Hyperuricaemia
C0365228|T201|DN|3084-1|LNC2HPO|Hyperuricaemia|Hyperuricaemia
C0365228|T201|OSN|3084-1|LNC2HPO|Hyperuricaemia|Hyperuricaemia
C0365228|T201|LC|3084-1|LNC2HPO|Hypouricemia|Hypouricemia
C0365228|T201|MTH_LN|3084-1|LNC2HPO|Hypouricemia|Hypouricemia
C0365228|T201|LN|3084-1|LNC2HPO|Hypouricemia|Hypouricemia
C0365228|T201|DN|3084-1|LNC2HPO|Hypouricemia|Hypouricemia
C0365228|T201|OSN|3084-1|LNC2HPO|Hypouricemia|Hypouricemia
C0942419|T201|LN|26449-9|LNC2HPO|Eosinophilia|Eosinophilia
C0942419|T201|DN|26449-9|LNC2HPO|Eosinophilia|Eosinophilia
C0942419|T201|OSN|26449-9|LNC2HPO|Eosinophilia|Eosinophilia
C0942419|T201|MTH_LN|26449-9|LNC2HPO|Eosinophilia|Eosinophilia
C0942419|T201|LC|26449-9|LNC2HPO|Eosinophilia|Eosinophilia
C0942440|T201|LN|26478-8|LNC2HPO|Lymphocytosis|Lymphocytosis
C0942440|T201|OSN|26478-8|LNC2HPO|Lymphocytosis|Lymphocytosis
C0942440|T201|DN|26478-8|LNC2HPO|Lymphocytosis|Lymphocytosis
C0942440|T201|MTH_LN|26478-8|LNC2HPO|Lymphocytosis|Lymphocytosis
C0942440|T201|LC|26478-8|LNC2HPO|Lymphocytosis|Lymphocytosis
C0942440|T201|LN|26478-8|LNC2HPO|Lymphopenia|Lymphopenia
C0942440|T201|OSN|26478-8|LNC2HPO|Lymphopenia|Lymphopenia
C0942440|T201|DN|26478-8|LNC2HPO|Lymphopenia|Lymphopenia
C0942440|T201|MTH_LN|26478-8|LNC2HPO|Lymphopenia|Lymphopenia
C0942440|T201|LC|26478-8|LNC2HPO|Lymphopenia|Lymphopenia
C0942440|T201|LN|26478-8|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0942440|T201|OSN|26478-8|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0942440|T201|DN|26478-8|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0942440|T201|MTH_LN|26478-8|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0942440|T201|LC|26478-8|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0942440|T201|LN|26478-8|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0942440|T201|OSN|26478-8|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0942440|T201|DN|26478-8|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0942440|T201|MTH_LN|26478-8|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0942440|T201|LC|26478-8|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0550259|T201|LN|12772-0|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0550259|T201|MTH_LN|12772-0|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0550259|T201|DN|12772-0|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0550259|T201|OSN|12772-0|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0550259|T201|LC|12772-0|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0550259|T201|LN|12772-0|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0550259|T201|MTH_LN|12772-0|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0550259|T201|DN|12772-0|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0550259|T201|OSN|12772-0|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0550259|T201|LC|12772-0|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0797821|T201|LN|14646-4|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0797821|T201|MTH_LN|14646-4|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0797821|T201|DN|14646-4|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0797821|T201|OSN|14646-4|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0797821|T201|LC|14646-4|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0797821|T201|LN|14646-4|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0797821|T201|MTH_LN|14646-4|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0797821|T201|DN|14646-4|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0797821|T201|OSN|14646-4|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0797821|T201|LC|14646-4|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0801309|T201|LN|18263-4|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0801309|T201|MTH_LN|18263-4|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0801309|T201|DN|18263-4|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0801309|T201|OSN|18263-4|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0801309|T201|LC|18263-4|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0801309|T201|LN|18263-4|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0801309|T201|MTH_LN|18263-4|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0801309|T201|DN|18263-4|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0801309|T201|OSN|18263-4|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0801309|T201|LC|18263-4|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0364221|T201|LC|2085-9|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0364221|T201|DN|2085-9|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0364221|T201|MTH_LN|2085-9|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0364221|T201|LN|2085-9|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0364221|T201|OSN|2085-9|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0364221|T201|LC|2085-9|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0364221|T201|DN|2085-9|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0364221|T201|MTH_LN|2085-9|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0364221|T201|LN|2085-9|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0364221|T201|OSN|2085-9|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C2713261|T201|OLC|2086-7|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C2713261|T201|DN|2086-7|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C2713261|T201|MTH_LO|2086-7|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C2713261|T201|LO|2086-7|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C2713261|T201|OOSN|2086-7|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C2713261|T201|OLC|2086-7|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C2713261|T201|DN|2086-7|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C2713261|T201|MTH_LO|2086-7|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C2713261|T201|LO|2086-7|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C2713261|T201|OOSN|2086-7|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C2603387|T201|DN|35197-3|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C2603387|T201|MTH_LN|35197-3|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C2603387|T201|LN|35197-3|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C2603387|T201|OSN|35197-3|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C2603387|T201|LC|35197-3|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C2603387|T201|DN|35197-3|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C2603387|T201|MTH_LN|35197-3|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C2603387|T201|LN|35197-3|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C2603387|T201|OSN|35197-3|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C2603387|T201|LC|35197-3|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C1954893|T201|LN|49130-8|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C1954893|T201|DN|49130-8|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C1954893|T201|MTH_LN|49130-8|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C1954893|T201|OSN|49130-8|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C1954893|T201|LC|49130-8|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C1954893|T201|LN|49130-8|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C1954893|T201|DN|49130-8|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C1954893|T201|MTH_LN|49130-8|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C1954893|T201|OSN|49130-8|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C1954893|T201|LC|49130-8|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C1315880|T201|LN|33411-0|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C1315880|T201|MTH_LN|33411-0|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C1315880|T201|DN|33411-0|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C1315880|T201|OSN|33411-0|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C1315880|T201|LC|33411-0|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C1316637|T201|LN|34174-3|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C1316637|T201|MTH_LN|34174-3|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C1316637|T201|DN|34174-3|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C1316637|T201|OSN|34174-3|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C1316637|T201|LC|34174-3|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0368020|T201|LN|5794-3|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0368020|T201|MTH_LN|5794-3|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0368020|T201|DN|5794-3|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0368020|T201|OSN|5794-3|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0368020|T201|LC|5794-3|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0362930|T201|LN|725-2|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0362930|T201|MTH_LN|725-2|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0362930|T201|DN|725-2|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0362930|T201|OSN|725-2|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0362930|T201|LC|725-2|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0797471|T201|OLC|14290-1|LNC2HPO|Hematuria|Hematuria
C0797471|T201|MTH_LO|14290-1|LNC2HPO|Hematuria|Hematuria
C0797471|T201|DN|14290-1|LNC2HPO|Hematuria|Hematuria
C0797471|T201|LO|14290-1|LNC2HPO|Hematuria|Hematuria
C0797471|T201|OOSN|14290-1|LNC2HPO|Hematuria|Hematuria
C0803224|T201|LN|20409-9|LNC2HPO|Hematuria|Hematuria
C0803224|T201|DN|20409-9|LNC2HPO|Hematuria|Hematuria
C0803224|T201|OSN|20409-9|LNC2HPO|Hematuria|Hematuria
C0803224|T201|MTH_LN|20409-9|LNC2HPO|Hematuria|Hematuria
C0803224|T201|LC|20409-9|LNC2HPO|Hematuria|Hematuria
C1114250|T201|LN|30391-7|LNC2HPO|Hematuria|Hematuria
C1114250|T201|DN|30391-7|LNC2HPO|Hematuria|Hematuria
C1114250|T201|OSN|30391-7|LNC2HPO|Hematuria|Hematuria
C1114250|T201|MTH_LN|30391-7|LNC2HPO|Hematuria|Hematuria
C1114250|T201|LC|30391-7|LNC2HPO|Hematuria|Hematuria
C1830308|T201|LN|46419-8|LNC2HPO|Hematuria|Hematuria
C1830308|T201|OSN|46419-8|LNC2HPO|Hematuria|Hematuria
C1830308|T201|MTH_LN|46419-8|LNC2HPO|Hematuria|Hematuria
C1830308|T201|LC|46419-8|LNC2HPO|Hematuria|Hematuria
C1830308|T201|DN|46419-8|LNC2HPO|Hematuria|Hematuria
C2736161|T201|LN|57747-8|LNC2HPO|Hematuria|Hematuria
C2736161|T201|DN|57747-8|LNC2HPO|Hematuria|Hematuria
C2736161|T201|LC|57747-8|LNC2HPO|Hematuria|Hematuria
C2736161|T201|MTH_LN|57747-8|LNC2HPO|Hematuria|Hematuria
C2736161|T201|OSN|57747-8|LNC2HPO|Hematuria|Hematuria
C3262756|T201|LN|68902-6|LNC2HPO|Hematuria|Hematuria
C3262756|T201|OSN|68902-6|LNC2HPO|Hematuria|Hematuria
C3262756|T201|MTH_LN|68902-6|LNC2HPO|Hematuria|Hematuria
C3262756|T201|LC|68902-6|LNC2HPO|Hematuria|Hematuria
C3262756|T201|DN|68902-6|LNC2HPO|Hematuria|Hematuria
C3262757|T201|LN|68903-4|LNC2HPO|Hematuria|Hematuria
C3262757|T201|OSN|68903-4|LNC2HPO|Hematuria|Hematuria
C3262757|T201|MTH_LN|68903-4|LNC2HPO|Hematuria|Hematuria
C3262757|T201|LC|68903-4|LNC2HPO|Hematuria|Hematuria
C3262757|T201|DN|68903-4|LNC2HPO|Hematuria|Hematuria
C0362919|T201|LN|798-9|LNC2HPO|Hematuria|Hematuria
C0362919|T201|DN|798-9|LNC2HPO|Hematuria|Hematuria
C0362919|T201|OSN|798-9|LNC2HPO|Hematuria|Hematuria
C0362919|T201|MTH_LN|798-9|LNC2HPO|Hematuria|Hematuria
C0362919|T201|LC|798-9|LNC2HPO|Hematuria|Hematuria
C0362920|T201|LN|799-7|LNC2HPO|Hematuria|Hematuria
C0362920|T201|DN|799-7|LNC2HPO|Hematuria|Hematuria
C0362920|T201|OSN|799-7|LNC2HPO|Hematuria|Hematuria
C0362920|T201|MTH_LN|799-7|LNC2HPO|Hematuria|Hematuria
C0362920|T201|LC|799-7|LNC2HPO|Hematuria|Hematuria
C1315522|T201|LN|33051-4|LNC2HPO|Hematuria|Hematuria
C1315522|T201|MTH_LN|33051-4|LNC2HPO|Hematuria|Hematuria
C1315522|T201|DN|33051-4|LNC2HPO|Hematuria|Hematuria
C1315522|T201|OSN|33051-4|LNC2HPO|Hematuria|Hematuria
C1315522|T201|LC|33051-4|LNC2HPO|Hematuria|Hematuria
C2361818|T201|LN|53292-9|LNC2HPO|Hematuria|Hematuria
C2361818|T201|MTH_LN|53292-9|LNC2HPO|Hematuria|Hematuria
C2361818|T201|DN|53292-9|LNC2HPO|Hematuria|Hematuria
C2361818|T201|OSN|53292-9|LNC2HPO|Hematuria|Hematuria
C2361818|T201|LC|53292-9|LNC2HPO|Hematuria|Hematuria
C0797133|T201|LN|13945-1|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C0797133|T201|DN|13945-1|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C0797133|T201|MTH_LN|13945-1|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C0797133|T201|OSN|13945-1|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C0797133|T201|LC|13945-1|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C0797133|T201|LN|13945-1|LNC2HPO|Microhematuria|Microhematuria
C0797133|T201|DN|13945-1|LNC2HPO|Microhematuria|Microhematuria
C0797133|T201|MTH_LN|13945-1|LNC2HPO|Microhematuria|Microhematuria
C0797133|T201|OSN|13945-1|LNC2HPO|Microhematuria|Microhematuria
C0797133|T201|LC|13945-1|LNC2HPO|Microhematuria|Microhematuria
C0797133|T201|LN|13945-1|LNC2HPO|Occult hematuria|Occult hematuria
C0797133|T201|DN|13945-1|LNC2HPO|Occult hematuria|Occult hematuria
C0797133|T201|MTH_LN|13945-1|LNC2HPO|Occult hematuria|Occult hematuria
C0797133|T201|OSN|13945-1|LNC2HPO|Occult hematuria|Occult hematuria
C0797133|T201|LC|13945-1|LNC2HPO|Occult hematuria|Occult hematuria
C0368013|T201|LN|5808-1|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C0368013|T201|DN|5808-1|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C0368013|T201|OSN|5808-1|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C0368013|T201|MTH_LN|5808-1|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C0368013|T201|LC|5808-1|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C0368013|T201|LN|5808-1|LNC2HPO|Microhematuria|Microhematuria
C0368013|T201|DN|5808-1|LNC2HPO|Microhematuria|Microhematuria
C0368013|T201|OSN|5808-1|LNC2HPO|Microhematuria|Microhematuria
C0368013|T201|MTH_LN|5808-1|LNC2HPO|Microhematuria|Microhematuria
C0368013|T201|LC|5808-1|LNC2HPO|Microhematuria|Microhematuria
C0368013|T201|LN|5808-1|LNC2HPO|Occult hematuria|Occult hematuria
C0368013|T201|DN|5808-1|LNC2HPO|Occult hematuria|Occult hematuria
C0368013|T201|OSN|5808-1|LNC2HPO|Occult hematuria|Occult hematuria
C0368013|T201|MTH_LN|5808-1|LNC2HPO|Occult hematuria|Occult hematuria
C0368013|T201|LC|5808-1|LNC2HPO|Occult hematuria|Occult hematuria
C2925974|T201|LN|58449-0|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C2925974|T201|DN|58449-0|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C2925974|T201|LC|58449-0|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C2925974|T201|OSN|58449-0|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C2925974|T201|MTH_LN|58449-0|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C2925974|T201|LN|58449-0|LNC2HPO|Microhematuria|Microhematuria
C2925974|T201|DN|58449-0|LNC2HPO|Microhematuria|Microhematuria
C2925974|T201|LC|58449-0|LNC2HPO|Microhematuria|Microhematuria
C2925974|T201|OSN|58449-0|LNC2HPO|Microhematuria|Microhematuria
C2925974|T201|MTH_LN|58449-0|LNC2HPO|Microhematuria|Microhematuria
C2925974|T201|LN|58449-0|LNC2HPO|Occult hematuria|Occult hematuria
C2925974|T201|DN|58449-0|LNC2HPO|Occult hematuria|Occult hematuria
C2925974|T201|LC|58449-0|LNC2HPO|Occult hematuria|Occult hematuria
C2925974|T201|OSN|58449-0|LNC2HPO|Occult hematuria|Occult hematuria
C2925974|T201|MTH_LN|58449-0|LNC2HPO|Occult hematuria|Occult hematuria
C2924078|T201|LN|59830-0|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C2924078|T201|DN|59830-0|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C2924078|T201|LC|59830-0|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C2924078|T201|OSN|59830-0|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C2924078|T201|MTH_LN|59830-0|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C2924078|T201|LN|59830-0|LNC2HPO|Microhematuria|Microhematuria
C2924078|T201|DN|59830-0|LNC2HPO|Microhematuria|Microhematuria
C2924078|T201|LC|59830-0|LNC2HPO|Microhematuria|Microhematuria
C2924078|T201|OSN|59830-0|LNC2HPO|Microhematuria|Microhematuria
C2924078|T201|MTH_LN|59830-0|LNC2HPO|Microhematuria|Microhematuria
C2924078|T201|LN|59830-0|LNC2HPO|Occult hematuria|Occult hematuria
C2924078|T201|DN|59830-0|LNC2HPO|Occult hematuria|Occult hematuria
C2924078|T201|LC|59830-0|LNC2HPO|Occult hematuria|Occult hematuria
C2924078|T201|OSN|59830-0|LNC2HPO|Occult hematuria|Occult hematuria
C2924078|T201|MTH_LN|59830-0|LNC2HPO|Occult hematuria|Occult hematuria
C3262760|T201|LN|68912-5|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C3262760|T201|MTH_LN|68912-5|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C3262760|T201|OSN|68912-5|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C3262760|T201|LC|68912-5|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C3262760|T201|DN|68912-5|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C3262760|T201|LN|68912-5|LNC2HPO|Microhematuria|Microhematuria
C3262760|T201|MTH_LN|68912-5|LNC2HPO|Microhematuria|Microhematuria
C3262760|T201|OSN|68912-5|LNC2HPO|Microhematuria|Microhematuria
C3262760|T201|LC|68912-5|LNC2HPO|Microhematuria|Microhematuria
C3262760|T201|DN|68912-5|LNC2HPO|Microhematuria|Microhematuria
C3262760|T201|LN|68912-5|LNC2HPO|Occult hematuria|Occult hematuria
C3262760|T201|MTH_LN|68912-5|LNC2HPO|Occult hematuria|Occult hematuria
C3262760|T201|OSN|68912-5|LNC2HPO|Occult hematuria|Occult hematuria
C3262760|T201|LC|68912-5|LNC2HPO|Occult hematuria|Occult hematuria
C3262760|T201|DN|68912-5|LNC2HPO|Occult hematuria|Occult hematuria
C1315247|T201|LN|32776-7|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C1315247|T201|MTH_LN|32776-7|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C1315247|T201|DN|32776-7|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C1315247|T201|OSN|32776-7|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C1315247|T201|LC|32776-7|LNC2HPO|Microscopic hematuria|Microscopic hematuria
C1315247|T201|LN|32776-7|LNC2HPO|Microhematuria|Microhematuria
C1315247|T201|MTH_LN|32776-7|LNC2HPO|Microhematuria|Microhematuria
C1315247|T201|DN|32776-7|LNC2HPO|Microhematuria|Microhematuria
C1315247|T201|OSN|32776-7|LNC2HPO|Microhematuria|Microhematuria
C1315247|T201|LC|32776-7|LNC2HPO|Microhematuria|Microhematuria
C1315247|T201|LN|32776-7|LNC2HPO|Occult hematuria|Occult hematuria
C1315247|T201|MTH_LN|32776-7|LNC2HPO|Occult hematuria|Occult hematuria
C1315247|T201|DN|32776-7|LNC2HPO|Occult hematuria|Occult hematuria
C1315247|T201|OSN|32776-7|LNC2HPO|Occult hematuria|Occult hematuria
C1315247|T201|LC|32776-7|LNC2HPO|Occult hematuria|Occult hematuria
C3172449|T201|LN|63378-4|LNC2HPO|Gross hematuria|Gross hematuria
C3172449|T201|OSN|63378-4|LNC2HPO|Gross hematuria|Gross hematuria
C3172449|T201|LC|63378-4|LNC2HPO|Gross hematuria|Gross hematuria
C3172449|T201|MTH_LN|63378-4|LNC2HPO|Gross hematuria|Gross hematuria
C3172449|T201|DN|63378-4|LNC2HPO|Gross hematuria|Gross hematuria
C3172449|T201|LN|63378-4|LNC2HPO|Macroscopic hematuria|Macroscopic hematuria
C3172449|T201|OSN|63378-4|LNC2HPO|Macroscopic hematuria|Macroscopic hematuria
C3172449|T201|LC|63378-4|LNC2HPO|Macroscopic hematuria|Macroscopic hematuria
C3172449|T201|MTH_LN|63378-4|LNC2HPO|Macroscopic hematuria|Macroscopic hematuria
C3172449|T201|DN|63378-4|LNC2HPO|Macroscopic hematuria|Macroscopic hematuria
C2361881|T201|LN|53358-8|LNC2HPO|Gross hematuria|Gross hematuria
C2361881|T201|DN|53358-8|LNC2HPO|Gross hematuria|Gross hematuria
C2361881|T201|MTH_LN|53358-8|LNC2HPO|Gross hematuria|Gross hematuria
C2361881|T201|OSN|53358-8|LNC2HPO|Gross hematuria|Gross hematuria
C2361881|T201|LC|53358-8|LNC2HPO|Gross hematuria|Gross hematuria
C2361881|T201|LN|53358-8|LNC2HPO|Macroscopic hematuria|Macroscopic hematuria
C2361881|T201|DN|53358-8|LNC2HPO|Macroscopic hematuria|Macroscopic hematuria
C2361881|T201|MTH_LN|53358-8|LNC2HPO|Macroscopic hematuria|Macroscopic hematuria
C2361881|T201|OSN|53358-8|LNC2HPO|Macroscopic hematuria|Macroscopic hematuria
C2361881|T201|LC|53358-8|LNC2HPO|Macroscopic hematuria|Macroscopic hematuria
C2361883|T201|LN|53360-4|LNC2HPO|Gross hematuria|Gross hematuria
C2361883|T201|DN|53360-4|LNC2HPO|Gross hematuria|Gross hematuria
C2361883|T201|MTH_LN|53360-4|LNC2HPO|Gross hematuria|Gross hematuria
C2361883|T201|OSN|53360-4|LNC2HPO|Gross hematuria|Gross hematuria
C2361883|T201|LC|53360-4|LNC2HPO|Gross hematuria|Gross hematuria
C2361883|T201|LN|53360-4|LNC2HPO|Macroscopic hematuria|Macroscopic hematuria
C2361883|T201|DN|53360-4|LNC2HPO|Macroscopic hematuria|Macroscopic hematuria
C2361883|T201|MTH_LN|53360-4|LNC2HPO|Macroscopic hematuria|Macroscopic hematuria
C2361883|T201|OSN|53360-4|LNC2HPO|Macroscopic hematuria|Macroscopic hematuria
C2361883|T201|LC|53360-4|LNC2HPO|Macroscopic hematuria|Macroscopic hematuria
C1977255|T201|LN|49505-1|LNC2HPO|Hematuria|Hematuria
C1977255|T201|LC|49505-1|LNC2HPO|Hematuria|Hematuria
C1977255|T201|MTH_LN|49505-1|LNC2HPO|Hematuria|Hematuria
C1977255|T201|OSN|49505-1|LNC2HPO|Hematuria|Hematuria
C1977255|T201|DN|49505-1|LNC2HPO|Hematuria|Hematuria
C1978061|T201|LN|50226-0|LNC2HPO|Hematuria|Hematuria
C1978061|T201|MTH_LN|50226-0|LNC2HPO|Hematuria|Hematuria
C1978061|T201|DN|50226-0|LNC2HPO|Hematuria|Hematuria
C1978061|T201|OSN|50226-0|LNC2HPO|Hematuria|Hematuria
C1978061|T201|LC|50226-0|LNC2HPO|Hematuria|Hematuria
C0363002|T201|LN|800-3|LNC2HPO|Schistocytosis|Schistocytosis
C0363002|T201|MTH_LN|800-3|LNC2HPO|Schistocytosis|Schistocytosis
C0363002|T201|DN|800-3|LNC2HPO|Schistocytosis|Schistocytosis
C0363002|T201|OSN|800-3|LNC2HPO|Schistocytosis|Schistocytosis
C0363002|T201|LC|800-3|LNC2HPO|Schistocytosis|Schistocytosis
C0363002|T201|LN|800-3|LNC2HPO|Schistocytes|Schistocytes
C0363002|T201|MTH_LN|800-3|LNC2HPO|Schistocytes|Schistocytes
C0363002|T201|DN|800-3|LNC2HPO|Schistocytes|Schistocytes
C0363002|T201|OSN|800-3|LNC2HPO|Schistocytes|Schistocytes
C0363002|T201|LC|800-3|LNC2HPO|Schistocytes|Schistocytes
C1543030|T201|LN|38908-0|LNC2HPO|Poikilocytosis|Poikilocytosis
C1543030|T201|MTH_LN|38908-0|LNC2HPO|Poikilocytosis|Poikilocytosis
C1543030|T201|OSN|38908-0|LNC2HPO|Poikilocytosis|Poikilocytosis
C1543030|T201|DN|38908-0|LNC2HPO|Poikilocytosis|Poikilocytosis
C1543030|T201|LC|38908-0|LNC2HPO|Poikilocytosis|Poikilocytosis
C2363247|T201|LN|779-9|LNC2HPO|Poikilocytosis|Poikilocytosis
C2363247|T201|MTH_LN|779-9|LNC2HPO|Poikilocytosis|Poikilocytosis
C2363247|T201|DN|779-9|LNC2HPO|Poikilocytosis|Poikilocytosis
C2363247|T201|OSN|779-9|LNC2HPO|Poikilocytosis|Poikilocytosis
C2363247|T201|LC|779-9|LNC2HPO|Poikilocytosis|Poikilocytosis
C0943152|T201|LN|27340-9|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0943152|T201|MTH_LN|27340-9|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0943152|T201|DN|27340-9|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0943152|T201|OSN|27340-9|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0943152|T201|LC|27340-9|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0368025|T201|LN|5796-8|LNC2HPO|Hyaline casts|Hyaline casts
C0368025|T201|DN|5796-8|LNC2HPO|Hyaline casts|Hyaline casts
C0368025|T201|MTH_LN|5796-8|LNC2HPO|Hyaline casts|Hyaline casts
C0368025|T201|OSN|5796-8|LNC2HPO|Hyaline casts|Hyaline casts
C0368025|T201|LC|5796-8|LNC2HPO|Hyaline casts|Hyaline casts
C1315694|T201|LN|33223-9|LNC2HPO|Hyaline casts|Hyaline casts
C1315694|T201|MTH_LN|33223-9|LNC2HPO|Hyaline casts|Hyaline casts
C1315694|T201|LC|33223-9|LNC2HPO|Hyaline casts|Hyaline casts
C1315694|T201|OSN|33223-9|LNC2HPO|Hyaline casts|Hyaline casts
C1315694|T201|DN|33223-9|LNC2HPO|Hyaline casts|Hyaline casts
C1717156|T201|LN|46135-0|LNC2HPO|Hyaline casts|Hyaline casts
C1717156|T201|DN|46135-0|LNC2HPO|Hyaline casts|Hyaline casts
C1717156|T201|MTH_LN|46135-0|LNC2HPO|Hyaline casts|Hyaline casts
C1717156|T201|LC|46135-0|LNC2HPO|Hyaline casts|Hyaline casts
C1717156|T201|OSN|46135-0|LNC2HPO|Hyaline casts|Hyaline casts
C1979500|T201|LN|51484-4|LNC2HPO|Hyaline casts|Hyaline casts
C1979500|T201|DN|51484-4|LNC2HPO|Hyaline casts|Hyaline casts
C1979500|T201|MTH_LN|51484-4|LNC2HPO|Hyaline casts|Hyaline casts
C1979500|T201|OSN|51484-4|LNC2HPO|Hyaline casts|Hyaline casts
C1979500|T201|LC|51484-4|LNC2HPO|Hyaline casts|Hyaline casts
C0364417|T201|LN|2282-2|LNC2HPO|Folate deficiency|Folate deficiency
C0364417|T201|MTH_LN|2282-2|LNC2HPO|Folate deficiency|Folate deficiency
C0364417|T201|DN|2282-2|LNC2HPO|Folate deficiency|Folate deficiency
C0364417|T201|OSN|2282-2|LNC2HPO|Folate deficiency|Folate deficiency
C0364417|T201|LC|2282-2|LNC2HPO|Folate deficiency|Folate deficiency
C0364417|T201|LN|2282-2|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0364417|T201|MTH_LN|2282-2|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0364417|T201|DN|2282-2|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0364417|T201|OSN|2282-2|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0364417|T201|LC|2282-2|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0364419|T201|LC|2284-8|LNC2HPO|Folate deficiency|Folate deficiency
C0364419|T201|DN|2284-8|LNC2HPO|Folate deficiency|Folate deficiency
C0364419|T201|OSN|2284-8|LNC2HPO|Folate deficiency|Folate deficiency
C0364419|T201|LN|2284-8|LNC2HPO|Folate deficiency|Folate deficiency
C0364419|T201|MTH_LN|2284-8|LNC2HPO|Folate deficiency|Folate deficiency
C0364419|T201|LC|2284-8|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0364419|T201|DN|2284-8|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0364419|T201|OSN|2284-8|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0364419|T201|LN|2284-8|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0364419|T201|MTH_LN|2284-8|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0941562|T201|LN|25415-1|LNC2HPO|Folate deficiency|Folate deficiency
C0941562|T201|DN|25415-1|LNC2HPO|Folate deficiency|Folate deficiency
C0941562|T201|MTH_LN|25415-1|LNC2HPO|Folate deficiency|Folate deficiency
C0941562|T201|OSN|25415-1|LNC2HPO|Folate deficiency|Folate deficiency
C0941562|T201|LC|25415-1|LNC2HPO|Folate deficiency|Folate deficiency
C0941562|T201|LN|25415-1|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0941562|T201|DN|25415-1|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0941562|T201|MTH_LN|25415-1|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0941562|T201|OSN|25415-1|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0941562|T201|LC|25415-1|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C1544620|T201|LN|40665-2|LNC2HPO|Reticulocytosis|Reticulocytosis
C1544620|T201|LC|40665-2|LNC2HPO|Reticulocytosis|Reticulocytosis
C1544620|T201|MTH_LN|40665-2|LNC2HPO|Reticulocytosis|Reticulocytosis
C1544620|T201|DN|40665-2|LNC2HPO|Reticulocytosis|Reticulocytosis
C1544620|T201|OSN|40665-2|LNC2HPO|Reticulocytosis|Reticulocytosis
C1544620|T201|LN|40665-2|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C1544620|T201|LC|40665-2|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C1544620|T201|MTH_LN|40665-2|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C1544620|T201|DN|40665-2|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C1544620|T201|OSN|40665-2|LNC2HPO|Reticulocytopenia|Reticulocytopenia
C0941357|T201|LN|25162-9|LNC2HPO|Hyaline casts|Hyaline casts
C0941357|T201|MTH_LN|25162-9|LNC2HPO|Hyaline casts|Hyaline casts
C0941357|T201|DN|25162-9|LNC2HPO|Hyaline casts|Hyaline casts
C0941357|T201|OSN|25162-9|LNC2HPO|Hyaline casts|Hyaline casts
C0941357|T201|LC|25162-9|LNC2HPO|Hyaline casts|Hyaline casts
C1717334|T201|LN|44382-0|LNC2HPO|Hyaline casts|Hyaline casts
C1717334|T201|MTH_LN|44382-0|LNC2HPO|Hyaline casts|Hyaline casts
C1717334|T201|DN|44382-0|LNC2HPO|Hyaline casts|Hyaline casts
C1717334|T201|OSN|44382-0|LNC2HPO|Hyaline casts|Hyaline casts
C1717334|T201|LC|44382-0|LNC2HPO|Hyaline casts|Hyaline casts
C1978066|T201|LN|50231-0|LNC2HPO|Hyaline casts|Hyaline casts
C1978066|T201|MTH_LN|50231-0|LNC2HPO|Hyaline casts|Hyaline casts
C1978066|T201|DN|50231-0|LNC2HPO|Hyaline casts|Hyaline casts
C1978066|T201|OSN|50231-0|LNC2HPO|Hyaline casts|Hyaline casts
C1978066|T201|LC|50231-0|LNC2HPO|Hyaline casts|Hyaline casts
C1978482|T201|LN|50555-2|LNC2HPO|Glycosuria|Glycosuria
C1978482|T201|MTH_LN|50555-2|LNC2HPO|Glycosuria|Glycosuria
C1978482|T201|DN|50555-2|LNC2HPO|Glycosuria|Glycosuria
C1978482|T201|OSN|50555-2|LNC2HPO|Glycosuria|Glycosuria
C1978482|T201|LC|50555-2|LNC2HPO|Glycosuria|Glycosuria
C1978482|T201|LN|50555-2|LNC2HPO|Glucosuria|Glucosuria
C1978482|T201|MTH_LN|50555-2|LNC2HPO|Glucosuria|Glucosuria
C1978482|T201|DN|50555-2|LNC2HPO|Glucosuria|Glucosuria
C1978482|T201|OSN|50555-2|LNC2HPO|Glucosuria|Glucosuria
C1978482|T201|LC|50555-2|LNC2HPO|Glucosuria|Glucosuria
C0482705|T201|MTH_LN|3255-7|LNC2HPO|Hyperfibrinogenemia|Hyperfibrinogenemia
C0482705|T201|LN|3255-7|LNC2HPO|Hyperfibrinogenemia|Hyperfibrinogenemia
C0482705|T201|DN|3255-7|LNC2HPO|Hyperfibrinogenemia|Hyperfibrinogenemia
C0482705|T201|OSN|3255-7|LNC2HPO|Hyperfibrinogenemia|Hyperfibrinogenemia
C0482705|T201|LC|3255-7|LNC2HPO|Hyperfibrinogenemia|Hyperfibrinogenemia
C0482705|T201|MTH_LN|3255-7|LNC2HPO|Hypofibrinogenemia|Hypofibrinogenemia
C0482705|T201|LN|3255-7|LNC2HPO|Hypofibrinogenemia|Hypofibrinogenemia
C0482705|T201|DN|3255-7|LNC2HPO|Hypofibrinogenemia|Hypofibrinogenemia
C0482705|T201|OSN|3255-7|LNC2HPO|Hypofibrinogenemia|Hypofibrinogenemia
C0482705|T201|LC|3255-7|LNC2HPO|Hypofibrinogenemia|Hypofibrinogenemia
C2736165|T201|LN|57751-0|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C2736165|T201|MTH_LN|57751-0|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C2736165|T201|DN|57751-0|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C2736165|T201|OSN|57751-0|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C2736165|T201|LC|57751-0|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0362931|T201|LN|726-0|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0362931|T201|MTH_LN|726-0|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0362931|T201|DN|726-0|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0362931|T201|OSN|726-0|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0362931|T201|LC|726-0|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0366869|T201|LN|4636-7|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0366869|T201|MTH_LN|4636-7|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0366869|T201|DN|4636-7|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0366869|T201|OSN|4636-7|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0366869|T201|LC|4636-7|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C1954901|T201|LN|49137-3|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C1954901|T201|DN|49137-3|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C1954901|T201|MTH_LN|49137-3|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C1954901|T201|OSN|49137-3|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C1954901|T201|LC|49137-3|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C1978486|T201|LN|50559-4|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C1978486|T201|DN|50559-4|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C1978486|T201|OSN|50559-4|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C1978486|T201|MTH_LN|50559-4|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C1978486|T201|LC|50559-4|LNC2HPO|Hemoglobinuria|Hemoglobinuria
C0482602|T201|LN|2842-3|LNC2HPO|Hyperprolactinemia|Hyperprolactinemia
C0482602|T201|DN|2842-3|LNC2HPO|Hyperprolactinemia|Hyperprolactinemia
C0482602|T201|MTH_LN|2842-3|LNC2HPO|Hyperprolactinemia|Hyperprolactinemia
C0482602|T201|OSN|2842-3|LNC2HPO|Hyperprolactinemia|Hyperprolactinemia
C0482602|T201|LC|2842-3|LNC2HPO|Hyperprolactinemia|Hyperprolactinemia
C0482602|T201|LN|2842-3|LNC2HPO|Hyperprolactinaemia|Hyperprolactinaemia
C0482602|T201|DN|2842-3|LNC2HPO|Hyperprolactinaemia|Hyperprolactinaemia
C0482602|T201|MTH_LN|2842-3|LNC2HPO|Hyperprolactinaemia|Hyperprolactinaemia
C0482602|T201|OSN|2842-3|LNC2HPO|Hyperprolactinaemia|Hyperprolactinaemia
C0482602|T201|LC|2842-3|LNC2HPO|Hyperprolactinaemia|Hyperprolactinaemia
C0482602|T201|LN|2842-3|LNC2HPO|Prolactin excess|Prolactin excess
C0482602|T201|DN|2842-3|LNC2HPO|Prolactin excess|Prolactin excess
C0482602|T201|MTH_LN|2842-3|LNC2HPO|Prolactin excess|Prolactin excess
C0482602|T201|OSN|2842-3|LNC2HPO|Prolactin excess|Prolactin excess
C0482602|T201|LC|2842-3|LNC2HPO|Prolactin excess|Prolactin excess
C0482602|T201|LN|2842-3|LNC2HPO|Prolactin deficiency|Prolactin deficiency
C0482602|T201|DN|2842-3|LNC2HPO|Prolactin deficiency|Prolactin deficiency
C0482602|T201|MTH_LN|2842-3|LNC2HPO|Prolactin deficiency|Prolactin deficiency
C0482602|T201|OSN|2842-3|LNC2HPO|Prolactin deficiency|Prolactin deficiency
C0482602|T201|LC|2842-3|LNC2HPO|Prolactin deficiency|Prolactin deficiency
C0364111|T201|LN|1978-6|LNC2HPO|Bilirubinuria|Bilirubinuria
C0364111|T201|LC|1978-6|LNC2HPO|Bilirubinuria|Bilirubinuria
C0364111|T201|MTH_LN|1978-6|LNC2HPO|Bilirubinuria|Bilirubinuria
C0364111|T201|DN|1978-6|LNC2HPO|Bilirubinuria|Bilirubinuria
C0364111|T201|OSN|1978-6|LNC2HPO|Bilirubinuria|Bilirubinuria
C0803316|T201|LN|20505-4|LNC2HPO|Bilirubinuria|Bilirubinuria
C0803316|T201|LC|20505-4|LNC2HPO|Bilirubinuria|Bilirubinuria
C0803316|T201|MTH_LN|20505-4|LNC2HPO|Bilirubinuria|Bilirubinuria
C0803316|T201|DN|20505-4|LNC2HPO|Bilirubinuria|Bilirubinuria
C0803316|T201|OSN|20505-4|LNC2HPO|Bilirubinuria|Bilirubinuria
C0941345|T201|LN|25146-2|LNC2HPO|Bilirubinuria|Bilirubinuria
C0941345|T201|DN|25146-2|LNC2HPO|Bilirubinuria|Bilirubinuria
C0941345|T201|MTH_LN|25146-2|LNC2HPO|Bilirubinuria|Bilirubinuria
C0941345|T201|OSN|25146-2|LNC2HPO|Bilirubinuria|Bilirubinuria
C0941345|T201|LC|25146-2|LNC2HPO|Bilirubinuria|Bilirubinuria
C1526443|T201|LN|38442-0|LNC2HPO|Bilirubinuria|Bilirubinuria
C1526443|T201|DN|38442-0|LNC2HPO|Bilirubinuria|Bilirubinuria
C1526443|T201|MTH_LN|38442-0|LNC2HPO|Bilirubinuria|Bilirubinuria
C1526443|T201|LC|38442-0|LNC2HPO|Bilirubinuria|Bilirubinuria
C1526443|T201|OSN|38442-0|LNC2HPO|Bilirubinuria|Bilirubinuria
C1544963|T201|LN|41016-7|LNC2HPO|Bilirubinuria|Bilirubinuria
C1544963|T201|LC|41016-7|LNC2HPO|Bilirubinuria|Bilirubinuria
C1544963|T201|DN|41016-7|LNC2HPO|Bilirubinuria|Bilirubinuria
C1544963|T201|OSN|41016-7|LNC2HPO|Bilirubinuria|Bilirubinuria
C1544963|T201|MTH_LN|41016-7|LNC2HPO|Bilirubinuria|Bilirubinuria
C2361847|T201|LN|53327-3|LNC2HPO|Bilirubinuria|Bilirubinuria
C2361847|T201|LC|53327-3|LNC2HPO|Bilirubinuria|Bilirubinuria
C2361847|T201|DN|53327-3|LNC2HPO|Bilirubinuria|Bilirubinuria
C2361847|T201|OSN|53327-3|LNC2HPO|Bilirubinuria|Bilirubinuria
C2361847|T201|MTH_LN|53327-3|LNC2HPO|Bilirubinuria|Bilirubinuria
C3262266|T201|LN|68367-2|LNC2HPO|Bilirubinuria|Bilirubinuria
C3262266|T201|OSN|68367-2|LNC2HPO|Bilirubinuria|Bilirubinuria
C3262266|T201|LC|68367-2|LNC2HPO|Bilirubinuria|Bilirubinuria
C3262266|T201|MTH_LN|68367-2|LNC2HPO|Bilirubinuria|Bilirubinuria
C3262266|T201|DN|68367-2|LNC2HPO|Bilirubinuria|Bilirubinuria
C3481649|T201|LN|70199-5|LNC2HPO|Bilirubinuria|Bilirubinuria
C3481649|T201|OSN|70199-5|LNC2HPO|Bilirubinuria|Bilirubinuria
C3481649|T201|MTH_LN|70199-5|LNC2HPO|Bilirubinuria|Bilirubinuria
C3481649|T201|LC|70199-5|LNC2HPO|Bilirubinuria|Bilirubinuria
C3481649|T201|DN|70199-5|LNC2HPO|Bilirubinuria|Bilirubinuria
C2925975|T201|LN|58450-8|LNC2HPO|Bilirubinuria|Bilirubinuria
C2925975|T201|MTH_LN|58450-8|LNC2HPO|Bilirubinuria|Bilirubinuria
C2925975|T201|DN|58450-8|LNC2HPO|Bilirubinuria|Bilirubinuria
C2925975|T201|LC|58450-8|LNC2HPO|Bilirubinuria|Bilirubinuria
C2925975|T201|OSN|58450-8|LNC2HPO|Bilirubinuria|Bilirubinuria
C0367986|T201|LN|5771-1|LNC2HPO|Bilirubinuria|Bilirubinuria
C0367986|T201|MTH_LN|5771-1|LNC2HPO|Bilirubinuria|Bilirubinuria
C0367986|T201|DN|5771-1|LNC2HPO|Bilirubinuria|Bilirubinuria
C0367986|T201|OSN|5771-1|LNC2HPO|Bilirubinuria|Bilirubinuria
C0367986|T201|LC|5771-1|LNC2HPO|Bilirubinuria|Bilirubinuria
C1715351|T201|LN|44075-0|LNC2HPO|Bilirubinuria|Bilirubinuria
C1715351|T201|MTH_LN|44075-0|LNC2HPO|Bilirubinuria|Bilirubinuria
C1715351|T201|DN|44075-0|LNC2HPO|Bilirubinuria|Bilirubinuria
C1715351|T201|OSN|44075-0|LNC2HPO|Bilirubinuria|Bilirubinuria
C1715351|T201|LC|44075-0|LNC2HPO|Bilirubinuria|Bilirubinuria
C1315707|T201|LN|33236-1|LNC2HPO|Bilirubinuria|Bilirubinuria
C1315707|T201|MTH_LN|33236-1|LNC2HPO|Bilirubinuria|Bilirubinuria
C1315707|T201|DN|33236-1|LNC2HPO|Bilirubinuria|Bilirubinuria
C1315707|T201|OSN|33236-1|LNC2HPO|Bilirubinuria|Bilirubinuria
C1315707|T201|LC|33236-1|LNC2HPO|Bilirubinuria|Bilirubinuria
C0550041|T201|LN|10833-2|LNC2HPO|Hyperinsulinemia|Hyperinsulinemia
C0550041|T201|DN|10833-2|LNC2HPO|Hyperinsulinemia|Hyperinsulinemia
C0550041|T201|MTH_LN|10833-2|LNC2HPO|Hyperinsulinemia|Hyperinsulinemia
C0550041|T201|OSN|10833-2|LNC2HPO|Hyperinsulinemia|Hyperinsulinemia
C0550041|T201|LC|10833-2|LNC2HPO|Hyperinsulinemia|Hyperinsulinemia
C0550041|T201|LN|10833-2|LNC2HPO|Hypoinsulinemia|Hypoinsulinemia
C0550041|T201|DN|10833-2|LNC2HPO|Hypoinsulinemia|Hypoinsulinemia
C0550041|T201|MTH_LN|10833-2|LNC2HPO|Hypoinsulinemia|Hypoinsulinemia
C0550041|T201|OSN|10833-2|LNC2HPO|Hypoinsulinemia|Hypoinsulinemia
C0550041|T201|LC|10833-2|LNC2HPO|Hypoinsulinemia|Hypoinsulinemia
C0945357|T201|LN|26464-8|LNC2HPO|Leukocytosis|Leukocytosis
C0945357|T201|DN|26464-8|LNC2HPO|Leukocytosis|Leukocytosis
C0945357|T201|OSN|26464-8|LNC2HPO|Leukocytosis|Leukocytosis
C0945357|T201|MTH_LN|26464-8|LNC2HPO|Leukocytosis|Leukocytosis
C0945357|T201|LC|26464-8|LNC2HPO|Leukocytosis|Leukocytosis
C0945357|T201|LN|26464-8|LNC2HPO|Leukopenia|Leukopenia
C0945357|T201|DN|26464-8|LNC2HPO|Leukopenia|Leukopenia
C0945357|T201|OSN|26464-8|LNC2HPO|Leukopenia|Leukopenia
C0945357|T201|MTH_LN|26464-8|LNC2HPO|Leukopenia|Leukopenia
C0945357|T201|LC|26464-8|LNC2HPO|Leukopenia|Leukopenia
C0942947|T201|LN|27088-4|LNC2HPO|Folate deficiency|Folate deficiency
C0942947|T201|MTH_LN|27088-4|LNC2HPO|Folate deficiency|Folate deficiency
C0942947|T201|OSN|27088-4|LNC2HPO|Folate deficiency|Folate deficiency
C0942947|T201|DN|27088-4|LNC2HPO|Folate deficiency|Folate deficiency
C0942947|T201|LC|27088-4|LNC2HPO|Folate deficiency|Folate deficiency
C0942947|T201|LN|27088-4|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0942947|T201|MTH_LN|27088-4|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0942947|T201|OSN|27088-4|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0942947|T201|DN|27088-4|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0942947|T201|LC|27088-4|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0363850|T201|LN|1716-0|LNC2HPO|Aciduria|Aciduria
C0363850|T201|MTH_LN|1716-0|LNC2HPO|Aciduria|Aciduria
C0363850|T201|DN|1716-0|LNC2HPO|Aciduria|Aciduria
C0363850|T201|OSN|1716-0|LNC2HPO|Aciduria|Aciduria
C0363850|T201|LC|1716-0|LNC2HPO|Aciduria|Aciduria
C2734583|T201|LN|56489-8|LNC2HPO|Aciduria|Aciduria
C2734583|T201|OSN|56489-8|LNC2HPO|Aciduria|Aciduria
C2734583|T201|MTH_LN|56489-8|LNC2HPO|Aciduria|Aciduria
C2734583|T201|LC|56489-8|LNC2HPO|Aciduria|Aciduria
C2734583|T201|DN|56489-8|LNC2HPO|Aciduria|Aciduria
C3699474|T201|LN|74092-8|LNC2HPO|Aciduria|Aciduria
C3699474|T201|OSN|74092-8|LNC2HPO|Aciduria|Aciduria
C3699474|T201|MTH_LN|74092-8|LNC2HPO|Aciduria|Aciduria
C3699474|T201|LC|74092-8|LNC2HPO|Aciduria|Aciduria
C3699474|T201|DN|74092-8|LNC2HPO|Aciduria|Aciduria
C0549979|T201|LN|10966-0|LNC2HPO|Glycosuria|Glycosuria
C0549979|T201|MTH_LN|10966-0|LNC2HPO|Glycosuria|Glycosuria
C0549979|T201|DN|10966-0|LNC2HPO|Glycosuria|Glycosuria
C0549979|T201|OSN|10966-0|LNC2HPO|Glycosuria|Glycosuria
C0549979|T201|LC|10966-0|LNC2HPO|Glycosuria|Glycosuria
C0549979|T201|LN|10966-0|LNC2HPO|Glucosuria|Glucosuria
C0549979|T201|MTH_LN|10966-0|LNC2HPO|Glucosuria|Glucosuria
C0549979|T201|DN|10966-0|LNC2HPO|Glucosuria|Glucosuria
C0549979|T201|OSN|10966-0|LNC2HPO|Glucosuria|Glucosuria
C0549979|T201|LC|10966-0|LNC2HPO|Glucosuria|Glucosuria
C0549984|T201|LN|10967-8|LNC2HPO|Glycosuria|Glycosuria
C0549984|T201|MTH_LN|10967-8|LNC2HPO|Glycosuria|Glycosuria
C0549984|T201|DN|10967-8|LNC2HPO|Glycosuria|Glycosuria
C0549984|T201|OSN|10967-8|LNC2HPO|Glycosuria|Glycosuria
C0549984|T201|LC|10967-8|LNC2HPO|Glycosuria|Glycosuria
C0549984|T201|LN|10967-8|LNC2HPO|Glucosuria|Glucosuria
C0549984|T201|MTH_LN|10967-8|LNC2HPO|Glucosuria|Glucosuria
C0549984|T201|DN|10967-8|LNC2HPO|Glucosuria|Glucosuria
C0549984|T201|OSN|10967-8|LNC2HPO|Glucosuria|Glucosuria
C0549984|T201|LC|10967-8|LNC2HPO|Glucosuria|Glucosuria
C0549987|T201|LN|10968-6|LNC2HPO|Glycosuria|Glycosuria
C0549987|T201|MTH_LN|10968-6|LNC2HPO|Glycosuria|Glycosuria
C0549987|T201|DN|10968-6|LNC2HPO|Glycosuria|Glycosuria
C0549987|T201|OSN|10968-6|LNC2HPO|Glycosuria|Glycosuria
C0549987|T201|LC|10968-6|LNC2HPO|Glycosuria|Glycosuria
C0549987|T201|LN|10968-6|LNC2HPO|Glucosuria|Glucosuria
C0549987|T201|MTH_LN|10968-6|LNC2HPO|Glucosuria|Glucosuria
C0549987|T201|DN|10968-6|LNC2HPO|Glucosuria|Glucosuria
C0549987|T201|OSN|10968-6|LNC2HPO|Glucosuria|Glucosuria
C0549987|T201|LC|10968-6|LNC2HPO|Glucosuria|Glucosuria
C0550433|T201|LN|12239-0|LNC2HPO|Oligosacchariduria|Oligosacchariduria
C0550433|T201|MTH_LN|12239-0|LNC2HPO|Oligosacchariduria|Oligosacchariduria
C0550433|T201|DN|12239-0|LNC2HPO|Oligosacchariduria|Oligosacchariduria
C0550433|T201|OSN|12239-0|LNC2HPO|Oligosacchariduria|Oligosacchariduria
C0550433|T201|LC|12239-0|LNC2HPO|Oligosacchariduria|Oligosacchariduria
C0364661|T201|LN|2520-5|LNC2HPO|Hyperlactatorachia|Hyperlactatorachia
C0364661|T201|MTH_LN|2520-5|LNC2HPO|Hyperlactatorachia|Hyperlactatorachia
C0364661|T201|DN|2520-5|LNC2HPO|Hyperlactatorachia|Hyperlactatorachia
C0364661|T201|OSN|2520-5|LNC2HPO|Hyperlactatorachia|Hyperlactatorachia
C0364661|T201|LC|2520-5|LNC2HPO|Hyperlactatorachia|Hyperlactatorachia
C0364661|T201|LN|2520-5|LNC2HPO|Hypolactatorachia|Hypolactatorachia
C0364661|T201|MTH_LN|2520-5|LNC2HPO|Hypolactatorachia|Hypolactatorachia
C0364661|T201|DN|2520-5|LNC2HPO|Hypolactatorachia|Hypolactatorachia
C0364661|T201|OSN|2520-5|LNC2HPO|Hypolactatorachia|Hypolactatorachia
C0364661|T201|LC|2520-5|LNC2HPO|Hypolactatorachia|Hypolactatorachia
C0943617|T201|LN|27941-4|LNC2HPO|Hyperlactatorachia|Hyperlactatorachia
C0943617|T201|DN|27941-4|LNC2HPO|Hyperlactatorachia|Hyperlactatorachia
C0943617|T201|MTH_LN|27941-4|LNC2HPO|Hyperlactatorachia|Hyperlactatorachia
C0943617|T201|OSN|27941-4|LNC2HPO|Hyperlactatorachia|Hyperlactatorachia
C0943617|T201|LC|27941-4|LNC2HPO|Hyperlactatorachia|Hyperlactatorachia
C0943617|T201|LN|27941-4|LNC2HPO|Hypolactatorachia|Hypolactatorachia
C0943617|T201|DN|27941-4|LNC2HPO|Hypolactatorachia|Hypolactatorachia
C0943617|T201|MTH_LN|27941-4|LNC2HPO|Hypolactatorachia|Hypolactatorachia
C0943617|T201|OSN|27941-4|LNC2HPO|Hypolactatorachia|Hypolactatorachia
C0943617|T201|LC|27941-4|LNC2HPO|Hypolactatorachia|Hypolactatorachia
C2706875|T201|LN|54309-0|LNC2HPO|Hyperlactatorachia|Hyperlactatorachia
C2706875|T201|DN|54309-0|LNC2HPO|Hyperlactatorachia|Hyperlactatorachia
C2706875|T201|OSN|54309-0|LNC2HPO|Hyperlactatorachia|Hyperlactatorachia
C2706875|T201|LC|54309-0|LNC2HPO|Hyperlactatorachia|Hyperlactatorachia
C2706875|T201|MTH_LN|54309-0|LNC2HPO|Hyperlactatorachia|Hyperlactatorachia
C2706875|T201|LN|54309-0|LNC2HPO|Hypolactatorachia|Hypolactatorachia
C2706875|T201|DN|54309-0|LNC2HPO|Hypolactatorachia|Hypolactatorachia
C2706875|T201|OSN|54309-0|LNC2HPO|Hypolactatorachia|Hypolactatorachia
C2706875|T201|LC|54309-0|LNC2HPO|Hypolactatorachia|Hypolactatorachia
C2706875|T201|MTH_LN|54309-0|LNC2HPO|Hypolactatorachia|Hypolactatorachia
C3846945|T201|LN|75040-6|LNC2HPO|Hyperlactatorachia|Hyperlactatorachia
C3846945|T201|LC|75040-6|LNC2HPO|Hyperlactatorachia|Hyperlactatorachia
C3846945|T201|OSN|75040-6|LNC2HPO|Hyperlactatorachia|Hyperlactatorachia
C3846945|T201|MTH_LN|75040-6|LNC2HPO|Hyperlactatorachia|Hyperlactatorachia
C3846945|T201|DN|75040-6|LNC2HPO|Hyperlactatorachia|Hyperlactatorachia
C3846945|T201|LN|75040-6|LNC2HPO|Hypolactatorachia|Hypolactatorachia
C3846945|T201|LC|75040-6|LNC2HPO|Hypolactatorachia|Hypolactatorachia
C3846945|T201|OSN|75040-6|LNC2HPO|Hypolactatorachia|Hypolactatorachia
C3846945|T201|MTH_LN|75040-6|LNC2HPO|Hypolactatorachia|Hypolactatorachia
C3846945|T201|DN|75040-6|LNC2HPO|Hypolactatorachia|Hypolactatorachia
C0796899|T201|LN|13708-3|LNC2HPO|Argininuria|Argininuria
C0796899|T201|MTH_LN|13708-3|LNC2HPO|Argininuria|Argininuria
C0796899|T201|OSN|13708-3|LNC2HPO|Argininuria|Argininuria
C0796899|T201|DN|13708-3|LNC2HPO|Argininuria|Argininuria
C0796899|T201|LC|13708-3|LNC2HPO|Argininuria|Argininuria
C0364029|T201|LN|1894-5|LNC2HPO|Argininuria|Argininuria
C0364029|T201|MTH_LN|1894-5|LNC2HPO|Argininuria|Argininuria
C0364029|T201|DN|1894-5|LNC2HPO|Argininuria|Argininuria
C0364029|T201|OSN|1894-5|LNC2HPO|Argininuria|Argininuria
C0364029|T201|LC|1894-5|LNC2HPO|Argininuria|Argininuria
C0364030|T201|LN|1895-2|LNC2HPO|Argininuria|Argininuria
C0364030|T201|MTH_LN|1895-2|LNC2HPO|Argininuria|Argininuria
C0364030|T201|DN|1895-2|LNC2HPO|Argininuria|Argininuria
C0364030|T201|OSN|1895-2|LNC2HPO|Argininuria|Argininuria
C0364030|T201|LC|1895-2|LNC2HPO|Argininuria|Argininuria
C0882311|T201|LN|22697-7|LNC2HPO|Argininuria|Argininuria
C0882311|T201|DN|22697-7|LNC2HPO|Argininuria|Argininuria
C0882311|T201|OSN|22697-7|LNC2HPO|Argininuria|Argininuria
C0882311|T201|LC|22697-7|LNC2HPO|Argininuria|Argininuria
C0882311|T201|MTH_LN|22697-7|LNC2HPO|Argininuria|Argininuria
C0941489|T201|LN|25322-9|LNC2HPO|Argininuria|Argininuria
C0941489|T201|DN|25322-9|LNC2HPO|Argininuria|Argininuria
C0941489|T201|MTH_LN|25322-9|LNC2HPO|Argininuria|Argininuria
C0941489|T201|OSN|25322-9|LNC2HPO|Argininuria|Argininuria
C0941489|T201|LC|25322-9|LNC2HPO|Argininuria|Argininuria
C0941920|T201|LN|25860-8|LNC2HPO|Argininuria|Argininuria
C0941920|T201|DN|25860-8|LNC2HPO|Argininuria|Argininuria
C0941920|T201|MTH_LN|25860-8|LNC2HPO|Argininuria|Argininuria
C0941920|T201|OSN|25860-8|LNC2HPO|Argininuria|Argininuria
C0941920|T201|LC|25860-8|LNC2HPO|Argininuria|Argininuria
C0941921|T201|LN|25861-6|LNC2HPO|Argininuria|Argininuria
C0941921|T201|DN|25861-6|LNC2HPO|Argininuria|Argininuria
C0941921|T201|OSN|25861-6|LNC2HPO|Argininuria|Argininuria
C0941921|T201|LC|25861-6|LNC2HPO|Argininuria|Argininuria
C0941921|T201|MTH_LN|25861-6|LNC2HPO|Argininuria|Argininuria
C0943117|T201|LN|27296-3|LNC2HPO|Argininuria|Argininuria
C0943117|T201|DN|27296-3|LNC2HPO|Argininuria|Argininuria
C0943117|T201|MTH_LN|27296-3|LNC2HPO|Argininuria|Argininuria
C0943117|T201|OSN|27296-3|LNC2HPO|Argininuria|Argininuria
C0943117|T201|LC|27296-3|LNC2HPO|Argininuria|Argininuria
C1113962|T201|LN|30062-4|LNC2HPO|Argininuria|Argininuria
C1113962|T201|DN|30062-4|LNC2HPO|Argininuria|Argininuria
C1113962|T201|MTH_LN|30062-4|LNC2HPO|Argininuria|Argininuria
C1113962|T201|OSN|30062-4|LNC2HPO|Argininuria|Argininuria
C1113962|T201|LC|30062-4|LNC2HPO|Argininuria|Argininuria
C1715553|T201|LN|44299-6|LNC2HPO|Argininuria|Argininuria
C1715553|T201|MTH_LN|44299-6|LNC2HPO|Argininuria|Argininuria
C1715553|T201|OSN|44299-6|LNC2HPO|Argininuria|Argininuria
C1715553|T201|DN|44299-6|LNC2HPO|Argininuria|Argininuria
C1715553|T201|LC|44299-6|LNC2HPO|Argininuria|Argininuria
C2734826|T201|LN|56672-9|LNC2HPO|Argininuria|Argininuria
C2734826|T201|MTH_LN|56672-9|LNC2HPO|Argininuria|Argininuria
C2734826|T201|DN|56672-9|LNC2HPO|Argininuria|Argininuria
C2734826|T201|LC|56672-9|LNC2HPO|Argininuria|Argininuria
C2734826|T201|OSN|56672-9|LNC2HPO|Argininuria|Argininuria
C0799554|T201|LN|16401-2|LNC2HPO|Argininuria|Argininuria
C0799554|T201|MTH_LN|16401-2|LNC2HPO|Argininuria|Argininuria
C0799554|T201|DN|16401-2|LNC2HPO|Argininuria|Argininuria
C0799554|T201|OSN|16401-2|LNC2HPO|Argininuria|Argininuria
C0799554|T201|LC|16401-2|LNC2HPO|Argininuria|Argininuria
C2607831|T201|DN|35210-4|LNC2HPO|Folate deficiency|Folate deficiency
C2607831|T201|OSN|35210-4|LNC2HPO|Folate deficiency|Folate deficiency
C2607831|T201|LN|35210-4|LNC2HPO|Folate deficiency|Folate deficiency
C2607831|T201|MTH_LN|35210-4|LNC2HPO|Folate deficiency|Folate deficiency
C2607831|T201|LC|35210-4|LNC2HPO|Folate deficiency|Folate deficiency
C2607831|T201|DN|35210-4|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C2607831|T201|OSN|35210-4|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C2607831|T201|LN|35210-4|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C2607831|T201|MTH_LN|35210-4|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C2607831|T201|LC|35210-4|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0486101|T201|LN|10364-8|LNC2HPO|Hair xenobiotic|Hair xenobiotic
C0486101|T201|MTH_LN|10364-8|LNC2HPO|Hair xenobiotic|Hair xenobiotic
C0486101|T201|OSN|10364-8|LNC2HPO|Hair xenobiotic|Hair xenobiotic
C0486101|T201|LC|10364-8|LNC2HPO|Hair xenobiotic|Hair xenobiotic
C0486101|T201|DN|10364-8|LNC2HPO|Hair xenobiotic|Hair xenobiotic
C1544330|T201|LN|40355-0|LNC2HPO|Hair xenobiotic|Hair xenobiotic
C1544330|T201|MTH_LN|40355-0|LNC2HPO|Hair xenobiotic|Hair xenobiotic
C1544330|T201|OSN|40355-0|LNC2HPO|Hair xenobiotic|Hair xenobiotic
C1544330|T201|DN|40355-0|LNC2HPO|Hair xenobiotic|Hair xenobiotic
C1544330|T201|LC|40355-0|LNC2HPO|Hair xenobiotic|Hair xenobiotic
C1544393|T201|LN|40418-6|LNC2HPO|Meconium xenobiotic|Meconium xenobiotic
C1544393|T201|MTH_LN|40418-6|LNC2HPO|Meconium xenobiotic|Meconium xenobiotic
C1544393|T201|OSN|40418-6|LNC2HPO|Meconium xenobiotic|Meconium xenobiotic
C1544393|T201|DN|40418-6|LNC2HPO|Meconium xenobiotic|Meconium xenobiotic
C1544393|T201|LC|40418-6|LNC2HPO|Meconium xenobiotic|Meconium xenobiotic
C2969826|T201|LN|59892-0|LNC2HPO|Gastric fluid xenobiotic|Gastric fluid xenobiotic
C2969826|T201|DN|59892-0|LNC2HPO|Gastric fluid xenobiotic|Gastric fluid xenobiotic
C2969826|T201|LC|59892-0|LNC2HPO|Gastric fluid xenobiotic|Gastric fluid xenobiotic
C2969826|T201|OSN|59892-0|LNC2HPO|Gastric fluid xenobiotic|Gastric fluid xenobiotic
C2969826|T201|MTH_LN|59892-0|LNC2HPO|Gastric fluid xenobiotic|Gastric fluid xenobiotic
C0947495|T201|MTH_LN|14251-3|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C0947495|T201|DN|14251-3|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C0947495|T201|LN|14251-3|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C0947495|T201|OSN|14251-3|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C0947495|T201|LC|14251-3|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C0942080|T201|LN|26054-7|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C0942080|T201|MTH_LN|26054-7|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C0942080|T201|DN|26054-7|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C0942080|T201|OSN|26054-7|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C0942080|T201|LC|26054-7|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C1977524|T201|LN|49781-8|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C1977524|T201|DN|49781-8|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C1977524|T201|OSN|49781-8|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C1977524|T201|MTH_LN|49781-8|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C1977524|T201|LC|49781-8|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C2360395|T201|LN|51715-1|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C2360395|T201|OSN|51715-1|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C2360395|T201|DN|51715-1|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C2360395|T201|MTH_LN|51715-1|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C2360395|T201|LC|51715-1|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C2360498|T201|LN|51794-6|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C2360498|T201|DN|51794-6|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C2360498|T201|MTH_LN|51794-6|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C2360498|T201|OSN|51794-6|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C2360498|T201|LC|51794-6|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C2734787|T201|LN|56632-3|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C2734787|T201|DN|56632-3|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C2734787|T201|LC|56632-3|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C2734787|T201|MTH_LN|56632-3|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C2734787|T201|OSN|56632-3|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C2734953|T201|LN|56735-4|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C2734953|T201|MTH_LN|56735-4|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C2734953|T201|LC|56735-4|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C2734953|T201|DN|56735-4|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C2734953|T201|OSN|56735-4|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C3172373|T201|LN|63283-6|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C3172373|T201|LC|63283-6|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C3172373|T201|OSN|63283-6|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C3172373|T201|MTH_LN|63283-6|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C3172373|T201|DN|63283-6|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C4298342|T201|LN|82928-3|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C4298342|T201|MTH_LN|82928-3|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C4298342|T201|LC|82928-3|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C4298342|T201|OSN|82928-3|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C4298342|T201|DN|82928-3|LNC2HPO|AMA-M2 positive|AMA-M2 positive
C0368008|T201|LN|5784-4|LNC2HPO|Cystinuria|Cystinuria
C0368008|T201|MTH_LN|5784-4|LNC2HPO|Cystinuria|Cystinuria
C0368008|T201|DN|5784-4|LNC2HPO|Cystinuria|Cystinuria
C0368008|T201|OSN|5784-4|LNC2HPO|Cystinuria|Cystinuria
C0368008|T201|LC|5784-4|LNC2HPO|Cystinuria|Cystinuria
C0368008|T201|LN|5784-4|LNC2HPO|Aminoaciduria|Aminoaciduria
C0368008|T201|MTH_LN|5784-4|LNC2HPO|Aminoaciduria|Aminoaciduria
C0368008|T201|DN|5784-4|LNC2HPO|Aminoaciduria|Aminoaciduria
C0368008|T201|OSN|5784-4|LNC2HPO|Aminoaciduria|Aminoaciduria
C0368008|T201|LC|5784-4|LNC2HPO|Aminoaciduria|Aminoaciduria
C0368008|T201|LN|5784-4|LNC2HPO|Hyperaminoaciduria|Hyperaminoaciduria
C0368008|T201|MTH_LN|5784-4|LNC2HPO|Hyperaminoaciduria|Hyperaminoaciduria
C0368008|T201|DN|5784-4|LNC2HPO|Hyperaminoaciduria|Hyperaminoaciduria
C0368008|T201|OSN|5784-4|LNC2HPO|Hyperaminoaciduria|Hyperaminoaciduria
C0368008|T201|LC|5784-4|LNC2HPO|Hyperaminoaciduria|Hyperaminoaciduria
C0364490|T201|LC|2350-7|LNC2HPO|Glycosuria|Glycosuria
C0364490|T201|MTH_LN|2350-7|LNC2HPO|Glycosuria|Glycosuria
C0364490|T201|DN|2350-7|LNC2HPO|Glycosuria|Glycosuria
C0364490|T201|OSN|2350-7|LNC2HPO|Glycosuria|Glycosuria
C0364490|T201|LN|2350-7|LNC2HPO|Glycosuria|Glycosuria
C0364490|T201|LC|2350-7|LNC2HPO|Glucosuria|Glucosuria
C0364490|T201|MTH_LN|2350-7|LNC2HPO|Glucosuria|Glucosuria
C0364490|T201|DN|2350-7|LNC2HPO|Glucosuria|Glucosuria
C0364490|T201|OSN|2350-7|LNC2HPO|Glucosuria|Glucosuria
C0364490|T201|LN|2350-7|LNC2HPO|Glucosuria|Glucosuria
C0365100|T201|LN|2956-1|LNC2HPO|Hypernatriuria|Hypernatriuria
C0365100|T201|MTH_LN|2956-1|LNC2HPO|Hypernatriuria|Hypernatriuria
C0365100|T201|DN|2956-1|LNC2HPO|Hypernatriuria|Hypernatriuria
C0365100|T201|OSN|2956-1|LNC2HPO|Hypernatriuria|Hypernatriuria
C0365100|T201|LC|2956-1|LNC2HPO|Hypernatriuria|Hypernatriuria
C0365100|T201|LN|2956-1|LNC2HPO|Hyponatriuria|Hyponatriuria
C0365100|T201|MTH_LN|2956-1|LNC2HPO|Hyponatriuria|Hyponatriuria
C0365100|T201|DN|2956-1|LNC2HPO|Hyponatriuria|Hyponatriuria
C0365100|T201|OSN|2956-1|LNC2HPO|Hyponatriuria|Hyponatriuria
C0365100|T201|LC|2956-1|LNC2HPO|Hyponatriuria|Hyponatriuria
C0364972|T201|LN|2829-0|LNC2HPO|Hyperkaliuresis|Hyperkaliuresis
C0364972|T201|MTH_LN|2829-0|LNC2HPO|Hyperkaliuresis|Hyperkaliuresis
C0364972|T201|DN|2829-0|LNC2HPO|Hyperkaliuresis|Hyperkaliuresis
C0364972|T201|OSN|2829-0|LNC2HPO|Hyperkaliuresis|Hyperkaliuresis
C0364972|T201|LC|2829-0|LNC2HPO|Hyperkaliuresis|Hyperkaliuresis
C0364972|T201|LN|2829-0|LNC2HPO|Hypokaluria|Hypokaluria
C0364972|T201|MTH_LN|2829-0|LNC2HPO|Hypokaluria|Hypokaluria
C0364972|T201|DN|2829-0|LNC2HPO|Hypokaluria|Hypokaluria
C0364972|T201|OSN|2829-0|LNC2HPO|Hypokaluria|Hypokaluria
C0364972|T201|LC|2829-0|LNC2HPO|Hypokaluria|Hypokaluria
C0362902|T201|LN|713-8|LNC2HPO|Eosinophilia|Eosinophilia
C0362902|T201|MTH_LN|713-8|LNC2HPO|Eosinophilia|Eosinophilia
C0362902|T201|OSN|713-8|LNC2HPO|Eosinophilia|Eosinophilia
C0362902|T201|DN|713-8|LNC2HPO|Eosinophilia|Eosinophilia
C0362902|T201|LC|713-8|LNC2HPO|Eosinophilia|Eosinophilia
C0362903|T201|LN|714-6|LNC2HPO|Eosinophilia|Eosinophilia
C0362903|T201|MTH_LN|714-6|LNC2HPO|Eosinophilia|Eosinophilia
C0362903|T201|OSN|714-6|LNC2HPO|Eosinophilia|Eosinophilia
C0362903|T201|DN|714-6|LNC2HPO|Eosinophilia|Eosinophilia
C0362903|T201|LC|714-6|LNC2HPO|Eosinophilia|Eosinophilia
C0362895|T201|LN|707-0|LNC2HPO|Basophilia|Basophilia
C0362895|T201|MTH_LN|707-0|LNC2HPO|Basophilia|Basophilia
C0362895|T201|OSN|707-0|LNC2HPO|Basophilia|Basophilia
C0362895|T201|DN|707-0|LNC2HPO|Basophilia|Basophilia
C0362895|T201|LC|707-0|LNC2HPO|Basophilia|Basophilia
C0799763|T201|LN|16616-5|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0799763|T201|OSN|16616-5|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0799763|T201|MTH_LN|16616-5|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0799763|T201|DN|16616-5|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0799763|T201|LC|16616-5|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C0799763|T201|LN|16616-5|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0799763|T201|OSN|16616-5|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0799763|T201|MTH_LN|16616-5|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0799763|T201|DN|16616-5|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C0799763|T201|LC|16616-5|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C1953490|T201|LN|48090-5|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C1953490|T201|DN|48090-5|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C1953490|T201|OSN|48090-5|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C1953490|T201|MTH_LN|48090-5|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C1953490|T201|LC|48090-5|LNC2HPO|Hyperalphalipoproteinemia|Hyperalphalipoproteinemia
C1953490|T201|LN|48090-5|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C1953490|T201|DN|48090-5|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C1953490|T201|OSN|48090-5|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C1953490|T201|MTH_LN|48090-5|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C1953490|T201|LC|48090-5|LNC2HPO|Hypoalphalipoproteinemia|Hypoalphalipoproteinemia
C1714736|T201|LN|43392-0|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1714736|T201|OSN|43392-0|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1714736|T201|LC|43392-0|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1714736|T201|MTH_LN|43392-0|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1714736|T201|DN|43392-0|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1714737|T201|LN|43393-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1714737|T201|LC|43393-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1714737|T201|MTH_LN|43393-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1714737|T201|OSN|43393-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1714737|T201|DN|43393-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1714738|T201|LN|43394-6|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1714738|T201|DN|43394-6|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1714738|T201|OSN|43394-6|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1714738|T201|MTH_LN|43394-6|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1714738|T201|LC|43394-6|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1831079|T201|LN|46984-1|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1831079|T201|LC|46984-1|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1831079|T201|MTH_LN|46984-1|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1831079|T201|OSN|46984-1|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1831079|T201|DN|46984-1|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1831080|T201|LN|46985-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1831080|T201|MTH_LN|46985-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1831080|T201|OSN|46985-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1831080|T201|LC|46985-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1831080|T201|DN|46985-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1954746|T201|LN|49026-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1954746|T201|MTH_LN|49026-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1954746|T201|LC|49026-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1954746|T201|DN|49026-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1954746|T201|OSN|49026-8|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1954748|T201|LN|49027-6|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1954748|T201|MTH_LN|49027-6|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1954748|T201|OSN|49027-6|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1954748|T201|LC|49027-6|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1954748|T201|DN|49027-6|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2361616|T201|LN|53133-5|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2361616|T201|DN|53133-5|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2361616|T201|MTH_LN|53133-5|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2361616|T201|OSN|53133-5|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2361616|T201|LC|53133-5|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2734094|T201|LN|56136-5|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2734094|T201|LC|56136-5|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2734094|T201|OSN|56136-5|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2734094|T201|MTH_LN|56136-5|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2734094|T201|DN|56136-5|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2734095|T201|LN|56137-3|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2734095|T201|OSN|56137-3|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2734095|T201|LC|56137-3|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2734095|T201|MTH_LN|56137-3|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2734095|T201|DN|56137-3|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2734096|T201|LN|56138-1|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2734096|T201|LC|56138-1|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2734096|T201|MTH_LN|56138-1|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2734096|T201|OSN|56138-1|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2734096|T201|DN|56138-1|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2734097|T201|LN|56139-9|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2734097|T201|LC|56139-9|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2734097|T201|MTH_LN|56139-9|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2734097|T201|OSN|56139-9|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2734097|T201|DN|56139-9|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2735471|T201|LN|57938-3|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2735471|T201|LC|57938-3|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2735471|T201|OSN|57938-3|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2735471|T201|MTH_LN|57938-3|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2735471|T201|DN|57938-3|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2736108|T201|LN|57698-3|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2736108|T201|OSN|57698-3|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2736108|T201|DN|57698-3|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2736108|T201|MTH_LN|57698-3|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C2736108|T201|LC|57698-3|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C0799525|T201|LN|16362-6|LNC2HPO|Azotemia|Azotemia
C0799525|T201|MTH_LN|16362-6|LNC2HPO|Azotemia|Azotemia
C0799525|T201|DN|16362-6|LNC2HPO|Azotemia|Azotemia
C0799525|T201|OSN|16362-6|LNC2HPO|Azotemia|Azotemia
C0799525|T201|LC|16362-6|LNC2HPO|Azotemia|Azotemia
C0799525|T201|LN|16362-6|LNC2HPO|Azotaemia|Azotaemia
C0799525|T201|MTH_LN|16362-6|LNC2HPO|Azotaemia|Azotaemia
C0799525|T201|DN|16362-6|LNC2HPO|Azotaemia|Azotaemia
C0799525|T201|OSN|16362-6|LNC2HPO|Azotaemia|Azotaemia
C0799525|T201|LC|16362-6|LNC2HPO|Azotaemia|Azotaemia
C0799525|T201|LN|16362-6|LNC2HPO|Hyperammonemia|Hyperammonemia
C0799525|T201|MTH_LN|16362-6|LNC2HPO|Hyperammonemia|Hyperammonemia
C0799525|T201|DN|16362-6|LNC2HPO|Hyperammonemia|Hyperammonemia
C0799525|T201|OSN|16362-6|LNC2HPO|Hyperammonemia|Hyperammonemia
C0799525|T201|LC|16362-6|LNC2HPO|Hyperammonemia|Hyperammonemia
C0799525|T201|LN|16362-6|LNC2HPO|Hypoammonemia|Hypoammonemia
C0799525|T201|MTH_LN|16362-6|LNC2HPO|Hypoammonemia|Hypoammonemia
C0799525|T201|DN|16362-6|LNC2HPO|Hypoammonemia|Hypoammonemia
C0799525|T201|OSN|16362-6|LNC2HPO|Hypoammonemia|Hypoammonemia
C0799525|T201|LC|16362-6|LNC2HPO|Hypoammonemia|Hypoammonemia
C0363976|T201|LN|1841-6|LNC2HPO|Azotemia|Azotemia
C0363976|T201|MTH_LN|1841-6|LNC2HPO|Azotemia|Azotemia
C0363976|T201|DN|1841-6|LNC2HPO|Azotemia|Azotemia
C0363976|T201|OSN|1841-6|LNC2HPO|Azotemia|Azotemia
C0363976|T201|LC|1841-6|LNC2HPO|Azotemia|Azotemia
C0363976|T201|LN|1841-6|LNC2HPO|Azotaemia|Azotaemia
C0363976|T201|MTH_LN|1841-6|LNC2HPO|Azotaemia|Azotaemia
C0363976|T201|DN|1841-6|LNC2HPO|Azotaemia|Azotaemia
C0363976|T201|OSN|1841-6|LNC2HPO|Azotaemia|Azotaemia
C0363976|T201|LC|1841-6|LNC2HPO|Azotaemia|Azotaemia
C0363976|T201|LN|1841-6|LNC2HPO|Hyperammonemia|Hyperammonemia
C0363976|T201|MTH_LN|1841-6|LNC2HPO|Hyperammonemia|Hyperammonemia
C0363976|T201|DN|1841-6|LNC2HPO|Hyperammonemia|Hyperammonemia
C0363976|T201|OSN|1841-6|LNC2HPO|Hyperammonemia|Hyperammonemia
C0363976|T201|LC|1841-6|LNC2HPO|Hyperammonemia|Hyperammonemia
C0363976|T201|LN|1841-6|LNC2HPO|Hypoammonemia|Hypoammonemia
C0363976|T201|MTH_LN|1841-6|LNC2HPO|Hypoammonemia|Hypoammonemia
C0363976|T201|DN|1841-6|LNC2HPO|Hypoammonemia|Hypoammonemia
C0363976|T201|OSN|1841-6|LNC2HPO|Hypoammonemia|Hypoammonemia
C0363976|T201|LC|1841-6|LNC2HPO|Hypoammonemia|Hypoammonemia
C0803484|T201|LN|20684-7|LNC2HPO|Azotemia|Azotemia
C0803484|T201|MTH_LN|20684-7|LNC2HPO|Azotemia|Azotemia
C0803484|T201|DN|20684-7|LNC2HPO|Azotemia|Azotemia
C0803484|T201|OSN|20684-7|LNC2HPO|Azotemia|Azotemia
C0803484|T201|LC|20684-7|LNC2HPO|Azotemia|Azotemia
C0803484|T201|LN|20684-7|LNC2HPO|Azotaemia|Azotaemia
C0803484|T201|MTH_LN|20684-7|LNC2HPO|Azotaemia|Azotaemia
C0803484|T201|DN|20684-7|LNC2HPO|Azotaemia|Azotaemia
C0803484|T201|OSN|20684-7|LNC2HPO|Azotaemia|Azotaemia
C0803484|T201|LC|20684-7|LNC2HPO|Azotaemia|Azotaemia
C0803484|T201|LN|20684-7|LNC2HPO|Hyperammonemia|Hyperammonemia
C0803484|T201|MTH_LN|20684-7|LNC2HPO|Hyperammonemia|Hyperammonemia
C0803484|T201|DN|20684-7|LNC2HPO|Hyperammonemia|Hyperammonemia
C0803484|T201|OSN|20684-7|LNC2HPO|Hyperammonemia|Hyperammonemia
C0803484|T201|LC|20684-7|LNC2HPO|Hyperammonemia|Hyperammonemia
C0803484|T201|LN|20684-7|LNC2HPO|Hypoammonemia|Hypoammonemia
C0803484|T201|MTH_LN|20684-7|LNC2HPO|Hypoammonemia|Hypoammonemia
C0803484|T201|DN|20684-7|LNC2HPO|Hypoammonemia|Hypoammonemia
C0803484|T201|OSN|20684-7|LNC2HPO|Hypoammonemia|Hypoammonemia
C0803484|T201|LC|20684-7|LNC2HPO|Hypoammonemia|Hypoammonemia
C0880263|T201|LC|22763-7|LNC2HPO|Azotemia|Azotemia
C0880263|T201|DN|22763-7|LNC2HPO|Azotemia|Azotemia
C0880263|T201|MTH_LN|22763-7|LNC2HPO|Azotemia|Azotemia
C0880263|T201|LN|22763-7|LNC2HPO|Azotemia|Azotemia
C0880263|T201|OSN|22763-7|LNC2HPO|Azotemia|Azotemia
C0880263|T201|LC|22763-7|LNC2HPO|Azotaemia|Azotaemia
C0880263|T201|DN|22763-7|LNC2HPO|Azotaemia|Azotaemia
C0880263|T201|MTH_LN|22763-7|LNC2HPO|Azotaemia|Azotaemia
C0880263|T201|LN|22763-7|LNC2HPO|Azotaemia|Azotaemia
C0880263|T201|OSN|22763-7|LNC2HPO|Azotaemia|Azotaemia
C0880263|T201|LC|22763-7|LNC2HPO|Hyperammonemia|Hyperammonemia
C0880263|T201|DN|22763-7|LNC2HPO|Hyperammonemia|Hyperammonemia
C0880263|T201|MTH_LN|22763-7|LNC2HPO|Hyperammonemia|Hyperammonemia
C0880263|T201|LN|22763-7|LNC2HPO|Hyperammonemia|Hyperammonemia
C0880263|T201|OSN|22763-7|LNC2HPO|Hyperammonemia|Hyperammonemia
C0880263|T201|LC|22763-7|LNC2HPO|Hypoammonemia|Hypoammonemia
C0880263|T201|DN|22763-7|LNC2HPO|Hypoammonemia|Hypoammonemia
C0880263|T201|MTH_LN|22763-7|LNC2HPO|Hypoammonemia|Hypoammonemia
C0880263|T201|LN|22763-7|LNC2HPO|Hypoammonemia|Hypoammonemia
C0880263|T201|OSN|22763-7|LNC2HPO|Hypoammonemia|Hypoammonemia
C1315138|T201|LN|32664-5|LNC2HPO|Azotemia|Azotemia
C1315138|T201|DN|32664-5|LNC2HPO|Azotemia|Azotemia
C1315138|T201|OSN|32664-5|LNC2HPO|Azotemia|Azotemia
C1315138|T201|MTH_LN|32664-5|LNC2HPO|Azotemia|Azotemia
C1315138|T201|LC|32664-5|LNC2HPO|Azotemia|Azotemia
C1315138|T201|LN|32664-5|LNC2HPO|Azotaemia|Azotaemia
C1315138|T201|DN|32664-5|LNC2HPO|Azotaemia|Azotaemia
C1315138|T201|OSN|32664-5|LNC2HPO|Azotaemia|Azotaemia
C1315138|T201|MTH_LN|32664-5|LNC2HPO|Azotaemia|Azotaemia
C1315138|T201|LC|32664-5|LNC2HPO|Azotaemia|Azotaemia
C1315138|T201|LN|32664-5|LNC2HPO|Hyperammonemia|Hyperammonemia
C1315138|T201|DN|32664-5|LNC2HPO|Hyperammonemia|Hyperammonemia
C1315138|T201|OSN|32664-5|LNC2HPO|Hyperammonemia|Hyperammonemia
C1315138|T201|MTH_LN|32664-5|LNC2HPO|Hyperammonemia|Hyperammonemia
C1315138|T201|LC|32664-5|LNC2HPO|Hyperammonemia|Hyperammonemia
C1315138|T201|LN|32664-5|LNC2HPO|Hypoammonemia|Hypoammonemia
C1315138|T201|DN|32664-5|LNC2HPO|Hypoammonemia|Hypoammonemia
C1315138|T201|OSN|32664-5|LNC2HPO|Hypoammonemia|Hypoammonemia
C1315138|T201|MTH_LN|32664-5|LNC2HPO|Hypoammonemia|Hypoammonemia
C1315138|T201|LC|32664-5|LNC2HPO|Hypoammonemia|Hypoammonemia
C5201101|T201|LC|35254-2|LNC2HPO|Azotemia|Azotemia
C5201101|T201|DN|35254-2|LNC2HPO|Azotemia|Azotemia
C5201101|T201|MTH_LN|35254-2|LNC2HPO|Azotemia|Azotemia
C5201101|T201|OSN|35254-2|LNC2HPO|Azotemia|Azotemia
C5201101|T201|LN|35254-2|LNC2HPO|Azotemia|Azotemia
C5201101|T201|LC|35254-2|LNC2HPO|Azotaemia|Azotaemia
C5201101|T201|DN|35254-2|LNC2HPO|Azotaemia|Azotaemia
C5201101|T201|MTH_LN|35254-2|LNC2HPO|Azotaemia|Azotaemia
C5201101|T201|OSN|35254-2|LNC2HPO|Azotaemia|Azotaemia
C5201101|T201|LN|35254-2|LNC2HPO|Azotaemia|Azotaemia
C5201101|T201|LC|35254-2|LNC2HPO|Hyperammonemia|Hyperammonemia
C5201101|T201|DN|35254-2|LNC2HPO|Hyperammonemia|Hyperammonemia
C5201101|T201|MTH_LN|35254-2|LNC2HPO|Hyperammonemia|Hyperammonemia
C5201101|T201|OSN|35254-2|LNC2HPO|Hyperammonemia|Hyperammonemia
C5201101|T201|LN|35254-2|LNC2HPO|Hyperammonemia|Hyperammonemia
C5201101|T201|LC|35254-2|LNC2HPO|Hypoammonemia|Hypoammonemia
C5201101|T201|DN|35254-2|LNC2HPO|Hypoammonemia|Hypoammonemia
C5201101|T201|MTH_LN|35254-2|LNC2HPO|Hypoammonemia|Hypoammonemia
C5201101|T201|OSN|35254-2|LNC2HPO|Hypoammonemia|Hypoammonemia
C5201101|T201|LN|35254-2|LNC2HPO|Hypoammonemia|Hypoammonemia
C0484632|T201|LN|9318-7|LNC2HPO|Albuminuria|Albuminuria
C0484632|T201|MTH_LN|9318-7|LNC2HPO|Albuminuria|Albuminuria
C0484632|T201|OSN|9318-7|LNC2HPO|Albuminuria|Albuminuria
C0484632|T201|DN|9318-7|LNC2HPO|Albuminuria|Albuminuria
C0484632|T201|LC|9318-7|LNC2HPO|Albuminuria|Albuminuria
C0363893|T201|LN|1759-0|LNC2HPO|Hyperalbuminemia|Hyperalbuminemia
C0363893|T201|OSN|1759-0|LNC2HPO|Hyperalbuminemia|Hyperalbuminemia
C0363893|T201|MTH_LN|1759-0|LNC2HPO|Hyperalbuminemia|Hyperalbuminemia
C0363893|T201|DN|1759-0|LNC2HPO|Hyperalbuminemia|Hyperalbuminemia
C0363893|T201|LC|1759-0|LNC2HPO|Hyperalbuminemia|Hyperalbuminemia
C0363893|T201|LN|1759-0|LNC2HPO|Hyperalbuminaemia|Hyperalbuminaemia
C0363893|T201|OSN|1759-0|LNC2HPO|Hyperalbuminaemia|Hyperalbuminaemia
C0363893|T201|MTH_LN|1759-0|LNC2HPO|Hyperalbuminaemia|Hyperalbuminaemia
C0363893|T201|DN|1759-0|LNC2HPO|Hyperalbuminaemia|Hyperalbuminaemia
C0363893|T201|LC|1759-0|LNC2HPO|Hyperalbuminaemia|Hyperalbuminaemia
C0363893|T201|LN|1759-0|LNC2HPO|Hypoalbuminemia|Hypoalbuminemia
C0363893|T201|OSN|1759-0|LNC2HPO|Hypoalbuminemia|Hypoalbuminemia
C0363893|T201|MTH_LN|1759-0|LNC2HPO|Hypoalbuminemia|Hypoalbuminemia
C0363893|T201|DN|1759-0|LNC2HPO|Hypoalbuminemia|Hypoalbuminemia
C0363893|T201|LC|1759-0|LNC2HPO|Hypoalbuminemia|Hypoalbuminemia
C0363893|T201|LN|1759-0|LNC2HPO|Hypoalbuminaemia|Hypoalbuminaemia
C0363893|T201|OSN|1759-0|LNC2HPO|Hypoalbuminaemia|Hypoalbuminaemia
C0363893|T201|MTH_LN|1759-0|LNC2HPO|Hypoalbuminaemia|Hypoalbuminaemia
C0363893|T201|DN|1759-0|LNC2HPO|Hypoalbuminaemia|Hypoalbuminaemia
C0363893|T201|LC|1759-0|LNC2HPO|Hypoalbuminaemia|Hypoalbuminaemia
C0941344|T201|LN|25145-4|LNC2HPO|Bacteriuria|Bacteriuria
C0941344|T201|MTH_LN|25145-4|LNC2HPO|Bacteriuria|Bacteriuria
C0941344|T201|DN|25145-4|LNC2HPO|Bacteriuria|Bacteriuria
C0941344|T201|OSN|25145-4|LNC2HPO|Bacteriuria|Bacteriuria
C0941344|T201|LC|25145-4|LNC2HPO|Bacteriuria|Bacteriuria
C0368563|T201|LN|630-4|LNC2HPO|Bacteriuria|Bacteriuria
C0368563|T201|DN|630-4|LNC2HPO|Bacteriuria|Bacteriuria
C0368563|T201|MTH_LN|630-4|LNC2HPO|Bacteriuria|Bacteriuria
C0368563|T201|OSN|630-4|LNC2HPO|Bacteriuria|Bacteriuria
C0368563|T201|LC|630-4|LNC2HPO|Bacteriuria|Bacteriuria
C0484511|T201|LN|10438-0|LNC2HPO|Increase in B cell count|Increase in B cell count
C0484511|T201|MTH_LN|10438-0|LNC2HPO|Increase in B cell count|Increase in B cell count
C0484511|T201|DN|10438-0|LNC2HPO|Increase in B cell count|Increase in B cell count
C0484511|T201|OSN|10438-0|LNC2HPO|Increase in B cell count|Increase in B cell count
C0484511|T201|LC|10438-0|LNC2HPO|Increase in B cell count|Increase in B cell count
C0363783|T201|LN|1649-3|LNC2HPO|Hypercalciuria|Hypercalciuria
C0363783|T201|DN|1649-3|LNC2HPO|Hypercalciuria|Hypercalciuria
C0363783|T201|MTH_LN|1649-3|LNC2HPO|Hypercalciuria|Hypercalciuria
C0363783|T201|LC|1649-3|LNC2HPO|Hypercalciuria|Hypercalciuria
C0363783|T201|OSN|1649-3|LNC2HPO|Hypercalciuria|Hypercalciuria
C0363783|T201|LN|1649-3|LNC2HPO|Hypercalcinuria|Hypercalcinuria
C0363783|T201|DN|1649-3|LNC2HPO|Hypercalcinuria|Hypercalcinuria
C0363783|T201|MTH_LN|1649-3|LNC2HPO|Hypercalcinuria|Hypercalcinuria
C0363783|T201|LC|1649-3|LNC2HPO|Hypercalcinuria|Hypercalcinuria
C0363783|T201|OSN|1649-3|LNC2HPO|Hypercalcinuria|Hypercalcinuria
C0363783|T201|LN|1649-3|LNC2HPO|Hypocalciuria|Hypocalciuria
C0363783|T201|DN|1649-3|LNC2HPO|Hypocalciuria|Hypocalciuria
C0363783|T201|MTH_LN|1649-3|LNC2HPO|Hypocalciuria|Hypocalciuria
C0363783|T201|LC|1649-3|LNC2HPO|Hypocalciuria|Hypocalciuria
C0363783|T201|OSN|1649-3|LNC2HPO|Hypocalciuria|Hypocalciuria
C0484673|T201|LN|6874-2|LNC2HPO|Hypercalciuria|Hypercalciuria
C0484673|T201|MTH_LN|6874-2|LNC2HPO|Hypercalciuria|Hypercalciuria
C0484673|T201|DN|6874-2|LNC2HPO|Hypercalciuria|Hypercalciuria
C0484673|T201|OSN|6874-2|LNC2HPO|Hypercalciuria|Hypercalciuria
C0484673|T201|LC|6874-2|LNC2HPO|Hypercalciuria|Hypercalciuria
C0484673|T201|LN|6874-2|LNC2HPO|Hypercalcinuria|Hypercalcinuria
C0484673|T201|MTH_LN|6874-2|LNC2HPO|Hypercalcinuria|Hypercalcinuria
C0484673|T201|DN|6874-2|LNC2HPO|Hypercalcinuria|Hypercalcinuria
C0484673|T201|OSN|6874-2|LNC2HPO|Hypercalcinuria|Hypercalcinuria
C0484673|T201|LC|6874-2|LNC2HPO|Hypercalcinuria|Hypercalcinuria
C0484673|T201|LN|6874-2|LNC2HPO|Hypocalciuria|Hypocalciuria
C0484673|T201|MTH_LN|6874-2|LNC2HPO|Hypocalciuria|Hypocalciuria
C0484673|T201|DN|6874-2|LNC2HPO|Hypocalciuria|Hypocalciuria
C0484673|T201|OSN|6874-2|LNC2HPO|Hypocalciuria|Hypocalciuria
C0484673|T201|LC|6874-2|LNC2HPO|Hypocalciuria|Hypocalciuria
C0800969|T201|LC|17862-4|LNC2HPO|Hypercalciuria|Hypercalciuria
C0800969|T201|MTH_LN|17862-4|LNC2HPO|Hypercalciuria|Hypercalciuria
C0800969|T201|DN|17862-4|LNC2HPO|Hypercalciuria|Hypercalciuria
C0800969|T201|OSN|17862-4|LNC2HPO|Hypercalciuria|Hypercalciuria
C0800969|T201|LN|17862-4|LNC2HPO|Hypercalciuria|Hypercalciuria
C0800969|T201|LC|17862-4|LNC2HPO|Hypercalcinuria|Hypercalcinuria
C0800969|T201|MTH_LN|17862-4|LNC2HPO|Hypercalcinuria|Hypercalcinuria
C0800969|T201|DN|17862-4|LNC2HPO|Hypercalcinuria|Hypercalcinuria
C0800969|T201|OSN|17862-4|LNC2HPO|Hypercalcinuria|Hypercalcinuria
C0800969|T201|LN|17862-4|LNC2HPO|Hypercalcinuria|Hypercalcinuria
C0800969|T201|LC|17862-4|LNC2HPO|Hypocalciuria|Hypocalciuria
C0800969|T201|MTH_LN|17862-4|LNC2HPO|Hypocalciuria|Hypocalciuria
C0800969|T201|DN|17862-4|LNC2HPO|Hypocalciuria|Hypocalciuria
C0800969|T201|OSN|17862-4|LNC2HPO|Hypocalciuria|Hypocalciuria
C0800969|T201|LN|17862-4|LNC2HPO|Hypocalciuria|Hypocalciuria
C0800971|T201|LN|17864-0|LNC2HPO|Hypercalcemia|Hypercalcemia
C0800971|T201|DN|17864-0|LNC2HPO|Hypercalcemia|Hypercalcemia
C0800971|T201|MTH_LN|17864-0|LNC2HPO|Hypercalcemia|Hypercalcemia
C0800971|T201|OSN|17864-0|LNC2HPO|Hypercalcemia|Hypercalcemia
C0800971|T201|LC|17864-0|LNC2HPO|Hypercalcemia|Hypercalcemia
C0800971|T201|LN|17864-0|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0800971|T201|DN|17864-0|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0800971|T201|MTH_LN|17864-0|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0800971|T201|OSN|17864-0|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0800971|T201|LC|17864-0|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0800971|T201|LN|17864-0|LNC2HPO|Hypocalcemia|Hypocalcemia
C0800971|T201|DN|17864-0|LNC2HPO|Hypocalcemia|Hypocalcemia
C0800971|T201|MTH_LN|17864-0|LNC2HPO|Hypocalcemia|Hypocalcemia
C0800971|T201|OSN|17864-0|LNC2HPO|Hypocalcemia|Hypocalcemia
C0800971|T201|LC|17864-0|LNC2HPO|Hypocalcemia|Hypocalcemia
C0800971|T201|LN|17864-0|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0800971|T201|DN|17864-0|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0800971|T201|MTH_LN|17864-0|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0800971|T201|OSN|17864-0|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0800971|T201|LC|17864-0|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364153|T201|LN|2021-4|LNC2HPO|Hypercapnia|Hypercapnia
C0364153|T201|MTH_LN|2021-4|LNC2HPO|Hypercapnia|Hypercapnia
C0364153|T201|DN|2021-4|LNC2HPO|Hypercapnia|Hypercapnia
C0364153|T201|OSN|2021-4|LNC2HPO|Hypercapnia|Hypercapnia
C0364153|T201|LC|2021-4|LNC2HPO|Hypercapnia|Hypercapnia
C0364153|T201|LN|2021-4|LNC2HPO|Hypercarbia|Hypercarbia
C0364153|T201|MTH_LN|2021-4|LNC2HPO|Hypercarbia|Hypercarbia
C0364153|T201|DN|2021-4|LNC2HPO|Hypercarbia|Hypercarbia
C0364153|T201|OSN|2021-4|LNC2HPO|Hypercarbia|Hypercarbia
C0364153|T201|LC|2021-4|LNC2HPO|Hypercarbia|Hypercarbia
C0364153|T201|LN|2021-4|LNC2HPO|Hypocapnia|Hypocapnia
C0364153|T201|MTH_LN|2021-4|LNC2HPO|Hypocapnia|Hypocapnia
C0364153|T201|DN|2021-4|LNC2HPO|Hypocapnia|Hypocapnia
C0364153|T201|OSN|2021-4|LNC2HPO|Hypocapnia|Hypocapnia
C0364153|T201|LC|2021-4|LNC2HPO|Hypocapnia|Hypocapnia
C0364153|T201|LN|2021-4|LNC2HPO|Hypocarbia|Hypocarbia
C0364153|T201|MTH_LN|2021-4|LNC2HPO|Hypocarbia|Hypocarbia
C0364153|T201|DN|2021-4|LNC2HPO|Hypocarbia|Hypocarbia
C0364153|T201|OSN|2021-4|LNC2HPO|Hypocarbia|Hypocarbia
C0364153|T201|LC|2021-4|LNC2HPO|Hypocarbia|Hypocarbia
C1315242|T201|LN|32771-8|LNC2HPO|Hypercapnia|Hypercapnia
C1315242|T201|DN|32771-8|LNC2HPO|Hypercapnia|Hypercapnia
C1315242|T201|MTH_LN|32771-8|LNC2HPO|Hypercapnia|Hypercapnia
C1315242|T201|LC|32771-8|LNC2HPO|Hypercapnia|Hypercapnia
C1315242|T201|OSN|32771-8|LNC2HPO|Hypercapnia|Hypercapnia
C1315242|T201|LN|32771-8|LNC2HPO|Hypercarbia|Hypercarbia
C1315242|T201|DN|32771-8|LNC2HPO|Hypercarbia|Hypercarbia
C1315242|T201|MTH_LN|32771-8|LNC2HPO|Hypercarbia|Hypercarbia
C1315242|T201|LC|32771-8|LNC2HPO|Hypercarbia|Hypercarbia
C1315242|T201|OSN|32771-8|LNC2HPO|Hypercarbia|Hypercarbia
C1315242|T201|LN|32771-8|LNC2HPO|Hypocapnia|Hypocapnia
C1315242|T201|DN|32771-8|LNC2HPO|Hypocapnia|Hypocapnia
C1315242|T201|MTH_LN|32771-8|LNC2HPO|Hypocapnia|Hypocapnia
C1315242|T201|LC|32771-8|LNC2HPO|Hypocapnia|Hypocapnia
C1315242|T201|OSN|32771-8|LNC2HPO|Hypocapnia|Hypocapnia
C1315242|T201|LN|32771-8|LNC2HPO|Hypocarbia|Hypocarbia
C1315242|T201|DN|32771-8|LNC2HPO|Hypocarbia|Hypocarbia
C1315242|T201|MTH_LN|32771-8|LNC2HPO|Hypocarbia|Hypocarbia
C1315242|T201|LC|32771-8|LNC2HPO|Hypocarbia|Hypocarbia
C1315242|T201|OSN|32771-8|LNC2HPO|Hypocarbia|Hypocarbia
C0482544|T201|MTH_LN|1558-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482544|T201|LN|1558-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482544|T201|DN|1558-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482544|T201|OSN|1558-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482544|T201|LC|1558-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0482544|T201|MTH_LN|1558-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482544|T201|LN|1558-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482544|T201|DN|1558-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482544|T201|OSN|1558-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482544|T201|LC|1558-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0482544|T201|MTH_LN|1558-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482544|T201|LN|1558-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482544|T201|DN|1558-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482544|T201|OSN|1558-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0482544|T201|LC|1558-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0796934|T201|LN|13744-8|LNC2HPO|Galactosuria|Galactosuria
C0796934|T201|OSN|13744-8|LNC2HPO|Galactosuria|Galactosuria
C0796934|T201|MTH_LN|13744-8|LNC2HPO|Galactosuria|Galactosuria
C0796934|T201|DN|13744-8|LNC2HPO|Galactosuria|Galactosuria
C0796934|T201|LC|13744-8|LNC2HPO|Galactosuria|Galactosuria
C0363617|T201|LN|1483-7|LNC2HPO|Galactosuria|Galactosuria
C0363617|T201|MTH_LN|1483-7|LNC2HPO|Galactosuria|Galactosuria
C0363617|T201|DN|1483-7|LNC2HPO|Galactosuria|Galactosuria
C0363617|T201|OSN|1483-7|LNC2HPO|Galactosuria|Galactosuria
C0363617|T201|LC|1483-7|LNC2HPO|Galactosuria|Galactosuria
C0798243|T201|LN|15071-4|LNC2HPO|Galactosuria|Galactosuria
C0798243|T201|MTH_LN|15071-4|LNC2HPO|Galactosuria|Galactosuria
C0798243|T201|DN|15071-4|LNC2HPO|Galactosuria|Galactosuria
C0798243|T201|OSN|15071-4|LNC2HPO|Galactosuria|Galactosuria
C0798243|T201|LC|15071-4|LNC2HPO|Galactosuria|Galactosuria
C0941310|T201|LN|25102-5|LNC2HPO|Galactosuria|Galactosuria
C0941310|T201|DN|25102-5|LNC2HPO|Galactosuria|Galactosuria
C0941310|T201|OSN|25102-5|LNC2HPO|Galactosuria|Galactosuria
C0941310|T201|LC|25102-5|LNC2HPO|Galactosuria|Galactosuria
C0941310|T201|MTH_LN|25102-5|LNC2HPO|Galactosuria|Galactosuria
C1316773|T201|LN|34310-3|LNC2HPO|Galactosuria|Galactosuria
C1316773|T201|DN|34310-3|LNC2HPO|Galactosuria|Galactosuria
C1316773|T201|MTH_LN|34310-3|LNC2HPO|Galactosuria|Galactosuria
C1316773|T201|OSN|34310-3|LNC2HPO|Galactosuria|Galactosuria
C1316773|T201|LC|34310-3|LNC2HPO|Galactosuria|Galactosuria
C0363613|T201|LN|1479-5|LNC2HPO|Galactosemia|Galactosemia
C0363613|T201|DN|1479-5|LNC2HPO|Galactosemia|Galactosemia
C0363613|T201|OSN|1479-5|LNC2HPO|Galactosemia|Galactosemia
C0363613|T201|MTH_LN|1479-5|LNC2HPO|Galactosemia|Galactosemia
C0363613|T201|LC|1479-5|LNC2HPO|Galactosemia|Galactosemia
C0363613|T201|LN|1479-5|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0363613|T201|DN|1479-5|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0363613|T201|OSN|1479-5|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0363613|T201|MTH_LN|1479-5|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0363613|T201|LC|1479-5|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0363614|T201|LN|1480-3|LNC2HPO|Galactosemia|Galactosemia
C0363614|T201|MTH_LN|1480-3|LNC2HPO|Galactosemia|Galactosemia
C0363614|T201|DN|1480-3|LNC2HPO|Galactosemia|Galactosemia
C0363614|T201|OSN|1480-3|LNC2HPO|Galactosemia|Galactosemia
C0363614|T201|LC|1480-3|LNC2HPO|Galactosemia|Galactosemia
C0363614|T201|LN|1480-3|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0363614|T201|MTH_LN|1480-3|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0363614|T201|DN|1480-3|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0363614|T201|OSN|1480-3|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0363614|T201|LC|1480-3|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0363615|T201|LN|1481-1|LNC2HPO|Galactosemia|Galactosemia
C0363615|T201|MTH_LN|1481-1|LNC2HPO|Galactosemia|Galactosemia
C0363615|T201|DN|1481-1|LNC2HPO|Galactosemia|Galactosemia
C0363615|T201|OSN|1481-1|LNC2HPO|Galactosemia|Galactosemia
C0363615|T201|LC|1481-1|LNC2HPO|Galactosemia|Galactosemia
C0363615|T201|LN|1481-1|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0363615|T201|MTH_LN|1481-1|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0363615|T201|DN|1481-1|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0363615|T201|OSN|1481-1|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0363615|T201|LC|1481-1|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0363616|T201|LN|1482-9|LNC2HPO|Galactosemia|Galactosemia
C0363616|T201|MTH_LN|1482-9|LNC2HPO|Galactosemia|Galactosemia
C0363616|T201|DN|1482-9|LNC2HPO|Galactosemia|Galactosemia
C0363616|T201|OSN|1482-9|LNC2HPO|Galactosemia|Galactosemia
C0363616|T201|LC|1482-9|LNC2HPO|Galactosemia|Galactosemia
C0363616|T201|LN|1482-9|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0363616|T201|MTH_LN|1482-9|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0363616|T201|DN|1482-9|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0363616|T201|OSN|1482-9|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0363616|T201|LC|1482-9|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0364441|T201|LN|2306-9|LNC2HPO|Galactosemia|Galactosemia
C0364441|T201|MTH_LN|2306-9|LNC2HPO|Galactosemia|Galactosemia
C0364441|T201|OSN|2306-9|LNC2HPO|Galactosemia|Galactosemia
C0364441|T201|DN|2306-9|LNC2HPO|Galactosemia|Galactosemia
C0364441|T201|LC|2306-9|LNC2HPO|Galactosemia|Galactosemia
C0364441|T201|LN|2306-9|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0364441|T201|MTH_LN|2306-9|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0364441|T201|OSN|2306-9|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0364441|T201|DN|2306-9|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0364441|T201|LC|2306-9|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0364442|T201|LN|2307-7|LNC2HPO|Galactosemia|Galactosemia
C0364442|T201|MTH_LN|2307-7|LNC2HPO|Galactosemia|Galactosemia
C0364442|T201|DN|2307-7|LNC2HPO|Galactosemia|Galactosemia
C0364442|T201|OSN|2307-7|LNC2HPO|Galactosemia|Galactosemia
C0364442|T201|LC|2307-7|LNC2HPO|Galactosemia|Galactosemia
C0364442|T201|LN|2307-7|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0364442|T201|MTH_LN|2307-7|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0364442|T201|DN|2307-7|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0364442|T201|OSN|2307-7|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0364442|T201|LC|2307-7|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0364443|T201|LN|2308-5|LNC2HPO|Galactosemia|Galactosemia
C0364443|T201|DN|2308-5|LNC2HPO|Galactosemia|Galactosemia
C0364443|T201|MTH_LN|2308-5|LNC2HPO|Galactosemia|Galactosemia
C0364443|T201|OSN|2308-5|LNC2HPO|Galactosemia|Galactosemia
C0364443|T201|LC|2308-5|LNC2HPO|Galactosemia|Galactosemia
C0364443|T201|LN|2308-5|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0364443|T201|DN|2308-5|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0364443|T201|MTH_LN|2308-5|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0364443|T201|OSN|2308-5|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0364443|T201|LC|2308-5|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0364444|T201|LN|2309-3|LNC2HPO|Galactosuria|Galactosuria
C0364444|T201|MTH_LN|2309-3|LNC2HPO|Galactosuria|Galactosuria
C0364444|T201|DN|2309-3|LNC2HPO|Galactosuria|Galactosuria
C0364444|T201|OSN|2309-3|LNC2HPO|Galactosuria|Galactosuria
C0364444|T201|LC|2309-3|LNC2HPO|Galactosuria|Galactosuria
C0364445|T201|LN|2310-1|LNC2HPO|Galactosuria|Galactosuria
C0364445|T201|MTH_LN|2310-1|LNC2HPO|Galactosuria|Galactosuria
C0364445|T201|DN|2310-1|LNC2HPO|Galactosuria|Galactosuria
C0364445|T201|OSN|2310-1|LNC2HPO|Galactosuria|Galactosuria
C0364445|T201|LC|2310-1|LNC2HPO|Galactosuria|Galactosuria
C0941571|T201|LN|25426-8|LNC2HPO|Galactosemia|Galactosemia
C0941571|T201|DN|25426-8|LNC2HPO|Galactosemia|Galactosemia
C0941571|T201|MTH_LN|25426-8|LNC2HPO|Galactosemia|Galactosemia
C0941571|T201|OSN|25426-8|LNC2HPO|Galactosemia|Galactosemia
C0941571|T201|LC|25426-8|LNC2HPO|Galactosemia|Galactosemia
C0941571|T201|LN|25426-8|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0941571|T201|DN|25426-8|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0941571|T201|MTH_LN|25426-8|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0941571|T201|OSN|25426-8|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0941571|T201|LC|25426-8|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C1954977|T201|LN|49219-9|LNC2HPO|Galactosemia|Galactosemia
C1954977|T201|DN|49219-9|LNC2HPO|Galactosemia|Galactosemia
C1954977|T201|OSN|49219-9|LNC2HPO|Galactosemia|Galactosemia
C1954977|T201|MTH_LN|49219-9|LNC2HPO|Galactosemia|Galactosemia
C1954977|T201|LC|49219-9|LNC2HPO|Galactosemia|Galactosemia
C1954977|T201|LN|49219-9|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C1954977|T201|DN|49219-9|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C1954977|T201|OSN|49219-9|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C1954977|T201|MTH_LN|49219-9|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C1954977|T201|LC|49219-9|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C2599398|T201|LN|54084-9|LNC2HPO|Galactosemia|Galactosemia
C2599398|T201|LC|54084-9|LNC2HPO|Galactosemia|Galactosemia
C2599398|T201|DN|54084-9|LNC2HPO|Galactosemia|Galactosemia
C2599398|T201|MTH_LN|54084-9|LNC2HPO|Galactosemia|Galactosemia
C2599398|T201|OSN|54084-9|LNC2HPO|Galactosemia|Galactosemia
C2599398|T201|LN|54084-9|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C2599398|T201|LC|54084-9|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C2599398|T201|DN|54084-9|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C2599398|T201|MTH_LN|54084-9|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C2599398|T201|OSN|54084-9|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C2599399|T201|LN|54085-6|LNC2HPO|Galactosemia|Galactosemia
C2599399|T201|LC|54085-6|LNC2HPO|Galactosemia|Galactosemia
C2599399|T201|DN|54085-6|LNC2HPO|Galactosemia|Galactosemia
C2599399|T201|MTH_LN|54085-6|LNC2HPO|Galactosemia|Galactosemia
C2599399|T201|OSN|54085-6|LNC2HPO|Galactosemia|Galactosemia
C2599399|T201|LN|54085-6|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C2599399|T201|LC|54085-6|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C2599399|T201|DN|54085-6|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C2599399|T201|MTH_LN|54085-6|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C2599399|T201|OSN|54085-6|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C3846901|T201|LN|75093-5|LNC2HPO|Galactosemia|Galactosemia
C3846901|T201|OSN|75093-5|LNC2HPO|Galactosemia|Galactosemia
C3846901|T201|MTH_LN|75093-5|LNC2HPO|Galactosemia|Galactosemia
C3846901|T201|LC|75093-5|LNC2HPO|Galactosemia|Galactosemia
C3846901|T201|DN|75093-5|LNC2HPO|Galactosemia|Galactosemia
C3846901|T201|LN|75093-5|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C3846901|T201|OSN|75093-5|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C3846901|T201|MTH_LN|75093-5|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C3846901|T201|LC|75093-5|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C3846901|T201|DN|75093-5|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C1316774|T201|LN|34311-1|LNC2HPO|Galactosuria|Galactosuria
C1316774|T201|DN|34311-1|LNC2HPO|Galactosuria|Galactosuria
C1316774|T201|MTH_LN|34311-1|LNC2HPO|Galactosuria|Galactosuria
C1316774|T201|OSN|34311-1|LNC2HPO|Galactosuria|Galactosuria
C1316774|T201|LC|34311-1|LNC2HPO|Galactosuria|Galactosuria
C0796799|T201|LN|13608-5|LNC2HPO|Hyperinsulinemia|Hyperinsulinemia
C0796799|T201|DN|13608-5|LNC2HPO|Hyperinsulinemia|Hyperinsulinemia
C0796799|T201|OSN|13608-5|LNC2HPO|Hyperinsulinemia|Hyperinsulinemia
C0796799|T201|MTH_LN|13608-5|LNC2HPO|Hyperinsulinemia|Hyperinsulinemia
C0796799|T201|LC|13608-5|LNC2HPO|Hyperinsulinemia|Hyperinsulinemia
C0796799|T201|LN|13608-5|LNC2HPO|Hypoinsulinemia|Hypoinsulinemia
C0796799|T201|DN|13608-5|LNC2HPO|Hypoinsulinemia|Hypoinsulinemia
C0796799|T201|OSN|13608-5|LNC2HPO|Hypoinsulinemia|Hypoinsulinemia
C0796799|T201|MTH_LN|13608-5|LNC2HPO|Hypoinsulinemia|Hypoinsulinemia
C0796799|T201|LC|13608-5|LNC2HPO|Hypoinsulinemia|Hypoinsulinemia
C0796800|T201|LN|13609-3|LNC2HPO|Hyperinsulinemia|Hyperinsulinemia
C0796800|T201|DN|13609-3|LNC2HPO|Hyperinsulinemia|Hyperinsulinemia
C0796800|T201|OSN|13609-3|LNC2HPO|Hyperinsulinemia|Hyperinsulinemia
C0796800|T201|MTH_LN|13609-3|LNC2HPO|Hyperinsulinemia|Hyperinsulinemia
C0796800|T201|LC|13609-3|LNC2HPO|Hyperinsulinemia|Hyperinsulinemia
C0796800|T201|LN|13609-3|LNC2HPO|Hypoinsulinemia|Hypoinsulinemia
C0796800|T201|DN|13609-3|LNC2HPO|Hypoinsulinemia|Hypoinsulinemia
C0796800|T201|OSN|13609-3|LNC2HPO|Hypoinsulinemia|Hypoinsulinemia
C0796800|T201|MTH_LN|13609-3|LNC2HPO|Hypoinsulinemia|Hypoinsulinemia
C0796800|T201|LC|13609-3|LNC2HPO|Hypoinsulinemia|Hypoinsulinemia
C0363625|T201|LN|1491-0|LNC2HPO|Glycosuria|Glycosuria
C0363625|T201|MTH_LN|1491-0|LNC2HPO|Glycosuria|Glycosuria
C0363625|T201|DN|1491-0|LNC2HPO|Glycosuria|Glycosuria
C0363625|T201|OSN|1491-0|LNC2HPO|Glycosuria|Glycosuria
C0363625|T201|LC|1491-0|LNC2HPO|Glycosuria|Glycosuria
C0363625|T201|LN|1491-0|LNC2HPO|Glucosuria|Glucosuria
C0363625|T201|MTH_LN|1491-0|LNC2HPO|Glucosuria|Glucosuria
C0363625|T201|DN|1491-0|LNC2HPO|Glucosuria|Glucosuria
C0363625|T201|OSN|1491-0|LNC2HPO|Glucosuria|Glucosuria
C0363625|T201|LC|1491-0|LNC2HPO|Glucosuria|Glucosuria
C0363629|T201|LN|1495-1|LNC2HPO|Glycosuria|Glycosuria
C0363629|T201|DN|1495-1|LNC2HPO|Glycosuria|Glycosuria
C0363629|T201|OSN|1495-1|LNC2HPO|Glycosuria|Glycosuria
C0363629|T201|MTH_LN|1495-1|LNC2HPO|Glycosuria|Glycosuria
C0363629|T201|LC|1495-1|LNC2HPO|Glycosuria|Glycosuria
C0363629|T201|LN|1495-1|LNC2HPO|Glucosuria|Glucosuria
C0363629|T201|DN|1495-1|LNC2HPO|Glucosuria|Glucosuria
C0363629|T201|OSN|1495-1|LNC2HPO|Glucosuria|Glucosuria
C0363629|T201|MTH_LN|1495-1|LNC2HPO|Glucosuria|Glucosuria
C0363629|T201|LC|1495-1|LNC2HPO|Glucosuria|Glucosuria
C0363639|T201|LN|1505-7|LNC2HPO|Glycosuria|Glycosuria
C0363639|T201|MTH_LN|1505-7|LNC2HPO|Glycosuria|Glycosuria
C0363639|T201|DN|1505-7|LNC2HPO|Glycosuria|Glycosuria
C0363639|T201|OSN|1505-7|LNC2HPO|Glycosuria|Glycosuria
C0363639|T201|LC|1505-7|LNC2HPO|Glycosuria|Glycosuria
C0363639|T201|LN|1505-7|LNC2HPO|Glucosuria|Glucosuria
C0363639|T201|MTH_LN|1505-7|LNC2HPO|Glucosuria|Glucosuria
C0363639|T201|DN|1505-7|LNC2HPO|Glucosuria|Glucosuria
C0363639|T201|OSN|1505-7|LNC2HPO|Glucosuria|Glucosuria
C0363639|T201|LC|1505-7|LNC2HPO|Glucosuria|Glucosuria
C0798248|T201|LN|15076-3|LNC2HPO|Glycosuria|Glycosuria
C0798248|T201|MTH_LN|15076-3|LNC2HPO|Glycosuria|Glycosuria
C0798248|T201|DN|15076-3|LNC2HPO|Glycosuria|Glycosuria
C0798248|T201|OSN|15076-3|LNC2HPO|Glycosuria|Glycosuria
C0798248|T201|LC|15076-3|LNC2HPO|Glycosuria|Glycosuria
C0798248|T201|LN|15076-3|LNC2HPO|Glucosuria|Glucosuria
C0798248|T201|MTH_LN|15076-3|LNC2HPO|Glucosuria|Glucosuria
C0798248|T201|DN|15076-3|LNC2HPO|Glucosuria|Glucosuria
C0798248|T201|OSN|15076-3|LNC2HPO|Glucosuria|Glucosuria
C0798248|T201|LC|15076-3|LNC2HPO|Glucosuria|Glucosuria
C0798249|T201|LN|15077-1|LNC2HPO|Glycosuria|Glycosuria
C0798249|T201|MTH_LN|15077-1|LNC2HPO|Glycosuria|Glycosuria
C0798249|T201|DN|15077-1|LNC2HPO|Glycosuria|Glycosuria
C0798249|T201|OSN|15077-1|LNC2HPO|Glycosuria|Glycosuria
C0798249|T201|LC|15077-1|LNC2HPO|Glycosuria|Glycosuria
C0798249|T201|LN|15077-1|LNC2HPO|Glucosuria|Glucosuria
C0798249|T201|MTH_LN|15077-1|LNC2HPO|Glucosuria|Glucosuria
C0798249|T201|DN|15077-1|LNC2HPO|Glucosuria|Glucosuria
C0798249|T201|OSN|15077-1|LNC2HPO|Glucosuria|Glucosuria
C0798249|T201|LC|15077-1|LNC2HPO|Glucosuria|Glucosuria
C0363643|T201|LN|1509-9|LNC2HPO|Glycosuria|Glycosuria
C0363643|T201|MTH_LN|1509-9|LNC2HPO|Glycosuria|Glycosuria
C0363643|T201|DN|1509-9|LNC2HPO|Glycosuria|Glycosuria
C0363643|T201|OSN|1509-9|LNC2HPO|Glycosuria|Glycosuria
C0363643|T201|LC|1509-9|LNC2HPO|Glycosuria|Glycosuria
C0363643|T201|LN|1509-9|LNC2HPO|Glucosuria|Glucosuria
C0363643|T201|MTH_LN|1509-9|LNC2HPO|Glucosuria|Glucosuria
C0363643|T201|DN|1509-9|LNC2HPO|Glucosuria|Glucosuria
C0363643|T201|OSN|1509-9|LNC2HPO|Glucosuria|Glucosuria
C0363643|T201|LC|1509-9|LNC2HPO|Glucosuria|Glucosuria
C0363686|T201|LN|1555-2|LNC2HPO|Glycosuria|Glycosuria
C0363686|T201|MTH_LN|1555-2|LNC2HPO|Glycosuria|Glycosuria
C0363686|T201|DN|1555-2|LNC2HPO|Glycosuria|Glycosuria
C0363686|T201|OSN|1555-2|LNC2HPO|Glycosuria|Glycosuria
C0363686|T201|LC|1555-2|LNC2HPO|Glycosuria|Glycosuria
C0363686|T201|LN|1555-2|LNC2HPO|Glucosuria|Glucosuria
C0363686|T201|MTH_LN|1555-2|LNC2HPO|Glucosuria|Glucosuria
C0363686|T201|DN|1555-2|LNC2HPO|Glucosuria|Glucosuria
C0363686|T201|OSN|1555-2|LNC2HPO|Glucosuria|Glucosuria
C0363686|T201|LC|1555-2|LNC2HPO|Glucosuria|Glucosuria
C0801273|T201|LN|18227-9|LNC2HPO|Glycosuria|Glycosuria
C0801273|T201|MTH_LN|18227-9|LNC2HPO|Glycosuria|Glycosuria
C0801273|T201|DN|18227-9|LNC2HPO|Glycosuria|Glycosuria
C0801273|T201|OSN|18227-9|LNC2HPO|Glycosuria|Glycosuria
C0801273|T201|LC|18227-9|LNC2HPO|Glycosuria|Glycosuria
C0801273|T201|LN|18227-9|LNC2HPO|Glucosuria|Glucosuria
C0801273|T201|MTH_LN|18227-9|LNC2HPO|Glucosuria|Glucosuria
C0801273|T201|DN|18227-9|LNC2HPO|Glucosuria|Glucosuria
C0801273|T201|OSN|18227-9|LNC2HPO|Glucosuria|Glucosuria
C0801273|T201|LC|18227-9|LNC2HPO|Glucosuria|Glucosuria
C0804099|T201|LN|21305-8|LNC2HPO|Glycosuria|Glycosuria
C0804099|T201|MTH_LN|21305-8|LNC2HPO|Glycosuria|Glycosuria
C0804099|T201|DN|21305-8|LNC2HPO|Glycosuria|Glycosuria
C0804099|T201|OSN|21305-8|LNC2HPO|Glycosuria|Glycosuria
C0804099|T201|LC|21305-8|LNC2HPO|Glycosuria|Glycosuria
C0804099|T201|LN|21305-8|LNC2HPO|Glucosuria|Glucosuria
C0804099|T201|MTH_LN|21305-8|LNC2HPO|Glucosuria|Glucosuria
C0804099|T201|DN|21305-8|LNC2HPO|Glucosuria|Glucosuria
C0804099|T201|OSN|21305-8|LNC2HPO|Glucosuria|Glucosuria
C0804099|T201|LC|21305-8|LNC2HPO|Glucosuria|Glucosuria
C0804100|T201|LN|21306-6|LNC2HPO|Glycosuria|Glycosuria
C0804100|T201|MTH_LN|21306-6|LNC2HPO|Glycosuria|Glycosuria
C0804100|T201|DN|21306-6|LNC2HPO|Glycosuria|Glycosuria
C0804100|T201|OSN|21306-6|LNC2HPO|Glycosuria|Glycosuria
C0804100|T201|LC|21306-6|LNC2HPO|Glycosuria|Glycosuria
C0804100|T201|LN|21306-6|LNC2HPO|Glucosuria|Glucosuria
C0804100|T201|MTH_LN|21306-6|LNC2HPO|Glucosuria|Glucosuria
C0804100|T201|DN|21306-6|LNC2HPO|Glucosuria|Glucosuria
C0804100|T201|OSN|21306-6|LNC2HPO|Glucosuria|Glucosuria
C0804100|T201|LC|21306-6|LNC2HPO|Glucosuria|Glucosuria
C0804101|T201|LN|21307-4|LNC2HPO|Glycosuria|Glycosuria
C0804101|T201|MTH_LN|21307-4|LNC2HPO|Glycosuria|Glycosuria
C0804101|T201|DN|21307-4|LNC2HPO|Glycosuria|Glycosuria
C0804101|T201|OSN|21307-4|LNC2HPO|Glycosuria|Glycosuria
C0804101|T201|LC|21307-4|LNC2HPO|Glycosuria|Glycosuria
C0804101|T201|LN|21307-4|LNC2HPO|Glucosuria|Glucosuria
C0804101|T201|MTH_LN|21307-4|LNC2HPO|Glucosuria|Glucosuria
C0804101|T201|DN|21307-4|LNC2HPO|Glucosuria|Glucosuria
C0804101|T201|OSN|21307-4|LNC2HPO|Glucosuria|Glucosuria
C0804101|T201|LC|21307-4|LNC2HPO|Glucosuria|Glucosuria
C0803801|T201|MTH_LN|21004-7|LNC2HPO|Glucose intolerance|Glucose intolerance
C0803801|T201|LN|21004-7|LNC2HPO|Glucose intolerance|Glucose intolerance
C0803801|T201|DN|21004-7|LNC2HPO|Glucose intolerance|Glucose intolerance
C0803801|T201|OSN|21004-7|LNC2HPO|Glucose intolerance|Glucose intolerance
C0803801|T201|LC|21004-7|LNC2HPO|Glucose intolerance|Glucose intolerance
C0803801|T201|MTH_LN|21004-7|LNC2HPO|Impaired glucose tolerance|Impaired glucose tolerance
C0803801|T201|LN|21004-7|LNC2HPO|Impaired glucose tolerance|Impaired glucose tolerance
C0803801|T201|DN|21004-7|LNC2HPO|Impaired glucose tolerance|Impaired glucose tolerance
C0803801|T201|OSN|21004-7|LNC2HPO|Impaired glucose tolerance|Impaired glucose tolerance
C0803801|T201|LC|21004-7|LNC2HPO|Impaired glucose tolerance|Impaired glucose tolerance
C0880214|T201|LN|22705-8|LNC2HPO|Glycosuria|Glycosuria
C0880214|T201|DN|22705-8|LNC2HPO|Glycosuria|Glycosuria
C0880214|T201|MTH_LN|22705-8|LNC2HPO|Glycosuria|Glycosuria
C0880214|T201|OSN|22705-8|LNC2HPO|Glycosuria|Glycosuria
C0880214|T201|LC|22705-8|LNC2HPO|Glycosuria|Glycosuria
C0880214|T201|LN|22705-8|LNC2HPO|Glucosuria|Glucosuria
C0880214|T201|DN|22705-8|LNC2HPO|Glucosuria|Glucosuria
C0880214|T201|MTH_LN|22705-8|LNC2HPO|Glucosuria|Glucosuria
C0880214|T201|OSN|22705-8|LNC2HPO|Glucosuria|Glucosuria
C0880214|T201|LC|22705-8|LNC2HPO|Glucosuria|Glucosuria
C0364491|T201|LN|2351-5|LNC2HPO|Glycosuria|Glycosuria
C0364491|T201|MTH_LN|2351-5|LNC2HPO|Glycosuria|Glycosuria
C0364491|T201|DN|2351-5|LNC2HPO|Glycosuria|Glycosuria
C0364491|T201|OSN|2351-5|LNC2HPO|Glycosuria|Glycosuria
C0364491|T201|LC|2351-5|LNC2HPO|Glycosuria|Glycosuria
C0364491|T201|LN|2351-5|LNC2HPO|Glucosuria|Glucosuria
C0364491|T201|MTH_LN|2351-5|LNC2HPO|Glucosuria|Glucosuria
C0364491|T201|DN|2351-5|LNC2HPO|Glucosuria|Glucosuria
C0364491|T201|OSN|2351-5|LNC2HPO|Glucosuria|Glucosuria
C0364491|T201|LC|2351-5|LNC2HPO|Glucosuria|Glucosuria
C0550203|T201|LN|12177-2|LNC2HPO|Aminoaciduria|Aminoaciduria
C0550203|T201|MTH_LN|12177-2|LNC2HPO|Aminoaciduria|Aminoaciduria
C0550203|T201|DN|12177-2|LNC2HPO|Aminoaciduria|Aminoaciduria
C0550203|T201|OSN|12177-2|LNC2HPO|Aminoaciduria|Aminoaciduria
C0550203|T201|LC|12177-2|LNC2HPO|Aminoaciduria|Aminoaciduria
C0550203|T201|LN|12177-2|LNC2HPO|Hyperaminoaciduria|Hyperaminoaciduria
C0550203|T201|MTH_LN|12177-2|LNC2HPO|Hyperaminoaciduria|Hyperaminoaciduria
C0550203|T201|DN|12177-2|LNC2HPO|Hyperaminoaciduria|Hyperaminoaciduria
C0550203|T201|OSN|12177-2|LNC2HPO|Hyperaminoaciduria|Hyperaminoaciduria
C0550203|T201|LC|12177-2|LNC2HPO|Hyperaminoaciduria|Hyperaminoaciduria
C0550202|T201|LN|12467-7|LNC2HPO|Aminoaciduria|Aminoaciduria
C0550202|T201|MTH_LN|12467-7|LNC2HPO|Aminoaciduria|Aminoaciduria
C0550202|T201|DN|12467-7|LNC2HPO|Aminoaciduria|Aminoaciduria
C0550202|T201|OSN|12467-7|LNC2HPO|Aminoaciduria|Aminoaciduria
C0550202|T201|LC|12467-7|LNC2HPO|Aminoaciduria|Aminoaciduria
C0550202|T201|LN|12467-7|LNC2HPO|Hyperaminoaciduria|Hyperaminoaciduria
C0550202|T201|MTH_LN|12467-7|LNC2HPO|Hyperaminoaciduria|Hyperaminoaciduria
C0550202|T201|DN|12467-7|LNC2HPO|Hyperaminoaciduria|Hyperaminoaciduria
C0550202|T201|OSN|12467-7|LNC2HPO|Hyperaminoaciduria|Hyperaminoaciduria
C0550202|T201|LC|12467-7|LNC2HPO|Hyperaminoaciduria|Hyperaminoaciduria
C0801239|T201|LN|18191-7|LNC2HPO|Aminoaciduria|Aminoaciduria
C0801239|T201|MTH_LN|18191-7|LNC2HPO|Aminoaciduria|Aminoaciduria
C0801239|T201|DN|18191-7|LNC2HPO|Aminoaciduria|Aminoaciduria
C0801239|T201|OSN|18191-7|LNC2HPO|Aminoaciduria|Aminoaciduria
C0801239|T201|LC|18191-7|LNC2HPO|Aminoaciduria|Aminoaciduria
C0801239|T201|LN|18191-7|LNC2HPO|Hyperaminoaciduria|Hyperaminoaciduria
C0801239|T201|MTH_LN|18191-7|LNC2HPO|Hyperaminoaciduria|Hyperaminoaciduria
C0801239|T201|DN|18191-7|LNC2HPO|Hyperaminoaciduria|Hyperaminoaciduria
C0801239|T201|OSN|18191-7|LNC2HPO|Hyperaminoaciduria|Hyperaminoaciduria
C0801239|T201|LC|18191-7|LNC2HPO|Hyperaminoaciduria|Hyperaminoaciduria
C0367978|T201|LN|5763-8|LNC2HPO|Hyperzincemia|Hyperzincemia
C0367978|T201|DN|5763-8|LNC2HPO|Hyperzincemia|Hyperzincemia
C0367978|T201|MTH_LN|5763-8|LNC2HPO|Hyperzincemia|Hyperzincemia
C0367978|T201|OSN|5763-8|LNC2HPO|Hyperzincemia|Hyperzincemia
C0367978|T201|LC|5763-8|LNC2HPO|Hyperzincemia|Hyperzincemia
C1114053|T201|LN|30166-3|LNC2HPO|TSH excess|TSH excess
C1114053|T201|DN|30166-3|LNC2HPO|TSH excess|TSH excess
C1114053|T201|MTH_LN|30166-3|LNC2HPO|TSH excess|TSH excess
C1114053|T201|OSN|30166-3|LNC2HPO|TSH excess|TSH excess
C1114053|T201|LC|30166-3|LNC2HPO|TSH excess|TSH excess
C1114402|T201|LN|30567-2|LNC2HPO|TSH excess|TSH excess
C1114402|T201|DN|30567-2|LNC2HPO|TSH excess|TSH excess
C1114402|T201|MTH_LN|30567-2|LNC2HPO|TSH excess|TSH excess
C1114402|T201|OSN|30567-2|LNC2HPO|TSH excess|TSH excess
C1114402|T201|LC|30567-2|LNC2HPO|TSH excess|TSH excess
C0485076|T201|LN|10613-8|LNC2HPO|Impaired spermatogenesis|Impaired spermatogenesis
C0485076|T201|DN|10613-8|LNC2HPO|Impaired spermatogenesis|Impaired spermatogenesis
C0485076|T201|MTH_LN|10613-8|LNC2HPO|Impaired spermatogenesis|Impaired spermatogenesis
C0485076|T201|LC|10613-8|LNC2HPO|Impaired spermatogenesis|Impaired spermatogenesis
C0485076|T201|OSN|10613-8|LNC2HPO|Impaired spermatogenesis|Impaired spermatogenesis
C0485076|T201|LN|10613-8|LNC2HPO|Oligospermia|Oligospermia
C0485076|T201|DN|10613-8|LNC2HPO|Oligospermia|Oligospermia
C0485076|T201|MTH_LN|10613-8|LNC2HPO|Oligospermia|Oligospermia
C0485076|T201|LC|10613-8|LNC2HPO|Oligospermia|Oligospermia
C0485076|T201|OSN|10613-8|LNC2HPO|Oligospermia|Oligospermia
C1315188|T201|LN|32717-1|LNC2HPO|Hypernatremia|Hypernatremia
C1315188|T201|DN|32717-1|LNC2HPO|Hypernatremia|Hypernatremia
C1315188|T201|MTH_LN|32717-1|LNC2HPO|Hypernatremia|Hypernatremia
C1315188|T201|OSN|32717-1|LNC2HPO|Hypernatremia|Hypernatremia
C1315188|T201|LC|32717-1|LNC2HPO|Hypernatremia|Hypernatremia
C1315188|T201|LN|32717-1|LNC2HPO|Hyponatremia|Hyponatremia
C1315188|T201|DN|32717-1|LNC2HPO|Hyponatremia|Hyponatremia
C1315188|T201|MTH_LN|32717-1|LNC2HPO|Hyponatremia|Hyponatremia
C1315188|T201|OSN|32717-1|LNC2HPO|Hyponatremia|Hyponatremia
C1315188|T201|LC|32717-1|LNC2HPO|Hyponatremia|Hyponatremia
C0804319|T201|LN|21525-1|LNC2HPO|Hypernatriuria|Hypernatriuria
C0804319|T201|MTH_LN|21525-1|LNC2HPO|Hypernatriuria|Hypernatriuria
C0804319|T201|DN|21525-1|LNC2HPO|Hypernatriuria|Hypernatriuria
C0804319|T201|OSN|21525-1|LNC2HPO|Hypernatriuria|Hypernatriuria
C0804319|T201|LC|21525-1|LNC2HPO|Hypernatriuria|Hypernatriuria
C0804319|T201|LN|21525-1|LNC2HPO|Hyponatriuria|Hyponatriuria
C0804319|T201|MTH_LN|21525-1|LNC2HPO|Hyponatriuria|Hyponatriuria
C0804319|T201|DN|21525-1|LNC2HPO|Hyponatriuria|Hyponatriuria
C0804319|T201|OSN|21525-1|LNC2HPO|Hyponatriuria|Hyponatriuria
C0804319|T201|LC|21525-1|LNC2HPO|Hyponatriuria|Hyponatriuria
C0364097|T201|LN|1964-6|LNC2HPO|Bicarbonaturia|Bicarbonaturia
C0364097|T201|MTH_LN|1964-6|LNC2HPO|Bicarbonaturia|Bicarbonaturia
C0364097|T201|DN|1964-6|LNC2HPO|Bicarbonaturia|Bicarbonaturia
C0364097|T201|OSN|1964-6|LNC2HPO|Bicarbonaturia|Bicarbonaturia
C0364097|T201|LC|1964-6|LNC2HPO|Bicarbonaturia|Bicarbonaturia
C1952809|T201|LN|47579-8|LNC2HPO|Bicarbonaturia|Bicarbonaturia
C1952809|T201|DN|47579-8|LNC2HPO|Bicarbonaturia|Bicarbonaturia
C1952809|T201|MTH_LN|47579-8|LNC2HPO|Bicarbonaturia|Bicarbonaturia
C1952809|T201|OSN|47579-8|LNC2HPO|Bicarbonaturia|Bicarbonaturia
C1952809|T201|LC|47579-8|LNC2HPO|Bicarbonaturia|Bicarbonaturia
C1952810|T201|LN|47580-6|LNC2HPO|Bicarbonaturia|Bicarbonaturia
C1952810|T201|DN|47580-6|LNC2HPO|Bicarbonaturia|Bicarbonaturia
C1952810|T201|OSN|47580-6|LNC2HPO|Bicarbonaturia|Bicarbonaturia
C1952810|T201|MTH_LN|47580-6|LNC2HPO|Bicarbonaturia|Bicarbonaturia
C1952810|T201|LC|47580-6|LNC2HPO|Bicarbonaturia|Bicarbonaturia
C0485074|T201|LN|10611-2|LNC2HPO|Asthenospermia|Asthenospermia
C0485074|T201|MTH_LN|10611-2|LNC2HPO|Asthenospermia|Asthenospermia
C0485074|T201|DN|10611-2|LNC2HPO|Asthenospermia|Asthenospermia
C0485074|T201|LC|10611-2|LNC2HPO|Asthenospermia|Asthenospermia
C0485074|T201|OSN|10611-2|LNC2HPO|Asthenospermia|Asthenospermia
C0803455|T201|LN|20651-6|LNC2HPO|Hypermethioninemia|Hypermethioninemia
C0803455|T201|MTH_LN|20651-6|LNC2HPO|Hypermethioninemia|Hypermethioninemia
C0803455|T201|DN|20651-6|LNC2HPO|Hypermethioninemia|Hypermethioninemia
C0803455|T201|OSN|20651-6|LNC2HPO|Hypermethioninemia|Hypermethioninemia
C0803455|T201|LC|20651-6|LNC2HPO|Hypermethioninemia|Hypermethioninemia
C0803455|T201|LN|20651-6|LNC2HPO|Methioninemia|Methioninemia
C0803455|T201|MTH_LN|20651-6|LNC2HPO|Methioninemia|Methioninemia
C0803455|T201|DN|20651-6|LNC2HPO|Methioninemia|Methioninemia
C0803455|T201|OSN|20651-6|LNC2HPO|Methioninemia|Methioninemia
C0803455|T201|LC|20651-6|LNC2HPO|Methioninemia|Methioninemia
C0803455|T201|LN|20651-6|LNC2HPO|Hypomethioninemia|Hypomethioninemia
C0803455|T201|MTH_LN|20651-6|LNC2HPO|Hypomethioninemia|Hypomethioninemia
C0803455|T201|DN|20651-6|LNC2HPO|Hypomethioninemia|Hypomethioninemia
C0803455|T201|OSN|20651-6|LNC2HPO|Hypomethioninemia|Hypomethioninemia
C0803455|T201|LC|20651-6|LNC2HPO|Hypomethioninemia|Hypomethioninemia
C0803448|T201|LN|20644-1|LNC2HPO|Hyperglycinemia|Hyperglycinemia
C0803448|T201|MTH_LN|20644-1|LNC2HPO|Hyperglycinemia|Hyperglycinemia
C0803448|T201|DN|20644-1|LNC2HPO|Hyperglycinemia|Hyperglycinemia
C0803448|T201|OSN|20644-1|LNC2HPO|Hyperglycinemia|Hyperglycinemia
C0803448|T201|LC|20644-1|LNC2HPO|Hyperglycinemia|Hyperglycinemia
C0803448|T201|LN|20644-1|LNC2HPO|Hyperglycinaemia|Hyperglycinaemia
C0803448|T201|MTH_LN|20644-1|LNC2HPO|Hyperglycinaemia|Hyperglycinaemia
C0803448|T201|DN|20644-1|LNC2HPO|Hyperglycinaemia|Hyperglycinaemia
C0803448|T201|OSN|20644-1|LNC2HPO|Hyperglycinaemia|Hyperglycinaemia
C0803448|T201|LC|20644-1|LNC2HPO|Hyperglycinaemia|Hyperglycinaemia
C0803448|T201|LN|20644-1|LNC2HPO|Hypoglycinemia|Hypoglycinemia
C0803448|T201|MTH_LN|20644-1|LNC2HPO|Hypoglycinemia|Hypoglycinemia
C0803448|T201|DN|20644-1|LNC2HPO|Hypoglycinemia|Hypoglycinemia
C0803448|T201|OSN|20644-1|LNC2HPO|Hypoglycinemia|Hypoglycinemia
C0803448|T201|LC|20644-1|LNC2HPO|Hypoglycinemia|Hypoglycinemia
C0942549|T201|LN|26607-2|LNC2HPO|Cystathioninemia|Cystathioninemia
C0942549|T201|DN|26607-2|LNC2HPO|Cystathioninemia|Cystathioninemia
C0942549|T201|MTH_LN|26607-2|LNC2HPO|Cystathioninemia|Cystathioninemia
C0942549|T201|OSN|26607-2|LNC2HPO|Cystathioninemia|Cystathioninemia
C0942549|T201|LC|26607-2|LNC2HPO|Cystathioninemia|Cystathioninemia
C0364133|T201|LN|2000-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C0364133|T201|MTH_LN|2000-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C0364133|T201|DN|2000-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C0364133|T201|OSN|2000-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C0364133|T201|LC|2000-8|LNC2HPO|Hypercalcemia|Hypercalcemia
C0364133|T201|LN|2000-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0364133|T201|MTH_LN|2000-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0364133|T201|DN|2000-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0364133|T201|OSN|2000-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0364133|T201|LC|2000-8|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0364133|T201|LN|2000-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C0364133|T201|MTH_LN|2000-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C0364133|T201|DN|2000-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C0364133|T201|OSN|2000-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C0364133|T201|LC|2000-8|LNC2HPO|Hypocalcemia|Hypocalcemia
C0364133|T201|LN|2000-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364133|T201|MTH_LN|2000-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364133|T201|DN|2000-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364133|T201|OSN|2000-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364133|T201|LC|2000-8|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0362894|T201|LN|706-2|LNC2HPO|Basophilia|Basophilia
C0362894|T201|MTH_LN|706-2|LNC2HPO|Basophilia|Basophilia
C0362894|T201|OSN|706-2|LNC2HPO|Basophilia|Basophilia
C0362894|T201|DN|706-2|LNC2HPO|Basophilia|Basophilia
C0362894|T201|LC|706-2|LNC2HPO|Basophilia|Basophilia
C0362960|T201|LN|5905-5|LNC2HPO|Monocytosis|Monocytosis
C0362960|T201|MTH_LN|5905-5|LNC2HPO|Monocytosis|Monocytosis
C0362960|T201|OSN|5905-5|LNC2HPO|Monocytosis|Monocytosis
C0362960|T201|DN|5905-5|LNC2HPO|Monocytosis|Monocytosis
C0362960|T201|LC|5905-5|LNC2HPO|Monocytosis|Monocytosis
C0362960|T201|LN|5905-5|LNC2HPO|Monocytopenia|Monocytopenia
C0362960|T201|MTH_LN|5905-5|LNC2HPO|Monocytopenia|Monocytopenia
C0362960|T201|OSN|5905-5|LNC2HPO|Monocytopenia|Monocytopenia
C0362960|T201|DN|5905-5|LNC2HPO|Monocytopenia|Monocytopenia
C0362960|T201|LC|5905-5|LNC2HPO|Monocytopenia|Monocytopenia
C1315725|T201|LN|33256-9|LNC2HPO|Leukocytosis|Leukocytosis
C1315725|T201|DN|33256-9|LNC2HPO|Leukocytosis|Leukocytosis
C1315725|T201|OSN|33256-9|LNC2HPO|Leukocytosis|Leukocytosis
C1315725|T201|MTH_LN|33256-9|LNC2HPO|Leukocytosis|Leukocytosis
C1315725|T201|LC|33256-9|LNC2HPO|Leukocytosis|Leukocytosis
C1315725|T201|LN|33256-9|LNC2HPO|Leukopenia|Leukopenia
C1315725|T201|DN|33256-9|LNC2HPO|Leukopenia|Leukopenia
C1315725|T201|OSN|33256-9|LNC2HPO|Leukopenia|Leukopenia
C1315725|T201|MTH_LN|33256-9|LNC2HPO|Leukopenia|Leukopenia
C1315725|T201|LC|33256-9|LNC2HPO|Leukopenia|Leukopenia
C0362961|T201|LN|744-3|LNC2HPO|Monocytosis|Monocytosis
C0362961|T201|MTH_LN|744-3|LNC2HPO|Monocytosis|Monocytosis
C0362961|T201|OSN|744-3|LNC2HPO|Monocytosis|Monocytosis
C0362961|T201|DN|744-3|LNC2HPO|Monocytosis|Monocytosis
C0362961|T201|LC|744-3|LNC2HPO|Monocytosis|Monocytosis
C0362961|T201|LN|744-3|LNC2HPO|Monocytopenia|Monocytopenia
C0362961|T201|MTH_LN|744-3|LNC2HPO|Monocytopenia|Monocytopenia
C0362961|T201|OSN|744-3|LNC2HPO|Monocytopenia|Monocytopenia
C0362961|T201|DN|744-3|LNC2HPO|Monocytopenia|Monocytopenia
C0362961|T201|LC|744-3|LNC2HPO|Monocytopenia|Monocytopenia
C0362952|T201|LN|736-9|LNC2HPO|Lymphocytosis|Lymphocytosis
C0362952|T201|MTH_LN|736-9|LNC2HPO|Lymphocytosis|Lymphocytosis
C0362952|T201|OSN|736-9|LNC2HPO|Lymphocytosis|Lymphocytosis
C0362952|T201|DN|736-9|LNC2HPO|Lymphocytosis|Lymphocytosis
C0362952|T201|LC|736-9|LNC2HPO|Lymphocytosis|Lymphocytosis
C0362952|T201|LN|736-9|LNC2HPO|Lymphopenia|Lymphopenia
C0362952|T201|MTH_LN|736-9|LNC2HPO|Lymphopenia|Lymphopenia
C0362952|T201|OSN|736-9|LNC2HPO|Lymphopenia|Lymphopenia
C0362952|T201|DN|736-9|LNC2HPO|Lymphopenia|Lymphopenia
C0362952|T201|LC|736-9|LNC2HPO|Lymphopenia|Lymphopenia
C0362952|T201|LN|736-9|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0362952|T201|MTH_LN|736-9|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0362952|T201|OSN|736-9|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0362952|T201|DN|736-9|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0362952|T201|LC|736-9|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0362952|T201|LN|736-9|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0362952|T201|MTH_LN|736-9|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0362952|T201|OSN|736-9|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0362952|T201|DN|736-9|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0362952|T201|LC|736-9|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0362953|T201|LN|737-7|LNC2HPO|Lymphocytosis|Lymphocytosis
C0362953|T201|MTH_LN|737-7|LNC2HPO|Lymphocytosis|Lymphocytosis
C0362953|T201|OSN|737-7|LNC2HPO|Lymphocytosis|Lymphocytosis
C0362953|T201|DN|737-7|LNC2HPO|Lymphocytosis|Lymphocytosis
C0362953|T201|LC|737-7|LNC2HPO|Lymphocytosis|Lymphocytosis
C0362953|T201|LN|737-7|LNC2HPO|Lymphopenia|Lymphopenia
C0362953|T201|MTH_LN|737-7|LNC2HPO|Lymphopenia|Lymphopenia
C0362953|T201|OSN|737-7|LNC2HPO|Lymphopenia|Lymphopenia
C0362953|T201|DN|737-7|LNC2HPO|Lymphopenia|Lymphopenia
C0362953|T201|LC|737-7|LNC2HPO|Lymphopenia|Lymphopenia
C0362953|T201|LN|737-7|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0362953|T201|MTH_LN|737-7|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0362953|T201|OSN|737-7|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0362953|T201|DN|737-7|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0362953|T201|LC|737-7|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0362953|T201|LN|737-7|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0362953|T201|MTH_LN|737-7|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0362953|T201|OSN|737-7|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0362953|T201|DN|737-7|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0362953|T201|LC|737-7|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0364481|T201|LN|2341-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0364481|T201|MTH_LN|2341-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0364481|T201|DN|2341-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0364481|T201|OSN|2341-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0364481|T201|LC|2341-6|LNC2HPO|Hyperglycemia|Hyperglycemia
C0364481|T201|LN|2341-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0364481|T201|MTH_LN|2341-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0364481|T201|DN|2341-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0364481|T201|OSN|2341-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0364481|T201|LC|2341-6|LNC2HPO|Hypoglycemia|Hypoglycemia
C0364481|T201|LN|2341-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0364481|T201|MTH_LN|2341-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0364481|T201|DN|2341-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0364481|T201|OSN|2341-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0364481|T201|LC|2341-6|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0365405|T201|LN|5964-2|LNC2HPO|Prolonged prothrombin time|Prolonged prothrombin time
C0365405|T201|DN|5964-2|LNC2HPO|Prolonged prothrombin time|Prolonged prothrombin time
C0365405|T201|MTH_LN|5964-2|LNC2HPO|Prolonged prothrombin time|Prolonged prothrombin time
C0365405|T201|OSN|5964-2|LNC2HPO|Prolonged prothrombin time|Prolonged prothrombin time
C0365405|T201|LC|5964-2|LNC2HPO|Prolonged prothrombin time|Prolonged prothrombin time
C0365405|T201|LN|5964-2|LNC2HPO|Prolonged PT|Prolonged PT
C0365405|T201|DN|5964-2|LNC2HPO|Prolonged PT|Prolonged PT
C0365405|T201|MTH_LN|5964-2|LNC2HPO|Prolonged PT|Prolonged PT
C0365405|T201|OSN|5964-2|LNC2HPO|Prolonged PT|Prolonged PT
C0365405|T201|LC|5964-2|LNC2HPO|Prolonged PT|Prolonged PT
C0365405|T201|LN|5964-2|LNC2HPO|increased international normalised ratio|increased international normalised ratio
C0365405|T201|DN|5964-2|LNC2HPO|increased international normalised ratio|increased international normalised ratio
C0365405|T201|MTH_LN|5964-2|LNC2HPO|increased international normalised ratio|increased international normalised ratio
C0365405|T201|OSN|5964-2|LNC2HPO|increased international normalised ratio|increased international normalised ratio
C0365405|T201|LC|5964-2|LNC2HPO|increased international normalised ratio|increased international normalised ratio
C0550431|T201|LN|11147-6|LNC2HPO|Myoglobinuria|Myoglobinuria
C0550431|T201|MTH_LN|11147-6|LNC2HPO|Myoglobinuria|Myoglobinuria
C0550431|T201|OSN|11147-6|LNC2HPO|Myoglobinuria|Myoglobinuria
C0550431|T201|DN|11147-6|LNC2HPO|Myoglobinuria|Myoglobinuria
C0550431|T201|LC|11147-6|LNC2HPO|Myoglobinuria|Myoglobinuria
C0550473|T201|LN|11148-4|LNC2HPO|Hyperkaliuresis|Hyperkaliuresis
C0550473|T201|OSN|11148-4|LNC2HPO|Hyperkaliuresis|Hyperkaliuresis
C0550473|T201|MTH_LN|11148-4|LNC2HPO|Hyperkaliuresis|Hyperkaliuresis
C0550473|T201|DN|11148-4|LNC2HPO|Hyperkaliuresis|Hyperkaliuresis
C0550473|T201|LC|11148-4|LNC2HPO|Hyperkaliuresis|Hyperkaliuresis
C0550473|T201|LN|11148-4|LNC2HPO|Hypokaluria|Hypokaluria
C0550473|T201|OSN|11148-4|LNC2HPO|Hypokaluria|Hypokaluria
C0550473|T201|MTH_LN|11148-4|LNC2HPO|Hypokaluria|Hypokaluria
C0550473|T201|DN|11148-4|LNC2HPO|Hypokaluria|Hypokaluria
C0550473|T201|LC|11148-4|LNC2HPO|Hypokaluria|Hypokaluria
C0550513|T201|LN|11149-2|LNC2HPO|Hyponatriuria|Hyponatriuria
C0550513|T201|MTH_LN|11149-2|LNC2HPO|Hyponatriuria|Hyponatriuria
C0550513|T201|OSN|11149-2|LNC2HPO|Hyponatriuria|Hyponatriuria
C0550513|T201|DN|11149-2|LNC2HPO|Hyponatriuria|Hyponatriuria
C0550513|T201|LC|11149-2|LNC2HPO|Hyponatriuria|Hyponatriuria
C0362933|T201|LN|728-6|LNC2HPO|Hypochromic anemia|Hypochromic anemia
C0362933|T201|MTH_LN|728-6|LNC2HPO|Hypochromic anemia|Hypochromic anemia
C0362933|T201|DN|728-6|LNC2HPO|Hypochromic anemia|Hypochromic anemia
C0362933|T201|OSN|728-6|LNC2HPO|Hypochromic anemia|Hypochromic anemia
C0362933|T201|LC|728-6|LNC2HPO|Hypochromic anemia|Hypochromic anemia
C0362933|T201|LN|728-6|LNC2HPO|Hypochromic anaemia|Hypochromic anaemia
C0362933|T201|MTH_LN|728-6|LNC2HPO|Hypochromic anaemia|Hypochromic anaemia
C0362933|T201|DN|728-6|LNC2HPO|Hypochromic anaemia|Hypochromic anaemia
C0362933|T201|OSN|728-6|LNC2HPO|Hypochromic anaemia|Hypochromic anaemia
C0362933|T201|LC|728-6|LNC2HPO|Hypochromic anaemia|Hypochromic anaemia
C0797497|T201|LN|14316-4|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0797497|T201|MTH_LN|14316-4|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0797497|T201|DN|14316-4|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0797497|T201|OSN|14316-4|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0797497|T201|LC|14316-4|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0799360|T201|LN|16195-0|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0799360|T201|LC|16195-0|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0799360|T201|MTH_LN|16195-0|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0799360|T201|DN|16195-0|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0799360|T201|OSN|16195-0|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802252|T201|LN|19359-9|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802252|T201|MTH_LN|19359-9|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802252|T201|DN|19359-9|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802252|T201|OSN|19359-9|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802252|T201|LC|19359-9|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C2361846|T201|MTH_LN|53326-5|LNC2HPO|Urine issues|Urine issues
C2361846|T201|DN|53326-5|LNC2HPO|Urine issues|Urine issues
C2361846|T201|LN|53326-5|LNC2HPO|Urine issues|Urine issues
C2361846|T201|OSN|53326-5|LNC2HPO|Urine issues|Urine issues
C2361846|T201|LC|53326-5|LNC2HPO|Urine issues|Urine issues
C2361846|T201|MTH_LN|53326-5|LNC2HPO|Pee issues|Pee issues
C2361846|T201|DN|53326-5|LNC2HPO|Pee issues|Pee issues
C2361846|T201|LN|53326-5|LNC2HPO|Pee issues|Pee issues
C2361846|T201|OSN|53326-5|LNC2HPO|Pee issues|Pee issues
C2361846|T201|LC|53326-5|LNC2HPO|Pee issues|Pee issues
C2361846|T201|MTH_LN|53326-5|LNC2HPO|Hyposthenuria|Hyposthenuria
C2361846|T201|DN|53326-5|LNC2HPO|Hyposthenuria|Hyposthenuria
C2361846|T201|LN|53326-5|LNC2HPO|Hyposthenuria|Hyposthenuria
C2361846|T201|OSN|53326-5|LNC2HPO|Hyposthenuria|Hyposthenuria
C2361846|T201|LC|53326-5|LNC2HPO|Hyposthenuria|Hyposthenuria
C0364101|T201|LC|1968-7|LNC2HPO|Hyperbilirubinemia|Hyperbilirubinemia
C0364101|T201|DN|1968-7|LNC2HPO|Hyperbilirubinemia|Hyperbilirubinemia
C0364101|T201|MTH_LN|1968-7|LNC2HPO|Hyperbilirubinemia|Hyperbilirubinemia
C0364101|T201|LN|1968-7|LNC2HPO|Hyperbilirubinemia|Hyperbilirubinemia
C0364101|T201|OSN|1968-7|LNC2HPO|Hyperbilirubinemia|Hyperbilirubinemia
C0364275|T201|LC|2143-6|LNC2HPO|Cushing syndrome|Cushing syndrome
C0364275|T201|LN|2143-6|LNC2HPO|Cushing syndrome|Cushing syndrome
C0364275|T201|MTH_LN|2143-6|LNC2HPO|Cushing syndrome|Cushing syndrome
C0364275|T201|DN|2143-6|LNC2HPO|Cushing syndrome|Cushing syndrome
C0364275|T201|OSN|2143-6|LNC2HPO|Cushing syndrome|Cushing syndrome
C0364275|T201|LC|2143-6|LNC2HPO|Hypercortisolism|Hypercortisolism
C0364275|T201|LN|2143-6|LNC2HPO|Hypercortisolism|Hypercortisolism
C0364275|T201|MTH_LN|2143-6|LNC2HPO|Hypercortisolism|Hypercortisolism
C0364275|T201|DN|2143-6|LNC2HPO|Hypercortisolism|Hypercortisolism
C0364275|T201|OSN|2143-6|LNC2HPO|Hypercortisolism|Hypercortisolism
C0364275|T201|LC|2143-6|LNC2HPO|Hypocortisolism|Hypocortisolism
C0364275|T201|LN|2143-6|LNC2HPO|Hypocortisolism|Hypocortisolism
C0364275|T201|MTH_LN|2143-6|LNC2HPO|Hypocortisolism|Hypocortisolism
C0364275|T201|DN|2143-6|LNC2HPO|Hypocortisolism|Hypocortisolism
C0364275|T201|OSN|2143-6|LNC2HPO|Hypocortisolism|Hypocortisolism
C0364275|T201|LC|2143-6|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0364275|T201|LN|2143-6|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0364275|T201|MTH_LN|2143-6|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0364275|T201|DN|2143-6|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0364275|T201|OSN|2143-6|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0364275|T201|LC|2143-6|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0364275|T201|LN|2143-6|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0364275|T201|MTH_LN|2143-6|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0364275|T201|DN|2143-6|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0364275|T201|OSN|2143-6|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0551356|T201|LN|11572-5|LNC2HPO|Rheumatoid factor positive|Rheumatoid factor positive
C0551356|T201|LC|11572-5|LNC2HPO|Rheumatoid factor positive|Rheumatoid factor positive
C0551356|T201|OSN|11572-5|LNC2HPO|Rheumatoid factor positive|Rheumatoid factor positive
C0551356|T201|MTH_LN|11572-5|LNC2HPO|Rheumatoid factor positive|Rheumatoid factor positive
C0551356|T201|DN|11572-5|LNC2HPO|Rheumatoid factor positive|Rheumatoid factor positive
C0364971|T201|LN|2828-2|LNC2HPO|Hyperkaliuresis|Hyperkaliuresis
C0364971|T201|MTH_LN|2828-2|LNC2HPO|Hyperkaliuresis|Hyperkaliuresis
C0364971|T201|DN|2828-2|LNC2HPO|Hyperkaliuresis|Hyperkaliuresis
C0364971|T201|OSN|2828-2|LNC2HPO|Hyperkaliuresis|Hyperkaliuresis
C0364971|T201|LC|2828-2|LNC2HPO|Hyperkaliuresis|Hyperkaliuresis
C0365111|T201|MTH_LN|2965-2|LNC2HPO|Urine issues|Urine issues
C0365111|T201|LC|2965-2|LNC2HPO|Urine issues|Urine issues
C0365111|T201|DN|2965-2|LNC2HPO|Urine issues|Urine issues
C0365111|T201|LN|2965-2|LNC2HPO|Urine issues|Urine issues
C0365111|T201|OSN|2965-2|LNC2HPO|Urine issues|Urine issues
C0365111|T201|MTH_LN|2965-2|LNC2HPO|Pee issues|Pee issues
C0365111|T201|LC|2965-2|LNC2HPO|Pee issues|Pee issues
C0365111|T201|DN|2965-2|LNC2HPO|Pee issues|Pee issues
C0365111|T201|LN|2965-2|LNC2HPO|Pee issues|Pee issues
C0365111|T201|OSN|2965-2|LNC2HPO|Pee issues|Pee issues
C0365111|T201|MTH_LN|2965-2|LNC2HPO|Hyposthenuria|Hyposthenuria
C0365111|T201|LC|2965-2|LNC2HPO|Hyposthenuria|Hyposthenuria
C0365111|T201|DN|2965-2|LNC2HPO|Hyposthenuria|Hyposthenuria
C0365111|T201|LN|2965-2|LNC2HPO|Hyposthenuria|Hyposthenuria
C0365111|T201|OSN|2965-2|LNC2HPO|Hyposthenuria|Hyposthenuria
C0365110|T201|LN|2966-0|LNC2HPO|Urine issues|Urine issues
C0365110|T201|MTH_LN|2966-0|LNC2HPO|Urine issues|Urine issues
C0365110|T201|DN|2966-0|LNC2HPO|Urine issues|Urine issues
C0365110|T201|OSN|2966-0|LNC2HPO|Urine issues|Urine issues
C0365110|T201|LC|2966-0|LNC2HPO|Urine issues|Urine issues
C0365110|T201|LN|2966-0|LNC2HPO|Pee issues|Pee issues
C0365110|T201|MTH_LN|2966-0|LNC2HPO|Pee issues|Pee issues
C0365110|T201|DN|2966-0|LNC2HPO|Pee issues|Pee issues
C0365110|T201|OSN|2966-0|LNC2HPO|Pee issues|Pee issues
C0365110|T201|LC|2966-0|LNC2HPO|Pee issues|Pee issues
C0365110|T201|LN|2966-0|LNC2HPO|Hyposthenuria|Hyposthenuria
C0365110|T201|MTH_LN|2966-0|LNC2HPO|Hyposthenuria|Hyposthenuria
C0365110|T201|DN|2966-0|LNC2HPO|Hyposthenuria|Hyposthenuria
C0365110|T201|OSN|2966-0|LNC2HPO|Hyposthenuria|Hyposthenuria
C0365110|T201|LC|2966-0|LNC2HPO|Hyposthenuria|Hyposthenuria
C1716137|T201|LN|44933-0|LNC2HPO|Urine issues|Urine issues
C1716137|T201|DN|44933-0|LNC2HPO|Urine issues|Urine issues
C1716137|T201|MTH_LN|44933-0|LNC2HPO|Urine issues|Urine issues
C1716137|T201|OSN|44933-0|LNC2HPO|Urine issues|Urine issues
C1716137|T201|LC|44933-0|LNC2HPO|Urine issues|Urine issues
C1716137|T201|LN|44933-0|LNC2HPO|Pee issues|Pee issues
C1716137|T201|DN|44933-0|LNC2HPO|Pee issues|Pee issues
C1716137|T201|MTH_LN|44933-0|LNC2HPO|Pee issues|Pee issues
C1716137|T201|OSN|44933-0|LNC2HPO|Pee issues|Pee issues
C1716137|T201|LC|44933-0|LNC2HPO|Pee issues|Pee issues
C1716137|T201|LN|44933-0|LNC2HPO|Hyposthenuria|Hyposthenuria
C1716137|T201|DN|44933-0|LNC2HPO|Hyposthenuria|Hyposthenuria
C1716137|T201|MTH_LN|44933-0|LNC2HPO|Hyposthenuria|Hyposthenuria
C1716137|T201|OSN|44933-0|LNC2HPO|Hyposthenuria|Hyposthenuria
C1716137|T201|LC|44933-0|LNC2HPO|Hyposthenuria|Hyposthenuria
C1977831|T201|LN|49959-0|LNC2HPO|Urine issues|Urine issues
C1977831|T201|DN|49959-0|LNC2HPO|Urine issues|Urine issues
C1977831|T201|MTH_LN|49959-0|LNC2HPO|Urine issues|Urine issues
C1977831|T201|LC|49959-0|LNC2HPO|Urine issues|Urine issues
C1977831|T201|OSN|49959-0|LNC2HPO|Urine issues|Urine issues
C1977831|T201|LN|49959-0|LNC2HPO|Pee issues|Pee issues
C1977831|T201|DN|49959-0|LNC2HPO|Pee issues|Pee issues
C1977831|T201|MTH_LN|49959-0|LNC2HPO|Pee issues|Pee issues
C1977831|T201|LC|49959-0|LNC2HPO|Pee issues|Pee issues
C1977831|T201|OSN|49959-0|LNC2HPO|Pee issues|Pee issues
C1977831|T201|LN|49959-0|LNC2HPO|Hyposthenuria|Hyposthenuria
C1977831|T201|DN|49959-0|LNC2HPO|Hyposthenuria|Hyposthenuria
C1977831|T201|MTH_LN|49959-0|LNC2HPO|Hyposthenuria|Hyposthenuria
C1977831|T201|LC|49959-0|LNC2HPO|Hyposthenuria|Hyposthenuria
C1977831|T201|OSN|49959-0|LNC2HPO|Hyposthenuria|Hyposthenuria
C1978489|T201|LN|50562-8|LNC2HPO|Urine issues|Urine issues
C1978489|T201|DN|50562-8|LNC2HPO|Urine issues|Urine issues
C1978489|T201|MTH_LN|50562-8|LNC2HPO|Urine issues|Urine issues
C1978489|T201|OSN|50562-8|LNC2HPO|Urine issues|Urine issues
C1978489|T201|LC|50562-8|LNC2HPO|Urine issues|Urine issues
C1978489|T201|LN|50562-8|LNC2HPO|Pee issues|Pee issues
C1978489|T201|DN|50562-8|LNC2HPO|Pee issues|Pee issues
C1978489|T201|MTH_LN|50562-8|LNC2HPO|Pee issues|Pee issues
C1978489|T201|OSN|50562-8|LNC2HPO|Pee issues|Pee issues
C1978489|T201|LC|50562-8|LNC2HPO|Pee issues|Pee issues
C1978489|T201|LN|50562-8|LNC2HPO|Hyposthenuria|Hyposthenuria
C1978489|T201|DN|50562-8|LNC2HPO|Hyposthenuria|Hyposthenuria
C1978489|T201|MTH_LN|50562-8|LNC2HPO|Hyposthenuria|Hyposthenuria
C1978489|T201|OSN|50562-8|LNC2HPO|Hyposthenuria|Hyposthenuria
C1978489|T201|LC|50562-8|LNC2HPO|Hyposthenuria|Hyposthenuria
C0368059|T201|LN|5810-7|LNC2HPO|Urine issues|Urine issues
C0368059|T201|MTH_LN|5810-7|LNC2HPO|Urine issues|Urine issues
C0368059|T201|DN|5810-7|LNC2HPO|Urine issues|Urine issues
C0368059|T201|LC|5810-7|LNC2HPO|Urine issues|Urine issues
C0368059|T201|OSN|5810-7|LNC2HPO|Urine issues|Urine issues
C0368059|T201|LN|5810-7|LNC2HPO|Pee issues|Pee issues
C0368059|T201|MTH_LN|5810-7|LNC2HPO|Pee issues|Pee issues
C0368059|T201|DN|5810-7|LNC2HPO|Pee issues|Pee issues
C0368059|T201|LC|5810-7|LNC2HPO|Pee issues|Pee issues
C0368059|T201|OSN|5810-7|LNC2HPO|Pee issues|Pee issues
C0368059|T201|LN|5810-7|LNC2HPO|Hyposthenuria|Hyposthenuria
C0368059|T201|MTH_LN|5810-7|LNC2HPO|Hyposthenuria|Hyposthenuria
C0368059|T201|DN|5810-7|LNC2HPO|Hyposthenuria|Hyposthenuria
C0368059|T201|LC|5810-7|LNC2HPO|Hyposthenuria|Hyposthenuria
C0368059|T201|OSN|5810-7|LNC2HPO|Hyposthenuria|Hyposthenuria
C0368061|T201|LN|5811-5|LNC2HPO|Urine issues|Urine issues
C0368061|T201|MTH_LN|5811-5|LNC2HPO|Urine issues|Urine issues
C0368061|T201|DN|5811-5|LNC2HPO|Urine issues|Urine issues
C0368061|T201|LC|5811-5|LNC2HPO|Urine issues|Urine issues
C0368061|T201|OSN|5811-5|LNC2HPO|Urine issues|Urine issues
C0368061|T201|LN|5811-5|LNC2HPO|Pee issues|Pee issues
C0368061|T201|MTH_LN|5811-5|LNC2HPO|Pee issues|Pee issues
C0368061|T201|DN|5811-5|LNC2HPO|Pee issues|Pee issues
C0368061|T201|LC|5811-5|LNC2HPO|Pee issues|Pee issues
C0368061|T201|OSN|5811-5|LNC2HPO|Pee issues|Pee issues
C0368061|T201|LN|5811-5|LNC2HPO|Hyposthenuria|Hyposthenuria
C0368061|T201|MTH_LN|5811-5|LNC2HPO|Hyposthenuria|Hyposthenuria
C0368061|T201|DN|5811-5|LNC2HPO|Hyposthenuria|Hyposthenuria
C0368061|T201|LC|5811-5|LNC2HPO|Hyposthenuria|Hyposthenuria
C0368061|T201|OSN|5811-5|LNC2HPO|Hyposthenuria|Hyposthenuria
C2363327|T201|MTH_LN|26513-2|LNC2HPO|Neutrophilia|Neutrophilia
C2363327|T201|OSN|26513-2|LNC2HPO|Neutrophilia|Neutrophilia
C2363327|T201|DN|26513-2|LNC2HPO|Neutrophilia|Neutrophilia
C2363327|T201|LN|26513-2|LNC2HPO|Neutrophilia|Neutrophilia
C2363327|T201|LC|26513-2|LNC2HPO|Neutrophilia|Neutrophilia
C2363327|T201|MTH_LN|26513-2|LNC2HPO|Neutropenia|Neutropenia
C2363327|T201|OSN|26513-2|LNC2HPO|Neutropenia|Neutropenia
C2363327|T201|DN|26513-2|LNC2HPO|Neutropenia|Neutropenia
C2363327|T201|LN|26513-2|LNC2HPO|Neutropenia|Neutropenia
C2363327|T201|LC|26513-2|LNC2HPO|Neutropenia|Neutropenia
C2363327|T201|MTH_LN|26513-2|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C2363327|T201|OSN|26513-2|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C2363327|T201|DN|26513-2|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C2363327|T201|LN|26513-2|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C2363327|T201|LC|26513-2|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0797129|T201|OSN|13941-0|LNC2HPO|Lymphocytosis|Lymphocytosis
C0797129|T201|DN|13941-0|LNC2HPO|Lymphocytosis|Lymphocytosis
C0797129|T201|LN|13941-0|LNC2HPO|Lymphocytosis|Lymphocytosis
C0797129|T201|MTH_LN|13941-0|LNC2HPO|Lymphocytosis|Lymphocytosis
C0797129|T201|LC|13941-0|LNC2HPO|Lymphocytosis|Lymphocytosis
C0797129|T201|OSN|13941-0|LNC2HPO|Lymphopenia|Lymphopenia
C0797129|T201|DN|13941-0|LNC2HPO|Lymphopenia|Lymphopenia
C0797129|T201|LN|13941-0|LNC2HPO|Lymphopenia|Lymphopenia
C0797129|T201|MTH_LN|13941-0|LNC2HPO|Lymphopenia|Lymphopenia
C0797129|T201|LC|13941-0|LNC2HPO|Lymphopenia|Lymphopenia
C0797129|T201|OSN|13941-0|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0797129|T201|DN|13941-0|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0797129|T201|LN|13941-0|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0797129|T201|MTH_LN|13941-0|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0797129|T201|LC|13941-0|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0797129|T201|OSN|13941-0|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0797129|T201|DN|13941-0|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0797129|T201|LN|13941-0|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0797129|T201|MTH_LN|13941-0|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0797129|T201|LC|13941-0|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0485832|T201|LN|8061-4|LNC2HPO|Antinuclear antibodies|Antinuclear antibodies
C0485832|T201|MTH_LN|8061-4|LNC2HPO|Antinuclear antibodies|Antinuclear antibodies
C0485832|T201|DN|8061-4|LNC2HPO|Antinuclear antibodies|Antinuclear antibodies
C0485832|T201|OSN|8061-4|LNC2HPO|Antinuclear antibodies|Antinuclear antibodies
C0485832|T201|LC|8061-4|LNC2HPO|Antinuclear antibodies|Antinuclear antibodies
C0485832|T201|LN|8061-4|LNC2HPO|Antinuclear antibody positive|Antinuclear antibody positive
C0485832|T201|MTH_LN|8061-4|LNC2HPO|Antinuclear antibody positive|Antinuclear antibody positive
C0485832|T201|DN|8061-4|LNC2HPO|Antinuclear antibody positive|Antinuclear antibody positive
C0485832|T201|OSN|8061-4|LNC2HPO|Antinuclear antibody positive|Antinuclear antibody positive
C0485832|T201|LC|8061-4|LNC2HPO|Antinuclear antibody positive|Antinuclear antibody positive
C0485832|T201|LN|8061-4|LNC2HPO|Serum antinuclear antibody|Serum antinuclear antibody
C0485832|T201|MTH_LN|8061-4|LNC2HPO|Serum antinuclear antibody|Serum antinuclear antibody
C0485832|T201|DN|8061-4|LNC2HPO|Serum antinuclear antibody|Serum antinuclear antibody
C0485832|T201|OSN|8061-4|LNC2HPO|Serum antinuclear antibody|Serum antinuclear antibody
C0485832|T201|LC|8061-4|LNC2HPO|Serum antinuclear antibody|Serum antinuclear antibody
C0942449|T201|LN|26487-9|LNC2HPO|Monocytosis|Monocytosis
C0942449|T201|OSN|26487-9|LNC2HPO|Monocytosis|Monocytosis
C0942449|T201|DN|26487-9|LNC2HPO|Monocytosis|Monocytosis
C0942449|T201|MTH_LN|26487-9|LNC2HPO|Monocytosis|Monocytosis
C0942449|T201|LC|26487-9|LNC2HPO|Monocytosis|Monocytosis
C0942449|T201|LN|26487-9|LNC2HPO|Monocytopenia|Monocytopenia
C0942449|T201|OSN|26487-9|LNC2HPO|Monocytopenia|Monocytopenia
C0942449|T201|DN|26487-9|LNC2HPO|Monocytopenia|Monocytopenia
C0942449|T201|MTH_LN|26487-9|LNC2HPO|Monocytopenia|Monocytopenia
C0942449|T201|LC|26487-9|LNC2HPO|Monocytopenia|Monocytopenia
C0802050|T201|LN|19113-0|LNC2HPO|IgE deficiency|IgE deficiency
C0802050|T201|LC|19113-0|LNC2HPO|IgE deficiency|IgE deficiency
C0802050|T201|OSN|19113-0|LNC2HPO|IgE deficiency|IgE deficiency
C0802050|T201|MTH_LN|19113-0|LNC2HPO|IgE deficiency|IgE deficiency
C0802050|T201|DN|19113-0|LNC2HPO|IgE deficiency|IgE deficiency
C0798132|T201|LN|14959-1|LNC2HPO|Microalbuminuria|Microalbuminuria
C0798132|T201|MTH_LN|14959-1|LNC2HPO|Microalbuminuria|Microalbuminuria
C0798132|T201|DN|14959-1|LNC2HPO|Microalbuminuria|Microalbuminuria
C0798132|T201|OSN|14959-1|LNC2HPO|Microalbuminuria|Microalbuminuria
C0798132|T201|LC|14959-1|LNC2HPO|Microalbuminuria|Microalbuminuria
C2598649|T201|LN|53531-0|LNC2HPO|Microalbuminuria|Microalbuminuria
C2598649|T201|DN|53531-0|LNC2HPO|Microalbuminuria|Microalbuminuria
C2598649|T201|MTH_LN|53531-0|LNC2HPO|Microalbuminuria|Microalbuminuria
C2598649|T201|OSN|53531-0|LNC2HPO|Microalbuminuria|Microalbuminuria
C2598649|T201|LC|53531-0|LNC2HPO|Microalbuminuria|Microalbuminuria
C1645723|T201|LN|41653-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C1645723|T201|DN|41653-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C1645723|T201|OSN|41653-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C1645723|T201|MTH_LN|41653-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C1645723|T201|LC|41653-7|LNC2HPO|Hyperglycemia|Hyperglycemia
C1645723|T201|LN|41653-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C1645723|T201|DN|41653-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C1645723|T201|OSN|41653-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C1645723|T201|MTH_LN|41653-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C1645723|T201|LC|41653-7|LNC2HPO|Hypoglycemia|Hypoglycemia
C1645723|T201|LN|41653-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1645723|T201|DN|41653-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1645723|T201|OSN|41653-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1645723|T201|MTH_LN|41653-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1645723|T201|LC|41653-7|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797944|T201|LN|14770-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797944|T201|MTH_LN|14770-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797944|T201|DN|14770-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797944|T201|OSN|14770-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797944|T201|LC|14770-2|LNC2HPO|Hyperglycemia|Hyperglycemia
C0797944|T201|LN|14770-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797944|T201|MTH_LN|14770-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797944|T201|DN|14770-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797944|T201|OSN|14770-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797944|T201|LC|14770-2|LNC2HPO|Hypoglycemia|Hypoglycemia
C0797944|T201|LN|14770-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797944|T201|MTH_LN|14770-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797944|T201|DN|14770-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797944|T201|OSN|14770-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C0797944|T201|LC|14770-2|LNC2HPO|Hypoglycaemia|Hypoglycaemia
C1830776|T201|LN|46702-7|LNC2HPO|Pyuria|Pyuria
C1830776|T201|MTH_LN|46702-7|LNC2HPO|Pyuria|Pyuria
C1830776|T201|OSN|46702-7|LNC2HPO|Pyuria|Pyuria
C1830776|T201|LC|46702-7|LNC2HPO|Pyuria|Pyuria
C1830776|T201|DN|46702-7|LNC2HPO|Pyuria|Pyuria
C1830776|T201|LN|46702-7|LNC2HPO|Leukocyturia|Leukocyturia
C1830776|T201|MTH_LN|46702-7|LNC2HPO|Leukocyturia|Leukocyturia
C1830776|T201|OSN|46702-7|LNC2HPO|Leukocyturia|Leukocyturia
C1830776|T201|LC|46702-7|LNC2HPO|Leukocyturia|Leukocyturia
C1830776|T201|DN|46702-7|LNC2HPO|Leukocyturia|Leukocyturia
C0803223|T201|LN|20408-1|LNC2HPO|Pyuria|Pyuria
C0803223|T201|DN|20408-1|LNC2HPO|Pyuria|Pyuria
C0803223|T201|OSN|20408-1|LNC2HPO|Pyuria|Pyuria
C0803223|T201|MTH_LN|20408-1|LNC2HPO|Pyuria|Pyuria
C0803223|T201|LC|20408-1|LNC2HPO|Pyuria|Pyuria
C0803223|T201|LN|20408-1|LNC2HPO|Leukocyturia|Leukocyturia
C0803223|T201|DN|20408-1|LNC2HPO|Leukocyturia|Leukocyturia
C0803223|T201|OSN|20408-1|LNC2HPO|Leukocyturia|Leukocyturia
C0803223|T201|MTH_LN|20408-1|LNC2HPO|Leukocyturia|Leukocyturia
C0803223|T201|LC|20408-1|LNC2HPO|Leukocyturia|Leukocyturia
C0803269|T201|LN|20455-2|LNC2HPO|Pyuria|Pyuria
C0803269|T201|MTH_LN|20455-2|LNC2HPO|Pyuria|Pyuria
C0803269|T201|DN|20455-2|LNC2HPO|Pyuria|Pyuria
C0803269|T201|OSN|20455-2|LNC2HPO|Pyuria|Pyuria
C0803269|T201|LC|20455-2|LNC2HPO|Pyuria|Pyuria
C0803269|T201|LN|20455-2|LNC2HPO|Leukocyturia|Leukocyturia
C0803269|T201|MTH_LN|20455-2|LNC2HPO|Leukocyturia|Leukocyturia
C0803269|T201|DN|20455-2|LNC2HPO|Leukocyturia|Leukocyturia
C0803269|T201|OSN|20455-2|LNC2HPO|Leukocyturia|Leukocyturia
C0803269|T201|LC|20455-2|LNC2HPO|Leukocyturia|Leukocyturia
C1114261|T201|LN|30405-5|LNC2HPO|Pyuria|Pyuria
C1114261|T201|DN|30405-5|LNC2HPO|Pyuria|Pyuria
C1114261|T201|OSN|30405-5|LNC2HPO|Pyuria|Pyuria
C1114261|T201|MTH_LN|30405-5|LNC2HPO|Pyuria|Pyuria
C1114261|T201|LC|30405-5|LNC2HPO|Pyuria|Pyuria
C1114261|T201|LN|30405-5|LNC2HPO|Leukocyturia|Leukocyturia
C1114261|T201|DN|30405-5|LNC2HPO|Leukocyturia|Leukocyturia
C1114261|T201|OSN|30405-5|LNC2HPO|Leukocyturia|Leukocyturia
C1114261|T201|MTH_LN|30405-5|LNC2HPO|Leukocyturia|Leukocyturia
C1114261|T201|LC|30405-5|LNC2HPO|Leukocyturia|Leukocyturia
C1744633|T201|LN|24122-4|LNC2HPO|Pyuria|Pyuria
C1744633|T201|DN|24122-4|LNC2HPO|Pyuria|Pyuria
C1744633|T201|OSN|24122-4|LNC2HPO|Pyuria|Pyuria
C1744633|T201|MTH_LN|24122-4|LNC2HPO|Pyuria|Pyuria
C1744633|T201|LC|24122-4|LNC2HPO|Pyuria|Pyuria
C1744633|T201|LN|24122-4|LNC2HPO|Leukocyturia|Leukocyturia
C1744633|T201|DN|24122-4|LNC2HPO|Leukocyturia|Leukocyturia
C1744633|T201|OSN|24122-4|LNC2HPO|Leukocyturia|Leukocyturia
C1744633|T201|MTH_LN|24122-4|LNC2HPO|Leukocyturia|Leukocyturia
C1744633|T201|LC|24122-4|LNC2HPO|Leukocyturia|Leukocyturia
C1315523|T201|LN|33052-2|LNC2HPO|Pyuria|Pyuria
C1315523|T201|MTH_LN|33052-2|LNC2HPO|Pyuria|Pyuria
C1315523|T201|DN|33052-2|LNC2HPO|Pyuria|Pyuria
C1315523|T201|OSN|33052-2|LNC2HPO|Pyuria|Pyuria
C1315523|T201|LC|33052-2|LNC2HPO|Pyuria|Pyuria
C1315523|T201|LN|33052-2|LNC2HPO|Leukocyturia|Leukocyturia
C1315523|T201|MTH_LN|33052-2|LNC2HPO|Leukocyturia|Leukocyturia
C1315523|T201|DN|33052-2|LNC2HPO|Leukocyturia|Leukocyturia
C1315523|T201|OSN|33052-2|LNC2HPO|Leukocyturia|Leukocyturia
C1315523|T201|LC|33052-2|LNC2HPO|Leukocyturia|Leukocyturia
C1716495|T201|LN|45383-7|LNC2HPO|Pyuria|Pyuria
C1716495|T201|DN|45383-7|LNC2HPO|Pyuria|Pyuria
C1716495|T201|MTH_LN|45383-7|LNC2HPO|Pyuria|Pyuria
C1716495|T201|OSN|45383-7|LNC2HPO|Pyuria|Pyuria
C1716495|T201|LC|45383-7|LNC2HPO|Pyuria|Pyuria
C1716495|T201|LN|45383-7|LNC2HPO|Leukocyturia|Leukocyturia
C1716495|T201|DN|45383-7|LNC2HPO|Leukocyturia|Leukocyturia
C1716495|T201|MTH_LN|45383-7|LNC2HPO|Leukocyturia|Leukocyturia
C1716495|T201|OSN|45383-7|LNC2HPO|Leukocyturia|Leukocyturia
C1716495|T201|LC|45383-7|LNC2HPO|Leukocyturia|Leukocyturia
C1979503|T201|LN|51487-7|LNC2HPO|Pyuria|Pyuria
C1979503|T201|DN|51487-7|LNC2HPO|Pyuria|Pyuria
C1979503|T201|MTH_LN|51487-7|LNC2HPO|Pyuria|Pyuria
C1979503|T201|OSN|51487-7|LNC2HPO|Pyuria|Pyuria
C1979503|T201|LC|51487-7|LNC2HPO|Pyuria|Pyuria
C1979503|T201|LN|51487-7|LNC2HPO|Leukocyturia|Leukocyturia
C1979503|T201|DN|51487-7|LNC2HPO|Leukocyturia|Leukocyturia
C1979503|T201|MTH_LN|51487-7|LNC2HPO|Leukocyturia|Leukocyturia
C1979503|T201|OSN|51487-7|LNC2HPO|Leukocyturia|Leukocyturia
C1979503|T201|LC|51487-7|LNC2HPO|Leukocyturia|Leukocyturia
C2361322|T201|LN|53316-6|LNC2HPO|Pyuria|Pyuria
C2361322|T201|MTH_LN|53316-6|LNC2HPO|Pyuria|Pyuria
C2361322|T201|DN|53316-6|LNC2HPO|Pyuria|Pyuria
C2361322|T201|OSN|53316-6|LNC2HPO|Pyuria|Pyuria
C2361322|T201|LC|53316-6|LNC2HPO|Pyuria|Pyuria
C2361322|T201|LN|53316-6|LNC2HPO|Leukocyturia|Leukocyturia
C2361322|T201|MTH_LN|53316-6|LNC2HPO|Leukocyturia|Leukocyturia
C2361322|T201|DN|53316-6|LNC2HPO|Leukocyturia|Leukocyturia
C2361322|T201|OSN|53316-6|LNC2HPO|Leukocyturia|Leukocyturia
C2361322|T201|LC|53316-6|LNC2HPO|Leukocyturia|Leukocyturia
C2598498|T201|LN|53964-3|LNC2HPO|Pyuria|Pyuria
C2598498|T201|MTH_LN|53964-3|LNC2HPO|Pyuria|Pyuria
C2598498|T201|DN|53964-3|LNC2HPO|Pyuria|Pyuria
C2598498|T201|LC|53964-3|LNC2HPO|Pyuria|Pyuria
C2598498|T201|OSN|53964-3|LNC2HPO|Pyuria|Pyuria
C2598498|T201|LN|53964-3|LNC2HPO|Leukocyturia|Leukocyturia
C2598498|T201|MTH_LN|53964-3|LNC2HPO|Leukocyturia|Leukocyturia
C2598498|T201|DN|53964-3|LNC2HPO|Leukocyturia|Leukocyturia
C2598498|T201|LC|53964-3|LNC2HPO|Leukocyturia|Leukocyturia
C2598498|T201|OSN|53964-3|LNC2HPO|Leukocyturia|Leukocyturia
C0368036|T201|LN|5821-4|LNC2HPO|Pyuria|Pyuria
C0368036|T201|DN|5821-4|LNC2HPO|Pyuria|Pyuria
C0368036|T201|MTH_LN|5821-4|LNC2HPO|Pyuria|Pyuria
C0368036|T201|LC|5821-4|LNC2HPO|Pyuria|Pyuria
C0368036|T201|OSN|5821-4|LNC2HPO|Pyuria|Pyuria
C0368036|T201|LN|5821-4|LNC2HPO|Leukocyturia|Leukocyturia
C0368036|T201|DN|5821-4|LNC2HPO|Leukocyturia|Leukocyturia
C0368036|T201|MTH_LN|5821-4|LNC2HPO|Leukocyturia|Leukocyturia
C0368036|T201|LC|5821-4|LNC2HPO|Leukocyturia|Leukocyturia
C0368036|T201|OSN|5821-4|LNC2HPO|Leukocyturia|Leukocyturia
C2923139|T201|LN|58805-3|LNC2HPO|Pyuria|Pyuria
C2923139|T201|DN|58805-3|LNC2HPO|Pyuria|Pyuria
C2923139|T201|MTH_LN|58805-3|LNC2HPO|Pyuria|Pyuria
C2923139|T201|LC|58805-3|LNC2HPO|Pyuria|Pyuria
C2923139|T201|OSN|58805-3|LNC2HPO|Pyuria|Pyuria
C2923139|T201|LN|58805-3|LNC2HPO|Leukocyturia|Leukocyturia
C2923139|T201|DN|58805-3|LNC2HPO|Leukocyturia|Leukocyturia
C2923139|T201|MTH_LN|58805-3|LNC2HPO|Leukocyturia|Leukocyturia
C2923139|T201|LC|58805-3|LNC2HPO|Leukocyturia|Leukocyturia
C2923139|T201|OSN|58805-3|LNC2HPO|Leukocyturia|Leukocyturia
C2924077|T201|LN|59829-2|LNC2HPO|Pyuria|Pyuria
C2924077|T201|DN|59829-2|LNC2HPO|Pyuria|Pyuria
C2924077|T201|LC|59829-2|LNC2HPO|Pyuria|Pyuria
C2924077|T201|OSN|59829-2|LNC2HPO|Pyuria|Pyuria
C2924077|T201|MTH_LN|59829-2|LNC2HPO|Pyuria|Pyuria
C2924077|T201|LN|59829-2|LNC2HPO|Leukocyturia|Leukocyturia
C2924077|T201|DN|59829-2|LNC2HPO|Leukocyturia|Leukocyturia
C2924077|T201|LC|59829-2|LNC2HPO|Leukocyturia|Leukocyturia
C2924077|T201|OSN|59829-2|LNC2HPO|Leukocyturia|Leukocyturia
C2924077|T201|MTH_LN|59829-2|LNC2HPO|Leukocyturia|Leukocyturia
C3172620|T201|LN|63554-0|LNC2HPO|Pyuria|Pyuria
C3172620|T201|MTH_LN|63554-0|LNC2HPO|Pyuria|Pyuria
C3172620|T201|OSN|63554-0|LNC2HPO|Pyuria|Pyuria
C3172620|T201|LC|63554-0|LNC2HPO|Pyuria|Pyuria
C3172620|T201|DN|63554-0|LNC2HPO|Pyuria|Pyuria
C3172620|T201|LN|63554-0|LNC2HPO|Leukocyturia|Leukocyturia
C3172620|T201|MTH_LN|63554-0|LNC2HPO|Leukocyturia|Leukocyturia
C3172620|T201|OSN|63554-0|LNC2HPO|Leukocyturia|Leukocyturia
C3172620|T201|LC|63554-0|LNC2HPO|Leukocyturia|Leukocyturia
C3172620|T201|DN|63554-0|LNC2HPO|Leukocyturia|Leukocyturia
C0801449|T201|LN|18407-7|LNC2HPO|Pyuria|Pyuria
C0801449|T201|DN|18407-7|LNC2HPO|Pyuria|Pyuria
C0801449|T201|OSN|18407-7|LNC2HPO|Pyuria|Pyuria
C0801449|T201|MTH_LN|18407-7|LNC2HPO|Pyuria|Pyuria
C0801449|T201|LC|18407-7|LNC2HPO|Pyuria|Pyuria
C0801449|T201|LN|18407-7|LNC2HPO|Leukocyturia|Leukocyturia
C0801449|T201|DN|18407-7|LNC2HPO|Leukocyturia|Leukocyturia
C0801449|T201|OSN|18407-7|LNC2HPO|Leukocyturia|Leukocyturia
C0801449|T201|MTH_LN|18407-7|LNC2HPO|Leukocyturia|Leukocyturia
C0801449|T201|LC|18407-7|LNC2HPO|Leukocyturia|Leukocyturia
C2361327|T201|LN|53321-6|LNC2HPO|Urine issues|Urine issues
C2361327|T201|MTH_LN|53321-6|LNC2HPO|Urine issues|Urine issues
C2361327|T201|DN|53321-6|LNC2HPO|Urine issues|Urine issues
C2361327|T201|OSN|53321-6|LNC2HPO|Urine issues|Urine issues
C2361327|T201|LC|53321-6|LNC2HPO|Urine issues|Urine issues
C2361327|T201|LN|53321-6|LNC2HPO|Pee issues|Pee issues
C2361327|T201|MTH_LN|53321-6|LNC2HPO|Pee issues|Pee issues
C2361327|T201|DN|53321-6|LNC2HPO|Pee issues|Pee issues
C2361327|T201|OSN|53321-6|LNC2HPO|Pee issues|Pee issues
C2361327|T201|LC|53321-6|LNC2HPO|Pee issues|Pee issues
C0486210|T201|LN|8247-9|LNC2HPO|Urine issues|Urine issues
C0486210|T201|MTH_LN|8247-9|LNC2HPO|Urine issues|Urine issues
C0486210|T201|DN|8247-9|LNC2HPO|Urine issues|Urine issues
C0486210|T201|OSN|8247-9|LNC2HPO|Urine issues|Urine issues
C0486210|T201|LC|8247-9|LNC2HPO|Urine issues|Urine issues
C0486210|T201|LN|8247-9|LNC2HPO|Pee issues|Pee issues
C0486210|T201|MTH_LN|8247-9|LNC2HPO|Pee issues|Pee issues
C0486210|T201|DN|8247-9|LNC2HPO|Pee issues|Pee issues
C0486210|T201|OSN|8247-9|LNC2HPO|Pee issues|Pee issues
C0486210|T201|LC|8247-9|LNC2HPO|Pee issues|Pee issues
C1979494|T201|LN|51478-6|LNC2HPO|Urine issues|Urine issues
C1979494|T201|DN|51478-6|LNC2HPO|Urine issues|Urine issues
C1979494|T201|OSN|51478-6|LNC2HPO|Urine issues|Urine issues
C1979494|T201|MTH_LN|51478-6|LNC2HPO|Urine issues|Urine issues
C1979494|T201|LC|51478-6|LNC2HPO|Urine issues|Urine issues
C1979494|T201|LN|51478-6|LNC2HPO|Pee issues|Pee issues
C1979494|T201|DN|51478-6|LNC2HPO|Pee issues|Pee issues
C1979494|T201|OSN|51478-6|LNC2HPO|Pee issues|Pee issues
C1979494|T201|MTH_LN|51478-6|LNC2HPO|Pee issues|Pee issues
C1979494|T201|LC|51478-6|LNC2HPO|Pee issues|Pee issues
C1978070|T201|LN|50235-1|LNC2HPO|Urine issues|Urine issues
C1978070|T201|MTH_LN|50235-1|LNC2HPO|Urine issues|Urine issues
C1978070|T201|OSN|50235-1|LNC2HPO|Urine issues|Urine issues
C1978070|T201|LC|50235-1|LNC2HPO|Urine issues|Urine issues
C1978070|T201|DN|50235-1|LNC2HPO|Urine issues|Urine issues
C1978070|T201|LN|50235-1|LNC2HPO|Pee issues|Pee issues
C1978070|T201|MTH_LN|50235-1|LNC2HPO|Pee issues|Pee issues
C1978070|T201|OSN|50235-1|LNC2HPO|Pee issues|Pee issues
C1978070|T201|LC|50235-1|LNC2HPO|Pee issues|Pee issues
C1978070|T201|DN|50235-1|LNC2HPO|Pee issues|Pee issues
C1830310|T201|LN|46421-4|LNC2HPO|Urine issues|Urine issues
C1830310|T201|DN|46421-4|LNC2HPO|Urine issues|Urine issues
C1830310|T201|MTH_LN|46421-4|LNC2HPO|Urine issues|Urine issues
C1830310|T201|LC|46421-4|LNC2HPO|Urine issues|Urine issues
C1830310|T201|OSN|46421-4|LNC2HPO|Urine issues|Urine issues
C1830310|T201|LN|46421-4|LNC2HPO|Pee issues|Pee issues
C1830310|T201|DN|46421-4|LNC2HPO|Pee issues|Pee issues
C1830310|T201|MTH_LN|46421-4|LNC2HPO|Pee issues|Pee issues
C1830310|T201|LC|46421-4|LNC2HPO|Pee issues|Pee issues
C1830310|T201|OSN|46421-4|LNC2HPO|Pee issues|Pee issues
C0944138|T201|LN|28545-2|LNC2HPO|Urine issues|Urine issues
C0944138|T201|DN|28545-2|LNC2HPO|Urine issues|Urine issues
C0944138|T201|MTH_LN|28545-2|LNC2HPO|Urine issues|Urine issues
C0944138|T201|OSN|28545-2|LNC2HPO|Urine issues|Urine issues
C0944138|T201|LC|28545-2|LNC2HPO|Urine issues|Urine issues
C0944138|T201|LN|28545-2|LNC2HPO|Pee issues|Pee issues
C0944138|T201|DN|28545-2|LNC2HPO|Pee issues|Pee issues
C0944138|T201|MTH_LN|28545-2|LNC2HPO|Pee issues|Pee issues
C0944138|T201|OSN|28545-2|LNC2HPO|Pee issues|Pee issues
C0944138|T201|LC|28545-2|LNC2HPO|Pee issues|Pee issues
C0944223|T201|LN|28642-7|LNC2HPO|Hyperoxemia|Hyperoxemia
C0944223|T201|DN|28642-7|LNC2HPO|Hyperoxemia|Hyperoxemia
C0944223|T201|LC|28642-7|LNC2HPO|Hyperoxemia|Hyperoxemia
C0944223|T201|MTH_LN|28642-7|LNC2HPO|Hyperoxemia|Hyperoxemia
C0944223|T201|OSN|28642-7|LNC2HPO|Hyperoxemia|Hyperoxemia
C0944223|T201|LN|28642-7|LNC2HPO|Hypoxemia|Hypoxemia
C0944223|T201|DN|28642-7|LNC2HPO|Hypoxemia|Hypoxemia
C0944223|T201|LC|28642-7|LNC2HPO|Hypoxemia|Hypoxemia
C0944223|T201|MTH_LN|28642-7|LNC2HPO|Hypoxemia|Hypoxemia
C0944223|T201|OSN|28642-7|LNC2HPO|Hypoxemia|Hypoxemia
C3483886|T201|LN|71847-8|LNC2HPO|Hyperoxemia|Hyperoxemia
C3483886|T201|LC|71847-8|LNC2HPO|Hyperoxemia|Hyperoxemia
C3483886|T201|MTH_LN|71847-8|LNC2HPO|Hyperoxemia|Hyperoxemia
C3483886|T201|OSN|71847-8|LNC2HPO|Hyperoxemia|Hyperoxemia
C3483886|T201|DN|71847-8|LNC2HPO|Hyperoxemia|Hyperoxemia
C3483886|T201|LN|71847-8|LNC2HPO|Hypoxemia|Hypoxemia
C3483886|T201|LC|71847-8|LNC2HPO|Hypoxemia|Hypoxemia
C3483886|T201|MTH_LN|71847-8|LNC2HPO|Hypoxemia|Hypoxemia
C3483886|T201|OSN|71847-8|LNC2HPO|Hypoxemia|Hypoxemia
C3483886|T201|DN|71847-8|LNC2HPO|Hypoxemia|Hypoxemia
C2733831|T201|LN|55859-3|LNC2HPO|Folate deficiency in cerebrospinal fluid|Folate deficiency in cerebrospinal fluid
C2733831|T201|DN|55859-3|LNC2HPO|Folate deficiency in cerebrospinal fluid|Folate deficiency in cerebrospinal fluid
C2733831|T201|OSN|55859-3|LNC2HPO|Folate deficiency in cerebrospinal fluid|Folate deficiency in cerebrospinal fluid
C2733831|T201|LC|55859-3|LNC2HPO|Folate deficiency in cerebrospinal fluid|Folate deficiency in cerebrospinal fluid
C2733831|T201|MTH_LN|55859-3|LNC2HPO|Folate deficiency in cerebrospinal fluid|Folate deficiency in cerebrospinal fluid
C0482617|T201|LN|3193-0|LNC2HPO|Factor V deficiency|Factor V deficiency
C0482617|T201|DN|3193-0|LNC2HPO|Factor V deficiency|Factor V deficiency
C0482617|T201|MTH_LN|3193-0|LNC2HPO|Factor V deficiency|Factor V deficiency
C0482617|T201|OSN|3193-0|LNC2HPO|Factor V deficiency|Factor V deficiency
C0482617|T201|LC|3193-0|LNC2HPO|Factor V deficiency|Factor V deficiency
C0550349|T201|LN|10834-0|LNC2HPO|Hypergammaglobulinemia|Hypergammaglobulinemia
C0550349|T201|MTH_LN|10834-0|LNC2HPO|Hypergammaglobulinemia|Hypergammaglobulinemia
C0550349|T201|DN|10834-0|LNC2HPO|Hypergammaglobulinemia|Hypergammaglobulinemia
C0550349|T201|OSN|10834-0|LNC2HPO|Hypergammaglobulinemia|Hypergammaglobulinemia
C0550349|T201|LC|10834-0|LNC2HPO|Hypergammaglobulinemia|Hypergammaglobulinemia
C0550349|T201|LN|10834-0|LNC2HPO|Hypergammaglobulinaemia|Hypergammaglobulinaemia
C0550349|T201|MTH_LN|10834-0|LNC2HPO|Hypergammaglobulinaemia|Hypergammaglobulinaemia
C0550349|T201|DN|10834-0|LNC2HPO|Hypergammaglobulinaemia|Hypergammaglobulinaemia
C0550349|T201|OSN|10834-0|LNC2HPO|Hypergammaglobulinaemia|Hypergammaglobulinaemia
C0550349|T201|LC|10834-0|LNC2HPO|Hypergammaglobulinaemia|Hypergammaglobulinaemia
C0550349|T201|LN|10834-0|LNC2HPO|Hyperglobulinemia|Hyperglobulinemia
C0550349|T201|MTH_LN|10834-0|LNC2HPO|Hyperglobulinemia|Hyperglobulinemia
C0550349|T201|DN|10834-0|LNC2HPO|Hyperglobulinemia|Hyperglobulinemia
C0550349|T201|OSN|10834-0|LNC2HPO|Hyperglobulinemia|Hyperglobulinemia
C0550349|T201|LC|10834-0|LNC2HPO|Hyperglobulinemia|Hyperglobulinemia
C0550349|T201|LN|10834-0|LNC2HPO|Hypogammaglobulinemia|Hypogammaglobulinemia
C0550349|T201|MTH_LN|10834-0|LNC2HPO|Hypogammaglobulinemia|Hypogammaglobulinemia
C0550349|T201|DN|10834-0|LNC2HPO|Hypogammaglobulinemia|Hypogammaglobulinemia
C0550349|T201|OSN|10834-0|LNC2HPO|Hypogammaglobulinemia|Hypogammaglobulinemia
C0550349|T201|LC|10834-0|LNC2HPO|Hypogammaglobulinemia|Hypogammaglobulinemia
C0550349|T201|LN|10834-0|LNC2HPO|Immunoglobulin deficiency|Immunoglobulin deficiency
C0550349|T201|MTH_LN|10834-0|LNC2HPO|Immunoglobulin deficiency|Immunoglobulin deficiency
C0550349|T201|DN|10834-0|LNC2HPO|Immunoglobulin deficiency|Immunoglobulin deficiency
C0550349|T201|OSN|10834-0|LNC2HPO|Immunoglobulin deficiency|Immunoglobulin deficiency
C0550349|T201|LC|10834-0|LNC2HPO|Immunoglobulin deficiency|Immunoglobulin deficiency
C0803440|T201|LN|20636-7|LNC2HPO|Hyperalaninemia|Hyperalaninemia
C0803440|T201|MTH_LN|20636-7|LNC2HPO|Hyperalaninemia|Hyperalaninemia
C0803440|T201|DN|20636-7|LNC2HPO|Hyperalaninemia|Hyperalaninemia
C0803440|T201|OSN|20636-7|LNC2HPO|Hyperalaninemia|Hyperalaninemia
C0803440|T201|LC|20636-7|LNC2HPO|Hyperalaninemia|Hyperalaninemia
C0803440|T201|LN|20636-7|LNC2HPO|Hypoalaninemia|Hypoalaninemia
C0803440|T201|MTH_LN|20636-7|LNC2HPO|Hypoalaninemia|Hypoalaninemia
C0803440|T201|DN|20636-7|LNC2HPO|Hypoalaninemia|Hypoalaninemia
C0803440|T201|OSN|20636-7|LNC2HPO|Hypoalaninemia|Hypoalaninemia
C0803440|T201|LC|20636-7|LNC2HPO|Hypoalaninemia|Hypoalaninemia
C0364028|T201|LN|1893-7|LNC2HPO|Hyperargininemia|Hyperargininemia
C0364028|T201|DN|1893-7|LNC2HPO|Hyperargininemia|Hyperargininemia
C0364028|T201|MTH_LN|1893-7|LNC2HPO|Hyperargininemia|Hyperargininemia
C0364028|T201|OSN|1893-7|LNC2HPO|Hyperargininemia|Hyperargininemia
C0364028|T201|LC|1893-7|LNC2HPO|Hyperargininemia|Hyperargininemia
C0364028|T201|LN|1893-7|LNC2HPO|Arginine deficiency|Arginine deficiency
C0364028|T201|DN|1893-7|LNC2HPO|Arginine deficiency|Arginine deficiency
C0364028|T201|MTH_LN|1893-7|LNC2HPO|Arginine deficiency|Arginine deficiency
C0364028|T201|OSN|1893-7|LNC2HPO|Arginine deficiency|Arginine deficiency
C0364028|T201|LC|1893-7|LNC2HPO|Arginine deficiency|Arginine deficiency
C0364028|T201|LN|1893-7|LNC2HPO|Hypoargininemia|Hypoargininemia
C0364028|T201|DN|1893-7|LNC2HPO|Hypoargininemia|Hypoargininemia
C0364028|T201|MTH_LN|1893-7|LNC2HPO|Hypoargininemia|Hypoargininemia
C0364028|T201|OSN|1893-7|LNC2HPO|Hypoargininemia|Hypoargininemia
C0364028|T201|LC|1893-7|LNC2HPO|Hypoargininemia|Hypoargininemia
C0803441|T201|LN|20637-5|LNC2HPO|Hyperargininemia|Hyperargininemia
C0803441|T201|MTH_LN|20637-5|LNC2HPO|Hyperargininemia|Hyperargininemia
C0803441|T201|DN|20637-5|LNC2HPO|Hyperargininemia|Hyperargininemia
C0803441|T201|OSN|20637-5|LNC2HPO|Hyperargininemia|Hyperargininemia
C0803441|T201|LC|20637-5|LNC2HPO|Hyperargininemia|Hyperargininemia
C0803441|T201|LN|20637-5|LNC2HPO|Arginine deficiency|Arginine deficiency
C0803441|T201|MTH_LN|20637-5|LNC2HPO|Arginine deficiency|Arginine deficiency
C0803441|T201|DN|20637-5|LNC2HPO|Arginine deficiency|Arginine deficiency
C0803441|T201|OSN|20637-5|LNC2HPO|Arginine deficiency|Arginine deficiency
C0803441|T201|LC|20637-5|LNC2HPO|Arginine deficiency|Arginine deficiency
C0803441|T201|LN|20637-5|LNC2HPO|Hypoargininemia|Hypoargininemia
C0803441|T201|MTH_LN|20637-5|LNC2HPO|Hypoargininemia|Hypoargininemia
C0803441|T201|DN|20637-5|LNC2HPO|Hypoargininemia|Hypoargininemia
C0803441|T201|OSN|20637-5|LNC2HPO|Hypoargininemia|Hypoargininemia
C0803441|T201|LC|20637-5|LNC2HPO|Hypoargininemia|Hypoargininemia
C0364043|T201|LN|1908-3|LNC2HPO|Hyperasparaginemia|Hyperasparaginemia
C0364043|T201|DN|1908-3|LNC2HPO|Hyperasparaginemia|Hyperasparaginemia
C0364043|T201|MTH_LN|1908-3|LNC2HPO|Hyperasparaginemia|Hyperasparaginemia
C0364043|T201|OSN|1908-3|LNC2HPO|Hyperasparaginemia|Hyperasparaginemia
C0364043|T201|LC|1908-3|LNC2HPO|Hyperasparaginemia|Hyperasparaginemia
C0364043|T201|LN|1908-3|LNC2HPO|Hypoasparaginemia|Hypoasparaginemia
C0364043|T201|DN|1908-3|LNC2HPO|Hypoasparaginemia|Hypoasparaginemia
C0364043|T201|MTH_LN|1908-3|LNC2HPO|Hypoasparaginemia|Hypoasparaginemia
C0364043|T201|OSN|1908-3|LNC2HPO|Hypoasparaginemia|Hypoasparaginemia
C0364043|T201|LC|1908-3|LNC2HPO|Hypoasparaginemia|Hypoasparaginemia
C0803442|T201|LN|20638-3|LNC2HPO|Hyperasparaginemia|Hyperasparaginemia
C0803442|T201|MTH_LN|20638-3|LNC2HPO|Hyperasparaginemia|Hyperasparaginemia
C0803442|T201|DN|20638-3|LNC2HPO|Hyperasparaginemia|Hyperasparaginemia
C0803442|T201|OSN|20638-3|LNC2HPO|Hyperasparaginemia|Hyperasparaginemia
C0803442|T201|LC|20638-3|LNC2HPO|Hyperasparaginemia|Hyperasparaginemia
C0803442|T201|LN|20638-3|LNC2HPO|Hypoasparaginemia|Hypoasparaginemia
C0803442|T201|MTH_LN|20638-3|LNC2HPO|Hypoasparaginemia|Hypoasparaginemia
C0803442|T201|DN|20638-3|LNC2HPO|Hypoasparaginemia|Hypoasparaginemia
C0803442|T201|OSN|20638-3|LNC2HPO|Hypoasparaginemia|Hypoasparaginemia
C0803442|T201|LC|20638-3|LNC2HPO|Hypoasparaginemia|Hypoasparaginemia
C0880190|T201|LN|22672-0|LNC2HPO|Hypercystinemia|Hypercystinemia
C0880190|T201|DN|22672-0|LNC2HPO|Hypercystinemia|Hypercystinemia
C0880190|T201|MTH_LN|22672-0|LNC2HPO|Hypercystinemia|Hypercystinemia
C0880190|T201|OSN|22672-0|LNC2HPO|Hypercystinemia|Hypercystinemia
C0880190|T201|LC|22672-0|LNC2HPO|Hypercystinemia|Hypercystinemia
C0880190|T201|LN|22672-0|LNC2HPO|Hypocystinemia|Hypocystinemia
C0880190|T201|DN|22672-0|LNC2HPO|Hypocystinemia|Hypocystinemia
C0880190|T201|MTH_LN|22672-0|LNC2HPO|Hypocystinemia|Hypocystinemia
C0880190|T201|OSN|22672-0|LNC2HPO|Hypocystinemia|Hypocystinemia
C0880190|T201|LC|22672-0|LNC2HPO|Hypocystinemia|Hypocystinemia
C0880187|T201|MTH_LN|20642-5|LNC2HPO|Hyperglutamatemia|Hyperglutamatemia
C0880187|T201|DN|20642-5|LNC2HPO|Hyperglutamatemia|Hyperglutamatemia
C0880187|T201|LN|20642-5|LNC2HPO|Hyperglutamatemia|Hyperglutamatemia
C0880187|T201|OSN|20642-5|LNC2HPO|Hyperglutamatemia|Hyperglutamatemia
C0880187|T201|LC|20642-5|LNC2HPO|Hyperglutamatemia|Hyperglutamatemia
C0880187|T201|MTH_LN|20642-5|LNC2HPO|Hypoglutamatemia|Hypoglutamatemia
C0880187|T201|DN|20642-5|LNC2HPO|Hypoglutamatemia|Hypoglutamatemia
C0880187|T201|LN|20642-5|LNC2HPO|Hypoglutamatemia|Hypoglutamatemia
C0880187|T201|OSN|20642-5|LNC2HPO|Hypoglutamatemia|Hypoglutamatemia
C0880187|T201|LC|20642-5|LNC2HPO|Hypoglutamatemia|Hypoglutamatemia
C0803447|T201|LN|20643-3|LNC2HPO|Hyperglutaminemia|Hyperglutaminemia
C0803447|T201|MTH_LN|20643-3|LNC2HPO|Hyperglutaminemia|Hyperglutaminemia
C0803447|T201|DN|20643-3|LNC2HPO|Hyperglutaminemia|Hyperglutaminemia
C0803447|T201|OSN|20643-3|LNC2HPO|Hyperglutaminemia|Hyperglutaminemia
C0803447|T201|LC|20643-3|LNC2HPO|Hyperglutaminemia|Hyperglutaminemia
C0803447|T201|LN|20643-3|LNC2HPO|Hypoglutaminemia|Hypoglutaminemia
C0803447|T201|MTH_LN|20643-3|LNC2HPO|Hypoglutaminemia|Hypoglutaminemia
C0803447|T201|DN|20643-3|LNC2HPO|Hypoglutaminemia|Hypoglutaminemia
C0803447|T201|OSN|20643-3|LNC2HPO|Hypoglutaminemia|Hypoglutaminemia
C0803447|T201|LC|20643-3|LNC2HPO|Hypoglutaminemia|Hypoglutaminemia
C0803449|T201|LN|20645-8|LNC2HPO|Histidinemia|Histidinemia
C0803449|T201|MTH_LN|20645-8|LNC2HPO|Histidinemia|Histidinemia
C0803449|T201|DN|20645-8|LNC2HPO|Histidinemia|Histidinemia
C0803449|T201|OSN|20645-8|LNC2HPO|Histidinemia|Histidinemia
C0803449|T201|LC|20645-8|LNC2HPO|Histidinemia|Histidinemia
C0803449|T201|LN|20645-8|LNC2HPO|Hyperhistidinemia|Hyperhistidinemia
C0803449|T201|MTH_LN|20645-8|LNC2HPO|Hyperhistidinemia|Hyperhistidinemia
C0803449|T201|DN|20645-8|LNC2HPO|Hyperhistidinemia|Hyperhistidinemia
C0803449|T201|OSN|20645-8|LNC2HPO|Hyperhistidinemia|Hyperhistidinemia
C0803449|T201|LC|20645-8|LNC2HPO|Hyperhistidinemia|Hyperhistidinemia
C0803449|T201|LN|20645-8|LNC2HPO|Hypohistidinemia|Hypohistidinemia
C0803449|T201|MTH_LN|20645-8|LNC2HPO|Hypohistidinemia|Hypohistidinemia
C0803449|T201|DN|20645-8|LNC2HPO|Hypohistidinemia|Hypohistidinemia
C0803449|T201|OSN|20645-8|LNC2HPO|Hypohistidinemia|Hypohistidinemia
C0803449|T201|LC|20645-8|LNC2HPO|Hypohistidinemia|Hypohistidinemia
C0797153|T201|LN|13965-9|LNC2HPO|Hyperhomocystinemia|Hyperhomocystinemia
C0797153|T201|OSN|13965-9|LNC2HPO|Hyperhomocystinemia|Hyperhomocystinemia
C0797153|T201|DN|13965-9|LNC2HPO|Hyperhomocystinemia|Hyperhomocystinemia
C0797153|T201|MTH_LN|13965-9|LNC2HPO|Hyperhomocystinemia|Hyperhomocystinemia
C0797153|T201|LC|13965-9|LNC2HPO|Hyperhomocystinemia|Hyperhomocystinemia
C0797153|T201|LN|13965-9|LNC2HPO|Homocystinemia|Homocystinemia
C0797153|T201|OSN|13965-9|LNC2HPO|Homocystinemia|Homocystinemia
C0797153|T201|DN|13965-9|LNC2HPO|Homocystinemia|Homocystinemia
C0797153|T201|MTH_LN|13965-9|LNC2HPO|Homocystinemia|Homocystinemia
C0797153|T201|LC|13965-9|LNC2HPO|Homocystinemia|Homocystinemia
C0803451|T201|LN|20647-4|LNC2HPO|Hydroxyprolinemia|Hydroxyprolinemia
C0803451|T201|MTH_LN|20647-4|LNC2HPO|Hydroxyprolinemia|Hydroxyprolinemia
C0803451|T201|DN|20647-4|LNC2HPO|Hydroxyprolinemia|Hydroxyprolinemia
C0803451|T201|OSN|20647-4|LNC2HPO|Hydroxyprolinemia|Hydroxyprolinemia
C0803451|T201|LC|20647-4|LNC2HPO|Hydroxyprolinemia|Hydroxyprolinemia
C0803452|T201|LN|20648-2|LNC2HPO|Hyperisoleucinemia|Hyperisoleucinemia
C0803452|T201|MTH_LN|20648-2|LNC2HPO|Hyperisoleucinemia|Hyperisoleucinemia
C0803452|T201|DN|20648-2|LNC2HPO|Hyperisoleucinemia|Hyperisoleucinemia
C0803452|T201|OSN|20648-2|LNC2HPO|Hyperisoleucinemia|Hyperisoleucinemia
C0803452|T201|LC|20648-2|LNC2HPO|Hyperisoleucinemia|Hyperisoleucinemia
C0803452|T201|LN|20648-2|LNC2HPO|Hypoisoleucinemia|Hypoisoleucinemia
C0803452|T201|MTH_LN|20648-2|LNC2HPO|Hypoisoleucinemia|Hypoisoleucinemia
C0803452|T201|DN|20648-2|LNC2HPO|Hypoisoleucinemia|Hypoisoleucinemia
C0803452|T201|OSN|20648-2|LNC2HPO|Hypoisoleucinemia|Hypoisoleucinemia
C0803452|T201|LC|20648-2|LNC2HPO|Hypoisoleucinemia|Hypoisoleucinemia
C0803453|T201|LN|20649-0|LNC2HPO|Hyperleucinemia|Hyperleucinemia
C0803453|T201|MTH_LN|20649-0|LNC2HPO|Hyperleucinemia|Hyperleucinemia
C0803453|T201|DN|20649-0|LNC2HPO|Hyperleucinemia|Hyperleucinemia
C0803453|T201|OSN|20649-0|LNC2HPO|Hyperleucinemia|Hyperleucinemia
C0803453|T201|LC|20649-0|LNC2HPO|Hyperleucinemia|Hyperleucinemia
C0803453|T201|LN|20649-0|LNC2HPO|Hypoleucinemia|Hypoleucinemia
C0803453|T201|MTH_LN|20649-0|LNC2HPO|Hypoleucinemia|Hypoleucinemia
C0803453|T201|DN|20649-0|LNC2HPO|Hypoleucinemia|Hypoleucinemia
C0803453|T201|OSN|20649-0|LNC2HPO|Hypoleucinemia|Hypoleucinemia
C0803453|T201|LC|20649-0|LNC2HPO|Hypoleucinemia|Hypoleucinemia
C0803454|T201|LN|20650-8|LNC2HPO|Hyperlysinemia|Hyperlysinemia
C0803454|T201|MTH_LN|20650-8|LNC2HPO|Hyperlysinemia|Hyperlysinemia
C0803454|T201|DN|20650-8|LNC2HPO|Hyperlysinemia|Hyperlysinemia
C0803454|T201|OSN|20650-8|LNC2HPO|Hyperlysinemia|Hyperlysinemia
C0803454|T201|LC|20650-8|LNC2HPO|Hyperlysinemia|Hyperlysinemia
C0803454|T201|LN|20650-8|LNC2HPO|Hypolysinemia|Hypolysinemia
C0803454|T201|MTH_LN|20650-8|LNC2HPO|Hypolysinemia|Hypolysinemia
C0803454|T201|DN|20650-8|LNC2HPO|Hypolysinemia|Hypolysinemia
C0803454|T201|OSN|20650-8|LNC2HPO|Hypolysinemia|Hypolysinemia
C0803454|T201|LC|20650-8|LNC2HPO|Hypolysinemia|Hypolysinemia
C0803456|T201|LN|20652-4|LNC2HPO|Hyperornithinemia|Hyperornithinemia
C0803456|T201|MTH_LN|20652-4|LNC2HPO|Hyperornithinemia|Hyperornithinemia
C0803456|T201|DN|20652-4|LNC2HPO|Hyperornithinemia|Hyperornithinemia
C0803456|T201|OSN|20652-4|LNC2HPO|Hyperornithinemia|Hyperornithinemia
C0803456|T201|LC|20652-4|LNC2HPO|Hyperornithinemia|Hyperornithinemia
C0803456|T201|LN|20652-4|LNC2HPO|Hypoornithinemia|Hypoornithinemia
C0803456|T201|MTH_LN|20652-4|LNC2HPO|Hypoornithinemia|Hypoornithinemia
C0803456|T201|DN|20652-4|LNC2HPO|Hypoornithinemia|Hypoornithinemia
C0803456|T201|OSN|20652-4|LNC2HPO|Hypoornithinemia|Hypoornithinemia
C0803456|T201|LC|20652-4|LNC2HPO|Hypoornithinemia|Hypoornithinemia
C1544784|T201|LN|40829-4|LNC2HPO|Hyperornithinemia|Hyperornithinemia
C1544784|T201|MTH_LN|40829-4|LNC2HPO|Hyperornithinemia|Hyperornithinemia
C1544784|T201|OSN|40829-4|LNC2HPO|Hyperornithinemia|Hyperornithinemia
C1544784|T201|DN|40829-4|LNC2HPO|Hyperornithinemia|Hyperornithinemia
C1544784|T201|LC|40829-4|LNC2HPO|Hyperornithinemia|Hyperornithinemia
C0798049|T201|MTH_LN|14875-9|LNC2HPO|Hyperphenylalaninemia|Hyperphenylalaninemia
C0798049|T201|LN|14875-9|LNC2HPO|Hyperphenylalaninemia|Hyperphenylalaninemia
C0798049|T201|DN|14875-9|LNC2HPO|Hyperphenylalaninemia|Hyperphenylalaninemia
C0798049|T201|OSN|14875-9|LNC2HPO|Hyperphenylalaninemia|Hyperphenylalaninemia
C0798049|T201|LC|14875-9|LNC2HPO|Hyperphenylalaninemia|Hyperphenylalaninemia
C0798049|T201|MTH_LN|14875-9|LNC2HPO|Hypophenylalaninemia|Hypophenylalaninemia
C0798049|T201|LN|14875-9|LNC2HPO|Hypophenylalaninemia|Hypophenylalaninemia
C0798049|T201|DN|14875-9|LNC2HPO|Hypophenylalaninemia|Hypophenylalaninemia
C0798049|T201|OSN|14875-9|LNC2HPO|Hypophenylalaninemia|Hypophenylalaninemia
C0798049|T201|LC|14875-9|LNC2HPO|Hypophenylalaninemia|Hypophenylalaninemia
C1543831|T201|LN|39789-3|LNC2HPO|Hyperkalemia|Hyperkalemia
C1543831|T201|DN|39789-3|LNC2HPO|Hyperkalemia|Hyperkalemia
C1543831|T201|OSN|39789-3|LNC2HPO|Hyperkalemia|Hyperkalemia
C1543831|T201|MTH_LN|39789-3|LNC2HPO|Hyperkalemia|Hyperkalemia
C1543831|T201|LC|39789-3|LNC2HPO|Hyperkalemia|Hyperkalemia
C1543831|T201|LN|39789-3|LNC2HPO|Hypokalemia|Hypokalemia
C1543831|T201|DN|39789-3|LNC2HPO|Hypokalemia|Hypokalemia
C1543831|T201|OSN|39789-3|LNC2HPO|Hypokalemia|Hypokalemia
C1543831|T201|MTH_LN|39789-3|LNC2HPO|Hypokalemia|Hypokalemia
C1543831|T201|LC|39789-3|LNC2HPO|Hypokalemia|Hypokalemia
C0803458|T201|LN|20655-7|LNC2HPO|Hyperprolinemia|Hyperprolinemia
C0803458|T201|MTH_LN|20655-7|LNC2HPO|Hyperprolinemia|Hyperprolinemia
C0803458|T201|DN|20655-7|LNC2HPO|Hyperprolinemia|Hyperprolinemia
C0803458|T201|OSN|20655-7|LNC2HPO|Hyperprolinemia|Hyperprolinemia
C0803458|T201|LC|20655-7|LNC2HPO|Hyperprolinemia|Hyperprolinemia
C0803458|T201|LN|20655-7|LNC2HPO|Prolinemia|Prolinemia
C0803458|T201|MTH_LN|20655-7|LNC2HPO|Prolinemia|Prolinemia
C0803458|T201|DN|20655-7|LNC2HPO|Prolinemia|Prolinemia
C0803458|T201|OSN|20655-7|LNC2HPO|Prolinemia|Prolinemia
C0803458|T201|LC|20655-7|LNC2HPO|Prolinemia|Prolinemia
C0803458|T201|LN|20655-7|LNC2HPO|Hypoprolinemia|Hypoprolinemia
C0803458|T201|MTH_LN|20655-7|LNC2HPO|Hypoprolinemia|Hypoprolinemia
C0803458|T201|DN|20655-7|LNC2HPO|Hypoprolinemia|Hypoprolinemia
C0803458|T201|OSN|20655-7|LNC2HPO|Hypoprolinemia|Hypoprolinemia
C0803458|T201|LC|20655-7|LNC2HPO|Hypoprolinemia|Hypoprolinemia
C0803459|T201|LN|20656-5|LNC2HPO|Hyperserinemia|Hyperserinemia
C0803459|T201|MTH_LN|20656-5|LNC2HPO|Hyperserinemia|Hyperserinemia
C0803459|T201|DN|20656-5|LNC2HPO|Hyperserinemia|Hyperserinemia
C0803459|T201|OSN|20656-5|LNC2HPO|Hyperserinemia|Hyperserinemia
C0803459|T201|LC|20656-5|LNC2HPO|Hyperserinemia|Hyperserinemia
C0803459|T201|LN|20656-5|LNC2HPO|Hyposerinemia|Hyposerinemia
C0803459|T201|MTH_LN|20656-5|LNC2HPO|Hyposerinemia|Hyposerinemia
C0803459|T201|DN|20656-5|LNC2HPO|Hyposerinemia|Hyposerinemia
C0803459|T201|OSN|20656-5|LNC2HPO|Hyposerinemia|Hyposerinemia
C0803459|T201|LC|20656-5|LNC2HPO|Hyposerinemia|Hyposerinemia
C0803461|T201|LN|20658-1|LNC2HPO|Hyperthreoninemia|Hyperthreoninemia
C0803461|T201|MTH_LN|20658-1|LNC2HPO|Hyperthreoninemia|Hyperthreoninemia
C0803461|T201|DN|20658-1|LNC2HPO|Hyperthreoninemia|Hyperthreoninemia
C0803461|T201|OSN|20658-1|LNC2HPO|Hyperthreoninemia|Hyperthreoninemia
C0803461|T201|LC|20658-1|LNC2HPO|Hyperthreoninemia|Hyperthreoninemia
C0803461|T201|LN|20658-1|LNC2HPO|Hypothreoninemia|Hypothreoninemia
C0803461|T201|MTH_LN|20658-1|LNC2HPO|Hypothreoninemia|Hypothreoninemia
C0803461|T201|DN|20658-1|LNC2HPO|Hypothreoninemia|Hypothreoninemia
C0803461|T201|OSN|20658-1|LNC2HPO|Hypothreoninemia|Hypothreoninemia
C0803461|T201|LC|20658-1|LNC2HPO|Hypothreoninemia|Hypothreoninemia
C0881709|T201|MTH_LN|20659-9|LNC2HPO|Hypertryptophanemia|Hypertryptophanemia
C0881709|T201|LN|20659-9|LNC2HPO|Hypertryptophanemia|Hypertryptophanemia
C0881709|T201|DN|20659-9|LNC2HPO|Hypertryptophanemia|Hypertryptophanemia
C0881709|T201|OSN|20659-9|LNC2HPO|Hypertryptophanemia|Hypertryptophanemia
C0881709|T201|LC|20659-9|LNC2HPO|Hypertryptophanemia|Hypertryptophanemia
C0881709|T201|MTH_LN|20659-9|LNC2HPO|Hypotryptophanemia|Hypotryptophanemia
C0881709|T201|LN|20659-9|LNC2HPO|Hypotryptophanemia|Hypotryptophanemia
C0881709|T201|DN|20659-9|LNC2HPO|Hypotryptophanemia|Hypotryptophanemia
C0881709|T201|OSN|20659-9|LNC2HPO|Hypotryptophanemia|Hypotryptophanemia
C0881709|T201|LC|20659-9|LNC2HPO|Hypotryptophanemia|Hypotryptophanemia
C0803463|T201|LN|20660-7|LNC2HPO|Hypertyrosinemia|Hypertyrosinemia
C0803463|T201|MTH_LN|20660-7|LNC2HPO|Hypertyrosinemia|Hypertyrosinemia
C0803463|T201|DN|20660-7|LNC2HPO|Hypertyrosinemia|Hypertyrosinemia
C0803463|T201|OSN|20660-7|LNC2HPO|Hypertyrosinemia|Hypertyrosinemia
C0803463|T201|LC|20660-7|LNC2HPO|Hypertyrosinemia|Hypertyrosinemia
C0803463|T201|LN|20660-7|LNC2HPO|Tyrosinemia|Tyrosinemia
C0803463|T201|MTH_LN|20660-7|LNC2HPO|Tyrosinemia|Tyrosinemia
C0803463|T201|DN|20660-7|LNC2HPO|Tyrosinemia|Tyrosinemia
C0803463|T201|OSN|20660-7|LNC2HPO|Tyrosinemia|Tyrosinemia
C0803463|T201|LC|20660-7|LNC2HPO|Tyrosinemia|Tyrosinemia
C0803463|T201|LN|20660-7|LNC2HPO|Hypotyrosinemia|Hypotyrosinemia
C0803463|T201|MTH_LN|20660-7|LNC2HPO|Hypotyrosinemia|Hypotyrosinemia
C0803463|T201|DN|20660-7|LNC2HPO|Hypotyrosinemia|Hypotyrosinemia
C0803463|T201|OSN|20660-7|LNC2HPO|Hypotyrosinemia|Hypotyrosinemia
C0803463|T201|LC|20660-7|LNC2HPO|Hypotyrosinemia|Hypotyrosinemia
C0803464|T201|LN|20661-5|LNC2HPO|Hypervalinemia|Hypervalinemia
C0803464|T201|MTH_LN|20661-5|LNC2HPO|Hypervalinemia|Hypervalinemia
C0803464|T201|DN|20661-5|LNC2HPO|Hypervalinemia|Hypervalinemia
C0803464|T201|OSN|20661-5|LNC2HPO|Hypervalinemia|Hypervalinemia
C0803464|T201|LC|20661-5|LNC2HPO|Hypervalinemia|Hypervalinemia
C0803464|T201|LN|20661-5|LNC2HPO|Hypovalinemia|Hypovalinemia
C0803464|T201|MTH_LN|20661-5|LNC2HPO|Hypovalinemia|Hypovalinemia
C0803464|T201|DN|20661-5|LNC2HPO|Hypovalinemia|Hypovalinemia
C0803464|T201|OSN|20661-5|LNC2HPO|Hypovalinemia|Hypovalinemia
C0803464|T201|LC|20661-5|LNC2HPO|Hypovalinemia|Hypovalinemia
C1114247|T201|LN|30386-7|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C1114247|T201|OSN|30386-7|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C1114247|T201|DN|30386-7|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C1114247|T201|MTH_LN|30386-7|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C1114247|T201|LC|30386-7|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C1114247|T201|LN|30386-7|LNC2HPO|Microcytosis|Microcytosis
C1114247|T201|OSN|30386-7|LNC2HPO|Microcytosis|Microcytosis
C1114247|T201|DN|30386-7|LNC2HPO|Microcytosis|Microcytosis
C1114247|T201|MTH_LN|30386-7|LNC2HPO|Microcytosis|Microcytosis
C1114247|T201|LC|30386-7|LNC2HPO|Microcytosis|Microcytosis
C0362905|T201|LN|784-9|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C0362905|T201|MTH_LN|784-9|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C0362905|T201|DN|784-9|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C0362905|T201|OSN|784-9|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C0362905|T201|LC|784-9|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C0362905|T201|LN|784-9|LNC2HPO|Microcytosis|Microcytosis
C0362905|T201|MTH_LN|784-9|LNC2HPO|Microcytosis|Microcytosis
C0362905|T201|DN|784-9|LNC2HPO|Microcytosis|Microcytosis
C0362905|T201|OSN|784-9|LNC2HPO|Microcytosis|Microcytosis
C0362905|T201|LC|784-9|LNC2HPO|Microcytosis|Microcytosis
C0364600|T201|LN|2460-4|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C0364600|T201|MTH_LN|2460-4|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C0364600|T201|DN|2460-4|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C0364600|T201|OSN|2460-4|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C0364600|T201|LC|2460-4|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C0364600|T201|LN|2460-4|LNC2HPO|IgD deficiency|IgD deficiency
C0364600|T201|MTH_LN|2460-4|LNC2HPO|IgD deficiency|IgD deficiency
C0364600|T201|DN|2460-4|LNC2HPO|IgD deficiency|IgD deficiency
C0364600|T201|OSN|2460-4|LNC2HPO|IgD deficiency|IgD deficiency
C0364600|T201|LC|2460-4|LNC2HPO|IgD deficiency|IgD deficiency
C0364601|T201|LN|2461-2|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C0364601|T201|MTH_LN|2461-2|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C0364601|T201|DN|2461-2|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C0364601|T201|OSN|2461-2|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C0364601|T201|LC|2461-2|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C0364601|T201|LN|2461-2|LNC2HPO|IgD deficiency|IgD deficiency
C0364601|T201|MTH_LN|2461-2|LNC2HPO|IgD deficiency|IgD deficiency
C0364601|T201|DN|2461-2|LNC2HPO|IgD deficiency|IgD deficiency
C0364601|T201|OSN|2461-2|LNC2HPO|IgD deficiency|IgD deficiency
C0364601|T201|LC|2461-2|LNC2HPO|IgD deficiency|IgD deficiency
C2733775|T201|LN|56688-5|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C2733775|T201|DN|56688-5|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C2733775|T201|LC|56688-5|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C2733775|T201|MTH_LN|56688-5|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C2733775|T201|OSN|56688-5|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C2733775|T201|LN|56688-5|LNC2HPO|IgD deficiency|IgD deficiency
C2733775|T201|DN|56688-5|LNC2HPO|IgD deficiency|IgD deficiency
C2733775|T201|LC|56688-5|LNC2HPO|IgD deficiency|IgD deficiency
C2733775|T201|MTH_LN|56688-5|LNC2HPO|IgD deficiency|IgD deficiency
C2733775|T201|OSN|56688-5|LNC2HPO|IgD deficiency|IgD deficiency
C1715862|T201|LN|44592-4|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C1715862|T201|MTH_LN|44592-4|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C1715862|T201|DN|44592-4|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C1715862|T201|OSN|44592-4|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C1715862|T201|LC|44592-4|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C2733880|T201|LN|55903-9|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C2733880|T201|MTH_LN|55903-9|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C2733880|T201|DN|55903-9|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C2733880|T201|LC|55903-9|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C2733880|T201|OSN|55903-9|LNC2HPO|IgD hypergammaglobulinemia|IgD hypergammaglobulinemia
C0797024|T201|LN|13834-7|LNC2HPO|IgE deficiency|IgE deficiency
C0797024|T201|MTH_LN|13834-7|LNC2HPO|IgE deficiency|IgE deficiency
C0797024|T201|OSN|13834-7|LNC2HPO|IgE deficiency|IgE deficiency
C0797024|T201|DN|13834-7|LNC2HPO|IgE deficiency|IgE deficiency
C0797024|T201|LC|13834-7|LNC2HPO|IgE deficiency|IgE deficiency
C0942471|T201|LN|26511-6|LNC2HPO|Neutrophilia|Neutrophilia
C0942471|T201|OSN|26511-6|LNC2HPO|Neutrophilia|Neutrophilia
C0942471|T201|DN|26511-6|LNC2HPO|Neutrophilia|Neutrophilia
C0942471|T201|MTH_LN|26511-6|LNC2HPO|Neutrophilia|Neutrophilia
C0942471|T201|LC|26511-6|LNC2HPO|Neutrophilia|Neutrophilia
C0942471|T201|LN|26511-6|LNC2HPO|Neutropenia|Neutropenia
C0942471|T201|OSN|26511-6|LNC2HPO|Neutropenia|Neutropenia
C0942471|T201|DN|26511-6|LNC2HPO|Neutropenia|Neutropenia
C0942471|T201|MTH_LN|26511-6|LNC2HPO|Neutropenia|Neutropenia
C0942471|T201|LC|26511-6|LNC2HPO|Neutropenia|Neutropenia
C0942471|T201|LN|26511-6|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0942471|T201|OSN|26511-6|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0942471|T201|DN|26511-6|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0942471|T201|MTH_LN|26511-6|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0942471|T201|LC|26511-6|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0364605|T201|LN|2465-3|LNC2HPO|IgG deficiency|IgG deficiency
C0364605|T201|LC|2465-3|LNC2HPO|IgG deficiency|IgG deficiency
C0364605|T201|OSN|2465-3|LNC2HPO|IgG deficiency|IgG deficiency
C0364605|T201|MTH_LN|2465-3|LNC2HPO|IgG deficiency|IgG deficiency
C0364605|T201|DN|2465-3|LNC2HPO|IgG deficiency|IgG deficiency
C0942474|T201|LN|26515-7|LNC2HPO|Thrombocytosis|Thrombocytosis
C0942474|T201|DN|26515-7|LNC2HPO|Thrombocytosis|Thrombocytosis
C0942474|T201|OSN|26515-7|LNC2HPO|Thrombocytosis|Thrombocytosis
C0942474|T201|MTH_LN|26515-7|LNC2HPO|Thrombocytosis|Thrombocytosis
C0942474|T201|LC|26515-7|LNC2HPO|Thrombocytosis|Thrombocytosis
C0942474|T201|LN|26515-7|LNC2HPO|Thrombocythemia|Thrombocythemia
C0942474|T201|DN|26515-7|LNC2HPO|Thrombocythemia|Thrombocythemia
C0942474|T201|OSN|26515-7|LNC2HPO|Thrombocythemia|Thrombocythemia
C0942474|T201|MTH_LN|26515-7|LNC2HPO|Thrombocythemia|Thrombocythemia
C0942474|T201|LC|26515-7|LNC2HPO|Thrombocythemia|Thrombocythemia
C0942474|T201|LN|26515-7|LNC2HPO|Thrombocythaemia|Thrombocythaemia
C0942474|T201|DN|26515-7|LNC2HPO|Thrombocythaemia|Thrombocythaemia
C0942474|T201|OSN|26515-7|LNC2HPO|Thrombocythaemia|Thrombocythaemia
C0942474|T201|MTH_LN|26515-7|LNC2HPO|Thrombocythaemia|Thrombocythaemia
C0942474|T201|LC|26515-7|LNC2HPO|Thrombocythaemia|Thrombocythaemia
C0942474|T201|LN|26515-7|LNC2HPO|Thrombocytopenia|Thrombocytopenia
C0942474|T201|DN|26515-7|LNC2HPO|Thrombocytopenia|Thrombocytopenia
C0942474|T201|OSN|26515-7|LNC2HPO|Thrombocytopenia|Thrombocytopenia
C0942474|T201|MTH_LN|26515-7|LNC2HPO|Thrombocytopenia|Thrombocytopenia
C0942474|T201|LC|26515-7|LNC2HPO|Thrombocytopenia|Thrombocytopenia
C0482691|T201|LN|6301-6|LNC2HPO|Prolonged prothrombin time|Prolonged prothrombin time
C0482691|T201|DN|6301-6|LNC2HPO|Prolonged prothrombin time|Prolonged prothrombin time
C0482691|T201|MTH_LN|6301-6|LNC2HPO|Prolonged prothrombin time|Prolonged prothrombin time
C0482691|T201|LC|6301-6|LNC2HPO|Prolonged prothrombin time|Prolonged prothrombin time
C0482691|T201|OSN|6301-6|LNC2HPO|Prolonged prothrombin time|Prolonged prothrombin time
C0482691|T201|LN|6301-6|LNC2HPO|Prolonged PT|Prolonged PT
C0482691|T201|DN|6301-6|LNC2HPO|Prolonged PT|Prolonged PT
C0482691|T201|MTH_LN|6301-6|LNC2HPO|Prolonged PT|Prolonged PT
C0482691|T201|LC|6301-6|LNC2HPO|Prolonged PT|Prolonged PT
C0482691|T201|OSN|6301-6|LNC2HPO|Prolonged PT|Prolonged PT
C0482691|T201|LN|6301-6|LNC2HPO|increased international normalised ratio|increased international normalised ratio
C0482691|T201|DN|6301-6|LNC2HPO|increased international normalised ratio|increased international normalised ratio
C0482691|T201|MTH_LN|6301-6|LNC2HPO|increased international normalised ratio|increased international normalised ratio
C0482691|T201|LC|6301-6|LNC2HPO|increased international normalised ratio|increased international normalised ratio
C0482691|T201|OSN|6301-6|LNC2HPO|increased international normalised ratio|increased international normalised ratio
C0368018|T201|LN|5792-7|LNC2HPO|Glycosuria|Glycosuria
C0368018|T201|MTH_LN|5792-7|LNC2HPO|Glycosuria|Glycosuria
C0368018|T201|DN|5792-7|LNC2HPO|Glycosuria|Glycosuria
C0368018|T201|OSN|5792-7|LNC2HPO|Glycosuria|Glycosuria
C0368018|T201|LC|5792-7|LNC2HPO|Glycosuria|Glycosuria
C0368018|T201|LN|5792-7|LNC2HPO|Glucosuria|Glucosuria
C0368018|T201|MTH_LN|5792-7|LNC2HPO|Glucosuria|Glucosuria
C0368018|T201|DN|5792-7|LNC2HPO|Glucosuria|Glucosuria
C0368018|T201|OSN|5792-7|LNC2HPO|Glucosuria|Glucosuria
C0368018|T201|LC|5792-7|LNC2HPO|Glucosuria|Glucosuria
C0368043|T201|LN|5804-0|LNC2HPO|Proteinuria|Proteinuria
C0368043|T201|MTH_LN|5804-0|LNC2HPO|Proteinuria|Proteinuria
C0368043|T201|DN|5804-0|LNC2HPO|Proteinuria|Proteinuria
C0368043|T201|OSN|5804-0|LNC2HPO|Proteinuria|Proteinuria
C0368043|T201|LC|5804-0|LNC2HPO|Proteinuria|Proteinuria
C0364745|T201|MTH_LN|2601-3|LNC2HPO|Hypermagnesemia|Hypermagnesemia
C0364745|T201|LN|2601-3|LNC2HPO|Hypermagnesemia|Hypermagnesemia
C0364745|T201|DN|2601-3|LNC2HPO|Hypermagnesemia|Hypermagnesemia
C0364745|T201|OSN|2601-3|LNC2HPO|Hypermagnesemia|Hypermagnesemia
C0364745|T201|LC|2601-3|LNC2HPO|Hypermagnesemia|Hypermagnesemia
C0364745|T201|MTH_LN|2601-3|LNC2HPO|Hypomagnesemia|Hypomagnesemia
C0364745|T201|LN|2601-3|LNC2HPO|Hypomagnesemia|Hypomagnesemia
C0364745|T201|DN|2601-3|LNC2HPO|Hypomagnesemia|Hypomagnesemia
C0364745|T201|OSN|2601-3|LNC2HPO|Hypomagnesemia|Hypomagnesemia
C0364745|T201|LC|2601-3|LNC2HPO|Hypomagnesemia|Hypomagnesemia
C0550246|T201|LN|11557-6|LNC2HPO|Hypercapnia|Hypercapnia
C0550246|T201|LC|11557-6|LNC2HPO|Hypercapnia|Hypercapnia
C0550246|T201|MTH_LN|11557-6|LNC2HPO|Hypercapnia|Hypercapnia
C0550246|T201|DN|11557-6|LNC2HPO|Hypercapnia|Hypercapnia
C0550246|T201|OSN|11557-6|LNC2HPO|Hypercapnia|Hypercapnia
C0550246|T201|LN|11557-6|LNC2HPO|Hypercarbia|Hypercarbia
C0550246|T201|LC|11557-6|LNC2HPO|Hypercarbia|Hypercarbia
C0550246|T201|MTH_LN|11557-6|LNC2HPO|Hypercarbia|Hypercarbia
C0550246|T201|DN|11557-6|LNC2HPO|Hypercarbia|Hypercarbia
C0550246|T201|OSN|11557-6|LNC2HPO|Hypercarbia|Hypercarbia
C0550246|T201|LN|11557-6|LNC2HPO|Hypocapnia|Hypocapnia
C0550246|T201|LC|11557-6|LNC2HPO|Hypocapnia|Hypocapnia
C0550246|T201|MTH_LN|11557-6|LNC2HPO|Hypocapnia|Hypocapnia
C0550246|T201|DN|11557-6|LNC2HPO|Hypocapnia|Hypocapnia
C0550246|T201|OSN|11557-6|LNC2HPO|Hypocapnia|Hypocapnia
C0550246|T201|LN|11557-6|LNC2HPO|Hypocarbia|Hypocarbia
C0550246|T201|LC|11557-6|LNC2HPO|Hypocarbia|Hypocarbia
C0550246|T201|MTH_LN|11557-6|LNC2HPO|Hypocarbia|Hypocarbia
C0550246|T201|DN|11557-6|LNC2HPO|Hypocarbia|Hypocarbia
C0550246|T201|OSN|11557-6|LNC2HPO|Hypocarbia|Hypocarbia
C0550440|T201|LN|11556-8|LNC2HPO|Hyperoxemia|Hyperoxemia
C0550440|T201|LC|11556-8|LNC2HPO|Hyperoxemia|Hyperoxemia
C0550440|T201|MTH_LN|11556-8|LNC2HPO|Hyperoxemia|Hyperoxemia
C0550440|T201|DN|11556-8|LNC2HPO|Hyperoxemia|Hyperoxemia
C0550440|T201|OSN|11556-8|LNC2HPO|Hyperoxemia|Hyperoxemia
C0550440|T201|LN|11556-8|LNC2HPO|Hypoxemia|Hypoxemia
C0550440|T201|LC|11556-8|LNC2HPO|Hypoxemia|Hypoxemia
C0550440|T201|MTH_LN|11556-8|LNC2HPO|Hypoxemia|Hypoxemia
C0550440|T201|DN|11556-8|LNC2HPO|Hypoxemia|Hypoxemia
C0550440|T201|OSN|11556-8|LNC2HPO|Hypoxemia|Hypoxemia
C0550447|T201|LN|11558-4|LNC2HPO|Acid base imbalance|Acid base imbalance
C0550447|T201|LC|11558-4|LNC2HPO|Acid base imbalance|Acid base imbalance
C0550447|T201|MTH_LN|11558-4|LNC2HPO|Acid base imbalance|Acid base imbalance
C0550447|T201|OSN|11558-4|LNC2HPO|Acid base imbalance|Acid base imbalance
C0550447|T201|DN|11558-4|LNC2HPO|Acid base imbalance|Acid base imbalance
C0550447|T201|LN|11558-4|LNC2HPO|Alkalemia|Alkalemia
C0550447|T201|LC|11558-4|LNC2HPO|Alkalemia|Alkalemia
C0550447|T201|MTH_LN|11558-4|LNC2HPO|Alkalemia|Alkalemia
C0550447|T201|OSN|11558-4|LNC2HPO|Alkalemia|Alkalemia
C0550447|T201|DN|11558-4|LNC2HPO|Alkalemia|Alkalemia
C0550447|T201|LN|11558-4|LNC2HPO|Acidemia|Acidemia
C0550447|T201|LC|11558-4|LNC2HPO|Acidemia|Acidemia
C0550447|T201|MTH_LN|11558-4|LNC2HPO|Acidemia|Acidemia
C0550447|T201|OSN|11558-4|LNC2HPO|Acidemia|Acidemia
C0550447|T201|DN|11558-4|LNC2HPO|Acidemia|Acidemia
C0364104|T201|LC|1971-1|LNC2HPO|Hyperbilirubinemia|Hyperbilirubinemia
C0364104|T201|MTH_LN|1971-1|LNC2HPO|Hyperbilirubinemia|Hyperbilirubinemia
C0364104|T201|LN|1971-1|LNC2HPO|Hyperbilirubinemia|Hyperbilirubinemia
C0364104|T201|DN|1971-1|LNC2HPO|Hyperbilirubinemia|Hyperbilirubinemia
C0364104|T201|OSN|1971-1|LNC2HPO|Hyperbilirubinemia|Hyperbilirubinemia
C0487995|T201|MTH_LN|8310-5|LNC2HPO|Body temperature changes|Body temperature changes
C0487995|T201|LC|8310-5|LNC2HPO|Body temperature changes|Body temperature changes
C0487995|T201|OSN|8310-5|LNC2HPO|Body temperature changes|Body temperature changes
C0487995|T201|LN|8310-5|LNC2HPO|Body temperature changes|Body temperature changes
C0487995|T201|MTH_LN|8310-5|LNC2HPO|Poor temperature regulation|Poor temperature regulation
C0487995|T201|LC|8310-5|LNC2HPO|Poor temperature regulation|Poor temperature regulation
C0487995|T201|OSN|8310-5|LNC2HPO|Poor temperature regulation|Poor temperature regulation
C0487995|T201|LN|8310-5|LNC2HPO|Poor temperature regulation|Poor temperature regulation
C0487995|T201|MTH_LN|8310-5|LNC2HPO|Fever|Fever
C0487995|T201|LC|8310-5|LNC2HPO|Fever|Fever
C0487995|T201|OSN|8310-5|LNC2HPO|Fever|Fever
C0487995|T201|LN|8310-5|LNC2HPO|Fever|Fever
C0487995|T201|MTH_LN|8310-5|LNC2HPO|Hyperthermia|Hyperthermia
C0487995|T201|LC|8310-5|LNC2HPO|Hyperthermia|Hyperthermia
C0487995|T201|OSN|8310-5|LNC2HPO|Hyperthermia|Hyperthermia
C0487995|T201|LN|8310-5|LNC2HPO|Hyperthermia|Hyperthermia
C0487995|T201|MTH_LN|8310-5|LNC2HPO|Pyrexia|Pyrexia
C0487995|T201|LC|8310-5|LNC2HPO|Pyrexia|Pyrexia
C0487995|T201|OSN|8310-5|LNC2HPO|Pyrexia|Pyrexia
C0487995|T201|LN|8310-5|LNC2HPO|Pyrexia|Pyrexia
C0487995|T201|MTH_LN|8310-5|LNC2HPO|Hypothermia|Hypothermia
C0487995|T201|LC|8310-5|LNC2HPO|Hypothermia|Hypothermia
C0487995|T201|OSN|8310-5|LNC2HPO|Hypothermia|Hypothermia
C0487995|T201|LN|8310-5|LNC2HPO|Hypothermia|Hypothermia
C0803374|T201|LN|20565-8|LNC2HPO|Hypercapnia|Hypercapnia
C0803374|T201|MTH_LN|20565-8|LNC2HPO|Hypercapnia|Hypercapnia
C0803374|T201|DN|20565-8|LNC2HPO|Hypercapnia|Hypercapnia
C0803374|T201|OSN|20565-8|LNC2HPO|Hypercapnia|Hypercapnia
C0803374|T201|LC|20565-8|LNC2HPO|Hypercapnia|Hypercapnia
C0803374|T201|LN|20565-8|LNC2HPO|Hypercarbia|Hypercarbia
C0803374|T201|MTH_LN|20565-8|LNC2HPO|Hypercarbia|Hypercarbia
C0803374|T201|DN|20565-8|LNC2HPO|Hypercarbia|Hypercarbia
C0803374|T201|OSN|20565-8|LNC2HPO|Hypercarbia|Hypercarbia
C0803374|T201|LC|20565-8|LNC2HPO|Hypercarbia|Hypercarbia
C0803374|T201|LN|20565-8|LNC2HPO|Hypocapnia|Hypocapnia
C0803374|T201|MTH_LN|20565-8|LNC2HPO|Hypocapnia|Hypocapnia
C0803374|T201|DN|20565-8|LNC2HPO|Hypocapnia|Hypocapnia
C0803374|T201|OSN|20565-8|LNC2HPO|Hypocapnia|Hypocapnia
C0803374|T201|LC|20565-8|LNC2HPO|Hypocapnia|Hypocapnia
C0803374|T201|LN|20565-8|LNC2HPO|Hypocarbia|Hypocarbia
C0803374|T201|MTH_LN|20565-8|LNC2HPO|Hypocarbia|Hypocarbia
C0803374|T201|DN|20565-8|LNC2HPO|Hypocarbia|Hypocarbia
C0803374|T201|OSN|20565-8|LNC2HPO|Hypocarbia|Hypocarbia
C0803374|T201|LC|20565-8|LNC2HPO|Hypocarbia|Hypocarbia
C0364896|T201|LN|2753-2|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364896|T201|DN|2753-2|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364896|T201|MTH_LN|2753-2|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364896|T201|OSN|2753-2|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364896|T201|LC|2753-2|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364896|T201|LN|2753-2|LNC2HPO|Alkalosis|Alkalosis
C0364896|T201|DN|2753-2|LNC2HPO|Alkalosis|Alkalosis
C0364896|T201|MTH_LN|2753-2|LNC2HPO|Alkalosis|Alkalosis
C0364896|T201|OSN|2753-2|LNC2HPO|Alkalosis|Alkalosis
C0364896|T201|LC|2753-2|LNC2HPO|Alkalosis|Alkalosis
C0364896|T201|LN|2753-2|LNC2HPO|Acidosis|Acidosis
C0364896|T201|DN|2753-2|LNC2HPO|Acidosis|Acidosis
C0364896|T201|MTH_LN|2753-2|LNC2HPO|Acidosis|Acidosis
C0364896|T201|OSN|2753-2|LNC2HPO|Acidosis|Acidosis
C0364896|T201|LC|2753-2|LNC2HPO|Acidosis|Acidosis
C1369580|T201|LN|34714-6|LNC2HPO|Impaired platelet aggregation|Impaired platelet aggregation
C1369580|T201|DN|34714-6|LNC2HPO|Impaired platelet aggregation|Impaired platelet aggregation
C1369580|T201|MTH_LN|34714-6|LNC2HPO|Impaired platelet aggregation|Impaired platelet aggregation
C1369580|T201|LC|34714-6|LNC2HPO|Impaired platelet aggregation|Impaired platelet aggregation
C1369580|T201|OSN|34714-6|LNC2HPO|Impaired platelet aggregation|Impaired platelet aggregation
C1369580|T201|LN|34714-6|LNC2HPO|Defective platelet aggregation|Defective platelet aggregation
C1369580|T201|DN|34714-6|LNC2HPO|Defective platelet aggregation|Defective platelet aggregation
C1369580|T201|MTH_LN|34714-6|LNC2HPO|Defective platelet aggregation|Defective platelet aggregation
C1369580|T201|LC|34714-6|LNC2HPO|Defective platelet aggregation|Defective platelet aggregation
C1369580|T201|OSN|34714-6|LNC2HPO|Defective platelet aggregation|Defective platelet aggregation
C1369580|T201|LN|34714-6|LNC2HPO|Deficient platelet aggregation|Deficient platelet aggregation
C1369580|T201|DN|34714-6|LNC2HPO|Deficient platelet aggregation|Deficient platelet aggregation
C1369580|T201|MTH_LN|34714-6|LNC2HPO|Deficient platelet aggregation|Deficient platelet aggregation
C1369580|T201|LC|34714-6|LNC2HPO|Deficient platelet aggregation|Deficient platelet aggregation
C1369580|T201|OSN|34714-6|LNC2HPO|Deficient platelet aggregation|Deficient platelet aggregation
C1369580|T201|LN|34714-6|LNC2HPO|Platelet aggregation defect|Platelet aggregation defect
C1369580|T201|DN|34714-6|LNC2HPO|Platelet aggregation defect|Platelet aggregation defect
C1369580|T201|MTH_LN|34714-6|LNC2HPO|Platelet aggregation defect|Platelet aggregation defect
C1369580|T201|LC|34714-6|LNC2HPO|Platelet aggregation defect|Platelet aggregation defect
C1369580|T201|OSN|34714-6|LNC2HPO|Platelet aggregation defect|Platelet aggregation defect
C0798351|T201|LN|15180-3|LNC2HPO|Hypochromic anemia|Hypochromic anemia
C0798351|T201|MTH_LN|15180-3|LNC2HPO|Hypochromic anemia|Hypochromic anemia
C0798351|T201|OSN|15180-3|LNC2HPO|Hypochromic anemia|Hypochromic anemia
C0798351|T201|DN|15180-3|LNC2HPO|Hypochromic anemia|Hypochromic anemia
C0798351|T201|LC|15180-3|LNC2HPO|Hypochromic anemia|Hypochromic anemia
C0798351|T201|LN|15180-3|LNC2HPO|Hypochromic anaemia|Hypochromic anaemia
C0798351|T201|MTH_LN|15180-3|LNC2HPO|Hypochromic anaemia|Hypochromic anaemia
C0798351|T201|OSN|15180-3|LNC2HPO|Hypochromic anaemia|Hypochromic anaemia
C0798351|T201|DN|15180-3|LNC2HPO|Hypochromic anaemia|Hypochromic anaemia
C0798351|T201|LC|15180-3|LNC2HPO|Hypochromic anaemia|Hypochromic anaemia
C0364598|T201|LN|2458-8|LNC2HPO|IgA hypergammaglobulinemia|IgA hypergammaglobulinemia
C0364598|T201|OSN|2458-8|LNC2HPO|IgA hypergammaglobulinemia|IgA hypergammaglobulinemia
C0364598|T201|LC|2458-8|LNC2HPO|IgA hypergammaglobulinemia|IgA hypergammaglobulinemia
C0364598|T201|MTH_LN|2458-8|LNC2HPO|IgA hypergammaglobulinemia|IgA hypergammaglobulinemia
C0364598|T201|DN|2458-8|LNC2HPO|IgA hypergammaglobulinemia|IgA hypergammaglobulinemia
C0364598|T201|LN|2458-8|LNC2HPO|IgA deficiency|IgA deficiency
C0364598|T201|OSN|2458-8|LNC2HPO|IgA deficiency|IgA deficiency
C0364598|T201|LC|2458-8|LNC2HPO|IgA deficiency|IgA deficiency
C0364598|T201|MTH_LN|2458-8|LNC2HPO|IgA deficiency|IgA deficiency
C0364598|T201|DN|2458-8|LNC2HPO|IgA deficiency|IgA deficiency
C0364598|T201|LN|2458-8|LNC2HPO|Gamma-A globulin deficiency|Gamma-A globulin deficiency
C0364598|T201|OSN|2458-8|LNC2HPO|Gamma-A globulin deficiency|Gamma-A globulin deficiency
C0364598|T201|LC|2458-8|LNC2HPO|Gamma-A globulin deficiency|Gamma-A globulin deficiency
C0364598|T201|MTH_LN|2458-8|LNC2HPO|Gamma-A globulin deficiency|Gamma-A globulin deficiency
C0364598|T201|DN|2458-8|LNC2HPO|Gamma-A globulin deficiency|Gamma-A globulin deficiency
C0365034|T201|LN|2890-2|LNC2HPO|Proteinuria|Proteinuria
C0365034|T201|OSN|2890-2|LNC2HPO|Proteinuria|Proteinuria
C0365034|T201|MTH_LN|2890-2|LNC2HPO|Proteinuria|Proteinuria
C0365034|T201|DN|2890-2|LNC2HPO|Proteinuria|Proteinuria
C0365034|T201|LC|2890-2|LNC2HPO|Proteinuria|Proteinuria
C0364655|T201|LN|2514-8|LNC2HPO|Ketonuria|Ketonuria
C0364655|T201|MTH_LN|2514-8|LNC2HPO|Ketonuria|Ketonuria
C0364655|T201|DN|2514-8|LNC2HPO|Ketonuria|Ketonuria
C0364655|T201|OSN|2514-8|LNC2HPO|Ketonuria|Ketonuria
C0364655|T201|LC|2514-8|LNC2HPO|Ketonuria|Ketonuria
C0364655|T201|LN|2514-8|LNC2HPO|Acetonuria|Acetonuria
C0364655|T201|MTH_LN|2514-8|LNC2HPO|Acetonuria|Acetonuria
C0364655|T201|DN|2514-8|LNC2HPO|Acetonuria|Acetonuria
C0364655|T201|OSN|2514-8|LNC2HPO|Acetonuria|Acetonuria
C0364655|T201|LC|2514-8|LNC2HPO|Acetonuria|Acetonuria
C0364655|T201|LN|2514-8|LNC2HPO|Ketoaciduria|Ketoaciduria
C0364655|T201|MTH_LN|2514-8|LNC2HPO|Ketoaciduria|Ketoaciduria
C0364655|T201|DN|2514-8|LNC2HPO|Ketoaciduria|Ketoaciduria
C0364655|T201|OSN|2514-8|LNC2HPO|Ketoaciduria|Ketoaciduria
C0364655|T201|LC|2514-8|LNC2HPO|Ketoaciduria|Ketoaciduria
C0364655|T201|LN|2514-8|LNC2HPO|Ketonaciduria|Ketonaciduria
C0364655|T201|MTH_LN|2514-8|LNC2HPO|Ketonaciduria|Ketonaciduria
C0364655|T201|DN|2514-8|LNC2HPO|Ketonaciduria|Ketonaciduria
C0364655|T201|OSN|2514-8|LNC2HPO|Ketonaciduria|Ketonaciduria
C0364655|T201|LC|2514-8|LNC2HPO|Ketonaciduria|Ketonaciduria
C0364127|T201|LN|1994-3|LNC2HPO|Hypercalcemia|Hypercalcemia
C0364127|T201|DN|1994-3|LNC2HPO|Hypercalcemia|Hypercalcemia
C0364127|T201|MTH_LN|1994-3|LNC2HPO|Hypercalcemia|Hypercalcemia
C0364127|T201|OSN|1994-3|LNC2HPO|Hypercalcemia|Hypercalcemia
C0364127|T201|LC|1994-3|LNC2HPO|Hypercalcemia|Hypercalcemia
C0364127|T201|LN|1994-3|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0364127|T201|DN|1994-3|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0364127|T201|MTH_LN|1994-3|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0364127|T201|OSN|1994-3|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0364127|T201|LC|1994-3|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0364127|T201|LN|1994-3|LNC2HPO|Hypocalcemia|Hypocalcemia
C0364127|T201|DN|1994-3|LNC2HPO|Hypocalcemia|Hypocalcemia
C0364127|T201|MTH_LN|1994-3|LNC2HPO|Hypocalcemia|Hypocalcemia
C0364127|T201|OSN|1994-3|LNC2HPO|Hypocalcemia|Hypocalcemia
C0364127|T201|LC|1994-3|LNC2HPO|Hypocalcemia|Hypocalcemia
C0364127|T201|LN|1994-3|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364127|T201|DN|1994-3|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364127|T201|MTH_LN|1994-3|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364127|T201|OSN|1994-3|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364127|T201|LC|1994-3|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364128|T201|LN|1995-0|LNC2HPO|Hypercalcemia|Hypercalcemia
C0364128|T201|DN|1995-0|LNC2HPO|Hypercalcemia|Hypercalcemia
C0364128|T201|MTH_LN|1995-0|LNC2HPO|Hypercalcemia|Hypercalcemia
C0364128|T201|OSN|1995-0|LNC2HPO|Hypercalcemia|Hypercalcemia
C0364128|T201|LC|1995-0|LNC2HPO|Hypercalcemia|Hypercalcemia
C0364128|T201|LN|1995-0|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0364128|T201|DN|1995-0|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0364128|T201|MTH_LN|1995-0|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0364128|T201|OSN|1995-0|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0364128|T201|LC|1995-0|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0364128|T201|LN|1995-0|LNC2HPO|Hypocalcemia|Hypocalcemia
C0364128|T201|DN|1995-0|LNC2HPO|Hypocalcemia|Hypocalcemia
C0364128|T201|MTH_LN|1995-0|LNC2HPO|Hypocalcemia|Hypocalcemia
C0364128|T201|OSN|1995-0|LNC2HPO|Hypocalcemia|Hypocalcemia
C0364128|T201|LC|1995-0|LNC2HPO|Hypocalcemia|Hypocalcemia
C0364128|T201|LN|1995-0|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364128|T201|DN|1995-0|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364128|T201|MTH_LN|1995-0|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364128|T201|OSN|1995-0|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364128|T201|LC|1995-0|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0944746|T201|LN|29265-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0944746|T201|DN|29265-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0944746|T201|MTH_LN|29265-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0944746|T201|OSN|29265-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0944746|T201|LC|29265-6|LNC2HPO|Hypercalcemia|Hypercalcemia
C0944746|T201|LN|29265-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0944746|T201|DN|29265-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0944746|T201|MTH_LN|29265-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0944746|T201|OSN|29265-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0944746|T201|LC|29265-6|LNC2HPO|Hypercalcaemia|Hypercalcaemia
C0944746|T201|LN|29265-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0944746|T201|DN|29265-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0944746|T201|MTH_LN|29265-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0944746|T201|OSN|29265-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0944746|T201|LC|29265-6|LNC2HPO|Hypocalcemia|Hypocalcemia
C0944746|T201|LN|29265-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0944746|T201|DN|29265-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0944746|T201|MTH_LN|29265-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0944746|T201|OSN|29265-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0944746|T201|LC|29265-6|LNC2HPO|Hypocalcaemia|Hypocalcaemia
C0364851|T201|LN|2708-6|LNC2HPO|Hyperoxemia|Hyperoxemia
C0364851|T201|DN|2708-6|LNC2HPO|Hyperoxemia|Hyperoxemia
C0364851|T201|LC|2708-6|LNC2HPO|Hyperoxemia|Hyperoxemia
C0364851|T201|MTH_LN|2708-6|LNC2HPO|Hyperoxemia|Hyperoxemia
C0364851|T201|OSN|2708-6|LNC2HPO|Hyperoxemia|Hyperoxemia
C0364851|T201|LN|2708-6|LNC2HPO|Hypoxemia|Hypoxemia
C0364851|T201|DN|2708-6|LNC2HPO|Hypoxemia|Hypoxemia
C0364851|T201|LC|2708-6|LNC2HPO|Hypoxemia|Hypoxemia
C0364851|T201|MTH_LN|2708-6|LNC2HPO|Hypoxemia|Hypoxemia
C0364851|T201|OSN|2708-6|LNC2HPO|Hypoxemia|Hypoxemia
C1145645|T201|LN|2703-7|LNC2HPO|Hyperoxemia|Hyperoxemia
C1145645|T201|MTH_LN|2703-7|LNC2HPO|Hyperoxemia|Hyperoxemia
C1145645|T201|DN|2703-7|LNC2HPO|Hyperoxemia|Hyperoxemia
C1145645|T201|LC|2703-7|LNC2HPO|Hyperoxemia|Hyperoxemia
C1145645|T201|OSN|2703-7|LNC2HPO|Hyperoxemia|Hyperoxemia
C1145645|T201|LN|2703-7|LNC2HPO|Hypoxemia|Hypoxemia
C1145645|T201|MTH_LN|2703-7|LNC2HPO|Hypoxemia|Hypoxemia
C1145645|T201|DN|2703-7|LNC2HPO|Hypoxemia|Hypoxemia
C1145645|T201|LC|2703-7|LNC2HPO|Hypoxemia|Hypoxemia
C1145645|T201|OSN|2703-7|LNC2HPO|Hypoxemia|Hypoxemia
C0362987|T201|LN|770-8|LNC2HPO|Neutrophilia|Neutrophilia
C0362987|T201|MTH_LN|770-8|LNC2HPO|Neutrophilia|Neutrophilia
C0362987|T201|OSN|770-8|LNC2HPO|Neutrophilia|Neutrophilia
C0362987|T201|DN|770-8|LNC2HPO|Neutrophilia|Neutrophilia
C0362987|T201|LC|770-8|LNC2HPO|Neutrophilia|Neutrophilia
C0362987|T201|LN|770-8|LNC2HPO|Neutropenia|Neutropenia
C0362987|T201|MTH_LN|770-8|LNC2HPO|Neutropenia|Neutropenia
C0362987|T201|OSN|770-8|LNC2HPO|Neutropenia|Neutropenia
C0362987|T201|DN|770-8|LNC2HPO|Neutropenia|Neutropenia
C0362987|T201|LC|770-8|LNC2HPO|Neutropenia|Neutropenia
C0362987|T201|LN|770-8|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0362987|T201|MTH_LN|770-8|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0362987|T201|OSN|770-8|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0362987|T201|DN|770-8|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0362987|T201|LC|770-8|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C1114281|T201|LN|30428-7|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C1114281|T201|OSN|30428-7|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C1114281|T201|LC|30428-7|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C1114281|T201|DN|30428-7|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C1114281|T201|MTH_LN|30428-7|LNC2HPO|Erythrocyte macrocytosis|Erythrocyte macrocytosis
C1114281|T201|LN|30428-7|LNC2HPO|Microcytosis|Microcytosis
C1114281|T201|OSN|30428-7|LNC2HPO|Microcytosis|Microcytosis
C1114281|T201|LC|30428-7|LNC2HPO|Microcytosis|Microcytosis
C1114281|T201|DN|30428-7|LNC2HPO|Microcytosis|Microcytosis
C1114281|T201|MTH_LN|30428-7|LNC2HPO|Microcytosis|Microcytosis
C0365392|T201|LN|3173-2|LNC2HPO|Haemorrhagic disorders|Haemorrhagic disorders
C0365392|T201|MTH_LN|3173-2|LNC2HPO|Haemorrhagic disorders|Haemorrhagic disorders
C0365392|T201|LC|3173-2|LNC2HPO|Haemorrhagic disorders|Haemorrhagic disorders
C0365392|T201|DN|3173-2|LNC2HPO|Haemorrhagic disorders|Haemorrhagic disorders
C0365392|T201|OSN|3173-2|LNC2HPO|Haemorrhagic disorders|Haemorrhagic disorders
C0365392|T201|LN|3173-2|LNC2HPO|Prolonged PTT|Prolonged PTT
C0365392|T201|MTH_LN|3173-2|LNC2HPO|Prolonged PTT|Prolonged PTT
C0365392|T201|LC|3173-2|LNC2HPO|Prolonged PTT|Prolonged PTT
C0365392|T201|DN|3173-2|LNC2HPO|Prolonged PTT|Prolonged PTT
C0365392|T201|OSN|3173-2|LNC2HPO|Prolonged PTT|Prolonged PTT
C0365392|T201|LN|3173-2|LNC2HPO|Prolonged partial thromboplastin time|Prolonged partial thromboplastin time
C0365392|T201|MTH_LN|3173-2|LNC2HPO|Prolonged partial thromboplastin time|Prolonged partial thromboplastin time
C0365392|T201|LC|3173-2|LNC2HPO|Prolonged partial thromboplastin time|Prolonged partial thromboplastin time
C0365392|T201|DN|3173-2|LNC2HPO|Prolonged partial thromboplastin time|Prolonged partial thromboplastin time
C0365392|T201|OSN|3173-2|LNC2HPO|Prolonged partial thromboplastin time|Prolonged partial thromboplastin time
C0365392|T201|LN|3173-2|LNC2HPO|Partial thromboplastin time prolonged|Partial thromboplastin time prolonged
C0365392|T201|MTH_LN|3173-2|LNC2HPO|Partial thromboplastin time prolonged|Partial thromboplastin time prolonged
C0365392|T201|LC|3173-2|LNC2HPO|Partial thromboplastin time prolonged|Partial thromboplastin time prolonged
C0365392|T201|DN|3173-2|LNC2HPO|Partial thromboplastin time prolonged|Partial thromboplastin time prolonged
C0365392|T201|OSN|3173-2|LNC2HPO|Partial thromboplastin time prolonged|Partial thromboplastin time prolonged
C0365392|T201|LN|3173-2|LNC2HPO|Delayed thromboplastin generation|Delayed thromboplastin generation
C0365392|T201|MTH_LN|3173-2|LNC2HPO|Delayed thromboplastin generation|Delayed thromboplastin generation
C0365392|T201|LC|3173-2|LNC2HPO|Delayed thromboplastin generation|Delayed thromboplastin generation
C0365392|T201|DN|3173-2|LNC2HPO|Delayed thromboplastin generation|Delayed thromboplastin generation
C0365392|T201|OSN|3173-2|LNC2HPO|Delayed thromboplastin generation|Delayed thromboplastin generation
C0365392|T201|LN|3173-2|LNC2HPO|Prolonged activated partial thromboplastin time|Prolonged activated partial thromboplastin time
C0365392|T201|MTH_LN|3173-2|LNC2HPO|Prolonged activated partial thromboplastin time|Prolonged activated partial thromboplastin time
C0365392|T201|LC|3173-2|LNC2HPO|Prolonged activated partial thromboplastin time|Prolonged activated partial thromboplastin time
C0365392|T201|DN|3173-2|LNC2HPO|Prolonged activated partial thromboplastin time|Prolonged activated partial thromboplastin time
C0365392|T201|OSN|3173-2|LNC2HPO|Prolonged activated partial thromboplastin time|Prolonged activated partial thromboplastin time
C0797906|T201|LN|14732-2|LNC2HPO|Folate deficiency|Folate deficiency
C0797906|T201|DN|14732-2|LNC2HPO|Folate deficiency|Folate deficiency
C0797906|T201|OSN|14732-2|LNC2HPO|Folate deficiency|Folate deficiency
C0797906|T201|MTH_LN|14732-2|LNC2HPO|Folate deficiency|Folate deficiency
C0797906|T201|LC|14732-2|LNC2HPO|Folate deficiency|Folate deficiency
C0797906|T201|LN|14732-2|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0797906|T201|DN|14732-2|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0797906|T201|OSN|14732-2|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0797906|T201|MTH_LN|14732-2|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0797906|T201|LC|14732-2|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0798076|T201|LN|14903-9|LNC2HPO|Folate deficiency|Folate deficiency
C0798076|T201|MTH_LN|14903-9|LNC2HPO|Folate deficiency|Folate deficiency
C0798076|T201|DN|14903-9|LNC2HPO|Folate deficiency|Folate deficiency
C0798076|T201|OSN|14903-9|LNC2HPO|Folate deficiency|Folate deficiency
C0798076|T201|LC|14903-9|LNC2HPO|Folate deficiency|Folate deficiency
C0798076|T201|LN|14903-9|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0798076|T201|MTH_LN|14903-9|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0798076|T201|DN|14903-9|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0798076|T201|OSN|14903-9|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0798076|T201|LC|14903-9|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0551446|T201|LN|11025-4|LNC2HPO|Meconium xenobiotic|Meconium xenobiotic
C0551446|T201|MTH_LN|11025-4|LNC2HPO|Meconium xenobiotic|Meconium xenobiotic
C0551446|T201|DN|11025-4|LNC2HPO|Meconium xenobiotic|Meconium xenobiotic
C0551446|T201|OSN|11025-4|LNC2HPO|Meconium xenobiotic|Meconium xenobiotic
C0551446|T201|LC|11025-4|LNC2HPO|Meconium xenobiotic|Meconium xenobiotic
C0944657|T201|LN|29159-1|LNC2HPO|Meconium xenobiotic|Meconium xenobiotic
C0944657|T201|DN|29159-1|LNC2HPO|Meconium xenobiotic|Meconium xenobiotic
C0944657|T201|MTH_LN|29159-1|LNC2HPO|Meconium xenobiotic|Meconium xenobiotic
C0944657|T201|OSN|29159-1|LNC2HPO|Meconium xenobiotic|Meconium xenobiotic
C0944657|T201|LC|29159-1|LNC2HPO|Meconium xenobiotic|Meconium xenobiotic
C1714972|T201|LN|43595-8|LNC2HPO|Meconium xenobiotic|Meconium xenobiotic
C1714972|T201|MTH_LN|43595-8|LNC2HPO|Meconium xenobiotic|Meconium xenobiotic
C1714972|T201|OSN|43595-8|LNC2HPO|Meconium xenobiotic|Meconium xenobiotic
C1714972|T201|DN|43595-8|LNC2HPO|Meconium xenobiotic|Meconium xenobiotic
C1714972|T201|LC|43595-8|LNC2HPO|Meconium xenobiotic|Meconium xenobiotic
C1978283|T201|LN|50410-0|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C1978283|T201|OSN|50410-0|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C1978283|T201|LC|50410-0|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C1978283|T201|DN|50410-0|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C1978283|T201|MTH_LN|50410-0|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C2736262|T201|LN|57838-5|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C2736262|T201|OSN|57838-5|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C2736262|T201|LC|57838-5|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C2736262|T201|DN|57838-5|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C2736262|T201|MTH_LN|57838-5|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C3262763|T201|LN|68916-6|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C3262763|T201|MTH_LN|68916-6|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C3262763|T201|OSN|68916-6|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C3262763|T201|LC|68916-6|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C3262763|T201|DN|68916-6|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C3870342|T201|LN|75511-6|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C3870342|T201|MTH_LN|75511-6|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C3870342|T201|LC|75511-6|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C3870342|T201|DN|75511-6|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C3870342|T201|OSN|75511-6|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C3870037|T201|LN|75883-9|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C3870037|T201|OSN|75883-9|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C3870037|T201|LC|75883-9|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C3870037|T201|MTH_LN|75883-9|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C3870037|T201|DN|75883-9|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C3870010|T201|LN|75913-4|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C3870010|T201|LC|75913-4|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C3870010|T201|MTH_LN|75913-4|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C3870010|T201|OSN|75913-4|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C3870010|T201|DN|75913-4|LNC2HPO|Lupus anticoagulant|Lupus anticoagulant
C0802017|T201|LN|19064-5|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802017|T201|MTH_LN|19064-5|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802017|T201|DN|19064-5|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802017|T201|OSN|19064-5|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802017|T201|LC|19064-5|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802179|T201|LN|19282-3|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802179|T201|LC|19282-3|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802179|T201|MTH_LN|19282-3|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802179|T201|DN|19282-3|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802179|T201|OSN|19282-3|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802180|T201|LN|19283-1|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802180|T201|MTH_LN|19283-1|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802180|T201|DN|19283-1|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802180|T201|OSN|19283-1|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802180|T201|LC|19283-1|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802181|T201|LN|19284-9|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802181|T201|LC|19284-9|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802181|T201|MTH_LN|19284-9|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802181|T201|DN|19284-9|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802181|T201|OSN|19284-9|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802182|T201|LN|19285-6|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802182|T201|MTH_LN|19285-6|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802182|T201|DN|19285-6|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802182|T201|OSN|19285-6|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802182|T201|LC|19285-6|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802183|T201|LN|19286-4|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802183|T201|LC|19286-4|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802183|T201|MTH_LN|19286-4|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802183|T201|DN|19286-4|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802183|T201|OSN|19286-4|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0365618|T201|MTH_LN|3387-8|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0365618|T201|DN|3387-8|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0365618|T201|OSN|3387-8|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0365618|T201|LN|3387-8|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0365618|T201|LC|3387-8|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C2361441|T201|LN|52955-2|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C2361441|T201|DN|52955-2|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C2361441|T201|OSN|52955-2|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C2361441|T201|MTH_LN|52955-2|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C2361441|T201|LC|52955-2|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C2598945|T201|LN|53736-5|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C2598945|T201|DN|53736-5|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C2598945|T201|MTH_LN|53736-5|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C2598945|T201|OSN|53736-5|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C2598945|T201|LC|53736-5|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C2598471|T201|LN|53745-6|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C2598471|T201|DN|53745-6|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C2598471|T201|LC|53745-6|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C2598471|T201|OSN|53745-6|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C2598471|T201|MTH_LN|53745-6|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C3481554|T201|LN|70140-9|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C3481554|T201|OSN|70140-9|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C3481554|T201|MTH_LN|70140-9|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C3481554|T201|LC|70140-9|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C3481554|T201|DN|70140-9|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C3482215|T201|LN|70142-5|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C3482215|T201|LC|70142-5|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C3482215|T201|OSN|70142-5|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C3482215|T201|MTH_LN|70142-5|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C3482215|T201|DN|70142-5|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0486032|T201|LN|9428-4|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0486032|T201|MTH_LN|9428-4|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0486032|T201|DN|9428-4|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0486032|T201|OSN|9428-4|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0486032|T201|LC|9428-4|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0797489|T201|LN|14308-1|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0797489|T201|MTH_LN|14308-1|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0797489|T201|DN|14308-1|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0797489|T201|OSN|14308-1|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0797489|T201|LC|14308-1|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0797490|T201|LN|14309-9|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0797490|T201|MTH_LN|14309-9|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0797490|T201|DN|14309-9|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0797490|T201|OSN|14309-9|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0797490|T201|LC|14309-9|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802163|T201|MTH_LN|19263-3|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802163|T201|DN|19263-3|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802163|T201|LN|19263-3|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802163|T201|OSN|19263-3|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0802163|T201|LC|19263-3|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0803225|T201|LN|20410-7|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0803225|T201|LC|20410-7|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0803225|T201|MTH_LN|20410-7|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0803225|T201|DN|20410-7|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0803225|T201|OSN|20410-7|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C3481552|T201|LN|70138-3|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C3481552|T201|OSN|70138-3|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C3481552|T201|MTH_LN|70138-3|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C3481552|T201|LC|70138-3|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C3481552|T201|DN|70138-3|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0486015|T201|LN|8150-5|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0486015|T201|MTH_LN|8150-5|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0486015|T201|DN|8150-5|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0486015|T201|OSN|8150-5|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0486015|T201|LC|8150-5|LNC2HPO|Urine xenobiotic|Urine xenobiotic
C0942465|T201|LN|26503-3|LNC2HPO|Neutrophilia|Neutrophilia
C0942465|T201|DN|26503-3|LNC2HPO|Neutrophilia|Neutrophilia
C0942465|T201|OSN|26503-3|LNC2HPO|Neutrophilia|Neutrophilia
C0942465|T201|MTH_LN|26503-3|LNC2HPO|Neutrophilia|Neutrophilia
C0942465|T201|LC|26503-3|LNC2HPO|Neutrophilia|Neutrophilia
C0942465|T201|LN|26503-3|LNC2HPO|Neutropenia|Neutropenia
C0942465|T201|DN|26503-3|LNC2HPO|Neutropenia|Neutropenia
C0942465|T201|OSN|26503-3|LNC2HPO|Neutropenia|Neutropenia
C0942465|T201|MTH_LN|26503-3|LNC2HPO|Neutropenia|Neutropenia
C0942465|T201|LC|26503-3|LNC2HPO|Neutropenia|Neutropenia
C0942465|T201|LN|26503-3|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0942465|T201|DN|26503-3|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0942465|T201|OSN|26503-3|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0942465|T201|MTH_LN|26503-3|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0942465|T201|LC|26503-3|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C3258971|T201|LN|66139-7|LNC2HPO|Neutrophilia|Neutrophilia
C3258971|T201|LC|66139-7|LNC2HPO|Neutrophilia|Neutrophilia
C3258971|T201|OSN|66139-7|LNC2HPO|Neutrophilia|Neutrophilia
C3258971|T201|MTH_LN|66139-7|LNC2HPO|Neutrophilia|Neutrophilia
C3258971|T201|DN|66139-7|LNC2HPO|Neutrophilia|Neutrophilia
C3258971|T201|LN|66139-7|LNC2HPO|Neutropenia|Neutropenia
C3258971|T201|LC|66139-7|LNC2HPO|Neutropenia|Neutropenia
C3258971|T201|OSN|66139-7|LNC2HPO|Neutropenia|Neutropenia
C3258971|T201|MTH_LN|66139-7|LNC2HPO|Neutropenia|Neutropenia
C3258971|T201|DN|66139-7|LNC2HPO|Neutropenia|Neutropenia
C3258971|T201|LN|66139-7|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C3258971|T201|LC|66139-7|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C3258971|T201|OSN|66139-7|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C3258971|T201|MTH_LN|66139-7|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C3258971|T201|DN|66139-7|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C3699844|T201|LN|74398-9|LNC2HPO|Neutrophilia|Neutrophilia
C3699844|T201|LC|74398-9|LNC2HPO|Neutrophilia|Neutrophilia
C3699844|T201|MTH_LN|74398-9|LNC2HPO|Neutrophilia|Neutrophilia
C3699844|T201|OSN|74398-9|LNC2HPO|Neutrophilia|Neutrophilia
C3699844|T201|DN|74398-9|LNC2HPO|Neutrophilia|Neutrophilia
C3699844|T201|LN|74398-9|LNC2HPO|Neutropenia|Neutropenia
C3699844|T201|LC|74398-9|LNC2HPO|Neutropenia|Neutropenia
C3699844|T201|MTH_LN|74398-9|LNC2HPO|Neutropenia|Neutropenia
C3699844|T201|OSN|74398-9|LNC2HPO|Neutropenia|Neutropenia
C3699844|T201|DN|74398-9|LNC2HPO|Neutropenia|Neutropenia
C3699844|T201|LN|74398-9|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C3699844|T201|LC|74398-9|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C3699844|T201|MTH_LN|74398-9|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C3699844|T201|OSN|74398-9|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C3699844|T201|DN|74398-9|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0362969|T201|LN|753-4|LNC2HPO|Neutrophilia|Neutrophilia
C0362969|T201|DN|753-4|LNC2HPO|Neutrophilia|Neutrophilia
C0362969|T201|OSN|753-4|LNC2HPO|Neutrophilia|Neutrophilia
C0362969|T201|MTH_LN|753-4|LNC2HPO|Neutrophilia|Neutrophilia
C0362969|T201|LC|753-4|LNC2HPO|Neutrophilia|Neutrophilia
C0362969|T201|LN|753-4|LNC2HPO|Neutropenia|Neutropenia
C0362969|T201|DN|753-4|LNC2HPO|Neutropenia|Neutropenia
C0362969|T201|OSN|753-4|LNC2HPO|Neutropenia|Neutropenia
C0362969|T201|MTH_LN|753-4|LNC2HPO|Neutropenia|Neutropenia
C0362969|T201|LC|753-4|LNC2HPO|Neutropenia|Neutropenia
C0362969|T201|LN|753-4|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0362969|T201|DN|753-4|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0362969|T201|OSN|753-4|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0362969|T201|MTH_LN|753-4|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C0362969|T201|LC|753-4|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C4482807|T201|LN|85369-7|LNC2HPO|Neutrophilia|Neutrophilia
C4482807|T201|MTH_LN|85369-7|LNC2HPO|Neutrophilia|Neutrophilia
C4482807|T201|OSN|85369-7|LNC2HPO|Neutrophilia|Neutrophilia
C4482807|T201|LC|85369-7|LNC2HPO|Neutrophilia|Neutrophilia
C4482807|T201|DN|85369-7|LNC2HPO|Neutrophilia|Neutrophilia
C4482807|T201|LN|85369-7|LNC2HPO|Neutropenia|Neutropenia
C4482807|T201|MTH_LN|85369-7|LNC2HPO|Neutropenia|Neutropenia
C4482807|T201|OSN|85369-7|LNC2HPO|Neutropenia|Neutropenia
C4482807|T201|LC|85369-7|LNC2HPO|Neutropenia|Neutropenia
C4482807|T201|DN|85369-7|LNC2HPO|Neutropenia|Neutropenia
C4482807|T201|LN|85369-7|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C4482807|T201|MTH_LN|85369-7|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C4482807|T201|OSN|85369-7|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C4482807|T201|LC|85369-7|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C4482807|T201|DN|85369-7|LNC2HPO|Peripheral neutropenia|Peripheral neutropenia
C1716121|T201|LN|44915-7|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1716121|T201|DN|44915-7|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1716121|T201|OSN|44915-7|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1716121|T201|LC|44915-7|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1716121|T201|MTH_LN|44915-7|LNC2HPO|Hyperbetalipoproteinemia|Hyperbetalipoproteinemia
C1716121|T201|LN|44915-7|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C1716121|T201|DN|44915-7|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C1716121|T201|OSN|44915-7|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C1716121|T201|LC|44915-7|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C1716121|T201|MTH_LN|44915-7|LNC2HPO|Hypobetalipoproteinemia|Hypobetalipoproteinemia
C0366794|T201|LN|4563-3|LNC2HPO|Hemoglobin C|Hemoglobin C
C0366794|T201|DN|4563-3|LNC2HPO|Hemoglobin C|Hemoglobin C
C0366794|T201|MTH_LN|4563-3|LNC2HPO|Hemoglobin C|Hemoglobin C
C0366794|T201|LC|4563-3|LNC2HPO|Hemoglobin C|Hemoglobin C
C0366794|T201|OSN|4563-3|LNC2HPO|Hemoglobin C|Hemoglobin C
C0366794|T201|LN|4563-3|LNC2HPO|HbC hemoglobin|HbC hemoglobin
C0366794|T201|DN|4563-3|LNC2HPO|HbC hemoglobin|HbC hemoglobin
C0366794|T201|MTH_LN|4563-3|LNC2HPO|HbC hemoglobin|HbC hemoglobin
C0366794|T201|LC|4563-3|LNC2HPO|HbC hemoglobin|HbC hemoglobin
C0366794|T201|OSN|4563-3|LNC2HPO|HbC hemoglobin|HbC hemoglobin
C0484423|T201|LN|10327-5|LNC2HPO|Sputum eosinophilia|Sputum eosinophilia
C0484423|T201|MTH_LN|10327-5|LNC2HPO|Sputum eosinophilia|Sputum eosinophilia
C0484423|T201|OSN|10327-5|LNC2HPO|Sputum eosinophilia|Sputum eosinophilia
C0484423|T201|DN|10327-5|LNC2HPO|Sputum eosinophilia|Sputum eosinophilia
C0484423|T201|LC|10327-5|LNC2HPO|Sputum eosinophilia|Sputum eosinophilia
C1113904|T201|LN|29993-3|LNC2HPO|Sputum eosinophilia|Sputum eosinophilia
C1113904|T201|MTH_LN|29993-3|LNC2HPO|Sputum eosinophilia|Sputum eosinophilia
C1113904|T201|DN|29993-3|LNC2HPO|Sputum eosinophilia|Sputum eosinophilia
C1113904|T201|OSN|29993-3|LNC2HPO|Sputum eosinophilia|Sputum eosinophilia
C1113904|T201|LC|29993-3|LNC2HPO|Sputum eosinophilia|Sputum eosinophilia
C1114243|T201|LN|30381-8|LNC2HPO|Sputum eosinophilia|Sputum eosinophilia
C1114243|T201|OSN|30381-8|LNC2HPO|Sputum eosinophilia|Sputum eosinophilia
C1114243|T201|DN|30381-8|LNC2HPO|Sputum eosinophilia|Sputum eosinophilia
C1114243|T201|MTH_LN|30381-8|LNC2HPO|Sputum eosinophilia|Sputum eosinophilia
C1114243|T201|LC|30381-8|LNC2HPO|Sputum eosinophilia|Sputum eosinophilia
C0365282|T201|LN|3137-7|LNC2HPO|Tall stature|Tall stature
C0365282|T201|MTH_LN|3137-7|LNC2HPO|Tall stature|Tall stature
C0365282|T201|LC|3137-7|LNC2HPO|Tall stature|Tall stature
C0365282|T201|OSN|3137-7|LNC2HPO|Tall stature|Tall stature
C0365282|T201|LN|3137-7|LNC2HPO|Accelerated linear growth|Accelerated linear growth
C0365282|T201|MTH_LN|3137-7|LNC2HPO|Accelerated linear growth|Accelerated linear growth
C0365282|T201|LC|3137-7|LNC2HPO|Accelerated linear growth|Accelerated linear growth
C0365282|T201|OSN|3137-7|LNC2HPO|Accelerated linear growth|Accelerated linear growth
C0365282|T201|LN|3137-7|LNC2HPO|Short stature|Short stature
C0365282|T201|MTH_LN|3137-7|LNC2HPO|Short stature|Short stature
C0365282|T201|LC|3137-7|LNC2HPO|Short stature|Short stature
C0365282|T201|OSN|3137-7|LNC2HPO|Short stature|Short stature
C0365282|T201|LN|3137-7|LNC2HPO|Small stature|Small stature
C0365282|T201|MTH_LN|3137-7|LNC2HPO|Small stature|Small stature
C0365282|T201|LC|3137-7|LNC2HPO|Small stature|Small stature
C0365282|T201|OSN|3137-7|LNC2HPO|Small stature|Small stature
C0365282|T201|LN|3137-7|LNC2HPO|Stature below 3rd percentile|Stature below 3rd percentile
C0365282|T201|MTH_LN|3137-7|LNC2HPO|Stature below 3rd percentile|Stature below 3rd percentile
C0365282|T201|LC|3137-7|LNC2HPO|Stature below 3rd percentile|Stature below 3rd percentile
C0365282|T201|OSN|3137-7|LNC2HPO|Stature below 3rd percentile|Stature below 3rd percentile
C0365282|T201|LN|3137-7|LNC2HPO|Height less than 3rd percentile|Height less than 3rd percentile
C0365282|T201|MTH_LN|3137-7|LNC2HPO|Height less than 3rd percentile|Height less than 3rd percentile
C0365282|T201|LC|3137-7|LNC2HPO|Height less than 3rd percentile|Height less than 3rd percentile
C0365282|T201|OSN|3137-7|LNC2HPO|Height less than 3rd percentile|Height less than 3rd percentile
C0365286|T201|LN|3141-9|LNC2HPO|Weight gain|Weight gain
C0365286|T201|LC|3141-9|LNC2HPO|Weight gain|Weight gain
C0365286|T201|OSN|3141-9|LNC2HPO|Weight gain|Weight gain
C0365286|T201|MTH_LN|3141-9|LNC2HPO|Weight gain|Weight gain
C0365286|T201|LN|3141-9|LNC2HPO|Weight less than 3rd percentile|Weight less than 3rd percentile
C0365286|T201|LC|3141-9|LNC2HPO|Weight less than 3rd percentile|Weight less than 3rd percentile
C0365286|T201|OSN|3141-9|LNC2HPO|Weight less than 3rd percentile|Weight less than 3rd percentile
C0365286|T201|MTH_LN|3141-9|LNC2HPO|Weight less than 3rd percentile|Weight less than 3rd percentile
C1369594|T201|LN|34728-6|LNC2HPO|Hypercapnia|Hypercapnia
C1369594|T201|DN|34728-6|LNC2HPO|Hypercapnia|Hypercapnia
C1369594|T201|OSN|34728-6|LNC2HPO|Hypercapnia|Hypercapnia
C1369594|T201|MTH_LN|34728-6|LNC2HPO|Hypercapnia|Hypercapnia
C1369594|T201|LC|34728-6|LNC2HPO|Hypercapnia|Hypercapnia
C1369594|T201|LN|34728-6|LNC2HPO|Hypercarbia|Hypercarbia
C1369594|T201|DN|34728-6|LNC2HPO|Hypercarbia|Hypercarbia
C1369594|T201|OSN|34728-6|LNC2HPO|Hypercarbia|Hypercarbia
C1369594|T201|MTH_LN|34728-6|LNC2HPO|Hypercarbia|Hypercarbia
C1369594|T201|LC|34728-6|LNC2HPO|Hypercarbia|Hypercarbia
C1369594|T201|LN|34728-6|LNC2HPO|Hypocapnia|Hypocapnia
C1369594|T201|DN|34728-6|LNC2HPO|Hypocapnia|Hypocapnia
C1369594|T201|OSN|34728-6|LNC2HPO|Hypocapnia|Hypocapnia
C1369594|T201|MTH_LN|34728-6|LNC2HPO|Hypocapnia|Hypocapnia
C1369594|T201|LC|34728-6|LNC2HPO|Hypocapnia|Hypocapnia
C1369594|T201|LN|34728-6|LNC2HPO|Hypocarbia|Hypocarbia
C1369594|T201|DN|34728-6|LNC2HPO|Hypocarbia|Hypocarbia
C1369594|T201|OSN|34728-6|LNC2HPO|Hypocarbia|Hypocarbia
C1369594|T201|MTH_LN|34728-6|LNC2HPO|Hypocarbia|Hypocarbia
C1369594|T201|LC|34728-6|LNC2HPO|Hypocarbia|Hypocarbia
C0484705|T201|LC|9813-7|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484705|T201|OSN|9813-7|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484705|T201|MTH_LN|9813-7|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484705|T201|LN|9813-7|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484705|T201|DN|9813-7|LNC2HPO|Cushing syndrome|Cushing syndrome
C0484705|T201|LC|9813-7|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484705|T201|OSN|9813-7|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484705|T201|MTH_LN|9813-7|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484705|T201|LN|9813-7|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484705|T201|DN|9813-7|LNC2HPO|Hypercortisolism|Hypercortisolism
C0484705|T201|LC|9813-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484705|T201|OSN|9813-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484705|T201|MTH_LN|9813-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484705|T201|LN|9813-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484705|T201|DN|9813-7|LNC2HPO|Hypocortisolism|Hypocortisolism
C0484705|T201|LC|9813-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484705|T201|OSN|9813-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484705|T201|MTH_LN|9813-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484705|T201|LN|9813-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484705|T201|DN|9813-7|LNC2HPO|Glucocorticoid insufficiency|Glucocorticoid insufficiency
C0484705|T201|LC|9813-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484705|T201|OSN|9813-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484705|T201|MTH_LN|9813-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484705|T201|LN|9813-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0484705|T201|DN|9813-7|LNC2HPO|Hypocortisolemia|Hypocortisolemia
C0363688|T201|LN|1557-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363688|T201|MTH_LN|1557-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363688|T201|DN|1557-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363688|T201|OSN|1557-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363688|T201|LC|1557-8|LNC2HPO|Hyperglycemia|Hyperglycemia
C0363688|T201|LN|1557-8|LNC2HPO|Fasting hypoglycemia|Fasting hypoglycemia
C0363688|T201|MTH_LN|1557-8|LNC2HPO|Fasting hypoglycemia|Fasting hypoglycemia
C0363688|T201|DN|1557-8|LNC2HPO|Fasting hypoglycemia|Fasting hypoglycemia
C0363688|T201|OSN|1557-8|LNC2HPO|Fasting hypoglycemia|Fasting hypoglycemia
C0363688|T201|LC|1557-8|LNC2HPO|Fasting hypoglycemia|Fasting hypoglycemia
C1953449|T201|LN|48065-7|LNC2HPO|Haemorrhagic disorders|Haemorrhagic disorders
C1953449|T201|DN|48065-7|LNC2HPO|Haemorrhagic disorders|Haemorrhagic disorders
C1953449|T201|OSN|48065-7|LNC2HPO|Haemorrhagic disorders|Haemorrhagic disorders
C1953449|T201|MTH_LN|48065-7|LNC2HPO|Haemorrhagic disorders|Haemorrhagic disorders
C1953449|T201|LC|48065-7|LNC2HPO|Haemorrhagic disorders|Haemorrhagic disorders
C0364418|T201|LN|2283-0|LNC2HPO|Folate deficiency|Folate deficiency
C0364418|T201|MTH_LN|2283-0|LNC2HPO|Folate deficiency|Folate deficiency
C0364418|T201|DN|2283-0|LNC2HPO|Folate deficiency|Folate deficiency
C0364418|T201|OSN|2283-0|LNC2HPO|Folate deficiency|Folate deficiency
C0364418|T201|LC|2283-0|LNC2HPO|Folate deficiency|Folate deficiency
C0364418|T201|LN|2283-0|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0364418|T201|MTH_LN|2283-0|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0364418|T201|DN|2283-0|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0364418|T201|OSN|2283-0|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0364418|T201|LC|2283-0|LNC2HPO|Vitamin B9 deficiency|Vitamin B9 deficiency
C0484652|T201|LN|1798-8|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0484652|T201|DN|1798-8|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0484652|T201|MTH_LN|1798-8|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0484652|T201|OSN|1798-8|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0484652|T201|LC|1798-8|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0484652|T201|LN|1798-8|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0484652|T201|DN|1798-8|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0484652|T201|MTH_LN|1798-8|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0484652|T201|OSN|1798-8|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0484652|T201|LC|1798-8|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0363939|T201|LN|1805-1|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0363939|T201|MTH_LN|1805-1|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0363939|T201|DN|1805-1|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0363939|T201|OSN|1805-1|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0363939|T201|LC|1805-1|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0363939|T201|LN|1805-1|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0363939|T201|MTH_LN|1805-1|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0363939|T201|DN|1805-1|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0363939|T201|OSN|1805-1|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0363939|T201|LC|1805-1|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0363940|T201|LN|1806-9|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0363940|T201|DN|1806-9|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0363940|T201|MTH_LN|1806-9|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0363940|T201|OSN|1806-9|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0363940|T201|LC|1806-9|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0363940|T201|LN|1806-9|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0363940|T201|DN|1806-9|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0363940|T201|MTH_LN|1806-9|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0363940|T201|OSN|1806-9|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0363940|T201|LC|1806-9|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0363941|T201|LN|1807-7|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0363941|T201|DN|1807-7|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0363941|T201|MTH_LN|1807-7|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0363941|T201|OSN|1807-7|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0363941|T201|LC|1807-7|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0363941|T201|LN|1807-7|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0363941|T201|DN|1807-7|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0363941|T201|MTH_LN|1807-7|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0363941|T201|OSN|1807-7|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0363941|T201|LC|1807-7|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0363942|T201|LN|1808-5|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0363942|T201|DN|1808-5|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0363942|T201|MTH_LN|1808-5|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0363942|T201|OSN|1808-5|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0363942|T201|LC|1808-5|LNC2HPO|Hyperamylasemia|Hyperamylasemia
C0363942|T201|LN|1808-5|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0363942|T201|DN|1808-5|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0363942|T201|MTH_LN|1808-5|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0363942|T201|OSN|1808-5|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0363942|T201|LC|1808-5|LNC2HPO|Hypoamylasemia|Hypoamylasemia
C0803262|T201|LN|20448-7|LNC2HPO|Hyperinsulinemia|Hyperinsulinemia
C0803262|T201|DN|20448-7|LNC2HPO|Hyperinsulinemia|Hyperinsulinemia
C0803262|T201|MTH_LN|20448-7|LNC2HPO|Hyperinsulinemia|Hyperinsulinemia
C0803262|T201|OSN|20448-7|LNC2HPO|Hyperinsulinemia|Hyperinsulinemia
C0803262|T201|LC|20448-7|LNC2HPO|Hyperinsulinemia|Hyperinsulinemia
C0803262|T201|LN|20448-7|LNC2HPO|Hypoinsulinemia|Hypoinsulinemia
C0803262|T201|DN|20448-7|LNC2HPO|Hypoinsulinemia|Hypoinsulinemia
C0803262|T201|MTH_LN|20448-7|LNC2HPO|Hypoinsulinemia|Hypoinsulinemia
C0803262|T201|OSN|20448-7|LNC2HPO|Hypoinsulinemia|Hypoinsulinemia
C0803262|T201|LC|20448-7|LNC2HPO|Hypoinsulinemia|Hypoinsulinemia
C0942441|T201|LN|26479-6|LNC2HPO|CSF lymphocytosis|CSF lymphocytosis
C0942441|T201|OSN|26479-6|LNC2HPO|CSF lymphocytosis|CSF lymphocytosis
C0942441|T201|DN|26479-6|LNC2HPO|CSF lymphocytosis|CSF lymphocytosis
C0942441|T201|MTH_LN|26479-6|LNC2HPO|CSF lymphocytosis|CSF lymphocytosis
C0942441|T201|LC|26479-6|LNC2HPO|CSF lymphocytosis|CSF lymphocytosis
C0942441|T201|LN|26479-6|LNC2HPO|CSF lymphocytic pleiocytosis|CSF lymphocytic pleiocytosis
C0942441|T201|OSN|26479-6|LNC2HPO|CSF lymphocytic pleiocytosis|CSF lymphocytic pleiocytosis
C0942441|T201|DN|26479-6|LNC2HPO|CSF lymphocytic pleiocytosis|CSF lymphocytic pleiocytosis
C0942441|T201|MTH_LN|26479-6|LNC2HPO|CSF lymphocytic pleiocytosis|CSF lymphocytic pleiocytosis
C0942441|T201|LC|26479-6|LNC2HPO|CSF lymphocytic pleiocytosis|CSF lymphocytic pleiocytosis
C0365160|T201|LN|3016-3|LNC2HPO|TSH excess|TSH excess
C0365160|T201|MTH_LN|3016-3|LNC2HPO|TSH excess|TSH excess
C0365160|T201|DN|3016-3|LNC2HPO|TSH excess|TSH excess
C0365160|T201|OSN|3016-3|LNC2HPO|TSH excess|TSH excess
C0365160|T201|LC|3016-3|LNC2HPO|TSH excess|TSH excess
C0489258|T201|MTH_LN|9279-1|LNC2HPO|Unusual breathing patterns|Unusual breathing patterns
C0489258|T201|LC|9279-1|LNC2HPO|Unusual breathing patterns|Unusual breathing patterns
C0489258|T201|LN|9279-1|LNC2HPO|Unusual breathing patterns|Unusual breathing patterns
C0489258|T201|OSN|9279-1|LNC2HPO|Unusual breathing patterns|Unusual breathing patterns
C0489258|T201|MTH_LN|9279-1|LNC2HPO|Tachypnea|Tachypnea
C0489258|T201|LC|9279-1|LNC2HPO|Tachypnea|Tachypnea
C0489258|T201|LN|9279-1|LNC2HPO|Tachypnea|Tachypnea
C0489258|T201|OSN|9279-1|LNC2HPO|Tachypnea|Tachypnea
C0489258|T201|MTH_LN|9279-1|LNC2HPO|Polypnea|Polypnea
C0489258|T201|LC|9279-1|LNC2HPO|Polypnea|Polypnea
C0489258|T201|LN|9279-1|LNC2HPO|Polypnea|Polypnea
C0489258|T201|OSN|9279-1|LNC2HPO|Polypnea|Polypnea
C0489258|T201|MTH_LN|9279-1|LNC2HPO|Hypopnea|Hypopnea
C0489258|T201|LC|9279-1|LNC2HPO|Hypopnea|Hypopnea
C0489258|T201|LN|9279-1|LNC2HPO|Hypopnea|Hypopnea
C0489258|T201|OSN|9279-1|LNC2HPO|Hypopnea|Hypopnea
C0550439|T201|LN|13483-3|LNC2HPO|Hyperoxaluria|Hyperoxaluria
C0550439|T201|OSN|13483-3|LNC2HPO|Hyperoxaluria|Hyperoxaluria
C0550439|T201|MTH_LN|13483-3|LNC2HPO|Hyperoxaluria|Hyperoxaluria
C0550439|T201|DN|13483-3|LNC2HPO|Hyperoxaluria|Hyperoxaluria
C0550439|T201|LC|13483-3|LNC2HPO|Hyperoxaluria|Hyperoxaluria
C0796977|T201|LN|13787-7|LNC2HPO|Orotic aciduria|Orotic aciduria
C0796977|T201|OSN|13787-7|LNC2HPO|Orotic aciduria|Orotic aciduria
C0796977|T201|MTH_LN|13787-7|LNC2HPO|Orotic aciduria|Orotic aciduria
C0796977|T201|DN|13787-7|LNC2HPO|Orotic aciduria|Orotic aciduria
C0796977|T201|LC|13787-7|LNC2HPO|Orotic aciduria|Orotic aciduria
C0796977|T201|LN|13787-7|LNC2HPO|Oroticaciduria|Oroticaciduria
C0796977|T201|OSN|13787-7|LNC2HPO|Oroticaciduria|Oroticaciduria
C0796977|T201|MTH_LN|13787-7|LNC2HPO|Oroticaciduria|Oroticaciduria
C0796977|T201|DN|13787-7|LNC2HPO|Oroticaciduria|Oroticaciduria
C0796977|T201|LC|13787-7|LNC2HPO|Oroticaciduria|Oroticaciduria
C0797152|T201|LN|13964-2|LNC2HPO|Methylmalonic acidemia|Methylmalonic acidemia
C0797152|T201|DN|13964-2|LNC2HPO|Methylmalonic acidemia|Methylmalonic acidemia
C0797152|T201|MTH_LN|13964-2|LNC2HPO|Methylmalonic acidemia|Methylmalonic acidemia
C0797152|T201|OSN|13964-2|LNC2HPO|Methylmalonic acidemia|Methylmalonic acidemia
C0797152|T201|LC|13964-2|LNC2HPO|Methylmalonic acidemia|Methylmalonic acidemia
C0797154|T201|LN|13966-7|LNC2HPO|Cystinuria|Cystinuria
C0797154|T201|MTH_LN|13966-7|LNC2HPO|Cystinuria|Cystinuria
C0797154|T201|DN|13966-7|LNC2HPO|Cystinuria|Cystinuria
C0797154|T201|OSN|13966-7|LNC2HPO|Cystinuria|Cystinuria
C0797154|T201|LC|13966-7|LNC2HPO|Cystinuria|Cystinuria
C0797321|T201|LN|14135-8|LNC2HPO|CD8+ T-cell lymphopenia|CD8+ T-cell lymphopenia
C0797321|T201|LC|14135-8|LNC2HPO|CD8+ T-cell lymphopenia|CD8+ T-cell lymphopenia
C0797321|T201|DN|14135-8|LNC2HPO|CD8+ T-cell lymphopenia|CD8+ T-cell lymphopenia
C0797321|T201|OSN|14135-8|LNC2HPO|CD8+ T-cell lymphopenia|CD8+ T-cell lymphopenia
C0797321|T201|MTH_LN|14135-8|LNC2HPO|CD8+ T-cell lymphopenia|CD8+ T-cell lymphopenia
C0798036|T201|LN|14862-7|LNC2HPO|Hyperoxaluria|Hyperoxaluria
C0798036|T201|MTH_LN|14862-7|LNC2HPO|Hyperoxaluria|Hyperoxaluria
C0798036|T201|DN|14862-7|LNC2HPO|Hyperoxaluria|Hyperoxaluria
C0798036|T201|OSN|14862-7|LNC2HPO|Hyperoxaluria|Hyperoxaluria
C0798036|T201|LC|14862-7|LNC2HPO|Hyperoxaluria|Hyperoxaluria
C0798152|T201|LN|14979-9|LNC2HPO|Haemorrhagic disorders|Haemorrhagic disorders
C0798152|T201|LC|14979-9|LNC2HPO|Haemorrhagic disorders|Haemorrhagic disorders
C0798152|T201|DN|14979-9|LNC2HPO|Haemorrhagic disorders|Haemorrhagic disorders
C0798152|T201|MTH_LN|14979-9|LNC2HPO|Haemorrhagic disorders|Haemorrhagic disorders
C0798152|T201|OSN|14979-9|LNC2HPO|Haemorrhagic disorders|Haemorrhagic disorders
C0798152|T201|LN|14979-9|LNC2HPO|Prolonged PTT|Prolonged PTT
C0798152|T201|LC|14979-9|LNC2HPO|Prolonged PTT|Prolonged PTT
C0798152|T201|DN|14979-9|LNC2HPO|Prolonged PTT|Prolonged PTT
C0798152|T201|MTH_LN|14979-9|LNC2HPO|Prolonged PTT|Prolonged PTT
C0798152|T201|OSN|14979-9|LNC2HPO|Prolonged PTT|Prolonged PTT
C0798152|T201|LN|14979-9|LNC2HPO|Prolonged partial thromboplastin time|Prolonged partial thromboplastin time
C0798152|T201|LC|14979-9|LNC2HPO|Prolonged partial thromboplastin time|Prolonged partial thromboplastin time
C0798152|T201|DN|14979-9|LNC2HPO|Prolonged partial thromboplastin time|Prolonged partial thromboplastin time
C0798152|T201|MTH_LN|14979-9|LNC2HPO|Prolonged partial thromboplastin time|Prolonged partial thromboplastin time
C0798152|T201|OSN|14979-9|LNC2HPO|Prolonged partial thromboplastin time|Prolonged partial thromboplastin time
C0798152|T201|LN|14979-9|LNC2HPO|Partial thromboplastin time prolonged|Partial thromboplastin time prolonged
C0798152|T201|LC|14979-9|LNC2HPO|Partial thromboplastin time prolonged|Partial thromboplastin time prolonged
C0798152|T201|DN|14979-9|LNC2HPO|Partial thromboplastin time prolonged|Partial thromboplastin time prolonged
C0798152|T201|MTH_LN|14979-9|LNC2HPO|Partial thromboplastin time prolonged|Partial thromboplastin time prolonged
C0798152|T201|OSN|14979-9|LNC2HPO|Partial thromboplastin time prolonged|Partial thromboplastin time prolonged
C0798152|T201|LN|14979-9|LNC2HPO|Delayed thromboplastin generation|Delayed thromboplastin generation
C0798152|T201|LC|14979-9|LNC2HPO|Delayed thromboplastin generation|Delayed thromboplastin generation
C0798152|T201|DN|14979-9|LNC2HPO|Delayed thromboplastin generation|Delayed thromboplastin generation
C0798152|T201|MTH_LN|14979-9|LNC2HPO|Delayed thromboplastin generation|Delayed thromboplastin generation
C0798152|T201|OSN|14979-9|LNC2HPO|Delayed thromboplastin generation|Delayed thromboplastin generation
C0798152|T201|LN|14979-9|LNC2HPO|Prolonged activated partial thromboplastin time|Prolonged activated partial thromboplastin time
C0798152|T201|LC|14979-9|LNC2HPO|Prolonged activated partial thromboplastin time|Prolonged activated partial thromboplastin time
C0798152|T201|DN|14979-9|LNC2HPO|Prolonged activated partial thromboplastin time|Prolonged activated partial thromboplastin time
C0798152|T201|MTH_LN|14979-9|LNC2HPO|Prolonged activated partial thromboplastin time|Prolonged activated partial thromboplastin time
C0798152|T201|OSN|14979-9|LNC2HPO|Prolonged activated partial thromboplastin time|Prolonged activated partial thromboplastin time
C0798254|T201|LN|15082-1|LNC2HPO|Methemoglobinemia|Methemoglobinemia
C0798254|T201|MTH_LN|15082-1|LNC2HPO|Methemoglobinemia|Methemoglobinemia
C0798254|T201|DN|15082-1|LNC2HPO|Methemoglobinemia|Methemoglobinemia
C0798254|T201|OSN|15082-1|LNC2HPO|Methemoglobinemia|Methemoglobinemia
C0798254|T201|LC|15082-1|LNC2HPO|Methemoglobinemia|Methemoglobinemia
C0799307|T201|LN|16142-2|LNC2HPO|Steatorrhea|Steatorrhea
C0799307|T201|MTH_LN|16142-2|LNC2HPO|Steatorrhea|Steatorrhea
C0799307|T201|DN|16142-2|LNC2HPO|Steatorrhea|Steatorrhea
C0799307|T201|OSN|16142-2|LNC2HPO|Steatorrhea|Steatorrhea
C0799307|T201|LC|16142-2|LNC2HPO|Steatorrhea|Steatorrhea
C0799307|T201|LN|16142-2|LNC2HPO|Fat in feces|Fat in feces
C0799307|T201|MTH_LN|16142-2|LNC2HPO|Fat in feces|Fat in feces
C0799307|T201|DN|16142-2|LNC2HPO|Fat in feces|Fat in feces
C0799307|T201|OSN|16142-2|LNC2HPO|Fat in feces|Fat in feces
C0799307|T201|LC|16142-2|LNC2HPO|Fat in feces|Fat in feces
C0799700|T201|LN|16551-4|LNC2HPO|Hypercapnia|Hypercapnia
C0799700|T201|MTH_LN|16551-4|LNC2HPO|Hypercapnia|Hypercapnia
C0799700|T201|DN|16551-4|LNC2HPO|Hypercapnia|Hypercapnia
C0799700|T201|OSN|16551-4|LNC2HPO|Hypercapnia|Hypercapnia
C0799700|T201|LC|16551-4|LNC2HPO|Hypercapnia|Hypercapnia
C0799700|T201|LN|16551-4|LNC2HPO|Hypercarbia|Hypercarbia
C0799700|T201|MTH_LN|16551-4|LNC2HPO|Hypercarbia|Hypercarbia
C0799700|T201|DN|16551-4|LNC2HPO|Hypercarbia|Hypercarbia
C0799700|T201|OSN|16551-4|LNC2HPO|Hypercarbia|Hypercarbia
C0799700|T201|LC|16551-4|LNC2HPO|Hypercarbia|Hypercarbia
C0799700|T201|LN|16551-4|LNC2HPO|Hypocapnia|Hypocapnia
C0799700|T201|MTH_LN|16551-4|LNC2HPO|Hypocapnia|Hypocapnia
C0799700|T201|DN|16551-4|LNC2HPO|Hypocapnia|Hypocapnia
C0799700|T201|OSN|16551-4|LNC2HPO|Hypocapnia|Hypocapnia
C0799700|T201|LC|16551-4|LNC2HPO|Hypocapnia|Hypocapnia
C0799700|T201|LN|16551-4|LNC2HPO|Hypocarbia|Hypocarbia
C0799700|T201|MTH_LN|16551-4|LNC2HPO|Hypocarbia|Hypocarbia
C0799700|T201|DN|16551-4|LNC2HPO|Hypocarbia|Hypocarbia
C0799700|T201|OSN|16551-4|LNC2HPO|Hypocarbia|Hypocarbia
C0799700|T201|LC|16551-4|LNC2HPO|Hypocarbia|Hypocarbia
C0363822|T201|LN|1688-1|LNC2HPO|Vitamin B6 deficiency|Vitamin B6 deficiency
C0363822|T201|DN|1688-1|LNC2HPO|Vitamin B6 deficiency|Vitamin B6 deficiency
C0363822|T201|MTH_LN|1688-1|LNC2HPO|Vitamin B6 deficiency|Vitamin B6 deficiency
C0363822|T201|OSN|1688-1|LNC2HPO|Vitamin B6 deficiency|Vitamin B6 deficiency
C0363822|T201|LC|1688-1|LNC2HPO|Vitamin B6 deficiency|Vitamin B6 deficiency
C0363897|T201|LC|1763-2|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C0363897|T201|DN|1763-2|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C0363897|T201|MTH_LN|1763-2|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C0363897|T201|LN|1763-2|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C0363897|T201|OSN|1763-2|LNC2HPO|Hypoaldosteronism|Hypoaldosteronism
C0363897|T201|LC|1763-2|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C0363897|T201|DN|1763-2|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C0363897|T201|MTH_LN|1763-2|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C0363897|T201|LN|1763-2|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C0363897|T201|OSN|1763-2|LNC2HPO|Mineralocorticoid insufficiency|Mineralocorticoid insufficiency
C0363897|T201|LC|1763-2|LNC2HPO|Hyperaldosteronism|Hyperaldosteronism
C0363897|T201|DN|1763-2|LNC2HPO|Hyperaldosteronism|Hyperaldosteronism
C0363897|T201|MTH_LN|1763-2|LNC2HPO|Hyperaldosteronism|Hyperaldosteronism
C0363897|T201|LN|1763-2|LNC2HPO|Hyperaldosteronism|Hyperaldosteronism
C0363897|T201|OSN|1763-2|LNC2HPO|Hyperaldosteronism|Hyperaldosteronism
C0363897|T201|LC|1763-2|LNC2HPO|Mineralocorticoid excess|Mineralocorticoid excess
C0363897|T201|DN|1763-2|LNC2HPO|Mineralocorticoid excess|Mineralocorticoid excess
C0363897|T201|MTH_LN|1763-2|LNC2HPO|Mineralocorticoid excess|Mineralocorticoid excess
C0363897|T201|LN|1763-2|LNC2HPO|Mineralocorticoid excess|Mineralocorticoid excess
C0363897|T201|OSN|1763-2|LNC2HPO|Mineralocorticoid excess|Mineralocorticoid excess
C0800964|T201|MTH_LN|17857-4|LNC2HPO|Rheumatoid factor positive|Rheumatoid factor positive
C0800964|T201|DN|17857-4|LNC2HPO|Rheumatoid factor positive|Rheumatoid factor positive
C0800964|T201|LN|17857-4|LNC2HPO|Rheumatoid factor positive|Rheumatoid factor positive
C0800964|T201|OSN|17857-4|LNC2HPO|Rheumatoid factor positive|Rheumatoid factor positive
C0800964|T201|LC|17857-4|LNC2HPO|Rheumatoid factor positive|Rheumatoid factor positive
C0802012|T201|LN|19023-1|LNC2HPO|Granulocytosis|Granulocytosis
C0802012|T201|OSN|19023-1|LNC2HPO|Granulocytosis|Granulocytosis
C0802012|T201|MTH_LN|19023-1|LNC2HPO|Granulocytosis|Granulocytosis
C0802012|T201|DN|19023-1|LNC2HPO|Granulocytosis|Granulocytosis
C0802012|T201|LC|19023-1|LNC2HPO|Granulocytosis|Granulocytosis
C0802012|T201|LN|19023-1|LNC2HPO|Granulocytopenia|Granulocytopenia
C0802012|T201|OSN|19023-1|LNC2HPO|Granulocytopenia|Granulocytopenia
C0802012|T201|MTH_LN|19023-1|LNC2HPO|Granulocytopenia|Granulocytopenia
C0802012|T201|DN|19023-1|LNC2HPO|Granulocytopenia|Granulocytopenia
C0802012|T201|LC|19023-1|LNC2HPO|Granulocytopenia|Granulocytopenia
C0484665|T201|MTH_LN|1903-4|LNC2HPO|Vitamin C deficiency|Vitamin C deficiency
C0484665|T201|LN|1903-4|LNC2HPO|Vitamin C deficiency|Vitamin C deficiency
C0484665|T201|DN|1903-4|LNC2HPO|Vitamin C deficiency|Vitamin C deficiency
C0484665|T201|OSN|1903-4|LNC2HPO|Vitamin C deficiency|Vitamin C deficiency
C0484665|T201|LC|1903-4|LNC2HPO|Vitamin C deficiency|Vitamin C deficiency
C1153749|T201|LN|19214-6|LNC2HPO|Hyperoxemia|Hyperoxemia
C1153749|T201|MTH_LN|19214-6|LNC2HPO|Hyperoxemia|Hyperoxemia
C1153749|T201|DN|19214-6|LNC2HPO|Hyperoxemia|Hyperoxemia
C1153749|T201|OSN|19214-6|LNC2HPO|Hyperoxemia|Hyperoxemia
C1153749|T201|LC|19214-6|LNC2HPO|Hyperoxemia|Hyperoxemia
C1153749|T201|LN|19214-6|LNC2HPO|Hypoxemia|Hypoxemia
C1153749|T201|MTH_LN|19214-6|LNC2HPO|Hypoxemia|Hypoxemia
C1153749|T201|DN|19214-6|LNC2HPO|Hypoxemia|Hypoxemia
C1153749|T201|OSN|19214-6|LNC2HPO|Hypoxemia|Hypoxemia
C1153749|T201|LC|19214-6|LNC2HPO|Hypoxemia|Hypoxemia
C0364846|T201|LN|19255-9|LNC2HPO|Hyperoxemia|Hyperoxemia
C0364846|T201|MTH_LN|19255-9|LNC2HPO|Hyperoxemia|Hyperoxemia
C0364846|T201|DN|19255-9|LNC2HPO|Hyperoxemia|Hyperoxemia
C0364846|T201|OSN|19255-9|LNC2HPO|Hyperoxemia|Hyperoxemia
C0364846|T201|LC|19255-9|LNC2HPO|Hyperoxemia|Hyperoxemia
C0364846|T201|LN|19255-9|LNC2HPO|Hypoxemia|Hypoxemia
C0364846|T201|MTH_LN|19255-9|LNC2HPO|Hypoxemia|Hypoxemia
C0364846|T201|DN|19255-9|LNC2HPO|Hypoxemia|Hypoxemia
C0364846|T201|OSN|19255-9|LNC2HPO|Hypoxemia|Hypoxemia
C0364846|T201|LC|19255-9|LNC2HPO|Hypoxemia|Hypoxemia
C0364086|T201|LN|1953-9|LNC2HPO|Beta 2-microglobulinuria|Beta 2-microglobulinuria
C0364086|T201|MTH_LN|1953-9|LNC2HPO|Beta 2-microglobulinuria|Beta 2-microglobulinuria
C0364086|T201|DN|1953-9|LNC2HPO|Beta 2-microglobulinuria|Beta 2-microglobulinuria
C0364086|T201|OSN|1953-9|LNC2HPO|Beta 2-microglobulinuria|Beta 2-microglobulinuria
C0364086|T201|LC|1953-9|LNC2HPO|Beta 2-microglobulinuria|Beta 2-microglobulinuria
C0364152|T201|LN|2020-6|LNC2HPO|Hypercapnia|Hypercapnia
C0364152|T201|MTH_LN|2020-6|LNC2HPO|Hypercapnia|Hypercapnia
C0364152|T201|DN|2020-6|LNC2HPO|Hypercapnia|Hypercapnia
C0364152|T201|LC|2020-6|LNC2HPO|Hypercapnia|Hypercapnia
C0364152|T201|OSN|2020-6|LNC2HPO|Hypercapnia|Hypercapnia
C0364152|T201|LN|2020-6|LNC2HPO|Hypercarbia|Hypercarbia
C0364152|T201|MTH_LN|2020-6|LNC2HPO|Hypercarbia|Hypercarbia
C0364152|T201|DN|2020-6|LNC2HPO|Hypercarbia|Hypercarbia
C0364152|T201|LC|2020-6|LNC2HPO|Hypercarbia|Hypercarbia
C0364152|T201|OSN|2020-6|LNC2HPO|Hypercarbia|Hypercarbia
C0364152|T201|LN|2020-6|LNC2HPO|Hypocapnia|Hypocapnia
C0364152|T201|MTH_LN|2020-6|LNC2HPO|Hypocapnia|Hypocapnia
C0364152|T201|DN|2020-6|LNC2HPO|Hypocapnia|Hypocapnia
C0364152|T201|LC|2020-6|LNC2HPO|Hypocapnia|Hypocapnia
C0364152|T201|OSN|2020-6|LNC2HPO|Hypocapnia|Hypocapnia
C0364152|T201|LN|2020-6|LNC2HPO|Hypocarbia|Hypocarbia
C0364152|T201|MTH_LN|2020-6|LNC2HPO|Hypocarbia|Hypocarbia
C0364152|T201|DN|2020-6|LNC2HPO|Hypocarbia|Hypocarbia
C0364152|T201|LC|2020-6|LNC2HPO|Hypocarbia|Hypocarbia
C0364152|T201|OSN|2020-6|LNC2HPO|Hypocarbia|Hypocarbia
C0364159|T201|LN|2027-1|LNC2HPO|Hypercapnia|Hypercapnia
C0364159|T201|MTH_LN|2027-1|LNC2HPO|Hypercapnia|Hypercapnia
C0364159|T201|DN|2027-1|LNC2HPO|Hypercapnia|Hypercapnia
C0364159|T201|OSN|2027-1|LNC2HPO|Hypercapnia|Hypercapnia
C0364159|T201|LC|2027-1|LNC2HPO|Hypercapnia|Hypercapnia
C0364159|T201|LN|2027-1|LNC2HPO|Hypercarbia|Hypercarbia
C0364159|T201|MTH_LN|2027-1|LNC2HPO|Hypercarbia|Hypercarbia
C0364159|T201|DN|2027-1|LNC2HPO|Hypercarbia|Hypercarbia
C0364159|T201|OSN|2027-1|LNC2HPO|Hypercarbia|Hypercarbia
C0364159|T201|LC|2027-1|LNC2HPO|Hypercarbia|Hypercarbia
C0364159|T201|LN|2027-1|LNC2HPO|Hypocapnia|Hypocapnia
C0364159|T201|MTH_LN|2027-1|LNC2HPO|Hypocapnia|Hypocapnia
C0364159|T201|DN|2027-1|LNC2HPO|Hypocapnia|Hypocapnia
C0364159|T201|OSN|2027-1|LNC2HPO|Hypocapnia|Hypocapnia
C0364159|T201|LC|2027-1|LNC2HPO|Hypocapnia|Hypocapnia
C0364159|T201|LN|2027-1|LNC2HPO|Hypocarbia|Hypocarbia
C0364159|T201|MTH_LN|2027-1|LNC2HPO|Hypocarbia|Hypocarbia
C0364159|T201|DN|2027-1|LNC2HPO|Hypocarbia|Hypocarbia
C0364159|T201|OSN|2027-1|LNC2HPO|Hypocarbia|Hypocarbia
C0364159|T201|LC|2027-1|LNC2HPO|Hypocarbia|Hypocarbia
C0803294|T201|LN|20482-6|LNC2HPO|Granulocytosis|Granulocytosis
C0803294|T201|DN|20482-6|LNC2HPO|Granulocytosis|Granulocytosis
C0803294|T201|OSN|20482-6|LNC2HPO|Granulocytosis|Granulocytosis
C0803294|T201|MTH_LN|20482-6|LNC2HPO|Granulocytosis|Granulocytosis
C0803294|T201|LC|20482-6|LNC2HPO|Granulocytosis|Granulocytosis
C0803294|T201|LN|20482-6|LNC2HPO|Granulocytopenia|Granulocytopenia
C0803294|T201|DN|20482-6|LNC2HPO|Granulocytopenia|Granulocytopenia
C0803294|T201|OSN|20482-6|LNC2HPO|Granulocytopenia|Granulocytopenia
C0803294|T201|MTH_LN|20482-6|LNC2HPO|Granulocytopenia|Granulocytopenia
C0803294|T201|LC|20482-6|LNC2HPO|Granulocytopenia|Granulocytopenia
C0880191|T201|MTH_LN|20646-6|LNC2HPO|Hyperhomocystinemia|Hyperhomocystinemia
C0880191|T201|OSN|20646-6|LNC2HPO|Hyperhomocystinemia|Hyperhomocystinemia
C0880191|T201|DN|20646-6|LNC2HPO|Hyperhomocystinemia|Hyperhomocystinemia
C0880191|T201|LN|20646-6|LNC2HPO|Hyperhomocystinemia|Hyperhomocystinemia
C0880191|T201|LC|20646-6|LNC2HPO|Hyperhomocystinemia|Hyperhomocystinemia
C0880191|T201|MTH_LN|20646-6|LNC2HPO|Homocystinemia|Homocystinemia
C0880191|T201|OSN|20646-6|LNC2HPO|Homocystinemia|Homocystinemia
C0880191|T201|DN|20646-6|LNC2HPO|Homocystinemia|Homocystinemia
C0880191|T201|LN|20646-6|LNC2HPO|Homocystinemia|Homocystinemia
C0880191|T201|LC|20646-6|LNC2HPO|Homocystinemia|Homocystinemia
C0364201|T201|LN|2069-3|LNC2HPO|Hyperchloremia|Hyperchloremia
C0364201|T201|MTH_LN|2069-3|LNC2HPO|Hyperchloremia|Hyperchloremia
C0364201|T201|DN|2069-3|LNC2HPO|Hyperchloremia|Hyperchloremia
C0364201|T201|OSN|2069-3|LNC2HPO|Hyperchloremia|Hyperchloremia
C0364201|T201|LC|2069-3|LNC2HPO|Hyperchloremia|Hyperchloremia
C0364201|T201|LN|2069-3|LNC2HPO|Hypochloremia|Hypochloremia
C0364201|T201|MTH_LN|2069-3|LNC2HPO|Hypochloremia|Hypochloremia
C0364201|T201|DN|2069-3|LNC2HPO|Hypochloremia|Hypochloremia
C0364201|T201|OSN|2069-3|LNC2HPO|Hypochloremia|Hypochloremia
C0364201|T201|LC|2069-3|LNC2HPO|Hypochloremia|Hypochloremia
C0364214|T201|LN|2082-6|LNC2HPO|Hypercholesterolemia|Hypercholesterolemia
C0364214|T201|DN|2082-6|LNC2HPO|Hypercholesterolemia|Hypercholesterolemia
C0364214|T201|MTH_LN|2082-6|LNC2HPO|Hypercholesterolemia|Hypercholesterolemia
C0364214|T201|OSN|2082-6|LNC2HPO|Hypercholesterolemia|Hypercholesterolemia
C0364214|T201|LC|2082-6|LNC2HPO|Hypercholesterolemia|Hypercholesterolemia
C0364214|T201|LN|2082-6|LNC2HPO|Hypocholesterolemia|Hypocholesterolemia
C0364214|T201|DN|2082-6|LNC2HPO|Hypocholesterolemia|Hypocholesterolemia
C0364214|T201|MTH_LN|2082-6|LNC2HPO|Hypocholesterolemia|Hypocholesterolemia
C0364214|T201|OSN|2082-6|LNC2HPO|Hypocholesterolemia|Hypocholesterolemia
C0364214|T201|LC|2082-6|LNC2HPO|Hypocholesterolemia|Hypocholesterolemia
C0880188|T201|LN|22670-4|LNC2HPO|Hyperisoleucinemia|Hyperisoleucinemia
C0880188|T201|DN|22670-4|LNC2HPO|Hyperisoleucinemia|Hyperisoleucinemia
C0880188|T201|MTH_LN|22670-4|LNC2HPO|Hyperisoleucinemia|Hyperisoleucinemia
C0880188|T201|OSN|22670-4|LNC2HPO|Hyperisoleucinemia|Hyperisoleucinemia
C0880188|T201|LC|22670-4|LNC2HPO|Hyperisoleucinemia|Hyperisoleucinemia
C0880188|T201|LN|22670-4|LNC2HPO|Hypoisoleucinemia|Hypoisoleucinemia
C0880188|T201|DN|22670-4|LNC2HPO|Hypoisoleucinemia|Hypoisoleucinemia
C0880188|T201|MTH_LN|22670-4|LNC2HPO|Hypoisoleucinemia|Hypoisoleucinemia
C0880188|T201|OSN|22670-4|LNC2HPO|Hypoisoleucinemia|Hypoisoleucinemia
C0880188|T201|LC|22670-4|LNC2HPO|Hypoisoleucinemia|Hypoisoleucinemia
C0881402|T201|LN|24082-0|LNC2HPO|Impairment of galactose metabolism|Impairment of galactose metabolism
C0881402|T201|DN|24082-0|LNC2HPO|Impairment of galactose metabolism|Impairment of galactose metabolism
C0881402|T201|MTH_LN|24082-0|LNC2HPO|Impairment of galactose metabolism|Impairment of galactose metabolism
C0881402|T201|OSN|24082-0|LNC2HPO|Impairment of galactose metabolism|Impairment of galactose metabolism
C0881402|T201|LC|24082-0|LNC2HPO|Impairment of galactose metabolism|Impairment of galactose metabolism
C0881402|T201|LN|24082-0|LNC2HPO|Impaired galactose metabolism|Impaired galactose metabolism
C0881402|T201|DN|24082-0|LNC2HPO|Impaired galactose metabolism|Impaired galactose metabolism
C0881402|T201|MTH_LN|24082-0|LNC2HPO|Impaired galactose metabolism|Impaired galactose metabolism
C0881402|T201|OSN|24082-0|LNC2HPO|Impaired galactose metabolism|Impaired galactose metabolism
C0881402|T201|LC|24082-0|LNC2HPO|Impaired galactose metabolism|Impaired galactose metabolism
C0881402|T201|LN|24082-0|LNC2HPO|Galactosemia|Galactosemia
C0881402|T201|DN|24082-0|LNC2HPO|Galactosemia|Galactosemia
C0881402|T201|MTH_LN|24082-0|LNC2HPO|Galactosemia|Galactosemia
C0881402|T201|OSN|24082-0|LNC2HPO|Galactosemia|Galactosemia
C0881402|T201|LC|24082-0|LNC2HPO|Galactosemia|Galactosemia
C0881402|T201|LN|24082-0|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0881402|T201|DN|24082-0|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0881402|T201|MTH_LN|24082-0|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0881402|T201|OSN|24082-0|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0881402|T201|LC|24082-0|LNC2HPO|Hypergalactosemia|Hypergalactosemia
C0881717|T201|MTH_LN|24467-3|LNC2HPO|CD4+ T-cell lymphopenia|CD4+ T-cell lymphopenia
C0881717|T201|LC|24467-3|LNC2HPO|CD4+ T-cell lymphopenia|CD4+ T-cell lymphopenia
C0881717|T201|DN|24467-3|LNC2HPO|CD4+ T-cell lymphopenia|CD4+ T-cell lymphopenia
C0881717|T201|LN|24467-3|LNC2HPO|CD4+ T-cell lymphopenia|CD4+ T-cell lymphopenia
C0881717|T201|OSN|24467-3|LNC2HPO|CD4+ T-cell lymphopenia|CD4+ T-cell lymphopenia
C0881717|T201|MTH_LN|24467-3|LNC2HPO|CD4 T cell lymphopenia|CD4 T cell lymphopenia
C0881717|T201|LC|24467-3|LNC2HPO|CD4 T cell lymphopenia|CD4 T cell lymphopenia
C0881717|T201|DN|24467-3|LNC2HPO|CD4 T cell lymphopenia|CD4 T cell lymphopenia
C0881717|T201|LN|24467-3|LNC2HPO|CD4 T cell lymphopenia|CD4 T cell lymphopenia
C0881717|T201|OSN|24467-3|LNC2HPO|CD4 T cell lymphopenia|CD4 T cell lymphopenia
C0364607|T201|LN|2467-9|LNC2HPO|Immunoglobulin IgG2 deficiency|Immunoglobulin IgG2 deficiency
C0364607|T201|MTH_LN|2467-9|LNC2HPO|Immunoglobulin IgG2 deficiency|Immunoglobulin IgG2 deficiency
C0364607|T201|DN|2467-9|LNC2HPO|Immunoglobulin IgG2 deficiency|Immunoglobulin IgG2 deficiency
C0364607|T201|OSN|2467-9|LNC2HPO|Immunoglobulin IgG2 deficiency|Immunoglobulin IgG2 deficiency
C0364607|T201|LC|2467-9|LNC2HPO|Immunoglobulin IgG2 deficiency|Immunoglobulin IgG2 deficiency
C0941297|T201|LN|25087-8|LNC2HPO|3-Methylglutaconic aciduria|3-Methylglutaconic aciduria
C0941297|T201|DN|25087-8|LNC2HPO|3-Methylglutaconic aciduria|3-Methylglutaconic aciduria
C0941297|T201|OSN|25087-8|LNC2HPO|3-Methylglutaconic aciduria|3-Methylglutaconic aciduria
C0941297|T201|LC|25087-8|LNC2HPO|3-Methylglutaconic aciduria|3-Methylglutaconic aciduria
C0941297|T201|MTH_LN|25087-8|LNC2HPO|3-Methylglutaconic aciduria|3-Methylglutaconic aciduria
C0941297|T201|LN|25087-8|LNC2HPO|3-Methylglutaconicaciduria|3-Methylglutaconicaciduria
C0941297|T201|DN|25087-8|LNC2HPO|3-Methylglutaconicaciduria|3-Methylglutaconicaciduria
C0941297|T201|OSN|25087-8|LNC2HPO|3-Methylglutaconicaciduria|3-Methylglutaconicaciduria
C0941297|T201|LC|25087-8|LNC2HPO|3-Methylglutaconicaciduria|3-Methylglutaconicaciduria
C0941297|T201|MTH_LN|25087-8|LNC2HPO|3-Methylglutaconicaciduria|3-Methylglutaconicaciduria
C0941601|T201|LN|25464-9|LNC2HPO|Hyperlysinuria|Hyperlysinuria
C0941601|T201|DN|25464-9|LNC2HPO|Hyperlysinuria|Hyperlysinuria
C0941601|T201|MTH_LN|25464-9|LNC2HPO|Hyperlysinuria|Hyperlysinuria
C0941601|T201|OSN|25464-9|LNC2HPO|Hyperlysinuria|Hyperlysinuria
C0941601|T201|LC|25464-9|LNC2HPO|Hyperlysinuria|Hyperlysinuria
C0941601|T201|LN|25464-9|LNC2HPO|Lysinuria|Lysinuria
C0941601|T201|DN|25464-9|LNC2HPO|Lysinuria|Lysinuria
C0941601|T201|MTH_LN|25464-9|LNC2HPO|Lysinuria|Lysinuria
C0941601|T201|OSN|25464-9|LNC2HPO|Lysinuria|Lysinuria
C0941601|T201|LC|25464-9|LNC2HPO|Lysinuria|Lysinuria
C0941624|T201|LN|25491-2|LNC2HPO|Ornithinuria|Ornithinuria
C0941624|T201|DN|25491-2|LNC2HPO|Ornithinuria|Ornithinuria
C0941624|T201|MTH_LN|25491-2|LNC2HPO|Ornithinuria|Ornithinuria
C0941624|T201|OSN|25491-2|LNC2HPO|Ornithinuria|Ornithinuria
C0941624|T201|LC|25491-2|LNC2HPO|Ornithinuria|Ornithinuria
C0364712|T201|LN|2569-2|LNC2HPO|Dyslipidemia|Dyslipidemia
C0364712|T201|MTH_LN|2569-2|LNC2HPO|Dyslipidemia|Dyslipidemia
C0364712|T201|DN|2569-2|LNC2HPO|Dyslipidemia|Dyslipidemia
C0364712|T201|OSN|2569-2|LNC2HPO|Dyslipidemia|Dyslipidemia
C0364712|T201|LC|2569-2|LNC2HPO|Dyslipidemia|Dyslipidemia
C0364712|T201|LN|2569-2|LNC2HPO|Hyperlipidemia|Hyperlipidemia
C0364712|T201|MTH_LN|2569-2|LNC2HPO|Hyperlipidemia|Hyperlipidemia
C0364712|T201|DN|2569-2|LNC2HPO|Hyperlipidemia|Hyperlipidemia
C0364712|T201|OSN|2569-2|LNC2HPO|Hyperlipidemia|Hyperlipidemia
C0364712|T201|LC|2569-2|LNC2HPO|Hyperlipidemia|Hyperlipidemia
C0364712|T201|LN|2569-2|LNC2HPO|Hypolipidemia|Hypolipidemia
C0364712|T201|MTH_LN|2569-2|LNC2HPO|Hypolipidemia|Hypolipidemia
C0364712|T201|DN|2569-2|LNC2HPO|Hypolipidemia|Hypolipidemia
C0364712|T201|OSN|2569-2|LNC2HPO|Hypolipidemia|Hypolipidemia
C0364712|T201|LC|2569-2|LNC2HPO|Hypolipidemia|Hypolipidemia
C0364774|T201|LN|2629-4|LNC2HPO|Methylmalonic acidemia|Methylmalonic acidemia
C0364774|T201|DN|2629-4|LNC2HPO|Methylmalonic acidemia|Methylmalonic acidemia
C0364774|T201|MTH_LN|2629-4|LNC2HPO|Methylmalonic acidemia|Methylmalonic acidemia
C0364774|T201|OSN|2629-4|LNC2HPO|Methylmalonic acidemia|Methylmalonic acidemia
C0364774|T201|LC|2629-4|LNC2HPO|Methylmalonic acidemia|Methylmalonic acidemia
C0942546|T201|LN|26604-9|LNC2HPO|Hyperbetaalaninemia|Hyperbetaalaninemia
C0942546|T201|DN|26604-9|LNC2HPO|Hyperbetaalaninemia|Hyperbetaalaninemia
C0942546|T201|MTH_LN|26604-9|LNC2HPO|Hyperbetaalaninemia|Hyperbetaalaninemia
C0942546|T201|OSN|26604-9|LNC2HPO|Hyperbetaalaninemia|Hyperbetaalaninemia
C0942546|T201|LC|26604-9|LNC2HPO|Hyperbetaalaninemia|Hyperbetaalaninemia
C0942546|T201|LN|26604-9|LNC2HPO|Hyperbeta-alaninemia|Hyperbeta-alaninemia
C0942546|T201|DN|26604-9|LNC2HPO|Hyperbeta-alaninemia|Hyperbeta-alaninemia
C0942546|T201|MTH_LN|26604-9|LNC2HPO|Hyperbeta-alaninemia|Hyperbeta-alaninemia
C0942546|T201|OSN|26604-9|LNC2HPO|Hyperbeta-alaninemia|Hyperbeta-alaninemia
C0942546|T201|LC|26604-9|LNC2HPO|Hyperbeta-alaninemia|Hyperbeta-alaninemia
C0942660|T201|LN|26740-1|LNC2HPO|Hydroxyprolinuria|Hydroxyprolinuria
C0942660|T201|DN|26740-1|LNC2HPO|Hydroxyprolinuria|Hydroxyprolinuria
C0942660|T201|MTH_LN|26740-1|LNC2HPO|Hydroxyprolinuria|Hydroxyprolinuria
C0942660|T201|OSN|26740-1|LNC2HPO|Hydroxyprolinuria|Hydroxyprolinuria
C0942660|T201|LC|26740-1|LNC2HPO|Hydroxyprolinuria|Hydroxyprolinuria
C0942745|T201|LN|26843-3|LNC2HPO|Cystinuria|Cystinuria
C0942745|T201|MTH_LN|26843-3|LNC2HPO|Cystinuria|Cystinuria
C0942745|T201|DN|26843-3|LNC2HPO|Cystinuria|Cystinuria
C0942745|T201|OSN|26843-3|LNC2HPO|Cystinuria|Cystinuria
C0942745|T201|LC|26843-3|LNC2HPO|Cystinuria|Cystinuria
C0945434|T201|LN|26971-2|LNC2HPO|Smooth muscle antibody positive|Smooth muscle antibody positive
C0945434|T201|MTH_LN|26971-2|LNC2HPO|Smooth muscle antibody positive|Smooth muscle antibody positive
C0945434|T201|DN|26971-2|LNC2HPO|Smooth muscle antibody positive|Smooth muscle antibody positive
C0945434|T201|OSN|26971-2|LNC2HPO|Smooth muscle antibody positive|Smooth muscle antibody positive
C0945434|T201|LC|26971-2|LNC2HPO|Smooth muscle antibody positive|Smooth muscle antibody positive
C0364844|T201|LN|2701-1|LNC2HPO|Hyperoxaluria|Hyperoxaluria
C0364844|T201|MTH_LN|2701-1|LNC2HPO|Hyperoxaluria|Hyperoxaluria
C0364844|T201|DN|2701-1|LNC2HPO|Hyperoxaluria|Hyperoxaluria
C0364844|T201|OSN|2701-1|LNC2HPO|Hyperoxaluria|Hyperoxaluria
C0364844|T201|LC|2701-1|LNC2HPO|Hyperoxaluria|Hyperoxaluria
C1145646|T201|LN|2704-5|LNC2HPO|Hyperoxemia|Hyperoxemia
C1145646|T201|MTH_LN|2704-5|LNC2HPO|Hyperoxemia|Hyperoxemia
C1145646|T201|DN|2704-5|LNC2HPO|Hyperoxemia|Hyperoxemia
C1145646|T201|LC|2704-5|LNC2HPO|Hyperoxemia|Hyperoxemia
C1145646|T201|OSN|2704-5|LNC2HPO|Hyperoxemia|Hyperoxemia
C1145646|T201|LN|2704-5|LNC2HPO|Hypoxemia|Hypoxemia
C1145646|T201|MTH_LN|2704-5|LNC2HPO|Hypoxemia|Hypoxemia
C1145646|T201|DN|2704-5|LNC2HPO|Hypoxemia|Hypoxemia
C1145646|T201|LC|2704-5|LNC2HPO|Hypoxemia|Hypoxemia
C1145646|T201|OSN|2704-5|LNC2HPO|Hypoxemia|Hypoxemia
C1145647|T201|LN|2705-2|LNC2HPO|Hyperoxemia|Hyperoxemia
C1145647|T201|MTH_LN|2705-2|LNC2HPO|Hyperoxemia|Hyperoxemia
C1145647|T201|DN|2705-2|LNC2HPO|Hyperoxemia|Hyperoxemia
C1145647|T201|LC|2705-2|LNC2HPO|Hyperoxemia|Hyperoxemia
C1145647|T201|OSN|2705-2|LNC2HPO|Hyperoxemia|Hyperoxemia
C1145647|T201|LN|2705-2|LNC2HPO|Hypoxemia|Hypoxemia
C1145647|T201|MTH_LN|2705-2|LNC2HPO|Hypoxemia|Hypoxemia
C1145647|T201|DN|2705-2|LNC2HPO|Hypoxemia|Hypoxemia
C1145647|T201|LC|2705-2|LNC2HPO|Hypoxemia|Hypoxemia
C1145647|T201|OSN|2705-2|LNC2HPO|Hypoxemia|Hypoxemia
C0364852|T201|LN|2709-4|LNC2HPO|Hyperoxemia|Hyperoxemia
C0364852|T201|LC|2709-4|LNC2HPO|Hyperoxemia|Hyperoxemia
C0364852|T201|MTH_LN|2709-4|LNC2HPO|Hyperoxemia|Hyperoxemia
C0364852|T201|OSN|2709-4|LNC2HPO|Hyperoxemia|Hyperoxemia
C0364852|T201|LN|2709-4|LNC2HPO|Hypoxemia|Hypoxemia
C0364852|T201|LC|2709-4|LNC2HPO|Hypoxemia|Hypoxemia
C0364852|T201|MTH_LN|2709-4|LNC2HPO|Hypoxemia|Hypoxemia
C0364852|T201|OSN|2709-4|LNC2HPO|Hypoxemia|Hypoxemia
C0943118|T201|LN|27298-9|LNC2HPO|Proteinuria|Proteinuria
C0943118|T201|DN|27298-9|LNC2HPO|Proteinuria|Proteinuria
C0943118|T201|MTH_LN|27298-9|LNC2HPO|Proteinuria|Proteinuria
C0943118|T201|OSN|27298-9|LNC2HPO|Proteinuria|Proteinuria
C0943118|T201|LC|27298-9|LNC2HPO|Proteinuria|Proteinuria
C0364874|T201|LC|2731-8|LNC2HPO|Parathyroid dysfunction|Parathyroid dysfunction
C0364874|T201|DN|2731-8|LNC2HPO|Parathyroid dysfunction|Parathyroid dysfunction
C0364874|T201|MTH_LN|2731-8|LNC2HPO|Parathyroid dysfunction|Parathyroid dysfunction
C0364874|T201|LN|2731-8|LNC2HPO|Parathyroid dysfunction|Parathyroid dysfunction
C0364874|T201|OSN|2731-8|LNC2HPO|Parathyroid dysfunction|Parathyroid dysfunction
C0364874|T201|LC|2731-8|LNC2HPO|Parathyroid issue|Parathyroid issue
C0364874|T201|DN|2731-8|LNC2HPO|Parathyroid issue|Parathyroid issue
C0364874|T201|MTH_LN|2731-8|LNC2HPO|Parathyroid issue|Parathyroid issue
C0364874|T201|LN|2731-8|LNC2HPO|Parathyroid issue|Parathyroid issue
C0364874|T201|OSN|2731-8|LNC2HPO|Parathyroid issue|Parathyroid issue
C0364874|T201|LC|2731-8|LNC2HPO|Hyperparathyroidism|Hyperparathyroidism
C0364874|T201|DN|2731-8|LNC2HPO|Hyperparathyroidism|Hyperparathyroidism
C0364874|T201|MTH_LN|2731-8|LNC2HPO|Hyperparathyroidism|Hyperparathyroidism
C0364874|T201|LN|2731-8|LNC2HPO|Hyperparathyroidism|Hyperparathyroidism
C0364874|T201|OSN|2731-8|LNC2HPO|Hyperparathyroidism|Hyperparathyroidism
C0364874|T201|LC|2731-8|LNC2HPO|Hypoparathyroidism|Hypoparathyroidism
C0364874|T201|DN|2731-8|LNC2HPO|Hypoparathyroidism|Hypoparathyroidism
C0364874|T201|MTH_LN|2731-8|LNC2HPO|Hypoparathyroidism|Hypoparathyroidism
C0364874|T201|LN|2731-8|LNC2HPO|Hypoparathyroidism|Hypoparathyroidism
C0364874|T201|OSN|2731-8|LNC2HPO|Hypoparathyroidism|Hypoparathyroidism
C0364887|T201|LN|2744-1|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364887|T201|LC|2744-1|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364887|T201|MTH_LN|2744-1|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364887|T201|OSN|2744-1|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364887|T201|DN|2744-1|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364887|T201|LN|2744-1|LNC2HPO|Alkalemia|Alkalemia
C0364887|T201|LC|2744-1|LNC2HPO|Alkalemia|Alkalemia
C0364887|T201|MTH_LN|2744-1|LNC2HPO|Alkalemia|Alkalemia
C0364887|T201|OSN|2744-1|LNC2HPO|Alkalemia|Alkalemia
C0364887|T201|DN|2744-1|LNC2HPO|Alkalemia|Alkalemia
C0364887|T201|LN|2744-1|LNC2HPO|Acidemia|Acidemia
C0364887|T201|LC|2744-1|LNC2HPO|Acidemia|Acidemia
C0364887|T201|MTH_LN|2744-1|LNC2HPO|Acidemia|Acidemia
C0364887|T201|OSN|2744-1|LNC2HPO|Acidemia|Acidemia
C0364887|T201|DN|2744-1|LNC2HPO|Acidemia|Acidemia
C0364888|T201|MTH_LN|2745-8|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364888|T201|LN|2745-8|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364888|T201|OSN|2745-8|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364888|T201|DN|2745-8|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364888|T201|LC|2745-8|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364888|T201|MTH_LN|2745-8|LNC2HPO|Alkalemia|Alkalemia
C0364888|T201|LN|2745-8|LNC2HPO|Alkalemia|Alkalemia
C0364888|T201|OSN|2745-8|LNC2HPO|Alkalemia|Alkalemia
C0364888|T201|DN|2745-8|LNC2HPO|Alkalemia|Alkalemia
C0364888|T201|LC|2745-8|LNC2HPO|Alkalemia|Alkalemia
C0364888|T201|MTH_LN|2745-8|LNC2HPO|Acidemia|Acidemia
C0364888|T201|LN|2745-8|LNC2HPO|Acidemia|Acidemia
C0364888|T201|OSN|2745-8|LNC2HPO|Acidemia|Acidemia
C0364888|T201|DN|2745-8|LNC2HPO|Acidemia|Acidemia
C0364888|T201|LC|2745-8|LNC2HPO|Acidemia|Acidemia
C0364889|T201|LN|2746-6|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364889|T201|LC|2746-6|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364889|T201|MTH_LN|2746-6|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364889|T201|OSN|2746-6|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364889|T201|DN|2746-6|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364889|T201|LN|2746-6|LNC2HPO|Alkalemia|Alkalemia
C0364889|T201|LC|2746-6|LNC2HPO|Alkalemia|Alkalemia
C0364889|T201|MTH_LN|2746-6|LNC2HPO|Alkalemia|Alkalemia
C0364889|T201|OSN|2746-6|LNC2HPO|Alkalemia|Alkalemia
C0364889|T201|DN|2746-6|LNC2HPO|Alkalemia|Alkalemia
C0364889|T201|LN|2746-6|LNC2HPO|Acidemia|Acidemia
C0364889|T201|LC|2746-6|LNC2HPO|Acidemia|Acidemia
C0364889|T201|MTH_LN|2746-6|LNC2HPO|Acidemia|Acidemia
C0364889|T201|OSN|2746-6|LNC2HPO|Acidemia|Acidemia
C0364889|T201|DN|2746-6|LNC2HPO|Acidemia|Acidemia
C0364899|T201|LN|2756-5|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364899|T201|LC|2756-5|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364899|T201|DN|2756-5|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364899|T201|MTH_LN|2756-5|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364899|T201|OSN|2756-5|LNC2HPO|Acid base imbalance|Acid base imbalance
C0364899|T201|LN|2756-5|LNC2HPO|Alkalemia|Alkalemia
C0364899|T201|LC|2756-5|LNC2HPO|Alkalemia|Alkalemia
C0364899|T201|DN|2756-5|LNC2HPO|Alkalemia|Alkalemia
C0364899|T201|MTH_LN|2756-5|LNC2HPO|Alkalemia|Alkalemia
C0364899|T201|OSN|2756-5|LNC2HPO|Alkalemia|Alkalemia
C0364899|T201|LN|2756-5|LNC2HPO|Acidemia|Acidemia
C0364899|T201|LC|2756-5|LNC2HPO|Acidemia|Acidemia
C0364899|T201|DN|2756-5|LNC2HPO|Acidemia|Acidemia
C0364899|T201|MTH_LN|2756-5|LNC2HPO|Acidemia|Acidemia
C0364899|T201|OSN|2756-5|LNC2HPO|Acidemia|Acidemia
C0364906|T201|LN|2765-6|LNC2HPO|Hyperphenylalaninemia|Hyperphenylalaninemia
C0364906|T201|MTH_LN|2765-6|LNC2HPO|Hyperphenylalaninemia|Hyperphenylalaninemia
C0364906|T201|DN|2765-6|LNC2HPO|Hyperphenylalaninemia|Hyperphenylalaninemia
C0364906|T201|OSN|2765-6|LNC2HPO|Hyperphenylalaninemia|Hyperphenylalaninemia
C0364906|T201|LC|2765-6|LNC2HPO|Hyperphenylalaninemia|Hyperphenylalaninemia
C0364906|T201|LN|2765-6|LNC2HPO|Hypophenylalaninemia|Hypophenylalaninemia
C0364906|T201|MTH_LN|2765-6|LNC2HPO|Hypophenylalaninemia|Hypophenylalaninemia
C0364906|T201|DN|2765-6|LNC2HPO|Hypophenylalaninemia|Hypophenylalaninemia
C0364906|T201|OSN|2765-6|LNC2HPO|Hypophenylalaninemia|Hypophenylalaninemia
C0364906|T201|LC|2765-6|LNC2HPO|Hypophenylalaninemia|Hypophenylalaninemia
C0943506|T201|LN|27811-9|LNC2HPO|Antithrombin III deficiency|Antithrombin III deficiency
C0943506|T201|DN|27811-9|LNC2HPO|Antithrombin III deficiency|Antithrombin III deficiency
C0943506|T201|OSN|27811-9|LNC2HPO|Antithrombin III deficiency|Antithrombin III deficiency
C0943506|T201|MTH_LN|27811-9|LNC2HPO|Antithrombin III deficiency|Antithrombin III deficiency
C0943506|T201|LC|27811-9|LNC2HPO|Antithrombin III deficiency|Antithrombin III deficiency
C0943506|T201|LN|27811-9|LNC2HPO|Anti-thrombin III deficiency|Anti-thrombin III deficiency
C0943506|T201|DN|27811-9|LNC2HPO|Anti-thrombin III deficiency|Anti-thrombin III deficiency
C0943506|T201|OSN|27811-9|LNC2HPO|Anti-thrombin III deficiency|Anti-thrombin III deficiency
C0943506|T201|MTH_LN|27811-9|LNC2HPO|Anti-thrombin III deficiency|Anti-thrombin III deficiency
C0943506|T201|LC|27811-9|LNC2HPO|Anti-thrombin III deficiency|Anti-thrombin III deficiency
C0944184|T201|LN|28597-3|LNC2HPO|Carnosinuria|Carnosinuria
C0944184|T201|DN|28597-3|LNC2HPO|Carnosinuria|Carnosinuria
C0944184|T201|MTH_LN|28597-3|LNC2HPO|Carnosinuria|Carnosinuria
C0944184|T201|OSN|28597-3|LNC2HPO|Carnosinuria|Carnosinuria
C0944184|T201|LC|28597-3|LNC2HPO|Carnosinuria|Carnosinuria
C0944185|T201|LN|28599-9|LNC2HPO|Cystathioninuria|Cystathioninuria
C0944185|T201|DN|28599-9|LNC2HPO|Cystathioninuria|Cystathioninuria
C0944185|T201|MTH_LN|28599-9|LNC2HPO|Cystathioninuria|Cystathioninuria
C0944185|T201|OSN|28599-9|LNC2HPO|Cystathioninuria|Cystathioninuria
C0944185|T201|LC|28599-9|LNC2HPO|Cystathioninuria|Cystathioninuria
C0945632|T201|LN|28601-3|LNC2HPO|Hydroxyprolinuria|Hydroxyprolinuria
C0945632|T201|DN|28601-3|LNC2HPO|Hydroxyprolinuria|Hydroxyprolinuria
C0945632|T201|MTH_LN|28601-3|LNC2HPO|Hydroxyprolinuria|Hydroxyprolinuria
C0945632|T201|OSN|28601-3|LNC2HPO|Hydroxyprolinuria|Hydroxyprolinuria
C0945632|T201|LC|28601-3|LNC2HPO|Hydroxyprolinuria|Hydroxyprolinuria
C0944189|T201|LN|28604-7|LNC2HPO|Phosphoethanolaminuria|Phosphoethanolaminuria
C0944189|T201|DN|28604-7|LNC2HPO|Phosphoethanolaminuria|Phosphoethanolaminuria
C0944189|T201|MTH_LN|28604-7|LNC2HPO|Phosphoethanolaminuria|Phosphoethanolaminuria
C0944189|T201|OSN|28604-7|LNC2HPO|Phosphoethanolaminuria|Phosphoethanolaminuria
C0944189|T201|LC|28604-7|LNC2HPO|Phosphoethanolaminuria|Phosphoethanolaminuria
C0944192|T201|LN|28608-8|LNC2HPO|Tryptophanuria|Tryptophanuria
C0944192|T201|DN|28608-8|LNC2HPO|Tryptophanuria|Tryptophanuria
C0944192|T201|MTH_LN|28608-8|LNC2HPO|Tryptophanuria|Tryptophanuria
C0944192|T201|OSN|28608-8|LNC2HPO|Tryptophanuria|Tryptophanuria
C0944192|T201|LC|28608-8|LNC2HPO|Tryptophanuria|Tryptophanuria
C0365005|T201|LN|2862-1|LNC2HPO|Hyperalbuminemia|Hyperalbuminemia
C0365005|T201|DN|2862-1|LNC2HPO|Hyperalbuminemia|Hyperalbuminemia
C0365005|T201|MTH_LN|2862-1|LNC2HPO|Hyperalbuminemia|Hyperalbuminemia
C0365005|T201|OSN|2862-1|LNC2HPO|Hyperalbuminemia|Hyperalbuminemia
C0365005|T201|LC|2862-1|LNC2HPO|Hyperalbuminemia|Hyperalbuminemia
C0365005|T201|LN|2862-1|LNC2HPO|Hyperalbuminaemia|Hyperalbuminaemia
C0365005|T201|DN|2862-1|LNC2HPO|Hyperalbuminaemia|Hyperalbuminaemia
C0365005|T201|MTH_LN|2862-1|LNC2HPO|Hyperalbuminaemia|Hyperalbuminaemia
C0365005|T201|OSN|2862-1|LNC2HPO|Hyperalbuminaemia|Hyperalbuminaemia
C0365005|T201|LC|2862-1|LNC2HPO|Hyperalbuminaemia|Hyperalbuminaemia
C0365005|T201|LN|2862-1|LNC2HPO|Hypoalbuminemia|Hypoalbuminemia
C0365005|T201|DN|2862-1|LNC2HPO|Hypoalbuminemia|Hypoalbuminemia
C0365005|T201|MTH_LN|2862-1|LNC2HPO|Hypoalbuminemia|Hypoalbuminemia
C0365005|T201|OSN|2862-1|LNC2HPO|Hypoalbuminemia|Hypoalbuminemia
C0365005|T201|LC|2862-1|LNC2HPO|Hypoalbuminemia|Hypoalbuminemia
C0365005|T201|LN|2862-1|LNC2HPO|Hypoalbuminaemia|Hypoalbuminaemia
C0365005|T201|DN|2862-1|LNC2HPO|Hypoalbuminaemia|Hypoalbuminaemia
C0365005|T201|MTH_LN|2862-1|LNC2HPO|Hypoalbuminaemia|Hypoalbuminaemia
C0365005|T201|OSN|2862-1|LNC2HPO|Hypoalbuminaemia|Hypoalbuminaemia
C0365005|T201|LC|2862-1|LNC2HPO|Hypoalbuminaemia|Hypoalbuminaemia
C0365059|T201|LN|2915-7|LNC2HPO|Hyperreninemia|Hyperreninemia
C0365059|T201|MTH_LN|2915-7|LNC2HPO|Hyperreninemia|Hyperreninemia
C0365059|T201|DN|2915-7|LNC2HPO|Hyperreninemia|Hyperreninemia
C0365059|T201|OSN|2915-7|LNC2HPO|Hyperreninemia|Hyperreninemia
C0365059|T201|LC|2915-7|LNC2HPO|Hyperreninemia|Hyperreninemia
C0944742|T201|LN|29261-5|LNC2HPO|Lymphocytosis|Lymphocytosis
C0944742|T201|OSN|29261-5|LNC2HPO|Lymphocytosis|Lymphocytosis
C0944742|T201|DN|29261-5|LNC2HPO|Lymphocytosis|Lymphocytosis
C0944742|T201|MTH_LN|29261-5|LNC2HPO|Lymphocytosis|Lymphocytosis
C0944742|T201|LC|29261-5|LNC2HPO|Lymphocytosis|Lymphocytosis
C0944742|T201|LN|29261-5|LNC2HPO|Lymphopenia|Lymphopenia
C0944742|T201|OSN|29261-5|LNC2HPO|Lymphopenia|Lymphopenia
C0944742|T201|DN|29261-5|LNC2HPO|Lymphopenia|Lymphopenia
C0944742|T201|MTH_LN|29261-5|LNC2HPO|Lymphopenia|Lymphopenia
C0944742|T201|LC|29261-5|LNC2HPO|Lymphopenia|Lymphopenia
C0944742|T201|LN|29261-5|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0944742|T201|OSN|29261-5|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0944742|T201|DN|29261-5|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0944742|T201|MTH_LN|29261-5|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0944742|T201|LC|29261-5|LNC2HPO|Lymphocytopenia|Lymphocytopenia
C0944742|T201|LN|29261-5|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0944742|T201|OSN|29261-5|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0944742|T201|DN|29261-5|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0944742|T201|MTH_LN|29261-5|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0944742|T201|LC|29261-5|LNC2HPO|Absolute lymphocyte count decrease|Absolute lymphocyte count decrease
C0945006|T201|LN|29572-5|LNC2HPO|Hyperphenylalaninemia|Hyperphenylalaninemia
C0945006|T201|LC|29572-5|LNC2HPO|Hyperphenylalaninemia|Hyperphenylalaninemia
C0945006|T201|DN|29572-5|LNC2HPO|Hyperphenylalaninemia|Hyperphenylalaninemia
C0945006|T201|MTH_LN|29572-5|LNC2HPO|Hyperphenylalaninemia|Hyperphenylalaninemia
C0945006|T201|OSN|29572-5|LNC2HPO|Hyperphenylalaninemia|Hyperphenylalaninemia
C0945006|T201|LN|29572-5|LNC2HPO|Hypophenylalaninemia|Hypophenylalaninemia
C0945006|T201|LC|29572-5|LNC2HPO|Hypophenylalaninemia|Hypophenylalaninemia
C0945006|T201|DN|29572-5|LNC2HPO|Hypophenylalaninemia|Hypophenylalaninemia
C0945006|T201|MTH_LN|29572-5|LNC2HPO|Hypophenylalaninemia|Hypophenylalaninemia
C0945006|T201|OSN|29572-5|LNC2HPO|Hypophenylalaninemia|Hypophenylalaninemia
C0945007|T201|LN|29573-3|LNC2HPO|Hyperphenylalaninemia|Hyperphenylalaninemia
C0945007|T201|LC|29573-3|LNC2HPO|Hyperphenylalaninemia|Hyperphenylalaninemia
C0945007|T201|DN|29573-3|LNC2HPO|Hyperphenylalaninemia|Hyperphenylalaninemia
C0945007|T201|MTH_LN|29573-3|LNC2HPO|Hyperphenylalaninemia|Hyperphenylalaninemia
C0945007|T201|OSN|29573-3|LNC2HPO|Hyperphenylalaninemia|Hyperphenylalaninemia
C0945007|T201|LN|29573-3|LNC2HPO|Hypophenylalaninemia|Hypophenylalaninemia
C0945007|T201|LC|29573-3|LNC2HPO|Hypophenylalaninemia|Hypophenylalaninemia
C0945007|T201|DN|29573-3|LNC2HPO|Hypophenylalaninemia|Hypophenylalaninemia
C0945007|T201|MTH_LN|29573-3|LNC2HPO|Hypophenylalaninemia|Hypophenylalaninemia
C0945007|T201|OSN|29573-3|LNC2HPO|Hypophenylalaninemia|Hypophenylalaninemia
C1114843|T201|LN|29953-7|LNC2HPO|Antinuclear antibodies|Antinuclear antibodies
C1114843|T201|DN|29953-7|LNC2HPO|Antinuclear antibodies|Antinuclear antibodies
C1114843|T201|MTH_LN|29953-7|LNC2HPO|Antinuclear antibodies|Antinuclear antibodies
C1114843|T201|OSN|29953-7|LNC2HPO|Antinuclear antibodies|Antinuclear antibodies
C1114843|T201|LC|29953-7|LNC2HPO|Antinuclear antibodies|Antinuclear antibodies
C1114843|T201|LN|29953-7|LNC2HPO|Antinuclear antibody positive|Antinuclear antibody positive
C1114843|T201|DN|29953-7|LNC2HPO|Antinuclear antibody positive|Antinuclear antibody positive
C1114843|T201|MTH_LN|29953-7|LNC2HPO|Antinuclear antibody positive|Antinuclear antibody positive
C1114843|T201|OSN|29953-7|LNC2HPO|Antinuclear antibody positive|Antinuclear antibody positive
C1114843|T201|LC|29953-7|LNC2HPO|Antinuclear antibody positive|Antinuclear antibody positive
C1114843|T201|LN|29953-7|LNC2HPO|Serum antinuclear antibody|Serum antinuclear antibody
C1114843|T201|DN|29953-7|LNC2HPO|Serum antinuclear antibody|Serum antinuclear antibody
C1114843|T201|MTH_LN|29953-7|LNC2HPO|Serum antinuclear antibody|Serum antinuclear antibody
C1114843|T201|OSN|29953-7|LNC2HPO|Serum antinuclear antibody|Serum antinuclear antibody
C1114843|T201|LC|29953-7|LNC2HPO|Serum antinuclear antibody|Serum antinuclear antibody
C1113951|T201|LN|30047-5|LNC2HPO|Histidinuria|Histidinuria
C1113951|T201|DN|30047-5|LNC2HPO|Histidinuria|Histidinuria
C1113951|T201|MTH_LN|30047-5|LNC2HPO|Histidinuria|Histidinuria
C1113951|T201|OSN|30047-5|LNC2HPO|Histidinuria|Histidinuria
C1113951|T201|LC|30047-5|LNC2HPO|Histidinuria|Histidinuria
C1114856|T201|LN|30048-3|LNC2HPO|Hyperlysinuria|Hyperlysinuria
C1114856|T201|DN|30048-3|LNC2HPO|Hyperlysinuria|Hyperlysinuria
C1114856|T201|MTH_LN|30048-3|LNC2HPO|Hyperlysinuria|Hyperlysinuria
C1114856|T201|OSN|30048-3|LNC2HPO|Hyperlysinuria|Hyperlysinuria
C1114856|T201|LC|30048-3|LNC2HPO|Hyperlysinuria|Hyperlysinuria
C1114856|T201|LN|30048-3|LNC2HPO|Lysinuria|Lysinuria
C1114856|T201|DN|30048-3|LNC2HPO|Lysinuria|Lysinuria
C1114856|T201|MTH_LN|30048-3|LNC2HPO|Lysinuria|Lysinuria
C1114856|T201|OSN|30048-3|LNC2HPO|Lysinuria|Lysinuria
C1114856|T201|LC|30048-3|LNC2HPO|Lysinuria|Lysinuria
C1113952|T201|LN|30049-1|LNC2HPO|Ornithinuria|Ornithinuria
C1113952|T201|DN|30049-1|LNC2HPO|Ornithinuria|Ornithinuria
C1113952|T201|MTH_LN|30049-1|LNC2HPO|Ornithinuria|Ornithinuria
C1113952|T201|OSN|30049-1|LNC2HPO|Ornithinuria|Ornithinuria
C1113952|T201|LC|30049-1|LNC2HPO|Ornithinuria|Ornithinuria
C1114857|T201|LN|30051-7|LNC2HPO|Homocystinuria|Homocystinuria
C1114857|T201|OSN|30051-7|LNC2HPO|Homocystinuria|Homocystinuria
C1114857|T201|DN|30051-7|LNC2HPO|Homocystinuria|Homocystinuria
C1114857|T201|MTH_LN|30051-7|LNC2HPO|Homocystinuria|Homocystinuria
C1114857|T201|LC|30051-7|LNC2HPO|Homocystinuria|Homocystinuria
C1114858|T201|LN|30052-5|LNC2HPO|Isoleucinuria|Isoleucinuria
C1114858|T201|DN|30052-5|LNC2HPO|Isoleucinuria|Isoleucinuria
C1114858|T201|MTH_LN|30052-5|LNC2HPO|Isoleucinuria|Isoleucinuria
C1114858|T201|OSN|30052-5|LNC2HPO|Isoleucinuria|Isoleucinuria
C1114858|T201|LC|30052-5|LNC2HPO|Isoleucinuria|Isoleucinuria
C1114858|T201|LN|30052-5|LNC2HPO|Hyperisoleucinuria|Hyperisoleucinuria
C1114858|T201|DN|30052-5|LNC2HPO|Hyperisoleucinuria|Hyperisoleucinuria
C1114858|T201|MTH_LN|30052-5|LNC2HPO|Hyperisoleucinuria|Hyperisoleucinuria
C1114858|T201|OSN|30052-5|LNC2HPO|Hyperisoleucinuria|Hyperisoleucinuria
C1114858|T201|LC|30052-5|LNC2HPO|Hyperisoleucinuria|Hyperisoleucinuria
C1113957|T201|LN|30057-4|LNC2HPO|Hyperthreoninuria|Hyperthreoninuria
C1113957|T201|DN|30057-4|LNC2HPO|Hyperthreoninuria|Hyperthreoninuria
C1113957|T201|MTH_LN|30057-4|LNC2HPO|Hyperthreoninuria|Hyperthreoninuria
C1113957|T201|OSN|30057-4|LNC2HPO|Hyperthreoninuria|Hyperthreoninuria
C1113957|T201|LC|30057-4|LNC2HPO|Hyperthreoninuria|Hyperthreoninuria
C1113959|T201|LN|30059-0|LNC2HPO|Glutaric aciduria|Glutaric aciduria
C1113959|T201|DN|30059-0|LNC2HPO|Glutaric aciduria|Glutaric aciduria
C1113959|T201|MTH_LN|30059-0|LNC2HPO|Glutaric aciduria|Glutaric aciduria
C1113959|T201|OSN|30059-0|LNC2HPO|Glutaric aciduria|Glutaric aciduria
C1113959|T201|LC|30059-0|LNC2HPO|Glutaric aciduria|Glutaric aciduria
C1113959|T201|LN|30059-0|LNC2HPO|Glutarate aciduria|Glutarate aciduria
C1113959|T201|DN|30059-0|LNC2HPO|Glutarate aciduria|Glutarate aciduria
C1113959|T201|MTH_LN|30059-0|LNC2HPO|Glutarate aciduria|Glutarate aciduria
C1113959|T201|OSN|30059-0|LNC2HPO|Glutarate aciduria|Glutarate aciduria
C1113959|T201|LC|30059-0|LNC2HPO|Glutarate aciduria|Glutarate aciduria
C1113959|T201|LN|30059-0|LNC2HPO|Glutaricaciduria|Glutaricaciduria
C1113959|T201|DN|30059-0|LNC2HPO|Glutaricaciduria|Glutaricaciduria
C1113959|T201|MTH_LN|30059-0|LNC2HPO|Glutaricaciduria|Glutaricaciduria
C1113959|T201|OSN|30059-0|LNC2HPO|Glutaricaciduria|Glutaricaciduria
C1113959|T201|LC|30059-0|LNC2HPO|Glutaricaciduria|Glutaricaciduria
C1113965|T201|LN|30065-7|LNC2HPO|Cystinuria|Cystinuria
C1113965|T201|DN|30065-7|LNC2HPO|Cystinuria|Cystinuria
C1113965|T201|MTH_LN|30065-7|LNC2HPO|Cystinuria|Cystinuria
C1113965|T201|OSN|30065-7|LNC2HPO|Cystinuria|Cystinuria
C1113965|T201|LC|30065-7|LNC2HPO|Cystinuria|Cystinuria
C1113966|T201|LN|30066-5|LNC2HPO|Glycinuria|Glycinuria
C1113966|T201|DN|30066-5|LNC2HPO|Glycinuria|Glycinuria
C1113966|T201|MTH_LN|30066-5|LNC2HPO|Glycinuria|Glycinuria
C1113966|T201|OSN|30066-5|LNC2HPO|Glycinuria|Glycinuria
C1113966|T201|LC|30066-5|LNC2HPO|Glycinuria|Glycinuria
C1113966|T201|LN|30066-5|LNC2HPO|Hyperglycinuria|Hyperglycinuria
C1113966|T201|DN|30066-5|LNC2HPO|Hyperglycinuria|Hyperglycinuria
C1113966|T201|MTH_LN|30066-5|LNC2HPO|Hyperglycinuria|Hyperglycinuria
C1113966|T201|OSN|30066-5|LNC2HPO|Hyperglycinuria|Hyperglycinuria
C1113966|T201|LC|30066-5|LNC2HPO|Hyperglycinuria|Hyperglycinuria
C1113967|T201|LN|30067-3|LNC2HPO|Prolinuria|Prolinuria
C1113967|T201|DN|30067-3|LNC2HPO|Prolinuria|Prolinuria
C1113967|T201|MTH_LN|30067-3|LNC2HPO|Prolinuria|Prolinuria
C1113967|T201|OSN|30067-3|LNC2HPO|Prolinuria|Prolinuria
C1113967|T201|LC|30067-3|LNC2HPO|Prolinuria|Prolinuria
C1114387|T201|LN|30552-4|LNC2HPO|Vitamin B6 deficiency|Vitamin B6 deficiency
C1114387|T201|DN|30552-4|LNC2HPO|Vitamin B6 deficiency|Vitamin B6 deficiency
C1114387|T201|MTH_LN|30552-4|LNC2HPO|Vitamin B6 deficiency|Vitamin B6 deficiency
C1114387|T201|OSN|30552-4|LNC2HPO|Vitamin B6 deficiency|Vitamin B6 deficiency
C1114387|T201|LC|30552-4|LNC2HPO|Vitamin B6 deficiency|Vitamin B6 deficiency
C0365213|T201|LN|3069-2|LNC2HPO|Hypertryptophanemia|Hypertryptophanemia
C0365213|T201|MTH_LN|3069-2|LNC2HPO|Hypertryptophanemia|Hypertryptophanemia
C0365213|T201|DN|3069-2|LNC2HPO|Hypertryptophanemia|Hypertryptophanemia
C0365213|T201|OSN|3069-2|LNC2HPO|Hypertryptophanemia|Hypertryptophanemia
C0365213|T201|LC|3069-2|LNC2HPO|Hypertryptophanemia|Hypertryptophanemia
C0365213|T201|LN|3069-2|LNC2HPO|Hypotryptophanemia|Hypotryptophanemia
C0365213|T201|MTH_LN|3069-2|LNC2HPO|Hypotryptophanemia|Hypotryptophanemia
C0365213|T201|DN|3069-2|LNC2HPO|Hypotryptophanemia|Hypotryptophanemia
C0365213|T201|OSN|3069-2|LNC2HPO|Hypotryptophanemia|Hypotryptophanemia
C0365213|T201|LC|3069-2|LNC2HPO|Hypotryptophanemia|Hypotryptophanemia
C0365223|T201|LN|3079-1|LNC2HPO|Hypertyrosinemia|Hypertyrosinemia
C0365223|T201|MTH_LN|3079-1|LNC2HPO|Hypertyrosinemia|Hypertyrosinemia
C0365223|T201|DN|3079-1|LNC2HPO|Hypertyrosinemia|Hypertyrosinemia
C0365223|T201|OSN|3079-1|LNC2HPO|Hypertyrosinemia|Hypertyrosinemia
C0365223|T201|LC|3079-1|LNC2HPO|Hypertyrosinemia|Hypertyrosinemia
C0365223|T201|LN|3079-1|LNC2HPO|Tyrosinemia|Tyrosinemia
C0365223|T201|MTH_LN|3079-1|LNC2HPO|Tyrosinemia|Tyrosinemia
C0365223|T201|DN|3079-1|LNC2HPO|Tyrosinemia|Tyrosinemia
C0365223|T201|OSN|3079-1|LNC2HPO|Tyrosinemia|Tyrosinemia
C0365223|T201|LC|3079-1|LNC2HPO|Tyrosinemia|Tyrosinemia
C0365223|T201|LN|3079-1|LNC2HPO|Hypotyrosinemia|Hypotyrosinemia
C0365223|T201|MTH_LN|3079-1|LNC2HPO|Hypotyrosinemia|Hypotyrosinemia
C0365223|T201|DN|3079-1|LNC2HPO|Hypotyrosinemia|Hypotyrosinemia
C0365223|T201|OSN|3079-1|LNC2HPO|Hypotyrosinemia|Hypotyrosinemia
C0365223|T201|LC|3079-1|LNC2HPO|Hypotyrosinemia|Hypotyrosinemia
C0482633|T201|MTH_LN|3209-4|LNC2HPO|Factor VIII deficiency|Factor VIII deficiency
C0482633|T201|DN|3209-4|LNC2HPO|Factor VIII deficiency|Factor VIII deficiency
C0482633|T201|LN|3209-4|LNC2HPO|Factor VIII deficiency|Factor VIII deficiency
C0482633|T201|OSN|3209-4|LNC2HPO|Factor VIII deficiency|Factor VIII deficiency
C0482633|T201|LC|3209-4|LNC2HPO|Factor VIII deficiency|Factor VIII deficiency
C1315089|T201|LN|32615-7|LNC2HPO|Hyperhomocystinemia|Hyperhomocystinemia
C1315089|T201|DN|32615-7|LNC2HPO|Hyperhomocystinemia|Hyperhomocystinemia
C1315089|T201|MTH_LN|32615-7|LNC2HPO|Hyperhomocystinemia|Hyperhomocystinemia
C1315089|T201|OSN|32615-7|LNC2HPO|Hyperhomocystinemia|Hyperhomocystinemia
C1315089|T201|LC|32615-7|LNC2HPO|Hyperhomocystinemia|Hyperhomocystinemia
C1315089|T201|LN|32615-7|LNC2HPO|Homocystinemia|Homocystinemia
C1315089|T201|DN|32615-7|LNC2HPO|Homocystinemia|Homocystinemia
C1315089|T201|MTH_LN|32615-7|LNC2HPO|Homocystinemia|Homocystinemia
C1315089|T201|OSN|32615-7|LNC2HPO|Homocystinemia|Homocystinemia
C1315089|T201|LC|32615-7|LNC2HPO|Homocystinemia|Homocystinemia
C1315156|T201|LN|32682-7|LNC2HPO|Persistence of hemoglobin F|Persistence of hemoglobin F
C1315156|T201|DN|32682-7|LNC2HPO|Persistence of hemoglobin F|Persistence of hemoglobin F
C1315156|T201|MTH_LN|32682-7|LNC2HPO|Persistence of hemoglobin F|Persistence of hemoglobin F
C1315156|T201|LC|32682-7|LNC2HPO|Persistence of hemoglobin F|Persistence of hemoglobin F
C1315156|T201|OSN|32682-7|LNC2HPO|Persistence of hemoglobin F|Persistence of hemoglobin F
C1315156|T201|LN|32682-7|LNC2HPO|Persistence of HbF|Persistence of HbF
C1315156|T201|DN|32682-7|LNC2HPO|Persistence of HbF|Persistence of HbF
C1315156|T201|MTH_LN|32682-7|LNC2HPO|Persistence of HbF|Persistence of HbF
C1315156|T201|LC|32682-7|LNC2HPO|Persistence of HbF|Persistence of HbF
C1315156|T201|OSN|32682-7|LNC2HPO|Persistence of HbF|Persistence of HbF
C1316828|T201|LN|34366-5|LNC2HPO|Proteinuria|Proteinuria
C1316828|T201|DN|34366-5|LNC2HPO|Proteinuria|Proteinuria
C1316828|T201|LC|34366-5|LNC2HPO|Proteinuria|Proteinuria
C1316828|T201|OSN|34366-5|LNC2HPO|Proteinuria|Proteinuria
C1316828|T201|MTH_LN|34366-5|LNC2HPO|Proteinuria|Proteinuria
C1507814|T201|LN|35663-4|LNC2HPO|Proteinuria|Proteinuria
C1507814|T201|LC|35663-4|LNC2HPO|Proteinuria|Proteinuria
C1507814|T201|DN|35663-4|LNC2HPO|Proteinuria|Proteinuria
C1507814|T201|MTH_LN|35663-4|LNC2HPO|Proteinuria|Proteinuria
C1507814|T201|OSN|35663-4|LNC2HPO|Proteinuria|Proteinuria
C1641515|T201|LN|41647-9|LNC2HPO|Hypercapnia|Hypercapnia
C1641515|T201|DN|41647-9|LNC2HPO|Hypercapnia|Hypercapnia
C1641515|T201|MTH_LN|41647-9|LNC2HPO|Hypercapnia|Hypercapnia
C1641515|T201|OSN|41647-9|LNC2HPO|Hypercapnia|Hypercapnia
C1641515|T201|LC|41647-9|LNC2HPO|Hypercapnia|Hypercapnia
C1641515|T201|LN|41647-9|LNC2HPO|Hypercarbia|Hypercarbia
C1641515|T201|DN|41647-9|LNC2HPO|Hypercarbia|Hypercarbia
C1641515|T201|MTH_LN|41647-9|LNC2HPO|Hypercarbia|Hypercarbia
C1641515|T201|OSN|41647-9|LNC2HPO|Hypercarbia|Hypercarbia
C1641515|T201|LC|41647-9|LNC2HPO|Hypercarbia|Hypercarbia
C1641515|T201|LN|41647-9|LNC2HPO|Hypocapnia|Hypocapnia
C1641515|T201|DN|41647-9|LNC2HPO|Hypocapnia|Hypocapnia
C1641515|T201|MTH_LN|41647-9|LNC2HPO|Hypocapnia|Hypocapnia
C1641515|T201|OSN|41647-9|LNC2HPO|Hypocapnia|Hypocapnia
C1641515|T201|LC|41647-9|LNC2HPO|Hypocapnia|Hypocapnia
C1641515|T201|LN|41647-9|LNC2HPO|Hypocarbia|Hypocarbia
C1641515|T201|DN|41647-9|LNC2HPO|Hypocarbia|Hypocarbia
C1641515|T201|MTH_LN|41647-9|LNC2HPO|Hypocarbia|Hypocarbia
C1641515|T201|OSN|41647-9|LNC2HPO|Hypocarbia|Hypocarbia
C1641515|T201|LC|41647-9|LNC2HPO|Hypocarbia|Hypocarbia
C1717305|T201|LN|44050-3|LNC2HPO|Glucosephosphate isomerase deficiency|Glucosephosphate isomerase deficiency
C1717305|T201|DN|44050-3|LNC2HPO|Glucosephosphate isomerase deficiency|Glucosephosphate isomerase deficiency
C1717305|T201|OSN|44050-3|LNC2HPO|Glucosephosphate isomerase deficiency|Glucosephosphate isomerase deficiency
C1717305|T201|MTH_LN|44050-3|LNC2HPO|Glucosephosphate isomerase deficiency|Glucosephosphate isomerase deficiency
C1717305|T201|LC|44050-3|LNC2HPO|Glucosephosphate isomerase deficiency|Glucosephosphate isomerase deficiency
C1717305|T201|LN|44050-3|LNC2HPO|Phosphohexose isomerase deficiency|Phosphohexose isomerase deficiency
C1717305|T201|DN|44050-3|LNC2HPO|Phosphohexose isomerase deficiency|Phosphohexose isomerase deficiency
C1717305|T201|OSN|44050-3|LNC2HPO|Phosphohexose isomerase deficiency|Phosphohexose isomerase deficiency
C1717305|T201|MTH_LN|44050-3|LNC2HPO|Phosphohexose isomerase deficiency|Phosphohexose isomerase deficiency
C1717305|T201|LC|44050-3|LNC2HPO|Phosphohexose isomerase deficiency|Phosphohexose isomerase deficiency
C1978568|T201|LN|50609-7|LNC2HPO|Impaired neutrophil bactericidal activity|Impaired neutrophil bactericidal activity
C1978568|T201|DN|50609-7|LNC2HPO|Impaired neutrophil bactericidal activity|Impaired neutrophil bactericidal activity
C1978568|T201|OSN|50609-7|LNC2HPO|Impaired neutrophil bactericidal activity|Impaired neutrophil bactericidal activity
C1978568|T201|MTH_LN|50609-7|LNC2HPO|Impaired neutrophil bactericidal activity|Impaired neutrophil bactericidal activity
C1978568|T201|LC|50609-7|LNC2HPO|Impaired neutrophil bactericidal activity|Impaired neutrophil bactericidal activity
C1978568|T201|LN|50609-7|LNC2HPO|Impaired oxidative burst|Impaired oxidative burst
C1978568|T201|DN|50609-7|LNC2HPO|Impaired oxidative burst|Impaired oxidative burst
C1978568|T201|OSN|50609-7|LNC2HPO|Impaired oxidative burst|Impaired oxidative burst
C1978568|T201|MTH_LN|50609-7|LNC2HPO|Impaired oxidative burst|Impaired oxidative burst
C1978568|T201|LC|50609-7|LNC2HPO|Impaired oxidative burst|Impaired oxidative burst
C2360416|T201|LN|51733-4|LNC2HPO|Hyperoxemia|Hyperoxemia
C2360416|T201|MTH_LN|51733-4|LNC2HPO|Hyperoxemia|Hyperoxemia
C2360416|T201|DN|51733-4|LNC2HPO|Hyperoxemia|Hyperoxemia
C2360416|T201|LC|51733-4|LNC2HPO|Hyperoxemia|Hyperoxemia
C2360416|T201|OSN|51733-4|LNC2HPO|Hyperoxemia|Hyperoxemia
C2360416|T201|LN|51733-4|LNC2HPO|Hypoxemia|Hypoxemia
C2360416|T201|MTH_LN|51733-4|LNC2HPO|Hypoxemia|Hypoxemia
C2360416|T201|DN|51733-4|LNC2HPO|Hypoxemia|Hypoxemia
C2360416|T201|LC|51733-4|LNC2HPO|Hypoxemia|Hypoxemia
C2360416|T201|OSN|51733-4|LNC2HPO|Hypoxemia|Hypoxemia
C0367788|T201|LN|5631-7|LNC2HPO|Hypercupremia|Hypercupremia
C0367788|T201|MTH_LN|5631-7|LNC2HPO|Hypercupremia|Hypercupremia
C0367788|T201|DN|5631-7|LNC2HPO|Hypercupremia|Hypercupremia
C0367788|T201|OSN|5631-7|LNC2HPO|Hypercupremia|Hypercupremia
C0367788|T201|LC|5631-7|LNC2HPO|Hypercupremia|Hypercupremia
C0367788|T201|LN|5631-7|LNC2HPO|Hypocupremia|Hypocupremia
C0367788|T201|MTH_LN|5631-7|LNC2HPO|Hypocupremia|Hypocupremia
C0367788|T201|DN|5631-7|LNC2HPO|Hypocupremia|Hypocupremia
C0367788|T201|OSN|5631-7|LNC2HPO|Hypocupremia|Hypocupremia
C0367788|T201|LC|5631-7|LNC2HPO|Hypocupremia|Hypocupremia
C0367788|T201|LN|5631-7|LNC2HPO|Copper deficiency|Copper deficiency
C0367788|T201|MTH_LN|5631-7|LNC2HPO|Copper deficiency|Copper deficiency
C0367788|T201|DN|5631-7|LNC2HPO|Copper deficiency|Copper deficiency
C0367788|T201|OSN|5631-7|LNC2HPO|Copper deficiency|Copper deficiency
C0367788|T201|LC|5631-7|LNC2HPO|Copper deficiency|Copper deficiency
C0367869|T201|LN|5683-8|LNC2HPO|Hypermagnesemia|Hypermagnesemia
C0367869|T201|MTH_LN|5683-8|LNC2HPO|Hypermagnesemia|Hypermagnesemia
C0367869|T201|DN|5683-8|LNC2HPO|Hypermagnesemia|Hypermagnesemia
C0367869|T201|OSN|5683-8|LNC2HPO|Hypermagnesemia|Hypermagnesemia
C0367869|T201|LC|5683-8|LNC2HPO|Hypermagnesemia|Hypermagnesemia
C0367869|T201|LN|5683-8|LNC2HPO|Hypomagnesemia|Hypomagnesemia
C0367869|T201|MTH_LN|5683-8|LNC2HPO|Hypomagnesemia|Hypomagnesemia
C0367869|T201|DN|5683-8|LNC2HPO|Hypomagnesemia|Hypomagnesemia
C0367869|T201|OSN|5683-8|LNC2HPO|Hypomagnesemia|Hypomagnesemia
C0367869|T201|LC|5683-8|LNC2HPO|Hypomagnesemia|Hypomagnesemia
C2923385|T201|LN|59069-5|LNC2HPO|Antinuclear antibodies|Antinuclear antibodies
C2923385|T201|MTH_LN|59069-5|LNC2HPO|Antinuclear antibodies|Antinuclear antibodies
C2923385|T201|DN|59069-5|LNC2HPO|Antinuclear antibodies|Antinuclear antibodies
C2923385|T201|LC|59069-5|LNC2HPO|Antinuclear antibodies|Antinuclear antibodies
C2923385|T201|OSN|59069-5|LNC2HPO|Antinuclear antibodies|Antinuclear antibodies
C2923385|T201|LN|59069-5|LNC2HPO|Antinuclear antibody positive|Antinuclear antibody positive
C2923385|T201|MTH_LN|59069-5|LNC2HPO|Antinuclear antibody positive|Antinuclear antibody positive
C2923385|T201|DN|59069-5|LNC2HPO|Antinuclear antibody positive|Antinuclear antibody positive
C2923385|T201|LC|59069-5|LNC2HPO|Antinuclear antibody positive|Antinuclear antibody positive
C2923385|T201|OSN|59069-5|LNC2HPO|Antinuclear antibody positive|Antinuclear antibody positive
C2923385|T201|LN|59069-5|LNC2HPO|Serum antinuclear antibody|Serum antinuclear antibody
C2923385|T201|MTH_LN|59069-5|LNC2HPO|Serum antinuclear antibody|Serum antinuclear antibody
C2923385|T201|DN|59069-5|LNC2HPO|Serum antinuclear antibody|Serum antinuclear antibody
C2923385|T201|LC|59069-5|LNC2HPO|Serum antinuclear antibody|Serum antinuclear antibody
C2923385|T201|OSN|59069-5|LNC2HPO|Serum antinuclear antibody|Serum antinuclear antibody
C2923805|T201|LN|59408-5|LNC2HPO|Hyperoxemia|Hyperoxemia
C2923805|T201|LC|59408-5|LNC2HPO|Hyperoxemia|Hyperoxemia
C2923805|T201|MTH_LN|59408-5|LNC2HPO|Hyperoxemia|Hyperoxemia
C2923805|T201|OSN|59408-5|LNC2HPO|Hyperoxemia|Hyperoxemia
C2923805|T201|LN|59408-5|LNC2HPO|Hypoxemia|Hypoxemia
C2923805|T201|LC|59408-5|LNC2HPO|Hypoxemia|Hypoxemia
C2923805|T201|MTH_LN|59408-5|LNC2HPO|Hypoxemia|Hypoxemia
C2923805|T201|OSN|59408-5|LNC2HPO|Hypoxemia|Hypoxemia
C0482677|T201|MTH_LN|5946-9|LNC2HPO|Haemorrhagic disorders|Haemorrhagic disorders
C0482677|T201|LC|5946-9|LNC2HPO|Haemorrhagic disorders|Haemorrhagic disorders
C0482677|T201|DN|5946-9|LNC2HPO|Haemorrhagic disorders|Haemorrhagic disorders
C0482677|T201|LN|5946-9|LNC2HPO|Haemorrhagic disorders|Haemorrhagic disorders
C0482677|T201|OSN|5946-9|LNC2HPO|Haemorrhagic disorders|Haemorrhagic disorders
C0482677|T201|MTH_LN|5946-9|LNC2HPO|Prolonged PTT|Prolonged PTT
C0482677|T201|LC|5946-9|LNC2HPO|Prolonged PTT|Prolonged PTT
C0482677|T201|DN|5946-9|LNC2HPO|Prolonged PTT|Prolonged PTT
C0482677|T201|LN|5946-9|LNC2HPO|Prolonged PTT|Prolonged PTT
C0482677|T201|OSN|5946-9|LNC2HPO|Prolonged PTT|Prolonged PTT
C0482677|T201|MTH_LN|5946-9|LNC2HPO|Prolonged partial thromboplastin time|Prolonged partial thromboplastin time
C0482677|T201|LC|5946-9|LNC2HPO|Prolonged partial thromboplastin time|Prolonged partial thromboplastin time
C0482677|T201|DN|5946-9|LNC2HPO|Prolonged partial thromboplastin time|Prolonged partial thromboplastin time
C0482677|T201|LN|5946-9|LNC2HPO|Prolonged partial thromboplastin time|Prolonged partial thromboplastin time
C0482677|T201|OSN|5946-9|LNC2HPO|Prolonged partial thromboplastin time|Prolonged partial thromboplastin time
C0482677|T201|MTH_LN|5946-9|LNC2HPO|Partial thromboplastin time prolonged|Partial thromboplastin time prolonged
C0482677|T201|LC|5946-9|LNC2HPO|Partial thromboplastin time prolonged|Partial thromboplastin time prolonged
C0482677|T201|DN|5946-9|LNC2HPO|Partial thromboplastin time prolonged|Partial thromboplastin time prolonged
C0482677|T201|LN|5946-9|LNC2HPO|Partial thromboplastin time prolonged|Partial thromboplastin time prolonged
C0482677|T201|OSN|5946-9|LNC2HPO|Partial thromboplastin time prolonged|Partial thromboplastin time prolonged
C0482677|T201|MTH_LN|5946-9|LNC2HPO|Delayed thromboplastin generation|Delayed thromboplastin generation
C0482677|T201|LC|5946-9|LNC2HPO|Delayed thromboplastin generation|Delayed thromboplastin generation
C0482677|T201|DN|5946-9|LNC2HPO|Delayed thromboplastin generation|Delayed thromboplastin generation
C0482677|T201|LN|5946-9|LNC2HPO|Delayed thromboplastin generation|Delayed thromboplastin generation
C0482677|T201|OSN|5946-9|LNC2HPO|Delayed thromboplastin generation|Delayed thromboplastin generation
C0482677|T201|MTH_LN|5946-9|LNC2HPO|Prolonged activated partial thromboplastin time|Prolonged activated partial thromboplastin time
C0482677|T201|LC|5946-9|LNC2HPO|Prolonged activated partial thromboplastin time|Prolonged activated partial thromboplastin time
C0482677|T201|DN|5946-9|LNC2HPO|Prolonged activated partial thromboplastin time|Prolonged activated partial thromboplastin time
C0482677|T201|LN|5946-9|LNC2HPO|Prolonged activated partial thromboplastin time|Prolonged activated partial thromboplastin time
C0482677|T201|OSN|5946-9|LNC2HPO|Prolonged activated partial thromboplastin time|Prolonged activated partial thromboplastin time
C0484692|T201|LN|6687-8|LNC2HPO|Hypercitraturia|Hypercitraturia
C0484692|T201|MTH_LN|6687-8|LNC2HPO|Hypercitraturia|Hypercitraturia
C0484692|T201|DN|6687-8|LNC2HPO|Hypercitraturia|Hypercitraturia
C0484692|T201|OSN|6687-8|LNC2HPO|Hypercitraturia|Hypercitraturia
C0484692|T201|LC|6687-8|LNC2HPO|Hypercitraturia|Hypercitraturia
C0484692|T201|LN|6687-8|LNC2HPO|Hypocitraturia|Hypocitraturia
C0484692|T201|MTH_LN|6687-8|LNC2HPO|Hypocitraturia|Hypocitraturia
C0484692|T201|DN|6687-8|LNC2HPO|Hypocitraturia|Hypocitraturia
C0484692|T201|OSN|6687-8|LNC2HPO|Hypocitraturia|Hypocitraturia
C0484692|T201|LC|6687-8|LNC2HPO|Hypocitraturia|Hypocitraturia
C3654405|T201|LN|73572-0|LNC2HPO|Hypermagnesemia|Hypermagnesemia
C3654405|T201|LC|73572-0|LNC2HPO|Hypermagnesemia|Hypermagnesemia
C3654405|T201|MTH_LN|73572-0|LNC2HPO|Hypermagnesemia|Hypermagnesemia
C3654405|T201|OSN|73572-0|LNC2HPO|Hypermagnesemia|Hypermagnesemia
C3654405|T201|DN|73572-0|LNC2HPO|Hypermagnesemia|Hypermagnesemia
C3654405|T201|LN|73572-0|LNC2HPO|Hypomagnesemia|Hypomagnesemia
C3654405|T201|LC|73572-0|LNC2HPO|Hypomagnesemia|Hypomagnesemia
C3654405|T201|MTH_LN|73572-0|LNC2HPO|Hypomagnesemia|Hypomagnesemia
C3654405|T201|OSN|73572-0|LNC2HPO|Hypomagnesemia|Hypomagnesemia
C3654405|T201|DN|73572-0|LNC2HPO|Hypomagnesemia|Hypomagnesemia
C0484521|T201|LN|8101-8|LNC2HPO|CD8+ T-cell lymphopenia|CD8+ T-cell lymphopenia
C0484521|T201|LC|8101-8|LNC2HPO|CD8+ T-cell lymphopenia|CD8+ T-cell lymphopenia
C0484521|T201|DN|8101-8|LNC2HPO|CD8+ T-cell lymphopenia|CD8+ T-cell lymphopenia
C0484521|T201|MTH_LN|8101-8|LNC2HPO|CD8+ T-cell lymphopenia|CD8+ T-cell lymphopenia
C0484521|T201|OSN|8101-8|LNC2HPO|CD8+ T-cell lymphopenia|CD8+ T-cell lymphopenia
C0484548|T201|LN|8123-2|LNC2HPO|CD4+ T-cell lymphopenia|CD4+ T-cell lymphopenia
C0484548|T201|LC|8123-2|LNC2HPO|CD4+ T-cell lymphopenia|CD4+ T-cell lymphopenia
C0484548|T201|DN|8123-2|LNC2HPO|CD4+ T-cell lymphopenia|CD4+ T-cell lymphopenia
C0484548|T201|MTH_LN|8123-2|LNC2HPO|CD4+ T-cell lymphopenia|CD4+ T-cell lymphopenia
C0484548|T201|OSN|8123-2|LNC2HPO|CD4+ T-cell lymphopenia|CD4+ T-cell lymphopenia
C0484548|T201|LN|8123-2|LNC2HPO|CD4 T cell lymphopenia|CD4 T cell lymphopenia
C0484548|T201|LC|8123-2|LNC2HPO|CD4 T cell lymphopenia|CD4 T cell lymphopenia
C0484548|T201|DN|8123-2|LNC2HPO|CD4 T cell lymphopenia|CD4 T cell lymphopenia
C0484548|T201|MTH_LN|8123-2|LNC2HPO|CD4 T cell lymphopenia|CD4 T cell lymphopenia
C0484548|T201|OSN|8123-2|LNC2HPO|CD4 T cell lymphopenia|CD4 T cell lymphopenia
C0488794|T201|LC|8867-4|LNC2HPO|Cardiac arrhythmia|Cardiac arrhythmia
C0488794|T201|OSN|8867-4|LNC2HPO|Cardiac arrhythmia|Cardiac arrhythmia
C0488794|T201|MTH_LN|8867-4|LNC2HPO|Cardiac arrhythmia|Cardiac arrhythmia
C0488794|T201|LN|8867-4|LNC2HPO|Cardiac arrhythmia|Cardiac arrhythmia
C0488794|T201|LC|8867-4|LNC2HPO|Cardiac arrhythmias|Cardiac arrhythmias
C0488794|T201|OSN|8867-4|LNC2HPO|Cardiac arrhythmias|Cardiac arrhythmias
C0488794|T201|MTH_LN|8867-4|LNC2HPO|Cardiac arrhythmias|Cardiac arrhythmias
C0488794|T201|LN|8867-4|LNC2HPO|Cardiac arrhythmias|Cardiac arrhythmias
C0488794|T201|LC|8867-4|LNC2HPO|Arrhythmia|Arrhythmia
C0488794|T201|OSN|8867-4|LNC2HPO|Arrhythmia|Arrhythmia
C0488794|T201|MTH_LN|8867-4|LNC2HPO|Arrhythmia|Arrhythmia
C0488794|T201|LN|8867-4|LNC2HPO|Arrhythmia|Arrhythmia
C0488794|T201|LC|8867-4|LNC2HPO|Arrhythmias|Arrhythmias
C0488794|T201|OSN|8867-4|LNC2HPO|Arrhythmias|Arrhythmias
C0488794|T201|MTH_LN|8867-4|LNC2HPO|Arrhythmias|Arrhythmias
C0488794|T201|LN|8867-4|LNC2HPO|Arrhythmias|Arrhythmias
C0488794|T201|LC|8867-4|LNC2HPO|Irregular heart beat|Irregular heart beat
C0488794|T201|OSN|8867-4|LNC2HPO|Irregular heart beat|Irregular heart beat
C0488794|T201|MTH_LN|8867-4|LNC2HPO|Irregular heart beat|Irregular heart beat
C0488794|T201|LN|8867-4|LNC2HPO|Irregular heart beat|Irregular heart beat
C0488794|T201|LC|8867-4|LNC2HPO|Heart rhythm disorders|Heart rhythm disorders
C0488794|T201|OSN|8867-4|LNC2HPO|Heart rhythm disorders|Heart rhythm disorders
C0488794|T201|MTH_LN|8867-4|LNC2HPO|Heart rhythm disorders|Heart rhythm disorders
C0488794|T201|LN|8867-4|LNC2HPO|Heart rhythm disorders|Heart rhythm disorders
C0488794|T201|LC|8867-4|LNC2HPO|Cardiac rhythm disturbances|Cardiac rhythm disturbances
C0488794|T201|OSN|8867-4|LNC2HPO|Cardiac rhythm disturbances|Cardiac rhythm disturbances
C0488794|T201|MTH_LN|8867-4|LNC2HPO|Cardiac rhythm disturbances|Cardiac rhythm disturbances
C0488794|T201|LN|8867-4|LNC2HPO|Cardiac rhythm disturbances|Cardiac rhythm disturbances
C0488794|T201|LC|8867-4|LNC2HPO|Irregular heartbeat|Irregular heartbeat
C0488794|T201|OSN|8867-4|LNC2HPO|Irregular heartbeat|Irregular heartbeat
C0488794|T201|MTH_LN|8867-4|LNC2HPO|Irregular heartbeat|Irregular heartbeat
C0488794|T201|LN|8867-4|LNC2HPO|Irregular heartbeat|Irregular heartbeat
C0488794|T201|LC|8867-4|LNC2HPO|Cardiac conduction defects|Cardiac conduction defects
C0488794|T201|OSN|8867-4|LNC2HPO|Cardiac conduction defects|Cardiac conduction defects
C0488794|T201|MTH_LN|8867-4|LNC2HPO|Cardiac conduction defects|Cardiac conduction defects
C0488794|T201|LN|8867-4|LNC2HPO|Cardiac conduction defects|Cardiac conduction defects
C0488794|T201|LC|8867-4|LNC2HPO|Tachycardia|Tachycardia
C0488794|T201|OSN|8867-4|LNC2HPO|Tachycardia|Tachycardia
C0488794|T201|MTH_LN|8867-4|LNC2HPO|Tachycardia|Tachycardia
C0488794|T201|LN|8867-4|LNC2HPO|Tachycardia|Tachycardia
C0488794|T201|LC|8867-4|LNC2HPO|Rapid heart beat|Rapid heart beat
C0488794|T201|OSN|8867-4|LNC2HPO|Rapid heart beat|Rapid heart beat
C0488794|T201|MTH_LN|8867-4|LNC2HPO|Rapid heart beat|Rapid heart beat
C0488794|T201|LN|8867-4|LNC2HPO|Rapid heart beat|Rapid heart beat
C0488794|T201|LC|8867-4|LNC2HPO|Fast heart rate|Fast heart rate
C0488794|T201|OSN|8867-4|LNC2HPO|Fast heart rate|Fast heart rate
C0488794|T201|MTH_LN|8867-4|LNC2HPO|Fast heart rate|Fast heart rate
C0488794|T201|LN|8867-4|LNC2HPO|Fast heart rate|Fast heart rate
C0488794|T201|LC|8867-4|LNC2HPO|Heart racing|Heart racing
C0488794|T201|OSN|8867-4|LNC2HPO|Heart racing|Heart racing
C0488794|T201|MTH_LN|8867-4|LNC2HPO|Heart racing|Heart racing
C0488794|T201|LN|8867-4|LNC2HPO|Heart racing|Heart racing
C0488794|T201|LC|8867-4|LNC2HPO|Racing heart|Racing heart
C0488794|T201|OSN|8867-4|LNC2HPO|Racing heart|Racing heart
C0488794|T201|MTH_LN|8867-4|LNC2HPO|Racing heart|Racing heart
C0488794|T201|LN|8867-4|LNC2HPO|Racing heart|Racing heart
C0488794|T201|LC|8867-4|LNC2HPO|Bradycardia|Bradycardia
C0488794|T201|OSN|8867-4|LNC2HPO|Bradycardia|Bradycardia
C0488794|T201|MTH_LN|8867-4|LNC2HPO|Bradycardia|Bradycardia
C0488794|T201|LN|8867-4|LNC2HPO|Bradycardia|Bradycardia
C0488794|T201|LC|8867-4|LNC2HPO|Brachycardia|Brachycardia
C0488794|T201|OSN|8867-4|LNC2HPO|Brachycardia|Brachycardia
C0488794|T201|MTH_LN|8867-4|LNC2HPO|Brachycardia|Brachycardia
C0488794|T201|LN|8867-4|LNC2HPO|Brachycardia|Brachycardia
C0488794|T201|LC|8867-4|LNC2HPO|Slow heartbeats|Slow heartbeats
C0488794|T201|OSN|8867-4|LNC2HPO|Slow heartbeats|Slow heartbeats
C0488794|T201|MTH_LN|8867-4|LNC2HPO|Slow heartbeats|Slow heartbeats
C0488794|T201|LN|8867-4|LNC2HPO|Slow heartbeats|Slow heartbeats
C0943173|T201|LN|27365-6|LNC2HPO|Kappa Bence Jones proteinuria|Kappa Bence Jones proteinuria
C0943173|T201|LC|27365-6|LNC2HPO|Kappa Bence Jones proteinuria|Kappa Bence Jones proteinuria
C0943173|T201|DN|27365-6|LNC2HPO|Kappa Bence Jones proteinuria|Kappa Bence Jones proteinuria
C0943173|T201|MTH_LN|27365-6|LNC2HPO|Kappa Bence Jones proteinuria|Kappa Bence Jones proteinuria
C0943173|T201|OSN|27365-6|LNC2HPO|Kappa Bence Jones proteinuria|Kappa Bence Jones proteinuria
