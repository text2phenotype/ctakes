C0009170|T131|LP16048-8|LNC|COCAINE|COCAINE
C0085163|T131||LNC|CRACK COCAINE
C2203924|T131||LNC|METHYLPHENIDATE ABUSE
C1456332|T131||LNC|STIMULANT ABUSE
C3509122|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED DISORDER
C2874625|T131||LNC|OTHER STIMULANT ABUSE
C2874626|T131||LNC|OTHER STIMULANT ABUSE, UNCOMPLICATED
C2874631|T131||LNC|OTHER STIMULANT ABUSE WITH INTOXICATION, UNSPECIFIED
C3494717|T131||LNC|CATHA EDULIS ABUSE
C3509117|T131||LNC|STIMULANT ABUSE - UNCOMPLICATED
C3509118|T131||LNC|STIMULANT ABUSE WITH INTOXICATION
C3509119|T131||LNC|STIMULANT ABUSE WITH INTOXICATION - UNCOMPLICATED
C3509120|T131||LNC|STIMULANT ABUSE WITH INTOXICATION DELIRIUM
C3662831|T131||LNC|NONDEPENDENT AMPHETAMINE ABUSE
C4481000|T131||LNC|OTHER STIMULANT ABUSE IN REMISSION
C2874632|T131||LNC|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED MOOD DISORDER
C2874636|T131||LNC|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED
C2874637|T131||LNC|OTHER STIMULANT ABUSE WITH OTHER STIMULANT-INDUCED DISORDER
C2874638|T131||LNC|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED ANXIETY DISORDER
C2874639|T131||LNC|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED SEXUAL DYSFUNCTION
C2874640|T131||LNC|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED SLEEP DISORDER
C2874641|T131||LNC|OTHER STIMULANT ABUSE WITH UNSPECIFIED STIMULANT-INDUCED DISORDER
C3509123|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED ANXIETY DISORDER
C3509124|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED SEXUAL FUNCTION
C3509125|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED SLEEP DISORDER
C3509126|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED MOOD DISORDER
C3509127|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER
C3509128|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS
C3509129|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS
C0553808|T131||LNC|NONDEPENDENT AMPHETAMINE OR OTHER PSYCHOSTIMULANT ABUSE
C2874628|T131||LNC|OTHER STIMULANT ABUSE WITH INTOXICATION, UNCOMPLICATED
C2874629|T131||LNC|OTHER STIMULANT ABUSE WITH INTOXICATION DELIRIUM
C3509121|T131||LNC|STIMULANT ABUSE WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE
C3836657|T131||LNC|NONDEPENDENT INTRAVENOUS AMPHETAMINE ABUSE
C2874634|T131||LNC|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS
C2874635|T131||LNC|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS
C0338682|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE, CONTINUOUS
C0338683|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE, EPISODIC
C0338684|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE IN REMISSION
C2874630|T131||LNC|OTHER STIMULANT ABUSE WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE
C0085163|T131||LNC|COCAINE, CRACK
C0085163|T131||LNC|CRACK COCAINE
C0085163|T131||LNC|FREE BASE COCAINE
C0085163|T131||LNC|CRACK COCAINE [CHEMICAL/INGREDIENT]
C0085163|T131||LNC|CRACK
C0085163|T131||LNC|COCAINE FREEBASE
C0085163|T131||LNC|ROCKS - COCAINE
C0085163|T131||LNC|COCAINE FREEBASE 
C0009169|T131||LNC|COCA
C0009169|T131||LNC|ERYTHROXYLUM COCA LAM.
C0009169|T131||LNC|ERYTHROXYLONS
C0009169|T131||LNC|ERYTHROXYLON
C0009169|T131||LNC|COCA PLANT
C0009169|T131||LNC|COCAINE PLANT
C0009169|T131||LNC|ERYTHROXYLUM COCA
C0009169|T131||LNC|ERYTHROXYLUM COCA 
C0009169|T131||LNC|HAYO
C0975799|T131||LNC|COCAINE HCL PWDR
C0975799|T131||LNC|COCAINE HCL POWDER
C0975799|T131||LNC|COCAINE HCL PWDR [VA PRODUCT]
C0009170|T131|LP16048-8|LNC|COCAINE|COCAINE
C0009170|T131|LP16048-8|LNC|8-AZABICYCLO(3.2.1)OCTANE-2-CARBOXYLIC ACID, 3-(BENZOYLOXY)-8-METHYL-, METHYL ESTER, (1R-(EXO,EXO))-|COCAINE
C0009170|T131|LP16048-8|LNC|(1R,2R,3S,5S)-2-METHOXYCARBONYLTROPAN-3-YL BENZOATE|COCAINE
C0009170|T131|LP16048-8|LNC|COCAINE [CHEMICAL/INGREDIENT]|COCAINE
C0009170|T131|LP16048-8|LNC|COCAINE (SCHEDULE I SUBSTANCE)|COCAINE
C0009170|T131|LP16048-8|LNC|SNOW|COCAINE
C0009170|T131|LP16048-8|LNC|COKE|COCAINE
C0009170|T131|LP16048-8|LNC|COCA|COCAINE
C0009170|T131|LP16048-8|LNC|COCAINE PRODUCT|COCAINE
C0009170|T131|LP16048-8|LNC|COCAINE |COCAINE
C0009170|T131|LP16048-8|LNC|COCAINE |COCAINE
C2315434|T131||LNC|NASAL FORM COCAINE 
C2315434|T131||LNC|NASAL FORM COCAINE
C2316909|T131||LNC|OROPHARYNGEAL FORM COCAINE 
C2316909|T131||LNC|OROPHARYNGEAL FORM COCAINE
C2316959|T131||LNC|ORAL FORM COCAINE
C2316959|T131||LNC|ORAL FORM COCAINE 
C0282108|T131||LNC|COCAINE HYDROCHLORIDE
C0282108|T131||LNC|HYDROCHLORIDE, COCAINE
C0282108|T131||LNC|COCAINE HYDROCHLORIDE 
C0282108|T131||LNC|METHYL 3-BETA-HYDROXY-1-ALPHA-H,5-ALPHA-H-TROPAN-2-BETA-CARBOXYLATE, BENZOATE (ESTER) HCL
C0282108|T131||LNC|COCAINE HYDROCHLORIDE [CHEMICAL/INGREDIENT]
C0282108|T131||LNC|COCAINE HCL
C0282108|T131||LNC|HCL, COCAINE
C0282108|T131||LNC|COCAINE HYDROCHLORIDE 
C0171681|T131||LNC|RTI-82
C0171681|T131||LNC|8-AZABICYCLO(3.2.1)OCTANE-2-CARBOXYLIC ACID, 3-(4-CHLOROPHENYL)-8-METHYL-, 2-(4-AZIDO-3-IODOPHENYL)ETHYL ESTER, (EXO,EXO)-
C0171681|T131||LNC|RTI 82
C0532637|T131||LNC|TRIMETHYLSTANNYL-(2-CARBOMETHOXY-3-(4-PHENYL)TROPANE)
C0532637|T131||LNC|TRIMETHYLSTANNYL-BETA-CT
C0350656|T131||LNC|MORPHINE + COCAINE ELIXIR
C0350656|T131||LNC|MORPHINE + COCAINE ELIXIR 
C0350656|T131||LNC|MORPHINE + COCAINE ELIXIR 
C0359982|T131||LNC|COCAINE HYDROCHLORIDE POWDER
C0359982|T131||LNC|COCAINE HYDROCHLORIDE POWDER BP
C0359982|T131||LNC|COCAINE HYDROCHLORIDE POWDER 
C0359982|T131||LNC|COCAINE HYDROCHLORIDE POWDER BP 
C0359982|T131||LNC|COCAINE HYDROCHLORIDE POWDER BP 
C0359981|T131||LNC|COCAINE POWDER BP 
C0359981|T131||LNC|COCAINE POWDER BP
C0359981|T131||LNC|COCAINE POWDER BP 
C0350555|T131||LNC|COCAINE [NO DRUGS HERE] 
C0350555|T131||LNC|COCAINE [NO DRUGS HERE]
C0350555|T131||LNC|COCAINE [NO DRUGS HERE] 
C1985612|T131|LP44749-7|LNC|COCAINE &#X7C; URINE|COCAINE &#X7C; URINE
C1985611|T131|LP54539-9|LNC|COCAINE &#X7C; UNKNOWN SUBSTANCE|COCAINE &#X7C; UNKNOWN SUBSTANCE
C0082060|T131||LNC|BENZOYLECGONINE ETHYL ESTER
C0082060|T131||LNC|COCA-ETHYLENE
C0082060|T131||LNC|COCAETHYLENE
C0082060|T131||LNC|ETHYLCOCAINE
C0082060|T131||LNC|COCAETHYLENE 
C0053258|T131|LP16047-0|LNC|BENZOYL ECGONINE|BENZOYLECGONINE
C0053258|T131|LP16047-0|LNC|BENZOYLECGONINE|BENZOYLECGONINE
C0053258|T131|LP16047-0|LNC|BENZOYLECGONINE |BENZOYLECGONINE
C1985608|T131|LP48571-1|LNC|COCAINE &#X7C; MECONIUM|COCAINE &#X7C; MECONIUM
C1985609|T131|LP52055-8|LNC|COCAINE &#X7C; SALIVA|COCAINE &#X7C; SALIVA
C1985613|T131|LP48688-3|LNC|COCAINE &#X7C; VITREOUS FLUID|COCAINE &#X7C; VITREOUS FLUID
C0058917|T131||LNC|ECGONINE METHYL ESTER
C0058917|T131||LNC|METHYL ECGONINE
C1985610|T131|LP48467-2|LNC|COCAINE &#X7C; STOOL|COCAINE &#X7C; STOOL
C1985607|T131|LP48647-9|LNC|COCAINE &#X7C; HAIR|COCAINE &#X7C; HAIR
C1985606|T131|LP49060-4|LNC|COCAINE &#X7C; GASTRIC FLUID|COCAINE &#X7C; GASTRIC FLUID
C1455816|T131||LNC|COCAINE METABOLITES
C1455816|T131||LNC|COCAINE METABOLITE
C1455816|T131||LNC|COCAINE METABOLITE 
C1985605|T131|LP44748-9|LNC|COCAINE &#X7C; BLD-SER-PLAS|COCAINE &#X7C; BLD-SER-PLAS
C1985604|T131|LP49617-1|LNC|COCAINE &#X7C; BILE FLUID|COCAINE &#X7C; BILE FLUID
C0565790|T131||LNC|COCAINE - NON-PHARMACEUTICAL
C0565790|T131||LNC|COCAINE - NON-PHARMACEUTICAL 
C0072534|T131||LNC|PSEUDOCOCAINE
C0075888|T131||LNC|8-AZABICYCLO(3.2.1)OCTANE-2-CARBOXYLIC ACID, 3-(BENZOYLOXY)-8-METHYL-, METHYL ESTER, (1R-(EXO,EXO))-, MIXT. WITH 2-(DIMETHYLAMINO)ETHYL 4-(BUTYLAMINO)BENZOATE AND (R)-4-(1-HYDROXY-2-(METHYLAMINO)ETHYL)-1,2-BENZENEDIOL
C0075888|T131||LNC|TAC COMBINATION
C0075888|T131||LNC|TEC SOLUTION
C0621633|T131||LNC|BAKER'S COCKTAIL
C0621633|T131||LNC|ALUMINUM HYDROXIDE - CIMETIDINE - COCAINE - HYDROXYZINE - MORPHINE
C0621633|T131||LNC|ALUMINUM HYDROXIDE, CIMETIDINE, COCAINE, HYDROXYZINE, MORPHINE DRUG COMBINATION
C0621633|T131||LNC|BAKER'S MIXTURE
C0053928|T131||LNC|BONAIN'S LIQUID
C0056054|T131||LNC|COCAINE-DIPICRYLAMINATE
C0056054|T131||LNC|COCAINE - DIPICRYLAMINATE
C0056054|T131||LNC|COCAINE, DIPICRYLAMINATE DRUG COMBINATION
C0757327|T131||LNC|COCAINE BENZOYL THIOESTER
C0770042|T131||LNC|ECGONIDINE
C1827575|T131||LNC|MORPHINE + COCAINE
C1827575|T131||LNC|MORPHINE + COCAINE 
C1827575|T131||LNC|COCAINE + MORPHINE
C0031890|T131||LNC|PICROTOXIN
C0031890|T131||LNC|3,6-METHANO-8H-1,5,7-TRIOXACYCLOPENTA(IJ)CYCLOPROP(A)AZULENE-4,8(3H)-DIONE, HEXAHYDRO-2A-HYDROXY-9-(1-HYDROXY-1-METHYLETHYL)-8B-METHYL-, (1AR-(1AALPHA,2ABETA,3BETA,6BETA,6ABETA,8AS*,8BBETA,9S*))-, COMPD. WITH (1AR-(1AALPHA,2ABETA,3BETA,6BETA,6ABETA,8AS*,8BBETA,9R*))-HEXAHYDRO-2A-HYDROXY-8B-METHYL-9-(1-METHYLETHENYL)-3,6-METHANO-8H-1,5,7-TRIOXACYCLOPENTA(IJ)CYCLOPROP(A)AZULENE-4,8(3H)-DIONE (1:1)
C0031890|T131||LNC|3,6-METHANO-8H-1,5,7-TRIOXACYCLOPENTA(IJ)CYCLOPROP(A)AZULENE-4,8(3H)-DIONE, HEXAHYDRO-2A-HYDROXY-9-(1-HYDROXY-1-METHYLETHYL)-8B-METHYL-, (1AR-(1AALPHA,2ABETA,3BETA,6BETA,6ABETA,8AS*,8BBETA,9S*))-, COMPD. WITH (1AR-(1AALPHA,2ABETA,3BETA,6BETA,6ABETA,8AS*,8
C0031890|T131||LNC|PICROTOXIN [CHEMICAL/INGREDIENT]
C0031890|T131||LNC|PICROTOXIN 
C0031974|T131||LNC|PIPRADROL
C0031974|T131||LNC|PYRIDROL
C0031974|T131||LNC|PIPRADOL
C0031974|T131||LNC|PIPRADROL 
C0014479|T131|LP16128-8|LNC|EPHEDRINE|EPHEDRINE
C0014479|T131|LP16128-8|LNC|[R-(R*,S*)]-ALPHA-[1-(METHYLAMINO)ETHYL]BENZENEMETHANOL|EPHEDRINE
C0014479|T131|LP16128-8|LNC|(-)-EPHEDRINE|EPHEDRINE
C0014479|T131|LP16128-8|LNC|(1R,2S)-2-METHYLAMINO-1-PHENYL-PROPAN-1-OL|EPHEDRINE
C0014479|T131|LP16128-8|LNC|EPHEDRINE ERYTHRO ISOMER|EPHEDRINE
C0014479|T131|LP16128-8|LNC|EPHEDRINE |EPHEDRINE
C0014479|T131|LP16128-8|LNC|EPHEDRINE [CHEMICAL/INGREDIENT]|EPHEDRINE
C0014479|T131|LP16128-8|LNC|ERYTHRO ISOMER OF EPHEDRINE|EPHEDRINE
C0014479|T131|LP16128-8|LNC|ANTIASTHMATICS EPHEDRINE |EPHEDRINE
C0014479|T131|LP16128-8|LNC|ANTIASTHMATICS EPHEDRINE|EPHEDRINE
C0014479|T131|LP16128-8|LNC|EPHEDRINE |EPHEDRINE
C0014479|T131|LP16128-8|LNC|EPHEDRINE |EPHEDRINE
C0018602|T131||LNC|HARMALINE
C0018602|T131||LNC|3H-PYRIDO(3,4-B)INDOLE, 4,9-DIHYDRO-7-METHOXY-1-METHYL-
C0018602|T131||LNC|HARMALINE [CHEMICAL/INGREDIENT]
C0018602|T131||LNC|DIHYDROHARMINE
C0018602|T131||LNC|HARMIDINE
C0018602|T131||LNC|HARMALINE 
C0025611|T131|LP16194-0|LNC|METHAMPHETAMINE|METHAMPHETAMINE
C0025611|T131|LP16194-0|LNC|N METHYLAMPHETAMINE|METHAMPHETAMINE
C0025611|T131|LP16194-0|LNC|BENZENEETHANAMINE, N,ALPHA-DIMETHYL-, (S)-|METHAMPHETAMINE
C0025611|T131|LP16194-0|LNC|METAMFETAMINE|METHAMPHETAMINE
C0025611|T131|LP16194-0|LNC|METHAMPHETAMINE [CHEMICAL/INGREDIENT]|METHAMPHETAMINE
C0025611|T131|LP16194-0|LNC|METHYLAMPHETAMINE|METHAMPHETAMINE
C0025611|T131|LP16194-0|LNC|N-METHYLAMPHETAMINE|METHAMPHETAMINE
# C0025611|T131|LP16194-0|LNC|SPEED|METHAMPHETAMINE
# C0025611|T131|LP16194-0|LNC|GLASS|METHAMPHETAMINE
# C0025611|T131|LP16194-0|LNC|CRYSTAL|METHAMPHETAMINE
# C0025611|T131|LP16194-0|LNC|CHALK|METHAMPHETAMINE
# C0025611|T131|LP16194-0|LNC|METH|METHAMPHETAMINE
C0025611|T131|LP16194-0|LNC|METH USER|METHAMPHETAMINE
C0025611|T131|LP16194-0|LNC|METH ADDICT|METHAMPHETAMINE
C0025611|T131|LP16194-0|LNC|METH ADDICTION|METHAMPHETAMINE
C0025611|T131|LP16194-0|LNC|USES METH|METHAMPHETAMINE
C0025611|T131|LP16194-0|LNC|METHAMPHETAMINE |METHAMPHETAMINE
C0025611|T131|LP16194-0|LNC|METHAMPHETAMINE |METHAMPHETAMINE
C0028089|T131|LP16220-3|LNC|DIETHYLAMIDE, NICOTINIC|NIKETHAMIDE
C0028089|T131|LP16220-3|LNC|NIKETHAMIDE|NIKETHAMIDE
C0028089|T131|LP16220-3|LNC|3-PYRIDINECARBOXAMIDE, N,N-DIETHYL-|NIKETHAMIDE
C0028089|T131|LP16220-3|LNC|NIKETHAMIDE |NIKETHAMIDE
C0028089|T131|LP16220-3|LNC|CORETHAMID|NIKETHAMIDE
C0028089|T131|LP16220-3|LNC|NICOTINIC DIETHYLAMIDE|NIKETHAMIDE
C0028089|T131|LP16220-3|LNC|DOPING DRUG|NIKETHAMIDE
C0028089|T131|LP16220-3|LNC|NICETHAMIDE|NIKETHAMIDE
C0028089|T131|LP16220-3|LNC|NIKETHAMIDE [CHEMICAL/INGREDIENT]|NIKETHAMIDE
C0028089|T131|LP16220-3|LNC|DIETHYLNICOTINAMID|NIKETHAMIDE
C0028089|T131|LP16220-3|LNC|NIKETHAMIDE |NIKETHAMIDE
C0028089|T131|LP16220-3|LNC|NIKETHAMIDE |NIKETHAMIDE
C0031411|T131|LP16247-6|LNC|PHENMETRAZINE|PHENMETRAZINE
C0031411|T131|LP16247-6|LNC|MORPHOLINE, 3-METHYL-2-PHENYL-|PHENMETRAZINE
C0031411|T131|LP16247-6|LNC|FENMETRAZIN|PHENMETRAZINE
C0031411|T131|LP16247-6|LNC|PHENMETRALINE|PHENMETRAZINE
C0031411|T131|LP16247-6|LNC|OXAZIMEDRINE|PHENMETRAZINE
C0031411|T131|LP16247-6|LNC|PHENMETRAZINE [CHEMICAL/INGREDIENT]|PHENMETRAZINE
C0031411|T131|LP16247-6|LNC|DEFENMETRAZIN|PHENMETRAZINE
C0031411|T131|LP16247-6|LNC|PHENMETRAZINE |PHENMETRAZINE
C0031411|T131|LP16247-6|LNC|PHENMETRAZINE |PHENMETRAZINE
C0031447|T131|LP16250-0|LNC|PHENTERMINE|PHENTERMINE
C0031447|T131|LP16250-0|LNC|BENZENEETHANAMINE, ALPHA,ALPHA-DIMETHYL-|PHENTERMINE
C0031447|T131|LP16250-0|LNC|PHENTERMINE [CHEMICAL/INGREDIENT]|PHENTERMINE
C0031447|T131|LP16250-0|LNC|1,1-DIMETHYL-2-PHENYLETHYLAMINE|PHENTERMINE
C0031447|T131|LP16250-0|LNC|2-PHENYL-TERT-BUTYLAMINE|PHENTERMINE
C0031447|T131|LP16250-0|LNC|2-AMINO-2-METHYL-1-PHENYLPROPANE|PHENTERMINE
C0031447|T131|LP16250-0|LNC|PHENYL-TERTIARY-BUTYLAMINE|PHENTERMINE
C0031447|T131|LP16250-0|LNC|PHENTERMINE |PHENTERMINE
C0031447|T131|LP16250-0|LNC|PHENTERMINE |PHENTERMINE
C0012201|T131|LP19505-4|LNC|DIETHYLPROPION|DIETHYLPROPION
C0012201|T131|LP19505-4|LNC|1-PROPANONE, 2-(DIETHYLAMINO)-1-PHENYL-|DIETHYLPROPION
C0012201|T131|LP19505-4|LNC|AMFEPRAMONE|DIETHYLPROPION
C0012201|T131|LP19505-4|LNC|2-DIETHYLAMINOPROPIOPHENONE|DIETHYLPROPION
C0012201|T131|LP19505-4|LNC|DIETHYLPROPION [CHEMICAL/INGREDIENT]|DIETHYLPROPION
C0012201|T131|LP19505-4|LNC|AMFEPRAMON|DIETHYLPROPION
C0012201|T131|LP19505-4|LNC|PHEPRANON|DIETHYLPROPION
C0012201|T131|LP19505-4|LNC|DIETHYLPROPION |DIETHYLPROPION
C0012201|T131|LP19505-4|LNC|DIETHYLPROPION |DIETHYLPROPION
C0282133|T131||LNC|DIETHYLPROPION HYDROCHLORIDE
C0282133|T131||LNC|HYDROCHLORIDE, DIETHYLPROPION
C0282133|T131||LNC|1-PHENYL-2-DIETHYL-AMINO-1-PROPANONE HYDROCHLORIDE
C0282133|T131||LNC|ANOREXICS DIETHYLPROPION HYDROCHLORIDE
C0282133|T131||LNC|DIETHYLPROPION HYDROCHLORIDE 
C0282133|T131||LNC|DIETHYLPROPION HYDROCHLORIDE [CHEMICAL/INGREDIENT]
C0282133|T131||LNC|DIETHYLPROPION HYDROCHLORIDE 
C0282133|T131||LNC|DIETHYLPROPION HYDROCHLORIDE 
C0282133|T131||LNC|AMFEPRAMONE HYDROCHLORIDE
C0282133|T131||LNC|DIETHYLPROPION HYDROCHLORIDE [DUP] 
C0767825|T131||LNC|IRAMPANEL
C0767825|T131||LNC|DIMETHYL-(2-(2-(3-PHENYL-(1,2,4)OXADIAZOL-5-YL)PHENOXY)ETHYL)AMINE HYDROCHLORIDE
C0767825|T131||LNC|5-(O-(2-(DIMETHYLAMINO)ETHOXY)PHENYL)-3-PHENYL-1,2,4-OXADIAZOLE
C1565316|T131||LNC|(S)-N-(2-(1,6,7,8-TETRAHYDRO-2H-INDENO-(5,4)FURAN-8-YL)ETHYL)PROPIONAMIDE
C2699993|T131||LNC|ENDOMIDE
C2698084|T131||LNC|AMFETAMINIL
C0051684|T131||LNC|2,4-DIAMINO-5-PHENYLTHIAZOLE
C0051684|T131||LNC|AMIPHENAZOLE
C0051684|T131||LNC|AMIPHENAZOLE 
C0034295|T131||LNC|PYRITHIOXIN
C0034295|T131||LNC|PYRITINOL 
C0034295|T131||LNC|PYRITINOL
C0034295|T131||LNC|4-PYRIDINEMETHANOL, 3,3'-(DITHIOBIS(METHYLENE))BIS(5-HYDROXY-6-METHYL- )
C0034295|T131||LNC|PYRITHIOXIN [CHEMICAL/INGREDIENT]
C0034295|T131||LNC|PYRITHIOXINE
C0034295|T131||LNC|PIRITINOL
C0034295|T131||LNC|DIPYRIDOXOLYLDISULFIDE
C0034295|T131||LNC|PYRIDOXINEDISULFIDE
C0034295|T131||LNC|PYRITINOL 
C2700197|T131||LNC|FLUBANILATE
C0056852|T131||LNC|CYPRODENATE
C0056852|T131||LNC|DIMETHYLAMINO- 2-ETHYL-BETA-CYCLOHEXYLPROPIONIC ACID MALEATE
C0056852|T131||LNC|CYPRODEMANOL
C0000379|T131|LP19292-9|LNC|MDA|METHYLENEDIOXYAMPHETAMINE
C0000379|T131|LP19292-9|LNC|1,3-BENZODIOXOLE-5-ETHANAMINE, ALPHA-METHYL-|METHYLENEDIOXYAMPHETAMINE
C0000379|T131|LP19292-9|LNC|METHYLENEDIOXYAMPHETAMINE 03 04|METHYLENEDIOXYAMPHETAMINE
C0000379|T131|LP19292-9|LNC|ALPHA-METHYL-1,3-BENZODIOXOLE-5-ETHANAMINE|METHYLENEDIOXYAMPHETAMINE
C0000379|T131|LP19292-9|LNC|TENAMFETAMINE|METHYLENEDIOXYAMPHETAMINE
C0000379|T131|LP19292-9|LNC|METHYLENEDIOXYAMPHETAMINE|METHYLENEDIOXYAMPHETAMINE
C0000379|T131|LP19292-9|LNC|3,4-METHYLENEDIOXYAMPHETAMINE [CHEMICAL/INGREDIENT]|METHYLENEDIOXYAMPHETAMINE
C0000379|T131|LP19292-9|LNC|METHYLENEDIOXYAMPHETAMINE |METHYLENEDIOXYAMPHETAMINE
C2825428|T131||LNC|CYCLAZODONE
C0059791|T131||LNC|ETHYLAMPHETAMINE
C0059791|T131||LNC|ETILAMFETAMINE
C0059791|T131||LNC|N-ETHYLAMPHETAMINE
C0060167|T131||LNC|7-(2-((ALPHA-METHYLPHENETHYL)AMINO)ETHYL)THEOPHYLLINE
C0060167|T131||LNC|7-ETHYLTHEOPHYLLINEAMPHETAMINE
C0060167|T131||LNC|FENETHYLLINE
C0060167|T131||LNC|FENETYLLINE
C0060167|T131||LNC|THEOPHYLLINE ETHYLAMPHETAMINE
C0060167|T131||LNC|FENETHYLLINE 
C2825430|T131||LNC|FENETHYLLINE HYDROCHLORIDE
C0301388|T131||LNC|2-AMINO-1,1-DIPHENYLHEPTAMOL
C0301388|T131||LNC|HEXAPRADOL
C0301388|T131||LNC|ALPHA-(1-AMINOHEXYL)BENZHYDROL
C0301388|T131||LNC|HEXAPRADOL 
C0771352|T131||LNC|1,3,7-TRIMETHYL-3,7-DIHYDRO-1H-PURINE-2,6-DIONE MONOHYDRATE
C0115471|T131|LA28418-4|LNC|MDMA|ECSTASY
C0115471|T131|LA28418-4|LNC|ECSTASY|ECSTASY
C0115471|T131|LA28418-4|LNC|N METHYL 3,4 METHYLENEDIOXYAMPHETAMINE|ECSTASY
C0115471|T131|LA28418-4|LNC|N-METHYL-3,4-METHYLENEDIOXYAMPHETAMINE|ECSTASY
C0115471|T131|LA28418-4|LNC|1,3-BENZODIOXOLE-5-ETHANAMINE, N,ALPHA-DIMETHYL-|ECSTASY
C0115471|T131|LA28418-4|LNC|3,4 METHYLENEDIOXYMETHAMPHETAMINE|ECSTASY
C0115471|T131|LA28418-4|LNC|MMDA|ECSTASY
C0115471|T131|LA28418-4|LNC|3-METHOXY-4,5- METHYLENEDIOXYAMPHETAMINE|ECSTASY
C0115471|T131|LA28418-4|LNC|3,4-METHYLENEDIOXYMETHAMPHETAMINE|ECSTASY
C0115471|T131|LA28418-4|LNC|METHYLMETHYLENEDIOXYAMPHETAMINE N 03 04|ECSTASY
C0115471|T131|LA28418-4|LNC|ECSTASY - DRUG|ECSTASY
C0115471|T131|LA28418-4|LNC|METHYLENE-DIOXYMETHAMPHETAMINE|ECSTASY
C0115471|T131|LA28418-4|LNC|ECSTASY |ECSTASY
C0115471|T131|LA28418-4|LNC|ECSTASY - AGENT|ECSTASY
C0115471|T131|LA28418-4|LNC|N-METHYL-3,4-METHYLENEDIOXYAMPHETAMINE [CHEMICAL/INGREDIENT]|ECSTASY
C0115471|T131|LA28418-4|LNC|METHYLENEDIOXYMETHAMPHETAMINE|ECSTASY
C0115471|T131|LA28418-4|LNC|XTC|ECSTASY
C0115471|T131|LA28418-4|LNC|N-METHYL-3, 4-METHYLENEDIOXYAMPHETAMINE |ECSTASY
C0115471|T131|LA28418-4|LNC|E - ECSTASY|ECSTASY
C0115471|T131|LA28418-4|LNC|N-METHYL-3, 4-METHYLENEDIOXYAMPHETAMINE|ECSTASY
C0115471|T131|LA28418-4|LNC|ECSTASY - AGENT |ECSTASY
C0115471|T131|LA28418-4|LNC|METHYLENE-DIOXYMETHAMPHETAMINE |ECSTASY
C0115471|T131|LA28418-4|LNC|MDM|ECSTASY
C0115471|T131|LA28418-4|LNC|MDMA - METHYLENEDIOXYMETHAMPHETAMINE|ECSTASY
C0115471|T131|LA28418-4|LNC|METHYLENE-DIOXYMETHAMPHETAMINE |ECSTASY
C0115471|T131|LA28418-4|LNC|METHYLENEDIOXYMETHAMPHETAMINE |ECSTASY
C0115471|T131|LA28418-4|LNC|ECSTASY - DRUG |ECSTASY
C0115471|T131|LA28418-4|LNC|METHYLENEDIOXYMETHAMFETAMINE|ECSTASY
C0553808|T131||LNC|NONDEPENDENT AMPHETAMINE OR OTHER PSYCHOSTIMULANT ABUSE
C0553808|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE
C0553808|T131||LNC|STIMULANT ABUSE NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT
C0553808|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE 
C0553808|T131||LNC|NONDEPENDENT AMPHETAMINE OR OTHER PSYCHOSTIMULANT ABUSE 
C0553808|T131||LNC|NONDEPENDENT AMFETAMINE OR OTHER PSYCHOSTIMULANT ABUSE
C3509117|T131||LNC|STIMULANT ABUSE - UNCOMPLICATED 
C3509117|T131||LNC|STIMULANT ABUSE - UNCOMPLICATED
C3509118|T131||LNC|STIMULANT ABUSE WITH INTOXICATION
C3509118|T131||LNC|STIMULANT ABUSE WITH INTOXICATION 
C3509119|T131||LNC|STIMULANT ABUSE WITH INTOXICATION - UNCOMPLICATED 
C3509119|T131||LNC|STIMULANT ABUSE WITH INTOXICATION - UNCOMPLICATED
C3509120|T131||LNC|STIMULANT ABUSE WITH INTOXICATION DELIRIUM 
C3509120|T131||LNC|STIMULANT ABUSE WITH INTOXICATION DELIRIUM
C3509121|T131||LNC|STIMULANT ABUSE WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE
C3509121|T131||LNC|STIMULANT ABUSE WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE 
C3509126|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED MOOD DISORDER 
C3509126|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED MOOD DISORDER
C3509127|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER
C3509127|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER 
C3509128|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS
C3509128|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS 
C3509129|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS
C3509129|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS 
C3509122|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED DISORDER 
C3509122|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED DISORDER
C3509123|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED ANXIETY DISORDER
C3509123|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED ANXIETY DISORDER 
C3509124|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED SEXUAL FUNCTION 
C3509124|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED SEXUAL FUNCTION
C3509125|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED SLEEP DISORDER 
C3509125|T131||LNC|STIMULANT ABUSE WITH STIMULANT-INDUCED SLEEP DISORDER
C1456332|T131||LNC|STIMULANT ABUSE 
C1456332|T131||LNC|STIMULANT ABUSE
C1456332|T131||LNC|STIMULANT ABUSE 
C1456332|T131||LNC|PSYCHOSTIMULANT ABUSE
C1456332|T131||LNC|ABUSE; STIMULANTS
C1456332|T131||LNC|STIMULANTS; ABUSE
C3494717|T131||LNC|MIRAA ABUSE
C3494717|T131||LNC|KHAT ABUSE
C3494717|T131||LNC|QAT ABUSE
C3494717|T131||LNC|CATHA EDULIS ABUSE 
C3494717|T131||LNC|GAT ABUSE
C3494717|T131||LNC|CATHA EDULIS ABUSE
C3494717|T131||LNC|STIMULANT ABUSE CATJA EDULIS
C3494717|T131||LNC|CATHA EDULIS ABUSE 
C2874626|T131||LNC|OTHER STIMULANT ABUSE, UNCOMPLICATED
C2874631|T131||LNC|OTHER STIMULANT ABUSE WITH INTOXICATION
C2874631|T131||LNC|OTHER STIMULANT ABUSE WITH INTOXICATION, UNSPECIFIED
C2874632|T131||LNC|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED MOOD DISORDER
C2874636|T131||LNC|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED
C2874636|T131||LNC|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER
C2874636|T131||LNC|OTH STIMULANT ABUSE W STIM-INDUCE PSYCHOTIC DISORDER, UNSP
C2874637|T131||LNC|OTHER STIMULANT ABUSE WITH OTHER STIMULANT-INDUCED DISORDER
C2874641|T131||LNC|OTHER STIMULANT ABUSE WITH UNSPECIFIED STIMULANT-INDUCED DISORDER
C2874641|T131||LNC|OTHER STIMULANT ABUSE WITH UNSP STIMULANT-INDUCED DISORDER
C2874628|T131||LNC|OTHER STIMULANT ABUSE WITH INTOXICATION, UNCOMPLICATED
C2874629|T131||LNC|OTHER STIMULANT ABUSE WITH INTOXICATION DELIRIUM
C2874630|T131||LNC|OTHER STIMULANT ABUSE WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE
C2874630|T131||LNC|OTH STIMULANT ABUSE W INTOXICATION W PERCEPTUAL DISTURBANCE
C3662854|T131||LNC|NONDEPENDENT INTRAVEOUS AMPHETAMINE ABUSE 
C3662854|T131||LNC|NONDEPENDENT INTRAVEOUS AMPHETAMINE ABUSE
C3662831|T131||LNC|NONDEPENDENT AMPHETAMINE ABUSE 
C3662831|T131||LNC|NONDEPENDENT AMPHETAMINE ABUSE
C3662831|T131||LNC|STIMULANT ABUSE NONDEPENDENT AMPHETAMINE
C3662831|T131||LNC|NONDEPENDENT AMPHETAMINE ABUSE 
C3836657|T131||LNC|STIMULANT ABUSE NONDEPENDENT AMPHETAMINE INTRAVENOUS
C3836657|T131||LNC|NONDEPENDENT INTRAVENOUS AMPHETAMINE ABUSE 
C3836657|T131||LNC|NONDEPENDENT INTRAVENOUS AMPHETAMINE ABUSE
C2874634|T131||LNC|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS
C2874634|T131||LNC|OTH STIMULANT ABUSE W STIM-INDUCE PSYCH DISORDER W DELUSIONS
C2874635|T131||LNC|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS
C2874635|T131||LNC|OTH STIMULANT ABUSE W STIM-INDUCE PSYCH DISORDER W HALLUCIN
C2874638|T131||LNC|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED ANXIETY DISORDER
C2874638|T131||LNC|OTH STIMULANT ABUSE WITH STIMULANT-INDUCED ANXIETY DISORDER
C2874639|T131||LNC|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED SEXUAL DYSFUNCTION
C2874639|T131||LNC|OTH STIMULANT ABUSE W STIMULANT-INDUCED SEXUAL DYSFUNCTION
C2874640|T131||LNC|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED SLEEP DISORDER
C0338685|T131||LNC|NONDEPENDENT AMFETAMINE OR PSYCHOSTIMULANT ABUSE NOS
C0338685|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE, UNSPECIFIED
C0338685|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE NOS
C0338685|T131||LNC|NONDEPENDENT AMFETAMINE OR PSYCHOSTIMULANT ABUSE, UNSPECIFIED
C0338685|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE, UNSPECIFIED 
C0338685|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE NOS 
C0338683|T131||LNC|STIMULANT ABUSE NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT - EPISODIC
C0338683|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE - EPISODIC
C0338683|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE - EPISODIC 
C0338683|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE, EPISODIC
C0338683|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE, EPISODIC 
C0338683|T131||LNC|NONDEPENDENT AMFETAMINE OR PSYCHOSTIMULANT ABUSE, EPISODIC
C0338683|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE, EPISODIC 
C0338683|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE, EPISODIC 
C0338684|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE IN REMISSION
C0338684|T131||LNC|NONDEPENDENT AMFETAMINE OR PSYCHOSTIMULANT ABUSE IN REMISSION
C0338684|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE IN REMISSION (QUALIFIER VALUE)
C0338684|T131||LNC|STIMULANT ABUSE NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT - IN REMISSION
C0338684|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE - IN REMISSION
C0338684|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE - IN REMISSION 
C0338684|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE IN REMISSION 
C0338684|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE IN REMISSION 
C0338682|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE - CONTINUOUS
C0338682|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE - CONTINUOUS 
C0338682|T131||LNC|STIMULANT ABUSE NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT - CONTINUOUS
C0338682|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE, CONTINUOUS
C0338682|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE, CONTINUOUS 
C0338682|T131||LNC|NONDEPENDENT AMFETAMINE OR PSYCHOSTIMULANT ABUSE, CONTINUOUS
C0338682|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE, CONTINUOUS 
C0338682|T131||LNC|NONDEPENDENT AMPHETAMINE OR PSYCHOSTIMULANT ABUSE, CONTINUOUS 
C2104574|T131||LNC|CONTINUOUS METHAMPHETAMINE ABUSE
C2104574|T131||LNC|CONTINUOUS METHAMPHETAMINE ABUSE 
C2104575|T131||LNC|EPISODIC METHAMPHETAMINE ABUSE 
C2104575|T131||LNC|EPISODIC METHAMPHETAMINE ABUSE
C2104576|T131||LNC|METHAMPHETAMINE ABUSE IN REMISSION 
C2104576|T131||LNC|METHAMPHETAMINE ABUSE IN REMISSION
