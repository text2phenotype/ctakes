C0551008|T034|11011-4|LNC|HEPATITIS C QUANTITATION|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C0551008|T034|11011-4|LNC|HEPATITIS C RNA|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C0551008|T034|11011-4|LNC|HCV LOG10|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C0551008|T034|11011-4|LNC|HCV RNA|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C0551008|T034|11011-4|LNC|HEPATITIS C VIRUS RNA|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C0551008|T034|11011-4|LNC|HEPATITIS C VIRUS RNA:ACNC:PT:SER/PLAS:QN:PROBE.AMP.TAR|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C0551008|T034|11011-4|LNC|LOINC 11011-4|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C0551008|T034|11011-4|LNC|LOINC 38180-6|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C1273338|T034||LNC|HEPATITIS C VIRAL LOAD
C1868902|T034||LNC|HCV VIRAL LOAD
C2697584|T034||LNC|HEPATITIS C VIRAL LOAD PCR MEASUREMENT
C0485398|T034|10676-5|LNC|HEPATITIS C VIRUS RNA|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE WITH AMPLIFICATION
C0485398|T034|10676-5|LNC|HEPATITIS C VIRUS RNA:ACNC:PT:SER/PLAS:QN:PROBE.AMP|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE WITH AMPLIFICATION
C0551008|T034|11011-4|LNC|HEPATITIS C VIRUS RNA:ACNC:PT:SER/PLAS:QN:PROBE.AMP.TAR|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C0803231|T034|20416-4|LNC|HEPATITIS C VIRUS RNA:NCNC:PT:SER/PLAS:QN:PROBE.AMP.TAR|HEPATITIS C VIRUS RIBONUCLEIC ACID:NUMBER CONCENTRATION (COUNT/VOL):POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C0803380|T034|20571-6|LNC|HEPATITIS C VIRUS RNA:NCNC:PT:SER/PLAS:QN:PROBE.AMP.SIG|HEPATITIS C VIRUS RIBONUCLEIC ACID:NUMBER CONCENTRATION (COUNT/VOL):POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.SIG
C0945037|T034|29609-5|LNC|HEPATITIS C VIRUS RNA:ACNC:PT:SER/PLAS:QN:PROBE.AMP.SIG|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.SIG
C1508112|T034|38180-6|LNC|HEPATITIS C VIRUS RNA:LACNC:PT:SER/PLAS:QN:PROBE.AMP.TAR|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C1623573|T034|42003-4|LNC|HEPATITIS C VIRUS RNA:LNCNC:PT:SER/PLAS:QN:PROBE.AMP.SIG|HCV RNA SERPL PROBE+SIG AMP-LOG#
C1643191|T034|42617-1|LNC|HEPATITIS C VIRUS RNA:LACNC:PT:SER/PLAS:QN:PROBE.AMP.SIG|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.SIG
C1831320|T034|47252-2|LNC|HEPATITIS C VIRUS RNA:LNCNC:PT:SER/PLAS:QN:PROBE.AMP.TAR|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG NUMBER CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C1977893|T034|50023-1|LNC|HEPATITIS C VIRUS RNA PANEL:-:PT:SER/PLAS:QN:PROBE.AMP.TAR|HEPATITIS C VIRUS RIBONUCLEIC ACID PANEL:-:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C4064960|T034||LNC|HEPATITIS C VIRUS RNA VIRAL LOAD IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION
C1369569|T034|34703-9|LNC|HEPATITIS C VIRUS RNA:ACNC:PT:SER/PLAS:QN:PROBE.AMP.TAR DETECTION LIMIT = 500 IU/ML|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD DETECTION LIMIT = 500 IU/ML
C1369570|T034|34704-7|LNC|HEPATITIS C VIRUS RNA:ACNC:PT:SER/PLAS:QN:PROBE.AMP.TAR DETECTION LIMIT = 50 IU/ML|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD DETECTION LIMIT = 50 IU/ML
C1977509|T034|49758-6|LNC|HEPATITIS C VIRUS RNA:ACNC:PT:SER/PLAS:QN:PROBE.AMP.TAR DETECTION LIMIT = 5 IU/ML|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD DETECTION LIMIT = 5 IU/ML
C0551008|T034|11011-4|LNC|HEPATITIS C VIRUS RNA:ACNC:PT:SER/PLAS:QN:PROBE.AMP.TAR|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C0551008|T034|11011-4|LNC|HCV RNA SERPL PCR-ACNC|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C0551008|T034|11011-4|LNC|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C0551008|T034|11011-4|LNC|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C1273338|T034||LNC|HEPATITIS C VIRAL LOAD
C1273338|T034||LNC|HEPATITIS C VIRAL LOAD 
C4064960|T034||LNC|PROBE & TARGET AMPLIF HEPATITIS C VIRUS RNA SERUM/PLASMA VIRAL LOAD
C4064960|T034||LNC|HEPATITIS C VIRUS RNA VIRAL LOAD IN SERUM OR PLASMA BY PROBE WITH TARGET AMPLIFICATION 
C4064960|T034||LNC|HEPATITIS C VIRUS RNA VIRAL LOAD IN SERUM OR PLASMA BY PROBE WITH TARGET AMPLIFICATION
C1868902|T034||LNC|HEPATITIS C VIRAL LOAD MEASUREMENT
C1868902|T034||LNC|HCV RNA
C1868902|T034||LNC|HEPATITIS C RNA
C1868902|T034||LNC|HCV VIRAL LOAD
C1868902|T034||LNC|HCVVLD
C0485398|T034|10676-5|LNC|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE WITH AMPLIFICATION|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE WITH AMPLIFICATION
C0485398|T034|10676-5|LNC|HCV RNA SERPL AMP PRB-ACNC|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE WITH AMPLIFICATION
C0485398|T034|10676-5|LNC|HEPATITIS C VIRUS RNA:ACNC:PT:SER/PLAS:QN:PROBE.AMP|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE WITH AMPLIFICATION
C0485398|T034|10676-5|LNC|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE WITH AMPLIFICATION
C0803231|T034|20416-4|LNC|HCV RNA # SERPL PCR|HEPATITIS C VIRUS RIBONUCLEIC ACID:NUMBER CONCENTRATION (COUNT/VOL):POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C0803231|T034|20416-4|LNC|HEPATITIS C VIRUS RNA:NCNC:PT:SER/PLAS:QN:PROBE.AMP.TAR|HEPATITIS C VIRUS RIBONUCLEIC ACID:NUMBER CONCENTRATION (COUNT/VOL):POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C0803231|T034|20416-4|LNC|HEPATITIS C VIRUS RIBONUCLEIC ACID:NUMBER CONCENTRATION (COUNT/VOL):POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR|HEPATITIS C VIRUS RIBONUCLEIC ACID:NUMBER CONCENTRATION (COUNT/VOL):POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C0803231|T034|20416-4|LNC|HEPATITIS C VIRUS RNA [#/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD|HEPATITIS C VIRUS RIBONUCLEIC ACID:NUMBER CONCENTRATION (COUNT/VOL):POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C0803380|T034|20571-6|LNC|HCV RNA # SERPL BDNA|HEPATITIS C VIRUS RIBONUCLEIC ACID:NUMBER CONCENTRATION (COUNT/VOL):POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.SIG
C0803380|T034|20571-6|LNC|HEPATITIS C VIRUS RNA:NCNC:PT:SER/PLAS:QN:PROBE.AMP.SIG|HEPATITIS C VIRUS RIBONUCLEIC ACID:NUMBER CONCENTRATION (COUNT/VOL):POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.SIG
C0803380|T034|20571-6|LNC|HEPATITIS C VIRUS RIBONUCLEIC ACID:NUMBER CONCENTRATION (COUNT/VOL):POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.SIG|HEPATITIS C VIRUS RIBONUCLEIC ACID:NUMBER CONCENTRATION (COUNT/VOL):POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.SIG
C0803380|T034|20571-6|LNC|HEPATITIS C VIRUS RNA [#/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND SIGNAL AMPLIFICATION METHOD|HEPATITIS C VIRUS RIBONUCLEIC ACID:NUMBER CONCENTRATION (COUNT/VOL):POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.SIG
C0945037|T034|29609-5|LNC|HCV RNA SERPL BDNA-ACNC|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.SIG
C0945037|T034|29609-5|LNC|HEPATITIS C VIRUS RNA:ACNC:PT:SER/PLAS:QN:PROBE.AMP.SIG|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.SIG
C0945037|T034|29609-5|LNC|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.SIG|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.SIG
C0945037|T034|29609-5|LNC|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND SIGNAL AMPLIFICATION METHOD|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.SIG
C1508112|T034|38180-6|LNC|HEPATITIS C VIRUS RNA:LACNC:PT:SER/PLAS:QN:PROBE.AMP.TAR|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C1508112|T034|38180-6|LNC|HCV RNA SERPL PCR-LOG IU|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C1508112|T034|38180-6|LNC|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C1508112|T034|38180-6|LNC|HEPATITIS C VIRUS RNA [LOG UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C1623573|T034|42003-4|LNC|HEPATITIS C VIRUS RNA:LNCNC:PT:SER/PLAS:QN:PROBE.AMP.SIG|HCV RNA SERPL PROBE+SIG AMP-LOG#
C1623573|T034|42003-4|LNC|HCV RNA SERPL BDNA-LOG#|HCV RNA SERPL PROBE+SIG AMP-LOG#
C1623573|T034|42003-4|LNC|HEPATITIS C VIRUS RNA [LOG #/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND SIGNAL AMPLIFICATION METHOD|HCV RNA SERPL PROBE+SIG AMP-LOG#
C1623573|T034|42003-4|LNC|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG NUMBER CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.SIG|HCV RNA SERPL PROBE+SIG AMP-LOG#
C1643191|T034|42617-1|LNC|HCV RNA SERPL BDNA-LOG IU|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.SIG
C1643191|T034|42617-1|LNC|HEPATITIS C VIRUS RNA:LACNC:PT:SER/PLAS:QN:PROBE.AMP.SIG|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.SIG
C1643191|T034|42617-1|LNC|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.SIG|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.SIG
C1643191|T034|42617-1|LNC|HEPATITIS C VIRUS RNA [LOG UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND SIGNAL AMPLIFICATION METHOD|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.SIG
C1831320|T034|47252-2|LNC|HEPATITIS C VIRUS RNA:LNCNC:PT:SER/PLAS:QN:PROBE.AMP.TAR|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG NUMBER CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C1831320|T034|47252-2|LNC|HCV RNA SERPL PCR-LOG#|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG NUMBER CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C1831320|T034|47252-2|LNC|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG NUMBER CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG NUMBER CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C1831320|T034|47252-2|LNC|HEPATITIS C VIRUS RNA [LOG #/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG NUMBER CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C1977157|T034|49371-8|LNC|HEPATITIS C VIRUS RNA [#/VOLUME] (VIRAL LOAD) IN TISSUE BY PROBE AND TARGET AMPLIFICATION METHOD|HEPATITIS C VIRUS RIBONUCLEIC ACID:NUMBER CONCENTRATION (COUNT/VOL):POINT IN TIME:TISSUE, UNSPECIFIED:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C1977158|T034|49372-6|LNC|HEPATITIS C VIRUS RNA:LNCNC:PT:XXX:QN:PROBE.AMP.TAR|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG NUMBER CONCENTRATION:POINT IN TIME:TO BE SPECIFIED IN ANOTHER PART OF THE MESSAGE:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C1977158|T034|49372-6|LNC|HCV RNA XXX PCR-LOG#|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG NUMBER CONCENTRATION:POINT IN TIME:TO BE SPECIFIED IN ANOTHER PART OF THE MESSAGE:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C1977158|T034|49372-6|LNC|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG NUMBER CONCENTRATION:POINT IN TIME:TO BE SPECIFIED IN ANOTHER PART OF THE MESSAGE:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG NUMBER CONCENTRATION:POINT IN TIME:TO BE SPECIFIED IN ANOTHER PART OF THE MESSAGE:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C1977158|T034|49372-6|LNC|HEPATITIS C VIRUS RNA [LOG #/VOLUME] (VIRAL LOAD) IN UNSPECIFIED SPECIMEN BY PROBE AND TARGET AMPLIFICATION METHOD|HEPATITIS C VIRUS RIBONUCLEIC ACID:LOG NUMBER CONCENTRATION:POINT IN TIME:TO BE SPECIFIED IN ANOTHER PART OF THE MESSAGE:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C1977893|T034|50023-1|LNC|HCV RNA PNL SERPL PCR|HEPATITIS C VIRUS RIBONUCLEIC ACID PANEL:-:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C1977893|T034|50023-1|LNC|HEPATITIS C VIRUS RNA PANEL:-:PT:SER/PLAS:QN:PROBE.AMP.TAR|HEPATITIS C VIRUS RIBONUCLEIC ACID PANEL:-:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C1977893|T034|50023-1|LNC|HEPATITIS C VIRUS RIBONUCLEIC ACID PANEL:-:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR|HEPATITIS C VIRUS RIBONUCLEIC ACID PANEL:-:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C1977893|T034|50023-1|LNC|HEPATITIS C VIRUS RNA PANEL (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD|HEPATITIS C VIRUS RIBONUCLEIC ACID PANEL:-:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR
C1369569|T034|34703-9|LNC|HEPATITIS C VIRUS RNA:ACNC:PT:SER/PLAS:QN:PROBE.AMP.TAR DETECTION LIMIT = 500 IU/ML|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD DETECTION LIMIT = 500 IU/ML
C1369569|T034|34703-9|LNC|HCV RNA SERPL PCR DL=500-ACNC|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD DETECTION LIMIT = 500 IU/ML
C1369569|T034|34703-9|LNC|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR DETECTION LIMIT = 500 IU/ML|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD DETECTION LIMIT = 500 IU/ML
C1369569|T034|34703-9|LNC|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD DETECTION LIMIT = 500 IU/ML|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD DETECTION LIMIT = 500 IU/ML
C1369570|T034|34704-7|LNC|HEPATITIS C VIRUS RNA:ACNC:PT:SER/PLAS:QN:PROBE.AMP.TAR DETECTION LIMIT = 50 IU/ML|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD DETECTION LIMIT = 50 IU/ML
C1369570|T034|34704-7|LNC|HCV RNA SERPL PCR DL=50-ACNC|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD DETECTION LIMIT = 50 IU/ML
C1369570|T034|34704-7|LNC|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR DETECTION LIMIT = 50 IU/ML|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD DETECTION LIMIT = 50 IU/ML
C1369570|T034|34704-7|LNC|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD DETECTION LIMIT = 50 IU/ML|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD DETECTION LIMIT = 50 IU/ML
C1977509|T034|49758-6|LNC|HEPATITIS C VIRUS RNA:ACNC:PT:SER/PLAS:QN:PROBE.AMP.TAR DETECTION LIMIT = 5 IU/ML|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD DETECTION LIMIT = 5 IU/ML
C1977509|T034|49758-6|LNC|HCV RNA SERPL PCR DL=5-ACNC|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD DETECTION LIMIT = 5 IU/ML
C1977509|T034|49758-6|LNC|HEPATITIS C VIRUS RIBONUCLEIC ACID:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DNA NUCLEIC ACID PROBE.AMP.TAR DETECTION LIMIT = 5 IU/ML|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD DETECTION LIMIT = 5 IU/ML
C1977509|T034|49758-6|LNC|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD DETECTION LIMIT = 5 IU/ML|HEPATITIS C VIRUS RNA [UNITS/VOLUME] (VIRAL LOAD) IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD DETECTION LIMIT = 5 IU/ML
