C1328839|T047||SNOMEDCT_US|AUTOIMMUNE INFLAMMATORY BOWEL DISEASE
C0400936|T047|235890007|SNOMEDCT_US|AUTOIMMUNE LIVER DISEASE|AUTOIMMUNE LIVER DISEASE (DISORDER)
C0400936|T047|235890007|SNOMEDCT_US|AUTOIMMUNE LIVER DISEASE |AUTOIMMUNE LIVER DISEASE (DISORDER)
C0854359|T047|408539000|SNOMEDCT_US|AUTOIMMUNE ENDOCRINE DISEASE INSULIN SYNDROME|INSULIN AUTOIMMUNE SYNDROME (DISORDER)
C1328839|T047||SNOMEDCT_US|AUTOIMMUNE INFLAMMATORY BOWEL DISEASE
C0854359|T047|408539000|SNOMEDCT_US|AUTOIMMUNE INSULIN SYNDROME|INSULIN AUTOIMMUNE SYNDROME (DISORDER)
C0854359|T047|408539000|SNOMEDCT_US|AUTOIMMUNE INSULIN SYNDROME |INSULIN AUTOIMMUNE SYNDROME (DISORDER)
C0400936|T047|235890007|SNOMEDCT_US|AUTOIMMUNE LIVER DISEASE|AUTOIMMUNE LIVER DISEASE (DISORDER)
C0400936|T047|235890007|SNOMEDCT_US|AUTOIMMUNE LIVER DISEASE |AUTOIMMUNE LIVER DISEASE (DISORDER)
C0004364|T047|85828009|SNOMEDCT_US|AUTOIMMUNE SYKDOMMER|AUTOIMMUNE DISEASE (DISORDER)
C0854359|T047|408539000|SNOMEDCT_US|INSULIN AUTOIMMUNE SYNDROME|INSULIN AUTOIMMUNE SYNDROME (DISORDER)
C0854359|T047|408539000|SNOMEDCT_US|INSULIN AUTOIMMUNE SYNDROME |INSULIN AUTOIMMUNE SYNDROME (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|CROHN DISEASE|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|CROHNS DISEASE|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|CROHN'S DISEASE|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|CROHN'S DISEASE [REGIONAL ENTERITIS]|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|CROHN'S DISEASE, UNSPECIFIED|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|INFLAMMATORY BOWEL DISEASE 1|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|IBD1|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|CROHN DIS|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|CROHNS DIS|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|ELEOCOLITIS|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|ENTERITIS (REGIONAL)|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|CROHN'S DISEASE, NOS|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|CROHN'S DISEASE |CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|CROHN'S ILEITIS|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|REGIONAL ENTERITIS|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|GRANULOMATOUS ENTERITIS|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|CROHN'S DISEASE NOS|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|CROHN DISEASE [DISEASE/FINDING]|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|DISEASE;CROHNS|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|REGIONAL ENTERITIS - CROHN'S DISEASE|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|REGIONAL ENTERITIS - CROHN|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|CROHN'S REGIONAL ENTERITIS|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|CROHN'S ENTERITIS|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|-- CROHN'S DISEASE|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|MORBUS CROHN|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|GRANULOMATOUS ENTERITIS AND COLITIS|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|DISEASE CROHNS|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|CROHN'S|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|CD - CROHN'S DISEASE|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|RE - REGIONAL ENTERITIS|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|CROHN'S DISEASE |CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|CROHN|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|GRANULOMATOUS ENTERITIS, NOS|CROHN'S DISEASE (DISORDER)
C0010346|T047|34000006|SNOMEDCT_US|REGIONAL ENTERITIS, NOS|CROHN'S DISEASE (DISORDER)
C0678202|T047|196984001|SNOMEDCT_US|REGIONAL ENTERITIS|REGIONAL ENTERITIS NOS (DISORDER)
C0678202|T047|196984001|SNOMEDCT_US|REGIONAL ENTERITIS |REGIONAL ENTERITIS NOS (DISORDER)
C0678202|T047|196984001|SNOMEDCT_US|REGIONAL ENTERITIS NOS|REGIONAL ENTERITIS NOS (DISORDER)
C0678202|T047|196984001|SNOMEDCT_US|ENTERITIS;REGIONAL|REGIONAL ENTERITIS NOS (DISORDER)
C0678202|T047|196984001|SNOMEDCT_US|GRANULOMATOUS ENTERITIS|REGIONAL ENTERITIS NOS (DISORDER)
C0678202|T047|196984001|SNOMEDCT_US|REGIONAL ENTERITIS |REGIONAL ENTERITIS NOS (DISORDER)
C0678202|T047|196984001|SNOMEDCT_US|ENTERITIS - REGIONAL|REGIONAL ENTERITIS NOS (DISORDER)
C0678202|T047|196984001|SNOMEDCT_US|REGIONAL ENTERITIS NOS |REGIONAL ENTERITIS NOS (DISORDER)
C0678202|T047|196984001|SNOMEDCT_US|GRANULOMATOUS ENTERITIS |REGIONAL ENTERITIS NOS (DISORDER)
C0678202|T047|196984001|SNOMEDCT_US|REGIONAL ENTERITIS OF UNSPECIFIED SITE|REGIONAL ENTERITIS NOS (DISORDER)
C0678202|T047|196984001|SNOMEDCT_US|ENTERITIS, REGIONAL|REGIONAL ENTERITIS NOS (DISORDER)
C0678202|T047|196984001|SNOMEDCT_US|BOWEL; REGIONAL ENTERITIS|REGIONAL ENTERITIS NOS (DISORDER)
C0678202|T047|196984001|SNOMEDCT_US|ENTERITIS, GRANULOMATOUS|REGIONAL ENTERITIS NOS (DISORDER)
C0267807|T047|19682006|SNOMEDCT_US|LUPUS HEPATITIS|LUPUS HEPATITIS (DISORDER)
C0267807|T047|19682006|SNOMEDCT_US|LUPOID HEPATITIS|LUPUS HEPATITIS (DISORDER)
C0267807|T047|19682006|SNOMEDCT_US|LUPUS HEPATITIS |LUPUS HEPATITIS (DISORDER)
C0267807|T047|19682006|SNOMEDCT_US|HEPATITIS; LUPOID|LUPUS HEPATITIS (DISORDER)
C0267807|T047|19682006|SNOMEDCT_US|LUPOID; HEPATITIS|LUPUS HEPATITIS (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|PRIMARY BILIARY CIRRHOSIS|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|PRIMARY BILIARY CIRRHOSIS |BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|BILIARY CIRRHOSIS PRIMARY|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|PBC|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|PBC1|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|BILIARY CIRRHOSIS, PRIMARY, 1|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|PRIMARY BILARY CIRRHOSIS (PBC)|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|CHRONIC NONSUPPURATIVE DESTRUCTIVE CHOLANGITIS|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|BILIARY CIRRHOSIS (& [PRIMARY]) |BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|BILIARY CIRRHOSIS|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|BILIARY CIRRHOSIS (& [PRIMARY])|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|CHRONIC NON-SUPPURATIVE DESTRUCTIVE CHOLANGITIS|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|CHOLANGITIS, CHRONIC NONSUPPURATIVE DESTRUCTIVE|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|PBC- PRIMARY BILIARY CIRRHOSIS|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|PRIMARY BILIARY CIRRHOSIS |BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|BILIARY; CIRRHOSIS, PRIMARY|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|HANOT|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|CHOLANGITIS; CHRONIC NONSUPPURATIVE DESTRUCTIVE|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|CHRONIC; CHOLANGITIS, CHRONIC NONSUPPURATIVE DESTRUCTIVE, DESTRUCTIVE|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|CIRRHOSIS; BILIARY, PRIMARY|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|BILIARY CIRRHOSIS, PRIMARY|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|CIRRHOSIS;BILIARY;PRIMARY|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0241910|T047|408335007|SNOMEDCT_US|AUTOIMMUNE HEPATITIDES|AUTOIMMUNE HEPATITIS (DISORDER)
C0241910|T047|408335007|SNOMEDCT_US|AUTOIMMUNE HEPATITIS|AUTOIMMUNE HEPATITIS (DISORDER)
C0241910|T047|408335007|SNOMEDCT_US|HEPATITIDES, AUTOIMMUNE|AUTOIMMUNE HEPATITIS (DISORDER)
C0241910|T047|408335007|SNOMEDCT_US|HEPATITIS, AUTOIMMUNE|AUTOIMMUNE HEPATITIS (DISORDER)
C0241910|T047|408335007|SNOMEDCT_US|AUTOIMMUNE HEPATITIS |AUTOIMMUNE HEPATITIS (DISORDER)
C0241910|T047|408335007|SNOMEDCT_US|HEPATITIS CHRONIC ACTIVE AUTOIMMUNE|AUTOIMMUNE HEPATITIS (DISORDER)
C0241910|T047|408335007|SNOMEDCT_US|CHRONIC ACTIVE AUTOIMMUNE HEPATITIS|AUTOIMMUNE HEPATITIS (DISORDER)
C0241910|T047|408335007|SNOMEDCT_US|CHRONIC ACTIVE AUTOIMMUNE HEPATITIS |AUTOIMMUNE HEPATITIS (DISORDER)
C0241910|T047|408335007|SNOMEDCT_US|HEPATITIDES, AUTOIMMUNE CHRONIC|AUTOIMMUNE HEPATITIS (DISORDER)
C0241910|T047|408335007|SNOMEDCT_US|HEPATITIS, AUTOIMMUNE CHRONIC|AUTOIMMUNE HEPATITIS (DISORDER)
C0241910|T047|408335007|SNOMEDCT_US|AUTOIMMUNE CHRONIC HEPATITIDES|AUTOIMMUNE HEPATITIS (DISORDER)
C0241910|T047|408335007|SNOMEDCT_US|CHRONIC HEPATITIDES, AUTOIMMUNE|AUTOIMMUNE HEPATITIS (DISORDER)
C0241910|T047|408335007|SNOMEDCT_US|CHRONIC HEPATITIS, AUTOIMMUNE|AUTOIMMUNE HEPATITIS (DISORDER)
C0241910|T047|408335007|SNOMEDCT_US|HEPATITIS, AUTOIMMUNE [DISEASE/FINDING]|AUTOIMMUNE HEPATITIS (DISORDER)
C0241910|T047|408335007|SNOMEDCT_US|AUTOIMMUNE CHRONIC HEPATITIS|AUTOIMMUNE HEPATITIS (DISORDER)
C0241910|T047|408335007|SNOMEDCT_US|HEPATITIS AUTOIMMUNE|AUTOIMMUNE HEPATITIS (DISORDER)
C0241910|T047|408335007|SNOMEDCT_US|AUTOIMMUNE CHRONIC ACTIVE HEPATITIS|AUTOIMMUNE HEPATITIS (DISORDER)
C0241910|T047|408335007|SNOMEDCT_US|AUTOIMMUNE HEPATITIS |AUTOIMMUNE HEPATITIS (DISORDER)
C0241910|T047|408335007|SNOMEDCT_US|AUTOIMMUNE; HEPATITIS|AUTOIMMUNE HEPATITIS (DISORDER)
C0241910|T047|408335007|SNOMEDCT_US|HEPATITIS; AUTOIMMUNE|AUTOIMMUNE HEPATITIS (DISORDER)
C0854359|T047|408539000|SNOMEDCT_US|INSULIN AUTOIMMUNE SYNDROME|INSULIN AUTOIMMUNE SYNDROME (DISORDER)
C0854359|T047|408539000|SNOMEDCT_US|AUTOIMMUNE ENDOCRINE DISEASE INSULIN SYNDROME|INSULIN AUTOIMMUNE SYNDROME (DISORDER)
C0854359|T047|408539000|SNOMEDCT_US|AUTOIMMUNE INSULIN SYNDROME|INSULIN AUTOIMMUNE SYNDROME (DISORDER)
C0854359|T047|408539000|SNOMEDCT_US|AUTOIMMUNE INSULIN SYNDROME |INSULIN AUTOIMMUNE SYNDROME (DISORDER)
C0854359|T047|408539000|SNOMEDCT_US|INSULIN AUTOIMMUNE SYNDROME |INSULIN AUTOIMMUNE SYNDROME (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|REITER'S SYNDROME|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|REITER'S DISEASE|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|REITERS DISEASE|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|REITER DIS|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|DISEASE, REITER'S|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|SYNDROME, REITER|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|DISEASE, REITER|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|REITERS DIS|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|FIESSINGER LEROY REITER SYNDROME|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|REITER'S SYNDROME WITH ARTHROPATHY|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|REITER'S SYNDROME WITH ARTHROPATHY |REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|REITER'S SYNDROME |REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|REITER SYNDROME|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|REITER DISEASE|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|REITER'S DISEASE, UNSPECIFIED SITE|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|REITERS SYNDROME|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|REITER'S DISEASE |REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|FIESSINGER-LEROY-REITER SYNDROME|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|URETHROOCULOARTICULAR SYNDROME|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|ARTHRITIS; URETHRITICA|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|REITER; TRIAD|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|REITER|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|SYNDROME; URETHRO-OCULO-ARTICULAR|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|TRIAD; REITER|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|URETHRITICA; ARTHRITIS|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|URETHRO-OCULO-ARTICULAR; SYNDROME|REITER'S DISEASE (DISORDER)
C0035012|T047|67224007|SNOMEDCT_US|UROARTHRITIS; INFECTIOUS|REITER'S DISEASE (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|ADDISONS DISEASE|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|DISEASE, ADDISON|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|ADDISON'S DISEASE|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|PRIMARY ADRENOCORTICAL INSUFFICIENCY|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|ADRENAL INSUFFICIENCY (ADDISON DISEASE)|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|ADDISON DISEASE|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|PRIMARY ADRENOCORTICAL FAILURE|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|ADDISONS DIS|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|ADDISON DIS|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|ADDISON'S DISEASE NOS|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|PRIMARY ADRENAL INSUFFICIENCY|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|PRIMARY ADRENAL INSUFFICIENCY |PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|ADDISON DISEASE [DISEASE/FINDING]|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|PRIMARY HYPOADRENALISM|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|DISEASE;ADDISONS|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|HYPOCORTISOLISM|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|ADDISON'S DISEASE, NOS|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|ADDISON'S DISEASE |PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|ADDISON'S DISEASE, NOS |PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|PRIMARY ADRENAL DEFICIENCY|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|CHRONIC PRIMARY ADRENAL INSUFFICIENCY|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|DISEASE ADDISON'S|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|PRIMARY ADRENOCORTICAL INSUFFICIENCY |PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|CORTICOADRENAL; DEFICIENCY, PRIMARY|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|DEFICIENCY; ADRENOCORTICAL, PRIMARY|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|DEFICIENCY; CORTICOADRENAL, PRIMARY|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|DISEASE (OR DISORDER); BRONZED SKIN (ADDISON) (BRONZE DISEASE)|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|HYPOADRENOCORTICISM; PRIMARY|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|INSUFFICIENCY; ADRENAL, PRIMARY|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|INSUFFICIENCY; SUPRARENAL, PRIMARY|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|ADRENAL CORTEX; DEFICIENCY, PRIMARY|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|ADRENAL CORTEX; HYPOFUNCTION, PRIMARY|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|ADRENAL; INSUFFICIENCY, PRIMARY|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|PRIMARY; HYPOADRENOCORTICISM|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|ADDISON; DISEASE OR SYNDROME|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|SUPRARENAL; INSUFFICIENCY, PRIMARY|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|SYNDROME; ADDISON|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|ADDISON'S DISEASE [AMBIGUOUS]|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|HYPOADRENALISM, PRIMARY|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|HYPOADRENALISMS, PRIMARY|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|INSUFFICIENCIES, PRIMARY ADRENOCORTICAL|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|INSUFFICIENCY, PRIMARY ADRENOCORTICAL|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|PRIMARY ADRENOCORTICAL INSUFFICIENCIES|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|ADRENAL INSUFFICIENCY, PRIMARY|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|ADRENOCORTICAL INSUFFICIENCIES, PRIMARY|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C0001403|T047|373662000|SNOMEDCT_US|ADRENOCORTICAL INSUFFICIENCY, PRIMARY|PRIMARY ADRENOCORTICAL INSUFFICIENCY (DISORDER)
C1527336|T047|201444003|SNOMEDCT_US|SJOGREN'S SYNDROME|SICCA (SJOGREN'S) SYNDROME
C1527336|T047|201444003|SNOMEDCT_US|SYNDROME, SJOGREN'S|SICCA (SJOGREN'S) SYNDROME
C1527336|T047|201444003|SNOMEDCT_US|SJOGRENS SYNDROME|SICCA (SJOGREN'S) SYNDROME
C1527336|T047|201444003|SNOMEDCT_US|SICCA SYNDROME [SJOGREN]|SICCA (SJOGREN'S) SYNDROME
C1527336|T047|201444003|SNOMEDCT_US|SJOGREN'S DISEASE|SICCA (SJOGREN'S) SYNDROME
C1527336|T047|201444003|SNOMEDCT_US|SJOGREN SYNDROME|SICCA (SJOGREN'S) SYNDROME
C1527336|T047|201444003|SNOMEDCT_US|SJOGREN'S SYNDROME [DISEASE/FINDING]|SICCA (SJOGREN'S) SYNDROME
C1527336|T047|201444003|SNOMEDCT_US|SICCA (SJOGREN'S) SYNDROME|SICCA (SJOGREN'S) SYNDROME
C1527336|T047|201444003|SNOMEDCT_US|SJOGREN SYNDROME |SICCA (SJOGREN'S) SYNDROME
C1527336|T047|201444003|SNOMEDCT_US|SJOGREN'S|SICCA (SJOGREN'S) SYNDROME
C1527336|T047|201444003|SNOMEDCT_US|GOUGEROT-MULOCK-HOUWER SYNDROME|SICCA (SJOGREN'S) SYNDROME
C1527336|T047|201444003|SNOMEDCT_US|SYNDROME SJOGREN'S|SICCA (SJOGREN'S) SYNDROME
C1527336|T047|201444003|SNOMEDCT_US|SJOEGREN'S SYNDROME|SICCA (SJOGREN'S) SYNDROME
C1527336|T047|201444003|SNOMEDCT_US|SJÖGREN'S SYNDROME |SICCA (SJOGREN'S) SYNDROME
C1527336|T047|201444003|SNOMEDCT_US|SJÖGREN|SICCA (SJOGREN'S) SYNDROME
C0002880|T047|413603009|SNOMEDCT_US|AUTOIMMUNE HEMOLYTIC ANEMIA|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|ANEMIA, HEMOLYTIC, AUTOIMMUNE|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|HEMOLYTIC ANEMIA, AUTOIMMUNE|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|ANEMIA, AUTOIMMUNE HEMOLYTIC|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|AUTOIMMUN HEMOLYTIC ANEM|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|ANEMIA, HEMOLYTIC, AUTOIMMUNE [DISEASE/FINDING]|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|AUTOIMMUNE HAEMOLYTIC ANAEMIAS|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|AIHA - AUTOIMMUNE HEMOLYTIC ANEMIA|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|AIHA - AUTOIMMUNE HAEMOLYTIC ANAEMIA|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|AUTOIMMUNE HAEMOLYTIC ANAEMIA |AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|AUTOIMMUNE HEMOLYTIC ANEMIA NOS |AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|AUTOIMMUNE HAEMOLYTIC ANAEMIA|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|HEMOLYTIC ANEMIA DUE TO ANTIBODY|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|AUTOIMMUNE HEMOLYTIC ANEMIA NOS|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|HAEMOLYTIC ANAEMIA DUE TO ANTIBODY|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|AUTOIMMUNE HEMOLYTIC ANEMIA |AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|AUTOIMMUNE HEMOLYTIC ANEMIAS|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|AUTOIMMUNE HAEMOLYTIC ANAEMIA NOS|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|IMMUNE MEDIATED HEMOLYTIC ANEMIA|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|ANEMIA HEMOLYTIC AUTOIMMUNE (NOS)|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|ANAEMIA HAEMOLYTIC AUTOIMMUNE|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|ANEMIA HEMOLYTIC AUTOIMMUNE|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|HEMOLYTIC; ANEMIA, AUTOIMMUNE|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|ANEMIA; HEMOLYTIC, AUTOIMMUNE|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|AUTOIMMUNE HEMOLYTIC ANEMIA, NOS|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|HEMOLYTIC ANEMIA DUE TO ANTIBODY, NOS|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|ANEMIAS, AUTOIMMUNE HEMOLYTIC|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0002880|T047|413603009|SNOMEDCT_US|HEMOLYTIC ANEMIAS, AUTOIMMUNE|AUTOIMMUNE HEMOLYTIC ANEMIA (DISORDER)
C0020951|T047||SNOMEDCT_US|GREY AREA TO ME. HYPERSENSITIVITY AND AUTOIMMUNITY ARE IN DIFFERENT BUCKETS IN MY HEAD, BUT I SUPPOSE A TYPE III IS PRETTY MUCH ALWAYS DUE TO AUTOIMMUNITY
C0020951|T047||SNOMEDCT_US|DISEASE, IMMUNE COMPLEX
C0020951|T047||SNOMEDCT_US|DISEASES, IMMUNE COMPLEX
C0020951|T047||SNOMEDCT_US|HYPERSENSITIVITIES, TYPE III
C0020951|T047||SNOMEDCT_US|TYPE III HYPERSENSITIVITIES
C0020951|T047||SNOMEDCT_US|IMMUNE COMPLEX DISEASE
C0020951|T047||SNOMEDCT_US|IMMUNE COMPLEX DIS
C0020951|T047||SNOMEDCT_US|IMMUNE COMPLEX DISEASES [DISEASE/FINDING]
C0020951|T047||SNOMEDCT_US|TYPE III HYPERSENSITIVITY
C0020951|T047||SNOMEDCT_US|HYPERSENSITIVITY, TYPE III
C0011854|T047|190362004|SNOMEDCT_US|BRITTLE DIABETES MELLITUS|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, JUVENILE ONSET|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, KETOSIS PRONE|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|JUVENILE-ONSET DIABETES MELLITUS|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|KETOSIS-PRONE DIABETES MELLITUS|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, SUDDEN ONSET|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|MELLITUS, SUDDEN-ONSET DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|SUDDEN-ONSET DIABETES MELLITUS|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|JOD|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|IDDM1|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|INSULIN-DEPENDENT DIABETES MELLITUS 1|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|INSULIN-DEPENDENT DIABETES MELLITUS (TYPE I)|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, INSULIN-DEPENDENT, 1|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS TYPE 01|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|TYPE I DIABETES MELLITUS|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|JUVENILE DIABETES MELLITUS|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|KETOSIS PRONE DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|TYPE 1 DIABETES MELLITUS|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|TYPE 1 DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|TYPE I DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|JUVENILE DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, KETOSIS-PRONE|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|KPD|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|BRITTLE DIABETES (MELLITUS)|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|JUVENILE ONSET DIABETES (MELLITUS)|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|KETOSIS-PRONE DIABETES (MELLITUS)|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, TYPE 1 [DISEASE/FINDING]|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, BRITTLE|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, TYPE 1|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, JUVENILE-ONSET|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, SUDDEN-ONSET|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, TYPE I|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES;TYPE 1|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES;INSULIN DEPENDENT|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES;JUVENILE ONSET|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|INSULIN DEPENDENT DIABETES MELLITUS 1|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|JUVENILE ONSET DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES, JUVENILE-ONSET|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|JUVENILE-ONSET DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES TYPE 1|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|INSULIN-DEPENDENT DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS: [JUVENILE] OR [INSULIN DEPENDENT]|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS - JUVENILE|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS: [JUVENILE] OR [INSULIN DEPENDENT] |TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS TYPE 1|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|JUVENILE ONSET DIABETES MELLITUS|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|TYPE I DIABETES MELLITUS |TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|IDDM - INSULIN-DEPENDENT DIABETES MELLITUS|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|INSULIN DEPENDENT DIABETES MEL|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|-- DIABETES TYPE 1|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS TYPE I|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|TYPE 1 DIABETES MELLITUS |TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS JUVENILE ONSET|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS INSULIN-DEPENDENT|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS TYPE 1 |TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES; JUVENILE-ONSET|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES; KETOSIS-PRONE|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES; TYPE I|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|JUVENILE-ONSET; DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|KETOSIS, PRONE; DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|TYPE I; DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|JUVENILE ONSET OF DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|MULTIPLE SCLEROSIS|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|DISSEMINATED SCLEROSIS|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|MS|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|SCLEROSIS, MULTIPLE|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|INSULAR SCLEROSIS|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|MULTIPLE SCLEROSIS |MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|GENERALIZED MULTIPLE SCLEROSIS|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|GENERALIZED MULTIPLE SCLEROSIS |MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|SCLEROSIS, DISSEMINATED|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|MS (MULTIPLE SCLEROSIS)|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|MULTIPLE SCLEROSIS [DISEASE/FINDING]|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|SCLEROSIS;DISSEMINATED|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|MULTIPLE SCLEROSIS NOS|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|MULTIPLE SCLEROSIS NOS |MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|MULTIPLE SCLEROSIS |MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|MULTIPLE SCLEROSIS - MS|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|GENERALISED MULTIPLE SCLEROSIS|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|SCLEROSIS MULTIPLE|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|NEURO: MULTIPLE SCLEROSIS|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|DS - DISSEMINATED SCLEROSIS|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|MS - MULTIPLE SCLEROSIS|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|GENERALIZED MULTIPLE SCLEROSIS |MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|CEREBROSPINAL; SCLEROSIS|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|DISSEMINATED; SCLEROSIS|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|INSULAR; SCLEROSIS|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|SCLEROSIS; CEREBROSPINAL|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|SCLEROSIS; DISSEMINATED|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|SCLEROSIS; INSULAR|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|SCLEROSIS; MULTIPLE|MULTIPLE SCLEROSIS (DISORDER)
C0026769|T047|24700007|SNOMEDCT_US|MULTIPLE SCLEROSIS, NOS|MULTIPLE SCLEROSIS (DISORDER)
C0026896|T047|91637004|SNOMEDCT_US|MYASTHENIA GRAVIS|MYASTHENIA GRAVIS (DISORDER)
# C0026896|T047|91637004|SNOMEDCT_US|MG|MYASTHENIA GRAVIS (DISORDER)
C0026896|T047|91637004|SNOMEDCT_US|MYASTHENIA GRAVIS |MYASTHENIA GRAVIS (DISORDER)
C0026896|T047|91637004|SNOMEDCT_US|MYASTHENIA GRAVIS NOS|MYASTHENIA GRAVIS (DISORDER)
C0026896|T047|91637004|SNOMEDCT_US|MYASTHENIA GRAVIS [DISEASE/FINDING]|MYASTHENIA GRAVIS (DISORDER)
C0026896|T047|91637004|SNOMEDCT_US|MYASTHENIA GRAVIS NOS |MYASTHENIA GRAVIS (DISORDER)
C0026896|T047|91637004|SNOMEDCT_US|MYASTHENIA GRAVIS |MYASTHENIA GRAVIS (DISORDER)
C0026896|T047|91637004|SNOMEDCT_US|MYASTHENIA GRAVIS PARALYTICA|MYASTHENIA GRAVIS (DISORDER)
C0026896|T047|91637004|SNOMEDCT_US|ERB-GOLDFLAM DISEASE|MYASTHENIA GRAVIS (DISORDER)
C0026896|T047|91637004|SNOMEDCT_US|MG - MYASTHENIA GRAVIS|MYASTHENIA GRAVIS (DISORDER)
C0026896|T047|91637004|SNOMEDCT_US|ERB-GOLDFLAM|MYASTHENIA GRAVIS (DISORDER)
C0026896|T047|91637004|SNOMEDCT_US|GOLDFLAM-ERB|MYASTHENIA GRAVIS (DISORDER)
C0026896|T047|91637004|SNOMEDCT_US|GRAVIS; MYASTHENIA|MYASTHENIA GRAVIS (DISORDER)
C0026896|T047|91637004|SNOMEDCT_US|MYASTHENIA; GRAVIS|MYASTHENIA GRAVIS (DISORDER)
C0026896|T047|91637004|SNOMEDCT_US|MYASTHENIA GRAVIS, NOS|MYASTHENIA GRAVIS (DISORDER)
C0030807|T047|65172003|SNOMEDCT_US|PEMPHIGUS|PEMPHIGUS (DISORDER)
C0030807|T047|65172003|SNOMEDCT_US|PEMPHIGUS, UNSPECIFIED|PEMPHIGUS (DISORDER)
C0030807|T047|65172003|SNOMEDCT_US|PEMPHIGUS |PEMPHIGUS (DISORDER)
C0030807|T047|65172003|SNOMEDCT_US|PEMPHIGUS [DISEASE/FINDING]|PEMPHIGUS (DISORDER)
C0030807|T047|65172003|SNOMEDCT_US|PEMPHIGUS NOS|PEMPHIGUS (DISORDER)
C0030807|T047|65172003|SNOMEDCT_US|PEMPHIGUS |PEMPHIGUS (DISORDER)
C0030807|T047|65172003|SNOMEDCT_US|PEMPHIGUS NOS |PEMPHIGUS (DISORDER)
C0030807|T047|65172003|SNOMEDCT_US|PEMPHIGUS, NOS|PEMPHIGUS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RHEUMATOID ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|ARTHRITIS, RHEUMATOID|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RHEUMATOID ARTHRITIS, UNSPECIFIED|RHEUMATOID ARTHRITIS (DISORDER)
# C0003873|T047|69896004|SNOMEDCT_US|RA|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RA (RHEUMATOID ARTHRITIS)|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RHEUMATOID ARTHRITIS |RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|R ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RH ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|ARTHRITIS, RHEUMATOID [DISEASE/FINDING]|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RHEUMATOID ARTHRITIS NOS |RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RHEUMATOID ARTHRITIS NOS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RHEUMATOID ARTHRITIS |RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|ARTHRITIS RHEUMATOID|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|ATROPHIC ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|SYSTEMIC RHEUMATOID ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|CHRONIC RHEUMATIC ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RHEUMATIC GOUT|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RA - RHEUMATOID ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RHA - RHEUMATOID ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RHEUMATOID DISEASE|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|ATROPHIC; ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RHEUMATOID; ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|ARTHRITIS; ATROPHIC|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|ARTHRITIS; RHEUMATOID|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|ARTHRITIS OR POLYARTHRITIS, ATROPHIC|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|ARTHRITIS OR POLYARTHRITIS, RHEUMATIC|RHEUMATOID ARTHRITIS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|SYSTEMIC LUPUS ERYTHEMATOSIS|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|LUPUS, ERYTHEMATOSUS, SYSTEMIC|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|LUPUS ERYTHEMATOSUS, SYSTEMIC|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|SLE|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|SYSTEMIC LUPUS ERYTHEMATOSUS|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|SYSTEMIC LUPUS ERYTHEMATOSUS, UNSPECIFIED|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|DISSEMINATED LUPUS ERYTHEMATOSUS|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|LUPUS|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|SYSTEMIC LUPUS ERYTHEMATOSUS |SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|SYSTEMIC LUPUS|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|SYST LUPUS ERYTHEMATOSUS|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|SYSTEMIC LUPUS ERYTHEMATOSUS (SLE)|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|SLE NOS|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|SYSTEMIC LUPUS ERYTHEMATOSUS NOS|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|LUPUS ERYTHEMATOSUS DISSEMINATUS|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|LUPUS ERYTHEMATOSUS, SYSTEMIC [DISEASE/FINDING]|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|SYSTEMIC LUPUS ERYTHEMATOSUS NOS |SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|SYSTEMIC LUPUS ERYTHEMATOSUS |SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|LUPUS ERYTHEMATOSIS DISSEMINATED|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|SYNDROME LUPUS|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|LUPUS SYNDROME|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|SYNDROME DISSEMINATED LUPUS ERYTHEMATOSIS|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|LUPUS ERYTHEMATOSUS SYSTEMIC|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|LE SYSTEMIC|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|SYSTEMIC LUPUS ERYTHEMATOSUS SYND|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|LE SYNDROME|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|SLE - SYSTEMIC LUPUS ERYTHEMATOSUS|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|ERYTHEMATOSUS; LUPUS, SYSTEMIC|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|LUPUS; ERYTHEMATOSUS, SYSTEMIC|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|SYSTEM; LUPUS ERYTHEMATOSUS|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0024141|T047|55464009|SNOMEDCT_US|SLE - LUPUS ERYTHEMATOSUS, SYSTEMIC|SYSTEMIC LUPUS ERYTHEMATOSUS (DISORDER)
C0157987|T047|201963008|SNOMEDCT_US|ALLERGIC ARTHRITIS|ALLERGIC ARTHRITIS OF UNSPECIFIED SITE (DISORDER)
C0157987|T047|201963008|SNOMEDCT_US|ALLERGIC ARTHRITIS |ALLERGIC ARTHRITIS OF UNSPECIFIED SITE (DISORDER)
C0157987|T047|201963008|SNOMEDCT_US|ALLERG ARTHRITIS-UNSPEC|ALLERGIC ARTHRITIS OF UNSPECIFIED SITE (DISORDER)
C0157987|T047|201963008|SNOMEDCT_US|ARTHRITIS;ALLERGIC|ALLERGIC ARTHRITIS OF UNSPECIFIED SITE (DISORDER)
C0157987|T047|201963008|SNOMEDCT_US|ALLERGIC ARTHRITIS |ALLERGIC ARTHRITIS OF UNSPECIFIED SITE (DISORDER)
C0157987|T047|201963008|SNOMEDCT_US|ALLERGIC ARTHRITIS NOS |ALLERGIC ARTHRITIS OF UNSPECIFIED SITE (DISORDER)
C0157987|T047|201963008|SNOMEDCT_US|ALLERGIC ARTHRITIS NOS|ALLERGIC ARTHRITIS OF UNSPECIFIED SITE (DISORDER)
C0157987|T047|201963008|SNOMEDCT_US|ALLERGIC ARTHRITIS OF UNSPECIFIED SITE |ALLERGIC ARTHRITIS OF UNSPECIFIED SITE (DISORDER)
C0157987|T047|201963008|SNOMEDCT_US|ALLERGIC ARTHRITIS OF UNSPECIFIED SITE|ALLERGIC ARTHRITIS OF UNSPECIFIED SITE (DISORDER)
C0157987|T047|201963008|SNOMEDCT_US|ALLERGIC ARTHRITIS, SITE UNSPECIFIED|ALLERGIC ARTHRITIS OF UNSPECIFIED SITE (DISORDER)
C0157987|T047|201963008|SNOMEDCT_US|ARTHRITIS ALLERGIC|ALLERGIC ARTHRITIS OF UNSPECIFIED SITE (DISORDER)
C0157987|T047|201963008|SNOMEDCT_US|ARTHRITIS ALLERGIC NOS|ALLERGIC ARTHRITIS OF UNSPECIFIED SITE (DISORDER)
C0157987|T047|201963008|SNOMEDCT_US|ALLERGIC; ARTHRITIS|ALLERGIC ARTHRITIS OF UNSPECIFIED SITE (DISORDER)
C0157987|T047|201963008|SNOMEDCT_US|ARTHRITIS; ALLERGIC|ALLERGIC ARTHRITIS OF UNSPECIFIED SITE (DISORDER)
C0920350|T047|66944004|SNOMEDCT_US|AUTOIMMUNE THYROIDITIDES|AUTOIMMUNE THYROIDITIS (DISORDER)
C0920350|T047|66944004|SNOMEDCT_US|LYMPHOCYTIC THYROIDITIDES|AUTOIMMUNE THYROIDITIS (DISORDER)
C0920350|T047|66944004|SNOMEDCT_US|LYMPHOMATOUS THYROIDITIDES|AUTOIMMUNE THYROIDITIS (DISORDER)
C0920350|T047|66944004|SNOMEDCT_US|LYMPHOMATOUS THYROIDITIS|AUTOIMMUNE THYROIDITIS (DISORDER)
C0920350|T047|66944004|SNOMEDCT_US|THYROIDITIDES, AUTOIMMUNE|AUTOIMMUNE THYROIDITIS (DISORDER)
C0920350|T047|66944004|SNOMEDCT_US|THYROIDITIDES, LYMPHOCYTIC|AUTOIMMUNE THYROIDITIS (DISORDER)
C0920350|T047|66944004|SNOMEDCT_US|THYROIDITIDES, LYMPHOMATOUS|AUTOIMMUNE THYROIDITIS (DISORDER)
C0920350|T047|66944004|SNOMEDCT_US|THYROIDITIS, AUTOIMMUNE|AUTOIMMUNE THYROIDITIS (DISORDER)
C0920350|T047|66944004|SNOMEDCT_US|LYMPHOCYTIC THYROIDITIS|AUTOIMMUNE THYROIDITIS (DISORDER)
C0920350|T047|66944004|SNOMEDCT_US|AUTOIMMUNE THYROIDITIS|AUTOIMMUNE THYROIDITIS (DISORDER)
C0920350|T047|66944004|SNOMEDCT_US|THYROIDITIS, AUTOIMMUNE [DISEASE/FINDING]|AUTOIMMUNE THYROIDITIS (DISORDER)
C0920350|T047|66944004|SNOMEDCT_US|THYROIDITIS, LYMPHOMATOUS|AUTOIMMUNE THYROIDITIS (DISORDER)
C0920350|T047|66944004|SNOMEDCT_US|THYROIDITIS, LYMPHOCYTIC|AUTOIMMUNE THYROIDITIS (DISORDER)
C0920350|T047|66944004|SNOMEDCT_US|THYROIDITIS AUTOIMMUNE|AUTOIMMUNE THYROIDITIS (DISORDER)
C0920350|T047|66944004|SNOMEDCT_US|AUTOIMMUNE THYROIDITIS |AUTOIMMUNE THYROIDITIS (DISORDER)
C0920350|T047|66944004|SNOMEDCT_US|LYMPHOCYTIC THYROIDITIS |AUTOIMMUNE THYROIDITIS (DISORDER)
C0920350|T047|66944004|SNOMEDCT_US|AUTOIMMUNE THYROIDITIS |AUTOIMMUNE THYROIDITIS (DISORDER)
C0920350|T047|66944004|SNOMEDCT_US|AUTOIMMUNE; THYROIDITIS|AUTOIMMUNE THYROIDITIS (DISORDER)
C0920350|T047|66944004|SNOMEDCT_US|THYROIDITIS; AUTOIMMUNE|AUTOIMMUNE THYROIDITIS (DISORDER)
C0920350|T047|66944004|SNOMEDCT_US|AUTOIMMUNE THYROIDITIS, NOS|AUTOIMMUNE THYROIDITIS (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|ANTI PHOSPHOLIPID SYNDROME|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|ANTIPHOSPHOLIPID SYNDROME|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|SYNDROME, ANTI-PHOSPHOLIPID|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|SYNDROME, ANTIPHOSPHOLIPID|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|ANTI PHOSPHOLIPID ANTIBODY SYNDROME|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|ANTIBODY SYNDROME, ANTI-PHOSPHOLIPID|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|ANTIBODY SYNDROME, ANTIPHOSPHOLIPID|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|ANTIPHOSPHOLIPID ANTIBODY SYNDROMES|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|SYNDROME, ANTI-PHOSPHOLIPID ANTIBODY|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|SYNDROME, ANTIPHOSPHOLIPID ANTIBODY|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|ANTIPHOSPHOLIPID SYNDROME |ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|ANTIPHOSPHOLIPID ANTIBODY SYNDROME|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|ANTI-PHOSPHOLIPID SYNDROME|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|ANTIPHOSPHOLIPID SYNDROME [DISEASE/FINDING]|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|ANTI-PHOSPHOLIPID ANTIBODY SYNDROME|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|ANTICARDIOLIPIN SYNDROME|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|ANTIPHOSPHOLIPID SYNDROME |ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|SYNDROME, HUGHES|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|HUGHES SYNDROME|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|APL - ANTIPHOSPHOLIPID SYNDROME|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|APS - ANTIPHOSPHOLIPID SYNDROME|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|SYNDROME; ANTICARDIOLIPIN|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|SYNDROME; ANTIPHOSPHOLIPID|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|ANTICARDIOLIPIN; SYNDROME|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0085278|T047|26843008|SNOMEDCT_US|ANTIPHOSPHOLIPID; SYNDROME|ANTIPHOSPHOLIPID SYNDROME (DISORDER)
C0031036|T047|155441006|SNOMEDCT_US|POLYARTERITIS NODOSA|POLYARTERITIS NODOSA (DISORDER)
C0031036|T047|155441006|SNOMEDCT_US|PERIARTERITIS NODOSA|POLYARTERITIS NODOSA (DISORDER)
C0031036|T047|155441006|SNOMEDCT_US|PANARTERITIS NODOSA |POLYARTERITIS NODOSA (DISORDER)
C0031036|T047|155441006|SNOMEDCT_US|PERIARTERITIS NODOSA |POLYARTERITIS NODOSA (DISORDER)
C0031036|T047|155441006|SNOMEDCT_US|PANARTERITIS NODOSA|POLYARTERITIS NODOSA (DISORDER)
C0031036|T047|155441006|SNOMEDCT_US|POLYARTERITIS NODOSA |POLYARTERITIS NODOSA (DISORDER)
C0031036|T047|155441006|SNOMEDCT_US|PAN|POLYARTERITIS NODOSA (DISORDER)
C0031036|T047|155441006|SNOMEDCT_US|POLYARTERITIS NODOSA [DISEASE/FINDING]|POLYARTERITIS NODOSA (DISORDER)
C0031036|T047|155441006|SNOMEDCT_US|CLASSICAL POLYARTERITIS NODOSA|POLYARTERITIS NODOSA (DISORDER)
C0031036|T047|155441006|SNOMEDCT_US|POLYARTERITIS NODOSA NOS|POLYARTERITIS NODOSA (DISORDER)
C0031036|T047|155441006|SNOMEDCT_US|SYSTEMIC PERIARTERITIS NODOSA|POLYARTERITIS NODOSA (DISORDER)
C0031036|T047|155441006|SNOMEDCT_US|PAN - POLYARTERITIS NODOSA|POLYARTERITIS NODOSA (DISORDER)
C0031036|T047|155441006|SNOMEDCT_US|POLYARTERITIS NODOSA |POLYARTERITIS NODOSA (DISORDER)
C0031036|T047|155441006|SNOMEDCT_US|POLYARTERITIS NODOSA NOS |POLYARTERITIS NODOSA (DISORDER)
C0031036|T047|155441006|SNOMEDCT_US|KUSSMAUL'S DISEASE|POLYARTERITIS NODOSA (DISORDER)
C0031036|T047|155441006|SNOMEDCT_US|CLASSIC POLYARTERITIS NODOSA|POLYARTERITIS NODOSA (DISORDER)
C0031036|T047|155441006|SNOMEDCT_US|POLYARTERITIS NODOSUM|POLYARTERITIS NODOSA (DISORDER)
C0031036|T047|155441006|SNOMEDCT_US|KUSSMAUL; DISEASE|POLYARTERITIS NODOSA (DISORDER)
C0031036|T047|155441006|SNOMEDCT_US|DISEASE; KUSSMAUL|POLYARTERITIS NODOSA (DISORDER)
C0342302|T047|11530004|SNOMEDCT_US|BRITTLE DIABETES|BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|BRITTLE DIABETES MELLITUS |BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|UNSTABLE DIABETES MELLITUS|BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|BRITTLE DIABETES MELLITUS |BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|BRITTLE DIABETES MELLITUS|BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|UNSTABLE DIABETES|BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|UNSTABLE DIABETES MELLITUS |BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|BRITTLE DIABETES MELLITUS |BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|DIABETES BRITTLE|BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|LABILE DIABETES|BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|BRITTLE; DIABETES|BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|DIABETES; BRITTLE|BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|DIABETES; UNSTABLE|BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|UNSTABLE; DIABETES|BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|BRITTLE DIABETES |BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|UNSTABLE DIABETES |BRITTLE DIABETES MELLITUS (FINDING)
C0178468|T047||SNOMEDCT_US|AUTOIMMUNE THYROID DISEASE
C0687719|T047||SNOMEDCT_US|AUTOIMMUNE DISEASE, NOT ELSEWHERE CLASSIFIED
C0687719|T047||SNOMEDCT_US|AUTOIMMUNE DISEASE NEC
C0687719|T047||SNOMEDCT_US|AUTOIMMUNE DISEASE NEC IN ICD9CM
C0409974|T047|200936003|SNOMEDCT_US|LUPUS ERYTHEMATOSUS|LUPUS ERYTHEMATOSUS (DISORDER)
C0409974|T047|200936003|SNOMEDCT_US|LUPUS ERYTHEMATOSIS (NOS)|LUPUS ERYTHEMATOSUS (DISORDER)
C0409974|T047|200936003|SNOMEDCT_US|LUPUS ERYTHEMATOSUS NOS|LUPUS ERYTHEMATOSUS (DISORDER)
C0409974|T047|200936003|SNOMEDCT_US|LUPUS|LUPUS ERYTHEMATOSUS (DISORDER)
C0409974|T047|200936003|SNOMEDCT_US|LUPUS ERYTHEMATOSUS NOS |LUPUS ERYTHEMATOSUS (DISORDER)
C0409974|T047|200936003|SNOMEDCT_US|LE - LUPUS ERYTHEMATOSUS|LUPUS ERYTHEMATOSUS (DISORDER)
C0409974|T047|200936003|SNOMEDCT_US|LUPUS ERYTHEMATOSUS |LUPUS ERYTHEMATOSUS (DISORDER)
C0409974|T047|200936003|SNOMEDCT_US|ERYTHEMATOSUS; LUPUS|LUPUS ERYTHEMATOSUS (DISORDER)
C0409974|T047|200936003|SNOMEDCT_US|LUPUS; ERYTHEMATOSUS|LUPUS ERYTHEMATOSUS (DISORDER)
C0011608|T047|111196000|SNOMEDCT_US|DERMATITIS HERPETIFORMIS|DERMATITIS HERPETIFORMIS (DISORDER)
C0011608|T047|111196000|SNOMEDCT_US|DUHRINGS DISEASE|DERMATITIS HERPETIFORMIS (DISORDER)
C0011608|T047|111196000|SNOMEDCT_US|DISEASE, DUHRING'S|DERMATITIS HERPETIFORMIS (DISORDER)
C0011608|T047|111196000|SNOMEDCT_US|DISEASE, DUHRING|DERMATITIS HERPETIFORMIS (DISORDER)
C0011608|T047|111196000|SNOMEDCT_US|DUHRING DIS|DERMATITIS HERPETIFORMIS (DISORDER)
C0011608|T047|111196000|SNOMEDCT_US|DUHRINGS DIS|DERMATITIS HERPETIFORMIS (DISORDER)
C0011608|T047|111196000|SNOMEDCT_US|DERMATITIS HERPETIFORMIS |DERMATITIS HERPETIFORMIS (DISORDER)
C0011608|T047|111196000|SNOMEDCT_US|DUHRING'S DISEASE|DERMATITIS HERPETIFORMIS (DISORDER)
C0011608|T047|111196000|SNOMEDCT_US|DUHRING DISEASE|DERMATITIS HERPETIFORMIS (DISORDER)
C0011608|T047|111196000|SNOMEDCT_US|DERMATITIS HERPETIFORMIS [DISEASE/FINDING]|DERMATITIS HERPETIFORMIS (DISORDER)
C0011608|T047|111196000|SNOMEDCT_US|DERMATITIS;HERPETIFORMIS|DERMATITIS HERPETIFORMIS (DISORDER)
C0011608|T047|111196000|SNOMEDCT_US|DUHRING-BROCQ DISEASE|DERMATITIS HERPETIFORMIS (DISORDER)
C0011608|T047|111196000|SNOMEDCT_US|DH - DERMATITIS HERPETIFORMIS|DERMATITIS HERPETIFORMIS (DISORDER)
C0011608|T047|111196000|SNOMEDCT_US|DERMATITIS HERPETIFORMIS |DERMATITIS HERPETIFORMIS (DISORDER)
C0011608|T047|111196000|SNOMEDCT_US|DERMATOSIS HERPETIFORMIS|DERMATITIS HERPETIFORMIS (DISORDER)
C0011608|T047|111196000|SNOMEDCT_US|DERMATITIS; HERPETIFORMIS|DERMATITIS HERPETIFORMIS (DISORDER)
C0011608|T047|111196000|SNOMEDCT_US|DERMATOSIS; HERPETIFORMIS|DERMATITIS HERPETIFORMIS (DISORDER)
C0011608|T047|111196000|SNOMEDCT_US|HERPETIFORMIS; DERMATITIS|DERMATITIS HERPETIFORMIS (DISORDER)
C0011608|T047|111196000|SNOMEDCT_US|HERPETIFORMIS; DERMATOSIS|DERMATITIS HERPETIFORMIS (DISORDER)
C0011608|T047|111196000|SNOMEDCT_US|DUHRING|DERMATITIS HERPETIFORMIS (DISORDER)
C0011608|T047|111196000|SNOMEDCT_US|DERMATITIS HERPETIFORMIS [DUP] |DERMATITIS HERPETIFORMIS (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|BERGERS DISEASE|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|GLOMERULONEPHRITIDES, IGA|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|GLOMERULONEPHRITIS, IGA|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|IGA NEPHROPATHY|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|NEPHROPATHY, IMMUNOGLOBULIN A|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|BERGERS DIS|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|BERGER DIS|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|FOCAL GLOMERULONEPHRITIS|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|SEGMENTAL GLOMERULONEPHRITIS|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|IGA GLOMERULONEPHRITIS|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|GLOMERULONEPHRITIS, IGA [DISEASE/FINDING]|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|BERGER DISEASE|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|BERGER'S DISEASE|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|NEPHROPATHY, IGA|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|IMMUNOGLOBULIN A NEPHROPATHY|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|IGA TYPE NEPHRITIS|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|NEPHRITIS, IGA TYPE|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|NEPHROPATHY 1, IGA|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|IGA NEPHROPATHY 1|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|IMMUNOGLOBULIN A NEPHROPATHY |IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|IGA NEPHROPATHY |IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|GLOMERULONEPHRITIS FOCAL|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|NEPHROPATHY IGA|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|IGA NEPHROPATHY |IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|IGAN - IGA NEPHROPATHY|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|IGA; NEPHROPATHY|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|GLOMERULONEPHRITIS; IGA|IGA NEPHROPATHY (DISORDER)
C0017661|T047|236407003|SNOMEDCT_US|NEPHROPATHY; IGA|IGA NEPHROPATHY (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|GRAVES DISEASE|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|BASEDOWS DISEASE|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|DISEASE, BASEDOW|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|EXOPHTHALMIC GOITERS|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|GOITERS, EXOPHTHALMIC|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|DISEASE, BASEDOW'S|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|DISEASE, GRAVES'|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|BASEDOW'S DISEASE|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|EXOPHTHALMIC GOITER|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|BASEDOW DIS|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|BASEDOWS DIS|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|GRAVES DIS|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|GRAVES' DISEASE |GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|GRAVES' DISEASE|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|GRAVES' DISEASE (DIFFUSE TOXIC GOITER)|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|DISEASE GRAVES'|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|GRAVES DISEASE [DISEASE/FINDING]|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|BASEDOW DISEASE|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|GOITER, EXOPHTHALMIC|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|DISEASE;BASEDOWS|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|DISEASE;GRAVES|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|EXOPHTHALMIC GOITRE|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|HYPERTHYROIDISM, AUTOIMMUNE|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|GRAVES' DISEASE |GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|GRAVES' DISEASE - HYPERTHYROIDISM|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|BASEDOW'S DISEASE |GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|MORBUS BASEDOW|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|GOITER EXOPHTHALMIC|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|GRAVES-BASEDOW DISEASE|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|AUTOIMMUNE HYPERTHYROIDISM|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|GOITRE EXOPHTHALMIC|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|GRAVES' DISEASE WITH EXOPHTHALMOS|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|TOXIC DIFFUSE GOITER WITH EXOPHTHALMOS|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|TOXIC DIFFUSE GOITRE WITH EXOPHTHALMOS|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|TOXIC DIFFUSE GOITER WITH EXOPHTHALMOS |GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|FLAJANI|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|GRAVES|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|BASEDOW|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|EXOPHTHALMIC; GOITER|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|EXOPHTHALMOS; GOITER (ETIOLOGY)|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|EXOPHTHALMOS; GOITER (MANIFESTATION)|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|GOITER; EXOPHTHALMOS (ETIOLOGY)|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|GOITER; EXOPHTHALMOS (MANIFESTATION)|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|STRUMA; EXOPHTHALMIC|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|GRAVES' DISEASE [AMBIGUOUS]|GRAVES' DISEASE (DISORDER)
C0018213|T047|353295004|SNOMEDCT_US|DISEASE, GRAVES|GRAVES' DISEASE (DISORDER)
C0029077|T047|75315001|SNOMEDCT_US|SYMPATHETIC OPHTHALMIA|SYMPATHETIC UVEITIS (DISORDER)
C0029077|T047|75315001|SNOMEDCT_US|OPHTHALMIA, SYMPATHETIC|SYMPATHETIC UVEITIS (DISORDER)
C0029077|T047|75315001|SNOMEDCT_US|OPHTHALMIAS, SYMPATHETIC|SYMPATHETIC UVEITIS (DISORDER)
C0029077|T047|75315001|SNOMEDCT_US|SYMPATHETIC OPHTHALMIAS|SYMPATHETIC UVEITIS (DISORDER)
C0029077|T047|75315001|SNOMEDCT_US|SYMPATHETIC UVEITIDES|SYMPATHETIC UVEITIS (DISORDER)
C0029077|T047|75315001|SNOMEDCT_US|UVEITIDES, SYMPATHETIC|SYMPATHETIC UVEITIS (DISORDER)
C0029077|T047|75315001|SNOMEDCT_US|SYMPATHETIC UVEITIS|SYMPATHETIC UVEITIS (DISORDER)
C0029077|T047|75315001|SNOMEDCT_US|SYMPATHETIC UVEITIS |SYMPATHETIC UVEITIS (DISORDER)
C0029077|T047|75315001|SNOMEDCT_US|UVEITIS, SYMPATHETIC|SYMPATHETIC UVEITIS (DISORDER)
C0029077|T047|75315001|SNOMEDCT_US|OPHTHALMIA, SYMPATHETIC [DISEASE/FINDING]|SYMPATHETIC UVEITIS (DISORDER)
C0029077|T047|75315001|SNOMEDCT_US|SYMPATHETIC OPHTHALMITIS|SYMPATHETIC UVEITIS (DISORDER)
C0029077|T047|75315001|SNOMEDCT_US|SYMPATHETIC UVEITIS |SYMPATHETIC UVEITIS (DISORDER)
C0029077|T047|75315001|SNOMEDCT_US|OPHTHALMIA; SYMPATHETIC|SYMPATHETIC UVEITIS (DISORDER)
C0029077|T047|75315001|SNOMEDCT_US|SYMPATHETIC; OPHTHALMIA|SYMPATHETIC UVEITIS (DISORDER)
C0029077|T047|75315001|SNOMEDCT_US|SYMPATHETIC; UVEITIS|SYMPATHETIC UVEITIS (DISORDER)
C0029077|T047|75315001|SNOMEDCT_US|UVEITIS; SYMPATHETIC|SYMPATHETIC UVEITIS (DISORDER)
C0030805|T047|86142006|SNOMEDCT_US|BULLOUS PEMPHIGOID|PEMPHIGOID (DISORDER)
C0030805|T047|86142006|SNOMEDCT_US|PEMPHIGOID|PEMPHIGOID (DISORDER)
C0030805|T047|86142006|SNOMEDCT_US|PEMPHIGOID, BULLOUS|PEMPHIGOID (DISORDER)
C0030805|T047|86142006|SNOMEDCT_US|PEMPHIGOID, UNSPECIFIED|PEMPHIGOID (DISORDER)
C0030805|T047|86142006|SNOMEDCT_US|PEMPHIGOIDS|PEMPHIGOID (DISORDER)
C0030805|T047|86142006|SNOMEDCT_US|PEMPHIGOID |PEMPHIGOID (DISORDER)
C0030805|T047|86142006|SNOMEDCT_US|BULLOUS PEMPHIGOID |PEMPHIGOID (DISORDER)
C0030805|T047|86142006|SNOMEDCT_US|PEMPHIGOID, BULLOUS [DISEASE/FINDING]|PEMPHIGOID (DISORDER)
C0030805|T047|86142006|SNOMEDCT_US|PEMPHIGOID NOS |PEMPHIGOID (DISORDER)
C0030805|T047|86142006|SNOMEDCT_US|PEMPHIGOID NOS|PEMPHIGOID (DISORDER)
C0030805|T047|86142006|SNOMEDCT_US|PEMPHIGOID |PEMPHIGOID (DISORDER)
C0030805|T047|86142006|SNOMEDCT_US|BULLOUS PEMPHIGOID NOS|PEMPHIGOID (DISORDER)
C0030805|T047|86142006|SNOMEDCT_US|BP - BULLOUS PEMPHIGOID|PEMPHIGOID (DISORDER)
C0030805|T047|86142006|SNOMEDCT_US|BULLOUS PEMPHIGOID |PEMPHIGOID (DISORDER)
C0030805|T047|86142006|SNOMEDCT_US|BULLOUS; PEMPHIGOID|PEMPHIGOID (DISORDER)
C0030805|T047|86142006|SNOMEDCT_US|PEMPHIGOID; BULLOUS|PEMPHIGOID (DISORDER)
C0030805|T047|86142006|SNOMEDCT_US|PEMPHIGOID, NOS|PEMPHIGOID (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|GLOMERULONEPHRITIDES, MEMBRANOUS|MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|GLOMERULONEPHRITIS, MEMBRANOUS|MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|GLOMERULONEPHROPATHY, MEMBRANOUS|MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|GLOMERULOPATHY, EXTRAMEMBRANOUS|MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|GLOMERULOPATHY, MEMBRANOUS|MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|MEMBRANOUS GLOMERULONEPHRITIDES|MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|MEMBRANOUS GLOMERULONEPHRITIS|MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|CHRONIC NEPHRITIC SYNDROME, DIFFUSE MEMBRANOUS GLOMERULONEPHRITIS|MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|MEMBRANOUS NEPHROPATHY|MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|MEMBRANOUS GLOMERULONEPHROPATHY|MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|NEPHROPATHY MEMBRANOUS|MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|MEMBRANOUS GLOMERULONEPHRITIS |MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|MEMBRANOUS NEPHROPATHY |MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|GLOMERULONEPHRITIS MEMBRANOUS|MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|CHRONIC NEPHRITIC SYNDROME WITH DIFFUSE MEMBRANOUS GLOMERULONEPHRITIS|MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|MEMBRANOUS GLOMERULOPATHY|MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|GLOMERULONEPHRITIS, MEMBRANOUS [DISEASE/FINDING]|MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|EXTRAMEMBRANOUS GLOMERULOPATHY|MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|NEPHROPATHY, MEMBRANOUS|MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|CHRONIC NEPHRITIC SYNDROME W DIFFUSE MEMBRANOUS GLOMRLNEPH|MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|CHRONIC NEPHRITIC SYNDROME WITH DIFFUSE MEMBRANOUS GLOMERULONEPHRITIS |MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|MEMBRANOUS GLOMERULONEPHRITIS |MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|MGN - MEMBRANOUS GLOMERULONEPHRITIS|MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|CHRONIC NEPHRITIC SYNDROME, DIFFUSE MEMBRANOUS GLOMERULONEPHRITIS |MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|MEMBRANOUS GLOMERULONEPHRITIS NOS|MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0017665|T047|77182004|SNOMEDCT_US|MEMBRANOUS NEPHROPATHY NOS|MEMBRANOUS GLOMERULONEPHRITIS (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|EATON LAMBERT MYASTHENIC SYNDROME|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|EATON LAMBERT SYNDROME|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|LAMBERT EATON MYASTHENIC SYNDROME|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|LAMBERT EATON SYNDROME|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|LAMBERT-EATON MYASTHENIC SYNDROME|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|MYASTHENIC SYNDROME, EATON-LAMBERT|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|SYNDROME, EATON-LAMBERT MYASTHENIC|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|SYNDROME, LAMBERT-EATON|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|SYNDROME, LAMBERT-EATON MYASTHENIC|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|SYNDROME, EATON-LAMBERT|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|EATON-LAMBERT SYNDROME|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|MYOPATHIC MYASTHENIC SYNDROME OF LAMBERT EATON|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|MYASTHENIC MYOPATHIC SYNDROME LAMBERT EATON|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|MYASTHENIC SYNDROME, LAMBERT EATON|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|EATON-LAMBERT SYNDROME |EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|EATON-LAMBERT MYASTHENIC-MYOPATHIC SYNDROME|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|EATON-LAMBERT MYOPATHIC-MYASTHENIC SYNDROME|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|LAMBERT-EATON MYASTHENIC-MYOPATHIC SYNDROME|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|LAMBERT-EATON MYOPATHIC-MYASTHENIC SYNDROME|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|MYOPATHIC-MYASTHENIC SYNDROME OF LAMBERT-EATON|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|LAMBERT-EATON MYASTHENIC SYNDROME [DISEASE/FINDING]|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|MYASTHENIC-MYOPATHIC SYNDROME OF LAMBERT-EATON|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|EATON-LAMBERT MYASTHENIC SYNDROME|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|MYASTHENIC SYNDROME, LAMBERT-EATON|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|LAMBERT-EATON SYNDROME|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|MYOPATHIC-MYASTHENIC SYNDROME OF EATON-LAMBERT|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|MYASTHENIC-MYOPATHIC SYNDROME OF EATON-LAMBERT|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|MYASTHENIC SYNDROME OF LAMBERT EATON|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|LAMBERT-EATON MYASTHENIC-MYOPATHIC SYNDROMES|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|MYASTHENIC MYOPATHIC SYNDROME OF EATON LAMBERT|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|MYASTHENIC MYOPATHIC SYNDROME OF LAMBERT EATON|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|MYOPATHIC MYASTHENIC SYNDROME OF EATON LAMBERT|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|LAMBERT-EATON SYNDROME NOS|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|LAMBERT-EATON MYOPATHIC-MYASTHENIC SYNDROMES|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|EATON-LAMBERT MYOPATHIC-MYASTHENIC SYNDROMES|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|EATON LAMBERT MYASTHENIC SYNDROME |EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|LEMS - LAMBERT-EATON MYASTHENIC SYNDROME|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|MYASTHENIC SYNDROME|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|EATON-LAMBERT SYNDROME |EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|LAMBERT-EATON (ETIOLOGY)|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|LAMBERT-EATON (MANIFESTATION)|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|EATON-LAMBERT (ETIOLOGY)|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0022972|T047|230688006|SNOMEDCT_US|EATON-LAMBERT (MANIFESTATION)|EATON LAMBERT MYASTHENIC SYNDROME (DISORDER)
C0398650|T047|32273002|SNOMEDCT_US|AUTOIMMUNE THROMBOCYTOPENIC PURPURAS|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|DISEASE, WERLHOF|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IDIOPATHIC THROMBOCYTOPENIC PURPURAS|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|PURPURA, AUTOIMMUNE THROMBOCYTOPENIC|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|PURPURA, IDIOPATHIC THROMBOCYTOPENIC|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|PURPURA, THROMBOCYTOPENIC, IDIOPATHIC|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|PURPURAS, AUTOIMMUNE THROMBOCYTOPENIC|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|PURPURAS, IDIOPATHIC THROMBOCYTOPENIC|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|THROMBOCYTOPENIC PURPURA, IDIOPATHIC|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|THROMBOCYTOPENIC PURPURAS, IDIOPATHIC|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|WERLHOFS DISEASE|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|DISEASE, WERLHOF'S|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IDIOPATHIC THROMBOCYTOPENIC PURPURA|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|ITP|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IDIOPATHIC THROMBOCYTOPENIC PURPURA (ITP)|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|THROMBOCYTOPENIC PURPURA, AUTOIMMUNE|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|WERLHOF DIS|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|WERLHOFS DIS|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IMMUNE THROMBOCYTOPENIC PURPURA |ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IMMUNE THROMBOCYTOPENIC PURPURA|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IDIOPATHIC THROMBOCYTOPENIC PURPURA |ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|ITP (IDIOPATHIC THROMBOCYTOPENIC PURPURA)|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|ITP (IMMUNE THROMBOCYTOPENIC PURPURA)|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IDIOPATHIC THROMBOCYTOPENIA PURPURA|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IDIOPATHIC THROMBOCYTOPENIA|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|AITP|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IMMUNE THROMBOCYT PURPRA|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|WERLHOF'S DISEASE|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|PURPURA, THROMBOCYTOPENIC, IDIOPATHIC [DISEASE/FINDING]|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|WERLHOF DISEASE|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|AUTOIMMUNE THROMBOCYTOPENIC PURPURA|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|PURPURA, THROMBOCYTOPENIC, AUTOIMMUNE|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|AUTOIMMUNE THROMBOCYTOPENIA|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IDIOPATHIC PURPURA (& THROMBOCYTOPENIC)|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IDEOPATH THROMBOCYTOPENIC PUR|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IDIOPATHIC PURPURA|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|ITP - IDIOPATHIC THROMBOCYTOPENIC PURPURA|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IDIOPATHIC PURPURA (& THROMBOCYTOPENIC) |ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IMMUNE THROMBOCYTOPENIAS|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|PURPURAS, IMMUNE THROMBOCYTOPENIC|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|THROMBOCYTOPENIC PURPURAS, IMMUNE|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|THROMBOCYTOPENIA, IMMUNE|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|PURPURA, IMMUNE THROMBOCYTOPENIC|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|THROMBOCYTOPENIAS, IMMUNE|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|THROMBOCYTOPENIAS, AUTOIMMUNE|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|THROMBOCYTOPENIC PURPURA, IMMUNE|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|THROMBOCYTOPENIA, AUTOIMMUNE|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IMMUNE THROMBOCYTOPENIC PURPURAS|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|AUTOIMMUNE THROMBOCYTOPENIAS|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IMMUNE THROMBOCYTOPENIA|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|WERLHOF'S SYNDROME|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IDIOPATHIC THROMBOCYTOPENIC PURPURA |ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IMMUNE THROMBOCYTOPENIC PURPURA |ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|FRANK|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|WERLHOF|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IDIOPATHIC; PURPURA|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|PURPURA; IDIOPATHIC|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|PURPURA; THROMBOCYTOPENIC, IDIOPATHIC|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|THROMBOCYTOPENIC; PURPURA, IDIOPATHIC|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|ITP, NOS|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IDIOPATHIC THROMBOCYTOPENIC PURPURA, NOS|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IDIOPATHIC PURPURA, NOS|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0398650|T047|32273002|SNOMEDCT_US|IDIOPATH THROMBOCYTOPENIC PURP|ITP - IMMUNE THROMBOCYTOPENIC PURPURA
C0085409|T047|18947001|SNOMEDCT_US|AUTOIMMUNE POLYENDOCRINOPATHY|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|POLYENDOCRINOPATHIES, AUTOIMMUNE|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|POLYENDOCRINOPATHY, AUTOIMMUNE|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|AUTOIMMUNE POLYGLANDULAR FAILURE|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|LLOYD'S SYNDROME |LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|LLOYD'S SYNDROME|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|POLYENDOCRINE FAILURE SYNDROME |LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|ENDOCRINE LLOYD'S SYNDROME|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|POLYENDOCRINE FAILURE SYNDROME|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|AUTOIMMUNE POLYENDOCRINOPATHY SYNDROME|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|POLYENDOCRINOPATHIES, AUTOIMMUNE [DISEASE/FINDING]|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|AUTOIMMUNE POLYENDOCRINE SYNDROME |LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|AUTOIMMUNE POLYENDOCRINE SYNDROME|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|LLOYD'S SYNDROME |LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|AUTOIMMUNE POLYGLANDULAR FAILURE |LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|PGA|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|APS|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|POLYENDOCRINE AUTOIMMUNITY SYNDROME|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|POLYGLANDULAR AUTOIMMUNE SYNDROME|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|AUTOIMMUNE POLYENDOCRINOPATHY |LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|AUTOIMMUNE POLYGLANDULAR SYNDROME|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|AUTOIMMUNE; POLYGLANDULAR SYNDROME|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|DEFICIENCY; POLYGLANDULAR, AUTOIMMUNE|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|POLYGLANDULAR; DEFICIENCY, AUTOIMMUNE|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|POLYGLANDULAR; SYNDROME, AUTOIMMUNE|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|SYNDROME; AUTOIMMUNE POLYGLANDULAR|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|SYNDROME; POLYGLANDULAR, AUTOIMMUNE|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|AUTOIMMUNE POLYENDOCRINOPATHY, NOS|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|AUTOIMMUNE POLYGLANDULAR SYNDROME, NOS|LLOYD'S SYNDROME (DISORDER)
C0085409|T047|18947001|SNOMEDCT_US|POLYGLANDULAR AUTOIMMUNE SYNDROME, NOS|LLOYD'S SYNDROME (DISORDER)
C0403529|T047|236506009|SNOMEDCT_US|GOODPASTURE'S SYNDROME|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|ANTI GBM DISEASE|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|ANTI-GLOMERULAR BASEMENT MEMBRANE DISEASE|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|SYNDROME, GOODPASTURE'S|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|GOODPASTURES SYNDROME|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|SYNDROME, GOODPASTURE|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|GOODPASTURE SYNDROME|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|ANTI GLOMERULAR BASEMENT MEMBRANE DIS|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|ANTIGBM DISEASE|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|ANTI GBM DIS|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|GOODPASTURE'S SYNDROME |ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|SYNDROME GOOD PASTURE|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|SYNDROME GOOD POSTURES|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|GOODPASTURE DISEASE|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|ANTI-GBM DISEASE|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|ANTI-GLOMERULAR BASEMENT MEMBRANE DISEASE [DISEASE/FINDING]|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|LUNG PURPURA WITH NEPHRITIS|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|ANTI GLOMERULAR BASEMENT MEMBRANE DISEASE|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|GOODPASTURE'S SYNDROME |ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|SYNDROME GOODPASTURE'S|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|PULMONARY-RENAL SYNDROME|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|LUNG PURPURA WITH NEPHRITIS SYNDROME|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|ANTI-GBM NEPHRITIS WITH PULMONARY HEMORRHAGE|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|PULMONARY HEMORRHAGE WITH GLOMERULONEPHRITIS|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|PULMONARY HEMOSIDEROSIS WITH GLOMERULONEPHRITIS|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|ANTI GBM - ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|ANTI-GBM NEPHRITIS WITH PULMONARY HAEMORRHAGE|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|GOODPASTURE'S DISEASE|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|PULMONARY HAEMORRHAGE WITH GLOMERULONEPHRITIS|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|PULMONARY HAEMOSIDEROSIS WITH GLOMERULONEPHRITIS|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|GOODPASTURE'S DISEASE |ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|HAEMORRHAGIC PNEUMONIA AND GLOMERULONEPHRITIS|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|HEMORRHAGIC PNEUMONIA AND GLOMERULONEPHRITIS|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|GOODPASTURE|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|PULMONARY; RENAL SYNDROME (GOODPASTURE)|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|SYNDROME; PULMONARY-RENAL (GOODPASTURE)|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|T047|236506009|SNOMEDCT_US|LUNG PURPURA WITH GLOMERULONEPHRITIS|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0751871|T047||SNOMEDCT_US|NEUROL AUTOIMMUNE DIS
C0751871|T047||SNOMEDCT_US|AUTOIMMUNE DIS NERVOUS SYSTEM
C0751871|T047||SNOMEDCT_US|AUTOIMMUNE NERVOUS SYSTEM DIS
C0751871|T047||SNOMEDCT_US|NERVOUS SYSTEM AUTOIMMUNE DIS
C0751871|T047||SNOMEDCT_US|AUTOIMMUNE DIS NEUROL
C0751871|T047||SNOMEDCT_US|AUTOIMMUNE DISEASES OF THE NERVOUS SYSTEM
C0751871|T047||SNOMEDCT_US|AUTOIMMUNE DISEASE, NEUROLOGIC
C0751871|T047||SNOMEDCT_US|DISEASE, NEUROLOGIC AUTOIMMUNE
C0751871|T047||SNOMEDCT_US|DISEASES, NEUROLOGIC AUTOIMMUNE
C0751871|T047||SNOMEDCT_US|NEUROLOGIC AUTOIMMUNE DISEASE
C0751871|T047||SNOMEDCT_US|AUTOIMMUNE DISEASES, NERVOUS SYSTEM
C0751871|T047||SNOMEDCT_US|NERVOUS SYSTEM AUTOIMMUNE DISEASES
C0751871|T047||SNOMEDCT_US|AUTOIMMUNE DISEASES OF THE NERVOUS SYSTEM [DISEASE/FINDING]
C0751871|T047||SNOMEDCT_US|AUTOIMMUNE DISEASES, NEUROLOGIC
C0751871|T047||SNOMEDCT_US|AUTOIMMUNE NERVOUS SYSTEM DISEASES
C0751871|T047||SNOMEDCT_US|AUTOIMMUNE DISORDERS, NERVOUS SYSTEM
C0751871|T047||SNOMEDCT_US|NEUROLOGIC AUTOIMMUNE DISEASES
C0751871|T047||SNOMEDCT_US|AUTOIMMUNE DISORDERS OF THE NERVOUS SYSTEM
C0751871|T047||SNOMEDCT_US|AUTOIMMUNE NERVOUS SYSTEM DISORDER
C0751871|T047||SNOMEDCT_US|NERVOUS SYSTEM AUTOIMMUNE DISORDERS
C0004364|T047|85828009|SNOMEDCT_US|AUTOIMMUNE DISEASES|AUTOIMMUNE DISEASE (DISORDER)
C0004364|T047|85828009|SNOMEDCT_US|DISEASE, AUTOIMMUNE|AUTOIMMUNE DISEASE (DISORDER)
C0004364|T047|85828009|SNOMEDCT_US|DISEASES, AUTOIMMUNE|AUTOIMMUNE DISEASE (DISORDER)
C0004364|T047|85828009|SNOMEDCT_US|AUTOIMMUNE DISORDER|AUTOIMMUNE DISEASE (DISORDER)
C0004364|T047|85828009|SNOMEDCT_US|AUTOIMMUNITY|AUTOIMMUNE DISEASE (DISORDER)
C0004364|T047|85828009|SNOMEDCT_US|AUTOIMMUNE DISEASE|AUTOIMMUNE DISEASE (DISORDER)
C0004364|T047|85828009|SNOMEDCT_US|AUTOIMMUNE DIS|AUTOIMMUNE DISEASE (DISORDER)
C0004364|T047|85828009|SNOMEDCT_US|SELF RECOGNITION (IMMUNE)|AUTOIMMUNE DISEASE (DISORDER)
C0004364|T047|85828009|SNOMEDCT_US|AUTOIMMUNE DISEASE |AUTOIMMUNE DISEASE (DISORDER)
C0004364|T047|85828009|SNOMEDCT_US|AUTOIMMUNE DISORDERS|AUTOIMMUNE DISEASE (DISORDER)
C0004364|T047|85828009|SNOMEDCT_US|AUTOIMMUNE DISEASE NOS|AUTOIMMUNE DISEASE (DISORDER)
C0004364|T047|85828009|SNOMEDCT_US|AUTOIMMUNE DISEASES [DISEASE/FINDING]|AUTOIMMUNE DISEASE (DISORDER)
C0004364|T047|85828009|SNOMEDCT_US|AUTOIMMUNE DISEASE NOS |AUTOIMMUNE DISEASE (DISORDER)
C0004364|T047|85828009|SNOMEDCT_US|AUTOIMMUNE DISORDER NOS|AUTOIMMUNE DISEASE (DISORDER)
C0004364|T047|85828009|SNOMEDCT_US|AUTOIMMUNE DISEASE |AUTOIMMUNE DISEASE (DISORDER)
C0004364|T047|85828009|SNOMEDCT_US|AUTOIMMUNE DISEASE, NOS|AUTOIMMUNE DISEASE (DISORDER)
C0004364|T047|85828009|SNOMEDCT_US|AUTOIMMUNE DISORDER, NOS|AUTOIMMUNE DISEASE (DISORDER)
C0847092|T047||SNOMEDCT_US|BLOOD AUTOIMMUNE DISORDERS
C0847092|T047||SNOMEDCT_US|AUTOIMMUNE HEMATOLOGIC DISORDER
C0342552|T047|237822008|SNOMEDCT_US|ENDOCRINE AUTOIMMUNE DISORDERS|AUTOIMMUNE ENDOCRINE DISEASE (DISORDER)
C0342552|T047|237822008|SNOMEDCT_US|AUTOIMMUNE ENDOCRINE DISEASE|AUTOIMMUNE ENDOCRINE DISEASE (DISORDER)
C0342552|T047|237822008|SNOMEDCT_US|AUTOIMMUNE ENDOCRINE DISEASE |AUTOIMMUNE ENDOCRINE DISEASE (DISORDER)
C0342552|T047|237822008|SNOMEDCT_US|AUTOIMMUNE ENDOCRINE DISEASE |AUTOIMMUNE ENDOCRINE DISEASE (DISORDER)
C0342552|T047|237822008|SNOMEDCT_US|AUTOIMMUNE ENDOCRINE DISORDER|AUTOIMMUNE ENDOCRINE DISEASE (DISORDER)
C0852003|T047||SNOMEDCT_US|HEPATIC AUTOIMMUNE DISORDERS
C0852004|T047||SNOMEDCT_US|MUSCULAR AUTOIMMUNE DISORDERS
C0852005|T047||SNOMEDCT_US|LUPUS ERYTHEMATOSUS AND ASSOCIATED CONDITIONS
C0851816|T047||SNOMEDCT_US|AUTOIMMUNE DISORDERS NEC
C0852006|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS AND ASSOCIATED CONDITIONS
C0852007|T047||SNOMEDCT_US|SCLERODERMA AND ASSOCIATED DISORDERS
C0949027|T047||SNOMEDCT_US|SKIN AUTOIMMUNE DISORDERS NEC
C0036421|T047|128457007|SNOMEDCT_US|PROGRESSIVE SYSTEMIC SCLEROSIS|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|SCLERODERMA, SYSTEMIC|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|SYSTEMIC SCLEROSIS|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|SYSTEMIC SCLERODERMA|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|SYSTEMIC SCLEROSIS, UNSPECIFIED|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|DIFFUSE SCLEROSIS|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|DIFFUSE SCLERODERMA|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|PSS - PROGRESSIVE SYSTEMIC SCLEROSIS|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|SCLERODERMA, DIFFUSE|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|SCLEROSIS, SYSTEMIC|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|SCLERODERMA, SYSTEMIC [DISEASE/FINDING]|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|SCLERODERMA;PROGRESSIVE|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|PROGRESSIVE SYSTEM SCLEROSIS|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|SCLERODERMA SYNDROME |SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|SCLERODERMA SYNDROME|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|SSC, DIFFUSE SCLEROSIS|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|SS - SYSTEMIC SCLEROSIS|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|SYSTEMIC SCLEROSIS |SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|PSS (PROGRESSIVE SYSTEMIC SCLEROSIS)|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|SCLEROSIS; SYSTEMIC, PROGRESSIVE|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|SCLEROSIS; SYSTEMIC|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|SCLEROSIS; SYSTEM|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|SYSTEM; SCLEROSIS|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|SYSTEMIC; SCLEROSIS, PROGRESSIVE|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|SYSTEMIC; SCLEROSIS|SCLERODERMA SYNDROME (DISORDER)
C0036421|T047|128457007|SNOMEDCT_US|PROGRESSIVE SCLERODERMA|SCLERODERMA SYNDROME (DISORDER)
C2717865|T047||SNOMEDCT_US|PAUCI IMMUNE VASCULITIS
C2717865|T047||SNOMEDCT_US|ANCA ASSOCIATED VASCULITIDES
C2717865|T047||SNOMEDCT_US|VASCULITIS, PAUCI-IMMUNE
C2717865|T047||SNOMEDCT_US|VASCULITIDES, ANCA-ASSOCIATED
C2717865|T047||SNOMEDCT_US|ANTI NEUTROPHIL CYTOPLASMIC ANTIBODY ASSOCIATED VASCULITIS
C2717865|T047||SNOMEDCT_US|VASCULITIS, ANCA-ASSOCIATED
C2717865|T047||SNOMEDCT_US|PAUCI-IMMUNE VASCULITIDES
C2717865|T047||SNOMEDCT_US|VASCULITIDE, ANCA-ASSOCIATED
C2717865|T047||SNOMEDCT_US|VASCULITIDES, PAUCI-IMMUNE
C2717865|T047||SNOMEDCT_US|ANCA-ASSOCIATED VASCULITIDE
C2717865|T047||SNOMEDCT_US|ANCA ASSOCIATED VASCULITIS
C2717865|T047||SNOMEDCT_US|ANTI-NEUTROPHIL CYTOPLASMIC ANTIBODY-ASSOCIATED VASCULITIS
C2717865|T047||SNOMEDCT_US|PAUCI-IMMUNE VASCULITIS
C2717865|T047||SNOMEDCT_US|ANCA-ASSOCIATED VASCULITIDES
C2717865|T047||SNOMEDCT_US|ANCA-ASSOCIATED VASCULITIS
C2717865|T047||SNOMEDCT_US|ANTI-NEUTROPHIL CYTOPLASMIC ANTIBODY-ASSOCIATED VASCULITIS [DISEASE/FINDING]
C1328840|T047|702444009|SNOMEDCT_US|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME (DISORDER)
C1328840|T047|702444009|SNOMEDCT_US|ALPS|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME (DISORDER)
C1328840|T047|702444009|SNOMEDCT_US|AUTOIMMUN LYMPHPROF SYND|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME (DISORDER)
C1328840|T047|702444009|SNOMEDCT_US|LYMPHOPROLIFERATIVE SYNDROMES, AUTOIMMUNE|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME (DISORDER)
C1328840|T047|702444009|SNOMEDCT_US|SYNDROMES, AUTOIMMUNE LYMPHOPROLIFERATIVE|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME (DISORDER)
C1328840|T047|702444009|SNOMEDCT_US|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROMES|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME (DISORDER)
C1328840|T047|702444009|SNOMEDCT_US|LYMPHOPROLIFERATIVE SYNDROME, AUTOIMMUNE|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME (DISORDER)
C1328840|T047|702444009|SNOMEDCT_US|SYNDROME, AUTOIMMUNE LYMPHOPROLIFERATIVE|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME (DISORDER)
C1328840|T047|702444009|SNOMEDCT_US|SYNDROME, CANALE SMITH|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME (DISORDER)
C1328840|T047|702444009|SNOMEDCT_US|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME [ALPS]|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME (DISORDER)
C1328840|T047|702444009|SNOMEDCT_US|CANALE SMITH SYNDROME|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME (DISORDER)
C1328840|T047|702444009|SNOMEDCT_US|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME [DISEASE/FINDING]|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME (DISORDER)
C1328840|T047|702444009|SNOMEDCT_US|SYNDROMES, CANALE-SMITH|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME (DISORDER)
C1328840|T047|702444009|SNOMEDCT_US|CANALE-SMITH SYNDROMES|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME (DISORDER)
C1328840|T047|702444009|SNOMEDCT_US|SYNDROME, CANALE-SMITH|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME (DISORDER)
C1328840|T047|702444009|SNOMEDCT_US|CANALE-SMITH SYNDROME|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME (DISORDER)
C1328840|T047|702444009|SNOMEDCT_US|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME, TYPE I, AUTOSOMAL DOMINANT|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME (DISORDER)
C1328840|T047|702444009|SNOMEDCT_US|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME |AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME (DISORDER)
C1328840|T047|702444009|SNOMEDCT_US|ALPS (AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME)|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANKYLOSING SPONDYLITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|BECHTEREWS DISEASE|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|MARIE STRUEMPELL DISEASE|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLITIS, ANKYLOSING|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLITIS, RHEUMATOID|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|BECHTEREW DIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|MARIE STRUEMPELL DIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|BECHTEREWS DIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANKYLOSING SPONDYLITIS |ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANK SPOND|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLOARTHRITIDES, ANKYLOSING|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANKYLOSING SPONDYLOARTHRITIDES|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLARTHRITIDES, ANKYLOSING|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLARTHRITIS, ANKYLOSING|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLOARTHRITIS, ANKYLOSING|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANKYLOSING SPONDYLARTHRITIDES|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF SPINE|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|RHEUMATOID SPONDYLITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLARTHRITIS ANKYLOPOIETICA|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|BECHTEREW'S DISEASE|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|BECHTEREW DISEASE|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|MARIE-STRUEMPELL DISEASE|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLITIS, ANKYLOSING [DISEASE/FINDING]|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANKYLOSING SPONDYLARTHRITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANKYLOSING SPONDYLOARTHRITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|DISEASE;BECHTEREWS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANKYLOSING SPONDYLITIS |ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLITIS ANKYLOPOIETICA|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLOARTHRITIS ANKYLOPOIETICA|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLITIS ANKYLOSING|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|BEKHTEREV'S DISEASE|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|AS - ANKYLOSING SPONDYLITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|IDIOPATHIC ANKYLOSING SPONDYLITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|MARIE-STRUMPELL SPONDYLITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|MARIE STRÜMPELL SPONDYLITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ARTHRITIS; SPINE OR VERTEBRA, MARIE-STRÜMPELL|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ARTHRITIS; SPINE OR VERTEBRA, ANKYLOSING|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|MARIE-STRÜMPELL; SPONDYLITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|MARIE-STRÜMPELL|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|STRÜMPELL-MARIE|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|VON BECHTEREW|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|BECHTEREW|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|RHEUMATOID; ARTHRITIS, SPINE|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|RHEUMATOID; SPONDYLITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPINE OR VERTEBRA; ARTHRITIS, MARIE-STRÜMPELL|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPINE OR VERTEBRA; ARTHRITIS, ANKYLOSING|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLITIS; MARIE-STRÜMPELL|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLITIS; ANKYLOPOIETICA|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLITIS; ANKYLOSING|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLITIS; RHEUMATOID|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANKYLOPOIETICA; SPONDYLITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANKYLOSING; SPONDYLITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ARTHRITIS; RHEUMATOID, SPINE|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANKYLOSING SPONDYLITIS, NOS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF SPINE, NOS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLITIS, MARIE-STRUMPELL|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|RHEUMATIOID ARTHRITIS OF SPINE NOS|ANKYLOSING SPONDYLITIS (DISORDER)
C0026272|T047|398021003|SNOMEDCT_US|MIXED CONNECTIVE TISSUE DISEASE|CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME (DISORDER)
C0026272|T047|398021003|SNOMEDCT_US|SYNDROME, SHARP|CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME (DISORDER)
C0026272|T047|398021003|SNOMEDCT_US|CONNECTIVE TISSUE DIS MIXED|CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME (DISORDER)
C0026272|T047|398021003|SNOMEDCT_US|MIXED CONNECTIVE TISSUE DIS|CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME (DISORDER)
C0026272|T047|398021003|SNOMEDCT_US|MIXED CONNECTIVE TISSUE DISEASE |CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME (DISORDER)
C0026272|T047|398021003|SNOMEDCT_US|MIXED CONNECTIVE TISSUE DISEASE [DISEASE/FINDING]|CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME (DISORDER)
C0026272|T047|398021003|SNOMEDCT_US|SHARP SYNDROME|CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME (DISORDER)
C0026272|T047|398021003|SNOMEDCT_US|MCTD|CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME (DISORDER)
C0026272|T047|398021003|SNOMEDCT_US|CONNECTIVE TISSUE DISEASE, MIXED|CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME (DISORDER)
C0026272|T047|398021003|SNOMEDCT_US|MIXED COLLAGEN VASCULAR DISEASE |CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME (DISORDER)
C0026272|T047|398021003|SNOMEDCT_US|CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME|CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME (DISORDER)
C0026272|T047|398021003|SNOMEDCT_US|SHARP'S SYNDROME|CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME (DISORDER)
C0026272|T047|398021003|SNOMEDCT_US|MIXED COLLAGEN VASCULAR DISEASE|CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME (DISORDER)
C0026272|T047|398021003|SNOMEDCT_US|MCTD - MIXED CONNECTIVE TISSUE DISEASE|CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME (DISORDER)
C0026272|T047|398021003|SNOMEDCT_US|CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME |CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME (DISORDER)
C0026272|T047|398021003|SNOMEDCT_US|DISEASE (OR DISORDER); MIXED CONNECTIVE TISSUE|CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME (DISORDER)
C0026272|T047|398021003|SNOMEDCT_US|DISEASE (OR DISORDER); MIXED, CONNECTIVE TISSUE|CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME (DISORDER)
C0026272|T047|398021003|SNOMEDCT_US|DISEASE; MIXED CONNECTIVE TISSUE|CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME (DISORDER)
C0026272|T047|398021003|SNOMEDCT_US|MIXED, CONNECTIVE TISSUE; DISORDER|CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME (DISORDER)
C0026272|T047|398021003|SNOMEDCT_US|MIXED COLLAGEN VASCULAR DISEASE, NOS|CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME (DISORDER)
C0026272|T047|398021003|SNOMEDCT_US|MIXED CONNECTIVE TISSUE DISEASE, NOS|CONNECTIVE TISSUE DISEASE OVERLAP SYNDROME (DISORDER)
C2609059|T047|445187004|SNOMEDCT_US|ANTISYNTHETASE SYNDROME|ANTISYNTHETASE SYNDROME (DISORDER)
C2609059|T047|445187004|SNOMEDCT_US|ANTISYNTHETASE SYNDROME |ANTISYNTHETASE SYNDROME (DISORDER)
C0554876|T047||SNOMEDCT_US|POORLY CONTROLLED DIABETES MELLITUS 
C0554876|T047||SNOMEDCT_US|DIABETES MELLITUS POORLY CONTROLLED
C0554876|T047||SNOMEDCT_US|POORLY CONTROLLED DIABETES MELLITUS
C2930824|T047||SNOMEDCT_US|AUTOIMMUNE LIMBIC ENCEPHALITIS
C1260879|T047|400009001|SNOMEDCT_US|AUTOIMMUNE PROGESTERONE DERMATITIS|AUTOIMMUNE PROGESTERONE DERMATITIS/URTICARIA
C1260879|T047|400009001|SNOMEDCT_US|PROGESTERONE DERMATITIS|AUTOIMMUNE PROGESTERONE DERMATITIS/URTICARIA
C1260879|T047|400009001|SNOMEDCT_US|AUTOIMMUNE PROGESTERONE URTICARIA|AUTOIMMUNE PROGESTERONE DERMATITIS/URTICARIA
C1260879|T047|400009001|SNOMEDCT_US|AUTOIMMUNE PROGESTERONE DERMATITIS/URTICARIA |AUTOIMMUNE PROGESTERONE DERMATITIS/URTICARIA
C1260879|T047|400009001|SNOMEDCT_US|AUTOIMMUNE PROGESTERONE DERMATITIS/URTICARIA|AUTOIMMUNE PROGESTERONE DERMATITIS/URTICARIA
C0301928|T047|275446004|SNOMEDCT_US|PSYCHOGENIC PURPURA|GARDNER-DIAMOND SYNDROME (DISORDER)
C0301928|T047|275446004|SNOMEDCT_US|AUTOERYTHROCYTE SENSITIZATION|GARDNER-DIAMOND SYNDROME (DISORDER)
C0301928|T047|275446004|SNOMEDCT_US|GARDNER-DIAMOND SYNDROME|GARDNER-DIAMOND SYNDROME (DISORDER)
C0301928|T047|275446004|SNOMEDCT_US|PAINFUL BRUISING SYNDROME|GARDNER-DIAMOND SYNDROME (DISORDER)
C0301928|T047|275446004|SNOMEDCT_US|AUTOERYTHROCYTE SENSITIVITY DISORDER|GARDNER-DIAMOND SYNDROME (DISORDER)
C0301928|T047|275446004|SNOMEDCT_US|AUTO-ERYTHROCYTE SENSITIZATION|GARDNER-DIAMOND SYNDROME (DISORDER)
C0301928|T047|275446004|SNOMEDCT_US|AUTO-ERYTHROCYTE SENSITISATION|GARDNER-DIAMOND SYNDROME (DISORDER)
C0301928|T047|275446004|SNOMEDCT_US|AUTOERYTHROCYTE SENSITIVITY DISORDER |GARDNER-DIAMOND SYNDROME (DISORDER)
C0301928|T047|275446004|SNOMEDCT_US|AUTOERYTHROCYTE SENSITIVITY|GARDNER-DIAMOND SYNDROME (DISORDER)
C0301928|T047|275446004|SNOMEDCT_US|GARDNER-DIAMOND SYNDROME |GARDNER-DIAMOND SYNDROME (DISORDER)
C0301928|T047|275446004|SNOMEDCT_US|AUTO-ERYTHROCYTE SENSITISATION SYNDROME|GARDNER-DIAMOND SYNDROME (DISORDER)
C0301928|T047|275446004|SNOMEDCT_US|AUTO-ERYTHROCYTE SENSITIZATION SYNDROME|GARDNER-DIAMOND SYNDROME (DISORDER)
C0301928|T047|275446004|SNOMEDCT_US|AUTOERYTHROCYTE SENSITIVITY |GARDNER-DIAMOND SYNDROME (DISORDER)
C0301928|T047|275446004|SNOMEDCT_US|AUTOERYTHROCYTE SENSITIZATION; SYNDROME|GARDNER-DIAMOND SYNDROME (DISORDER)
C0301928|T047|275446004|SNOMEDCT_US|SYNDROME; AUTOERYTHROCYTE SENSITIZATION|GARDNER-DIAMOND SYNDROME (DISORDER)
C0301928|T047|275446004|SNOMEDCT_US|GARDENER-DIAMOND SYNDROME|GARDNER-DIAMOND SYNDROME (DISORDER)
C0301928|T047|275446004|SNOMEDCT_US|AUTOERYTHROCYTE SENSITIVITY DISORDER, NOS|GARDNER-DIAMOND SYNDROME (DISORDER)
C2931429|T047|446682003|SNOMEDCT_US|PEDIATRIC AUTOIMMUNE NEUROPSYCHIATRIC DISORDERS ASSOCIATED WITH STREPTOCOCCAL INFECTIONS|PANDAS - PEDIATRIC AUTOIMMUNE NEUROPSYCHIATRIC DISORDER ASSOCIATED WITH STREPTOCOCCAL INFECTION
C2931429|T047|446682003|SNOMEDCT_US|PANDAS - PAEDIATRIC AUTOIMMUNE NEUROPSYCHIATRIC DISORDER ASSOCIATED WITH STREPTOCOCCAL INFECTION|PANDAS - PEDIATRIC AUTOIMMUNE NEUROPSYCHIATRIC DISORDER ASSOCIATED WITH STREPTOCOCCAL INFECTION
C2931429|T047|446682003|SNOMEDCT_US|PAEDIATRIC AUTOIMMUNE NEUROPSYCHIATRIC DISORDER ASSOCIATED WITH STREPTOCOCCAL INFECTION|PANDAS - PEDIATRIC AUTOIMMUNE NEUROPSYCHIATRIC DISORDER ASSOCIATED WITH STREPTOCOCCAL INFECTION
C2931429|T047|446682003|SNOMEDCT_US|PEDIATRIC AUTOIMMUNE NEUROPSYCHIATRIC DISORDER ASSOCIATED WITH STREPTOCOCCAL INFECTION|PANDAS - PEDIATRIC AUTOIMMUNE NEUROPSYCHIATRIC DISORDER ASSOCIATED WITH STREPTOCOCCAL INFECTION
C2931429|T047|446682003|SNOMEDCT_US|PEDIATRIC AUTOIMMUNE NEUROPSYCHIATRIC DISORDER ASSOCIATED WITH STREPTOCOCCAL INFECTION |PANDAS - PEDIATRIC AUTOIMMUNE NEUROPSYCHIATRIC DISORDER ASSOCIATED WITH STREPTOCOCCAL INFECTION
C2931429|T047|446682003|SNOMEDCT_US|PANDAS - PEDIATRIC AUTOIMMUNE NEUROPSYCHIATRIC DISORDER ASSOCIATED WITH STREPTOCOCCAL INFECTION|PANDAS - PEDIATRIC AUTOIMMUNE NEUROPSYCHIATRIC DISORDER ASSOCIATED WITH STREPTOCOCCAL INFECTION
C2931429|T047|446682003|SNOMEDCT_US|PAEDIATRIC AUTOIMMUNE NEUROPSYCHIATRIC DISORDERS ASSOCIATED WITH STREPTOCOCCAL INFECTION|PANDAS - PEDIATRIC AUTOIMMUNE NEUROPSYCHIATRIC DISORDER ASSOCIATED WITH STREPTOCOCCAL INFECTION
C2931429|T047|446682003|SNOMEDCT_US|PEDIATRIC AUTOIMMUNE NEUROPSYCHIATRIC DISORDERS ASSOCIATED WITH STREPTOCOCCAL INFECTION|PANDAS - PEDIATRIC AUTOIMMUNE NEUROPSYCHIATRIC DISORDER ASSOCIATED WITH STREPTOCOCCAL INFECTION
C2931429|T047|446682003|SNOMEDCT_US|PANDAS|PANDAS - PEDIATRIC AUTOIMMUNE NEUROPSYCHIATRIC DISORDER ASSOCIATED WITH STREPTOCOCCAL INFECTION
C0341305|T047|235728001|SNOMEDCT_US|AUTOIMMUNE ENTEROPATHY|AUTOIMMUNE ENTEROPATHY (DISORDER)
C0341305|T047|235728001|SNOMEDCT_US|AUTOIMMUNE ENTEROPATHY |AUTOIMMUNE ENTEROPATHY (DISORDER)
C0406650|T047|95330001|SNOMEDCT_US|LINEAR IGA DISEASE|LINEAR IGA DERMATOSIS (DISORDER)
C0406650|T047|95330001|SNOMEDCT_US|LINEAR IGA DERMATOSES |LINEAR IGA DERMATOSIS (DISORDER)
C0406650|T047|95330001|SNOMEDCT_US|LINEAR IGA DERMATOSES|LINEAR IGA DERMATOSIS (DISORDER)
C0406650|T047|95330001|SNOMEDCT_US|LINEAR IGA DERMATOSIS|LINEAR IGA DERMATOSIS (DISORDER)
C0406650|T047|95330001|SNOMEDCT_US|IGA DERMATOSES, LINEAR|LINEAR IGA DERMATOSIS (DISORDER)
C0406650|T047|95330001|SNOMEDCT_US|LINEAR IGA BULLOUS DERMATOSIS|LINEAR IGA DERMATOSIS (DISORDER)
C0406650|T047|95330001|SNOMEDCT_US|DERMATOSIS, LINEAR IGA|LINEAR IGA DERMATOSIS (DISORDER)
C0406650|T047|95330001|SNOMEDCT_US|IGA DERMATOSIS, LINEAR|LINEAR IGA DERMATOSIS (DISORDER)
C0406650|T047|95330001|SNOMEDCT_US|DERMATOSES, LINEAR IGA|LINEAR IGA DERMATOSIS (DISORDER)
C0406650|T047|95330001|SNOMEDCT_US|LINEAR IGA BULLOUS DERMATOSIS [DISEASE/FINDING]|LINEAR IGA DERMATOSIS (DISORDER)
C0406650|T047|95330001|SNOMEDCT_US|LINEAR IMMUNOGLOBULIN A DERMATOSIS |LINEAR IGA DERMATOSIS (DISORDER)
C0406650|T047|95330001|SNOMEDCT_US|LINEAR IGA DERMATOSIS |LINEAR IGA DERMATOSIS (DISORDER)
C0406650|T047|95330001|SNOMEDCT_US|LINEAR IMMUNOGLOBULIN A DERMATOSIS|LINEAR IGA DERMATOSIS (DISORDER)
C0406650|T047|95330001|SNOMEDCT_US|LINEAR IGA|LINEAR IGA DERMATOSIS (DISORDER)
C0406650|T047|95330001|SNOMEDCT_US|LINEAR IG A DISEASE|LINEAR IGA DERMATOSIS (DISORDER)
C0406650|T047|95330001|SNOMEDCT_US|IGA - LINEAR IMMUNOGLOBULIN A BULLOUS DERMATOSIS|LINEAR IGA DERMATOSIS (DISORDER)
C0406650|T047|95330001|SNOMEDCT_US|LAD - LINEAR IGA DISEASE|LINEAR IGA DERMATOSIS (DISORDER)
C0406650|T047|95330001|SNOMEDCT_US|LINEAR IMMUNOGLOBULIN A BULLOUS DERMATOSIS|LINEAR IGA DERMATOSIS (DISORDER)
C0342340|T047|190454008|SNOMEDCT_US|AUTOIMMUNE PARATHYROIDITIS|AUTOIMMUNE PARATHYROIDITIS (DISORDER)
C0342340|T047|190454008|SNOMEDCT_US|AUTOIMMUNE PARATHYROIDITIS |AUTOIMMUNE PARATHYROIDITIS (DISORDER)
C0034152|T047|246074004|SNOMEDCT_US|PURPURA, SCHOENLEIN HENOCH|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURA, SCHOENLEIN-HENOCH|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|SCHOENLEIN HENOCH PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|ALLERGIC PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|HENOCH-SCHONLEIN PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURA, ALLERGIC|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURA, ANAPHYLACTOID|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|HENOCH-SCHOENLEIN PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|HENOCH-SCHONLEIN PURPURA |HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|ANAPHYLACTOID PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURA, HENOCH|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|HENOCH-SCHOLEIN PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|HENOCH-SCH@NLEIN PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|ALLERGIC PURPURA |HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|ALLERGIC VASCULAR PURPURA |HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|HENOCH SCHOENLEIN PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURA, HENOCH-SCHOENLEIN|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|ALLERGIC VASCULAR PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|HENOCH SCHONLEIN PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|HENOCH SCHONLEIN PURPURA |HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|VASCULAR ALLERGIC PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURAS, SCHONLEIN-HENOCH|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|SCHONLEIN-HENOCH PURPURAS|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURAS, HENOCH-SCHONLEIN|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|HENOCH SCHONLEIN PURPURAS|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURA, SCHONLEIN HENOCH|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|HENOCH-SCHONLEIN PURPURAS|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURA, HENOCH SCHONLEIN|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|SCHONLEIN PURPURA, HENOCH|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|SCHONLEIN PURPURAS, HENOCH|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|SCHONLEIN-HENOCH PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURAS, HENOCH SCHONLEIN|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURA, HENOCH-SCHONLEIN|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|SCHOENLEIN-HENOCH PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURA HENOCH(-SCHÖNLEIN)|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURA ANAPHYLACTOID|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURA, SCHOENLEIN-HENOCH [DISEASE/FINDING]|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|HENOCH PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURA, SCHONLEIN-HENOCH|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|HENOCH-SCH?NLEIN PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|AUTOIMMUNE PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|ALLERGIC PURPURA |HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|AUTOIMMUNE PURPURA |HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|HENOCH-SCHONLEIN ALL. PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|ALLERGIC PURPURA NOS |HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURA: [ALLERGIC] OR [HENOCH-SCHONLEIN ALLERGY]|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURA: [ALLERGIC] OR [HENOCH-SCHONLEIN ALLERGY] |HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|HENOCH-SCH?NLEIN PURPURA |HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|ALLERGIC PURPURA NOS|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|ANAPHYLACTIC VASCULAR PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURA ALLERGIC|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURA VASCULAR ALLERGIC|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|ANAPHYLACTOID VASCULAR PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|HENOCH-SCHONLEIN|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|HENOCH SHONLEIN PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|HSP|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|HENOCH'S PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|ACUTE VASCULAR PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|HENOCH-SCHOENLEIN VASCULITIS|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|SPRING FEVER|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|HSP - HENOCH-SCHONLEIN PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|SCHÖNLEIN; PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|SCHÖNLEIN|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|ALLERGIC; PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURA; SCHÖNLEIN|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURA; ALLERGIC|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURA; ANAPHYLACTOID|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|ANAPHYLACTOID; PURPURA|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|AUTOIMMUNE PURPURA  [AMBIGUOUS]|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURA, AUTOIMMUNE|HENOCH-SCH?NLEIN PURPURA
C0034152|T047|246074004|SNOMEDCT_US|PURPURA;HENOCH-SCHONLEIN|HENOCH-SCH?NLEIN PURPURA
C0272177|T047|111585004|SNOMEDCT_US|NEUTROPENIA ASSOCIATED WITH AUTOIMMUNE DISEASE|NEUTROPENIA ASSOCIATED WITH AUTOIMMUNE DISEASE (DISORDER)
C0272177|T047|111585004|SNOMEDCT_US|NEUTROPENIA ASSOCIATED WITH AUTOIMMUNE DISEASE |NEUTROPENIA ASSOCIATED WITH AUTOIMMUNE DISEASE (DISORDER)
C0272177|T047|111585004|SNOMEDCT_US|NEUTROPENIA ASSOCIATED WITH AUTOIMMUNE DISEASE |NEUTROPENIA ASSOCIATED WITH AUTOIMMUNE DISEASE (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|CHRONIC ARTHRITIS, JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|RHEUMATOID ARTHRITIS, JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE ARTHRITIS|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE ARTHRITIS, UNSPECIFIED|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ARTHRITIS, JUVENILE CHRONIC|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE IDIOPATHIC ARTHRITIS|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE CHRONIC ARTHRITIS|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE RHEUMATOID ARTHRITIS|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ARTHRITIS, JUVENILE IDIOPATHIC|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE ARTHRITIS |JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ARTHRITIS, JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ENTHESITIS RELATED ARTHRITIS, JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE OLIGOARTHRITIS|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ARTHRITIS, JUVENILE SYSTEMIC|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE ENTHESITIS-RELATED ARTHRITIS|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE SYSTEMIC ARTHRITIS|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ARTHRITIS, JUVENILE PSORIATIC|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE PSORIATIC ARTHRITIS|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ARTHRITIS, JUVENILE ENTHESITIS-RELATED|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|OLIGOARTHRITIS, JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ARTHRITIS, JUVENILE RHEUMATOID|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ENTHESITIS-RELATED ARTHRITIS, JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|PSORIATIC ARTHRITIS, JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|SYSTEMIC ARTHRITIS, JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ARTHRITIS, JUVENILE [DISEASE/FINDING]|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JIA|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|POLYARTHRITIS, JUVENILE, RHEUMATOID FACTOR POSITIVE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|POLYARTHRITIS, JUVENILE, RHEUMATOID FACTOR NEGATIVE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JCA - JUVENILE CHRONIC ARTHRITIS|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE CHRONIC ARTHRITIS |JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE; ARTHRITIS|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ARTHRITIS; JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE CHRONIC ARTHRITIS, POLYARTICULAR SEROPOSITIVE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE IDIOPATHIC ARTHRITIS |JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE IDIOPATHIC ARTHRITIS, POLYARTHRITIS, RHEUMATOID FACTOR POSITIVE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|IDIOPATHIC ARTHRITIS, JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ARTHRITIS;JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C2732697|T047|443899007|SNOMEDCT_US|AUTOIMMUNE INFLAMMATION OF SKELETAL MUSCLE |AUTOIMMUNE INFLAMMATION OF SKELETAL MUSCLE (DISORDER)
C2732697|T047|443899007|SNOMEDCT_US|AUTOIMMUNE INFLAMMATION OF SKELETAL MUSCLE|AUTOIMMUNE INFLAMMATION OF SKELETAL MUSCLE (DISORDER)
C2732697|T047|443899007|SNOMEDCT_US|AUTOIMMUNE MYOSITIS|AUTOIMMUNE INFLAMMATION OF SKELETAL MUSCLE (DISORDER)
C1328843|T047|427213005|SNOMEDCT_US|AUTOIMMUNE VASCULITIS|AUTOIMMUNE VASCULITIS (DISORDER)
C1328843|T047|427213005|SNOMEDCT_US|AUTOIMMUNE VASCULITIS |AUTOIMMUNE VASCULITIS (DISORDER)
C1328843|T047|427213005|SNOMEDCT_US|IMMUNE MEDIATED VASCULITIS|AUTOIMMUNE VASCULITIS (DISORDER)
C2609129|T047|448542008|SNOMEDCT_US|AUTOIMMUNE PANCREATITIS|AUTOIMMUNE PANCREATITIS (DISORDER)
C2609129|T047|448542008|SNOMEDCT_US|AUTOIMMUNE PANCREATITIS |AUTOIMMUNE PANCREATITIS (DISORDER)
C0456037|T047|276575001|SNOMEDCT_US|ANT - AUTOIMMUNE NEONATAL THROMBOCYTOPENIA|AUTOIMMUNE NEONATAL THROMBOCYTOPENIA (DISORDER)
C0456037|T047|276575001|SNOMEDCT_US|AUTOIMMUNE NEONATAL THROMBOCYTOPENIA|AUTOIMMUNE NEONATAL THROMBOCYTOPENIA (DISORDER)
C0456037|T047|276575001|SNOMEDCT_US|AUTOIMMUNE NEONATAL THROMBOCYTOPENIA |AUTOIMMUNE NEONATAL THROMBOCYTOPENIA (DISORDER)
C0342337|T047|237652003|SNOMEDCT_US|INSULIN RESISTANCE - TYPE B|INSULIN RESISTANCE - TYPE B (DISORDER)
C0342337|T047|237652003|SNOMEDCT_US|INSULIN RESISTANCE - TYPE B |INSULIN RESISTANCE - TYPE B (DISORDER)
C0400936|T047|235890007|SNOMEDCT_US|AUTOIMMUNE LIVER DISEASE|AUTOIMMUNE LIVER DISEASE (DISORDER)
C0400936|T047|235890007|SNOMEDCT_US|AUTOIMMUNE LIVER DISEASE |AUTOIMMUNE LIVER DISEASE (DISORDER)
C1970472|T047|707443007|SNOMEDCT_US|PULMONARY ALVEOLAR PROTEINOSIS, ACQUIRED|AUTOIMMUNE PULMONARY ALVEOLAR PROTEINOSIS
C1970472|T047|707443007|SNOMEDCT_US|PULMONARY ALVEOLAR LIPOPROTEINOSIS, ACQUIRED|AUTOIMMUNE PULMONARY ALVEOLAR PROTEINOSIS
C1970472|T047|707443007|SNOMEDCT_US|PULMONARY ALVEOLAR PROTEINOSIS, AUTOIMMUNE|AUTOIMMUNE PULMONARY ALVEOLAR PROTEINOSIS
C1970472|T047|707443007|SNOMEDCT_US|AUTOIMMUNE PULMONARY ALVEOLAR PROTEINOSIS |AUTOIMMUNE PULMONARY ALVEOLAR PROTEINOSIS
C1970472|T047|707443007|SNOMEDCT_US|AUTOIMMUNE PULMONARY ALVEOLAR PROTEINOSIS|AUTOIMMUNE PULMONARY ALVEOLAR PROTEINOSIS
C1970472|T047|707443007|SNOMEDCT_US|PAP, ACQUIRED|AUTOIMMUNE PULMONARY ALVEOLAR PROTEINOSIS
C1842763|T047|703523004|SNOMEDCT_US|SPONDYLOENCHONDRODYSPLASIA WITH IMMUNE DYSREGULATION|SPONDYLOENCHONDRODYSPLASIA WITH IMMUNE DYSREGULATION (DISORDER)
C1842763|T047|703523004|SNOMEDCT_US|SPENCDI|SPONDYLOENCHONDRODYSPLASIA WITH IMMUNE DYSREGULATION (DISORDER)
C1842763|T047|703523004|SNOMEDCT_US|COMBINED IMMUNODEFICIENCY WITH AUTOIMMUNITY AND SPONDYLOMETAPHYSEAL DYSPLASIA|SPONDYLOENCHONDRODYSPLASIA WITH IMMUNE DYSREGULATION (DISORDER)
C1842763|T047|703523004|SNOMEDCT_US|SPONDYLOENCHONDRODYSPLASIA WITH IMMUNE DYSREGULATION |SPONDYLOENCHONDRODYSPLASIA WITH IMMUNE DYSREGULATION (DISORDER)
C1842763|T047|703523004|SNOMEDCT_US|ROIFMAN-MELAMED SYNDROME|SPONDYLOENCHONDRODYSPLASIA WITH IMMUNE DYSREGULATION (DISORDER)
C1842763|T047|703523004|SNOMEDCT_US|ROIFMAN-COSTA SYNDROME|SPONDYLOENCHONDRODYSPLASIA WITH IMMUNE DYSREGULATION (DISORDER)
C0272137|T047|40387008|SNOMEDCT_US|GALACTOSYLTRANSFERASE DEFICIENCY|POLYAGGLUTINABLE ERYTHROCYTE SYNDROME (DISORDER)
C0272137|T047|40387008|SNOMEDCT_US|TN SYNDROME|POLYAGGLUTINABLE ERYTHROCYTE SYNDROME (DISORDER)
C0272137|T047|40387008|SNOMEDCT_US|TN POLYAGGLUTINATION SYNDROME|POLYAGGLUTINABLE ERYTHROCYTE SYNDROME (DISORDER)
C0272137|T047|40387008|SNOMEDCT_US|TNPS|POLYAGGLUTINABLE ERYTHROCYTE SYNDROME (DISORDER)
C0272137|T047|40387008|SNOMEDCT_US|POLYAGGLUTINABLE ERYTHROCYTE SYNDROME|POLYAGGLUTINABLE ERYTHROCYTE SYNDROME (DISORDER)
C0272137|T047|40387008|SNOMEDCT_US|POLYAGGLUTINABLE ERYTHROCYTE SYNDROME |POLYAGGLUTINABLE ERYTHROCYTE SYNDROME (DISORDER)
C1835931|T047||SNOMEDCT_US|ALPHA/BETA T-CELL LYMPHOPENIA WITH GAMMA/DELTA T-CELL EXPANSION, SEVERE CYTOMEGALOVIRUS INFECTION, AND AUTOIMMUNITY
C1835931|T047||SNOMEDCT_US|ALPHA-BETA T-CELL LYMPHOPENIA WITH GAMMA-DELTA T-CELL EXPANSION, SEVERE CYTOMEGALOVIRUS INFECTION, AND AUTOIMMUNITY
C1857958|T047||SNOMEDCT_US|DIABETES MELLITUS, CONGENITAL AUTOIMMUNE
C0026103|T047|7826003|SNOMEDCT_US|MIKULICZ'S DISEASE|MIKULICZ'S DISEASE (DISORDER)
C0026103|T047|7826003|SNOMEDCT_US|MIKULICZ'S SYNDROME|MIKULICZ'S DISEASE (DISORDER)
C0026103|T047|7826003|SNOMEDCT_US|DISEASE, MIKULICZ|MIKULICZ'S DISEASE (DISORDER)
C0026103|T047|7826003|SNOMEDCT_US|DISEASE, MIKULICZ'|MIKULICZ'S DISEASE (DISORDER)
C0026103|T047|7826003|SNOMEDCT_US|MIKULICZ' DISEASE|MIKULICZ'S DISEASE (DISORDER)
C0026103|T047|7826003|SNOMEDCT_US|MIKULICZ DIS|MIKULICZ'S DISEASE (DISORDER)
C0026103|T047|7826003|SNOMEDCT_US|MIKULICZ'S DISEASE |MIKULICZ'S DISEASE (DISORDER)
C0026103|T047|7826003|SNOMEDCT_US|MIKULICZ DISEASE|MIKULICZ'S DISEASE (DISORDER)
C0026103|T047|7826003|SNOMEDCT_US|MIKULICZ' DISEASE [DISEASE/FINDING]|MIKULICZ'S DISEASE (DISORDER)
C0026103|T047|7826003|SNOMEDCT_US|MIKULICZ SYNDROME|MIKULICZ'S DISEASE (DISORDER)
C0026103|T047|7826003|SNOMEDCT_US|MIKULICZ'S DISEASE |MIKULICZ'S DISEASE (DISORDER)
C0026103|T047|7826003|SNOMEDCT_US|MIKULICZ|MIKULICZ'S DISEASE (DISORDER)
C2717757|T047|702575003|SNOMEDCT_US|SYNDROME, SUSAC|RETINOCOCHLEOCEREBRAL VASCULOPATHY (DISORDER)
C2717757|T047|702575003|SNOMEDCT_US|SUSACS SYNDROME|RETINOCOCHLEOCEREBRAL VASCULOPATHY (DISORDER)
C2717757|T047|702575003|SNOMEDCT_US|VASCULOPATHIES, RETINOCOCHLEOCEREBRAL|RETINOCOCHLEOCEREBRAL VASCULOPATHY (DISORDER)
C2717757|T047|702575003|SNOMEDCT_US|RETINOCOCHLEOCEREBRAL VASCULOPATHIES|RETINOCOCHLEOCEREBRAL VASCULOPATHY (DISORDER)
C2717757|T047|702575003|SNOMEDCT_US|SYNDROME, SUSAC'S|RETINOCOCHLEOCEREBRAL VASCULOPATHY (DISORDER)
C2717757|T047|702575003|SNOMEDCT_US|SUSAC SYNDROME|RETINOCOCHLEOCEREBRAL VASCULOPATHY (DISORDER)
C2717757|T047|702575003|SNOMEDCT_US|VASCULOPATHY, RETINOCOCHLEOCEREBRAL|RETINOCOCHLEOCEREBRAL VASCULOPATHY (DISORDER)
C2717757|T047|702575003|SNOMEDCT_US|SUSAC SYNDROME [DISEASE/FINDING]|RETINOCOCHLEOCEREBRAL VASCULOPATHY (DISORDER)
C2717757|T047|702575003|SNOMEDCT_US|RETINOCOCHLEOCEREBRAL VASCULOPATHY|RETINOCOCHLEOCEREBRAL VASCULOPATHY (DISORDER)
C2717757|T047|702575003|SNOMEDCT_US|SUSAC'S SYNDROME|RETINOCOCHLEOCEREBRAL VASCULOPATHY (DISORDER)
C2717757|T047|702575003|SNOMEDCT_US|RETINOCOCHLEOCEREBRAL VASCULOPATHY |RETINOCOCHLEOCEREBRAL VASCULOPATHY (DISORDER)
C0409999|T047|239918008|SNOMEDCT_US|UNDIFFERENTIATED CONNECTIVE TISSUE DISEASE|UNDIFFERENTIATED CONNECTIVE TISSUE DISEASE (DISORDER)
C0409999|T047|239918008|SNOMEDCT_US|UCTD|UNDIFFERENTIATED CONNECTIVE TISSUE DISEASE (DISORDER)
C0409999|T047|239918008|SNOMEDCT_US|UNDIFFERENTIATED CONNECTIVE TISSUE DISEASE |UNDIFFERENTIATED CONNECTIVE TISSUE DISEASE (DISORDER)
C1861303|T047|726078000|SNOMEDCT_US|ACUG|EARLY ONSET SARCOIDOSIS
C1861303|T047|726078000|SNOMEDCT_US|SYNOVITIS, GRANULOMATOUS, WITH UVEITIS AND CRANIAL NEUROPATHIES |EARLY ONSET SARCOIDOSIS
C1861303|T047|726078000|SNOMEDCT_US|SYNOVITIS, GRANULOMATOUS, WITH UVEITIS AND CRANIAL NEUROPATHIES|EARLY ONSET SARCOIDOSIS
C1861303|T047|726078000|SNOMEDCT_US|BLAU SYNDROME|EARLY ONSET SARCOIDOSIS
C1861303|T047|726078000|SNOMEDCT_US|GRANULOMATOUS INFLAMMATORY ARTHRITIS, DERMATITIS, AND UVEITIS, FAMILIAL|EARLY ONSET SARCOIDOSIS
C1861303|T047|726078000|SNOMEDCT_US|GRANULOMATOSIS, FAMILIAL, BLAU TYPE|EARLY ONSET SARCOIDOSIS
C1861303|T047|726078000|SNOMEDCT_US|ARTHROCUTANEOUVEAL GRANULOMATOSIS|EARLY ONSET SARCOIDOSIS
C1861303|T047|726078000|SNOMEDCT_US|GRANULOMATOSIS, FAMILIAL JUVENILE SYSTEMIC|EARLY ONSET SARCOIDOSIS
C1861303|T047|726078000|SNOMEDCT_US|JABS SYNDROME|EARLY ONSET SARCOIDOSIS
C1861303|T047|726078000|SNOMEDCT_US|FAMILIAL GRANULOMATOSIS, BLAU TYPE|EARLY ONSET SARCOIDOSIS
C1861303|T047|726078000|SNOMEDCT_US|ARTHROCUTANEOUVEAL GRANULAMOTOSIS|EARLY ONSET SARCOIDOSIS
C1861303|T047|726078000|SNOMEDCT_US|GRANULOMATOUS INFLAMMATORY ARTHRITIS, DERMATITIS AND UVEITIS, FAMILIAL|EARLY ONSET SARCOIDOSIS
C1861303|T047|726078000|SNOMEDCT_US|FAMILIAL JUVENILE SYSTEMIC GRANULOMATOSIS|EARLY ONSET SARCOIDOSIS
C1861303|T047|726078000|SNOMEDCT_US|EARLY ONSET SARCOIDOSIS|EARLY ONSET SARCOIDOSIS
C1861303|T047|726078000|SNOMEDCT_US|PEDIATRIC GRANULOMATOUS ARTHRITIS|EARLY ONSET SARCOIDOSIS
C1861303|T047|726078000|SNOMEDCT_US|FAMILIAL GRANULOMATOUS INFLAMMATORY ARTHRITIS, DERMATITIS AND UVEITIS |EARLY ONSET SARCOIDOSIS
C1861303|T047|726078000|SNOMEDCT_US|FAMILIAL GRANULOMATOUS INFLAMMATORY ARTHRITIS, DERMATITIS AND UVEITIS|EARLY ONSET SARCOIDOSIS
C1861303|T047|726078000|SNOMEDCT_US|EARLY-ONSET SARCOIDOSIS|EARLY ONSET SARCOIDOSIS
C1861303|T047|726078000|SNOMEDCT_US|BLAUS|EARLY ONSET SARCOIDOSIS
C1861303|T047|726078000|SNOMEDCT_US|SYNOVITIS GRANULOMATOUS WITH UVEITIS AND CRANIAL NEUROPATHIES|EARLY ONSET SARCOIDOSIS
C0410000|T047|276657008|SNOMEDCT_US|OVERLAP SYNDROME|OVERLAP SYNDROME (DISORDER)
C0410000|T047|276657008|SNOMEDCT_US|OVERLAP SYNDROME |OVERLAP SYNDROME (DISORDER)
C0393799|T047|193175006|SNOMEDCT_US|MILLER FISHER SYNDROME|MILLER-FISHER VARIANT OF GUILLAIN-BARRE SYNDROME (DISORDER)
C0393799|T047|193175006|SNOMEDCT_US|SYNDROME, FISHER|MILLER-FISHER VARIANT OF GUILLAIN-BARRE SYNDROME (DISORDER)
C0393799|T047|193175006|SNOMEDCT_US|SYNDROME, MILLER FISHER|MILLER-FISHER VARIANT OF GUILLAIN-BARRE SYNDROME (DISORDER)
C0393799|T047|193175006|SNOMEDCT_US|SYNDROME, MILLER-FISHER|MILLER-FISHER VARIANT OF GUILLAIN-BARRE SYNDROME (DISORDER)
C0393799|T047|193175006|SNOMEDCT_US|MILLER-FISHER SYNDROME |MILLER-FISHER VARIANT OF GUILLAIN-BARRE SYNDROME (DISORDER)
C0393799|T047|193175006|SNOMEDCT_US|MILLER-FISHER SYNDROME|MILLER-FISHER VARIANT OF GUILLAIN-BARRE SYNDROME (DISORDER)
C0393799|T047|193175006|SNOMEDCT_US|FISHER SYNDROME|MILLER-FISHER VARIANT OF GUILLAIN-BARRE SYNDROME (DISORDER)
C0393799|T047|193175006|SNOMEDCT_US|GUILLAIN-BARRE SYNDROME, MILLER FISHER VARIANT|MILLER-FISHER VARIANT OF GUILLAIN-BARRE SYNDROME (DISORDER)
C0393799|T047|193175006|SNOMEDCT_US|MILLER FISHER SYNDROME [DISEASE/FINDING]|MILLER-FISHER VARIANT OF GUILLAIN-BARRE SYNDROME (DISORDER)
C0393799|T047|193175006|SNOMEDCT_US|MILLER FISHER VARIANT OF GUILLAIN BARRE SYNDROME|MILLER-FISHER VARIANT OF GUILLAIN-BARRE SYNDROME (DISORDER)
C0393799|T047|193175006|SNOMEDCT_US|GUILLAIN BARRE SYNDROME, MILLER FISHER VARIANT|MILLER-FISHER VARIANT OF GUILLAIN-BARRE SYNDROME (DISORDER)
C0393799|T047|193175006|SNOMEDCT_US|OPHTHALMOPLEGIA, ATAXIA AND AREFLEXIA SYNDROME|MILLER-FISHER VARIANT OF GUILLAIN-BARRE SYNDROME (DISORDER)
C0393799|T047|193175006|SNOMEDCT_US|MILLER-FISHER VARIANT OF GUILLAIN-BARRE SYNDROME |MILLER-FISHER VARIANT OF GUILLAIN-BARRE SYNDROME (DISORDER)
C0393799|T047|193175006|SNOMEDCT_US|MILLER-FISHER VARIANT OF GUILLAIN-BARRE SYNDROME|MILLER-FISHER VARIANT OF GUILLAIN-BARRE SYNDROME (DISORDER)
C0393799|T047|193175006|SNOMEDCT_US|FISHER'S SYNDROME|MILLER-FISHER VARIANT OF GUILLAIN-BARRE SYNDROME (DISORDER)
C0393799|T047|193175006|SNOMEDCT_US|OPHTHALMOPLEGIA, ATAXIA, AREFLEXIA SYNDROME|MILLER-FISHER VARIANT OF GUILLAIN-BARRE SYNDROME (DISORDER)
C0393799|T047|193175006|SNOMEDCT_US|FISHER'S SYNDROME |MILLER-FISHER VARIANT OF GUILLAIN-BARRE SYNDROME (DISORDER)
C0265235|T047|33410002|SNOMEDCT_US|MARSHALL SYNDROME|MARSHALL SYNDROME (DISORDER)
C0265235|T047|33410002|SNOMEDCT_US|DEAFNESS, MYOPIA, CATARACT, SADDLE NOSE-MARSHALL TYPE|MARSHALL SYNDROME (DISORDER)
C0265235|T047|33410002|SNOMEDCT_US|PFAPA SYNDROME|MARSHALL SYNDROME (DISORDER)
C0265235|T047|33410002|SNOMEDCT_US|PFAPA SYNDROME |MARSHALL SYNDROME (DISORDER)
C0265235|T047|33410002|SNOMEDCT_US|MRSHS|MARSHALL SYNDROME (DISORDER)
C0265235|T047|33410002|SNOMEDCT_US|PERIODIC FEVER, APHTHOUS STOMATITIS, PHARYNGITIS, ADENITIS SYNDROME|MARSHALL SYNDROME (DISORDER)
C0265235|T047|33410002|SNOMEDCT_US|SYNDROME OF PERIODIC FEVER, APHTHOUS STOMATITIS, PHARYNGITIS, CERVICAL ADENITIS|MARSHALL SYNDROME (DISORDER)
C0265235|T047|33410002|SNOMEDCT_US|MARSHALL'S SYNDROME|MARSHALL SYNDROME (DISORDER)
C0265235|T047|33410002|SNOMEDCT_US|MARSHALL SYNDROME |MARSHALL SYNDROME (DISORDER)
C0340971|T047|234425008|SNOMEDCT_US|AUTOIMMUNE NEUTROPENIA|AUTOIMMUNE NEUTROPENIA (DISORDER)
C0340971|T047|234425008|SNOMEDCT_US|NEUTROPENIA AUTOIMMUNE|AUTOIMMUNE NEUTROPENIA (DISORDER)
C0340971|T047|234425008|SNOMEDCT_US|AUTOIMMUNE NEUTROPENIA |AUTOIMMUNE NEUTROPENIA (DISORDER)
C0340971|T047|234425008|SNOMEDCT_US|AUTOIMMUNE NEUTROPENIA |AUTOIMMUNE NEUTROPENIA (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|HASHIMOTO'S DISEASE|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|HASHIMOTO THYROIDITIS|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|LYMPHOMATOUS THYROIDITIS|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|HASHIMOTOS DIS|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|HASHIMOTO DIS|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|HASHIMOTO'S THYROIDITIS|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|HASHIMOTO'S THYROIDITIS |STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|CHR LYMPHOCYT THYROIDIT|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|HASHIMOTO'S SYNDROMES|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|HASHIMOTOS SYNDROME|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|SYNDROMES, HASHIMOTO'S|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|HASHIMOTO SYNDROME|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|SYNDROME, HASHIMOTO'S|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|STRUMA LYMPHOMATOSA|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|HASHIMOTO DISEASE [DISEASE/FINDING]|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|HASHIMOTO DISEASE|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|CHRONIC LYMPHOCYTIC THYROIDITIS|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|HASHIMOTO'S SYNDROME|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|DISEASE;HASHIMOTOS|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|HASHIMOTO STRUMA|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|STRUMA LYMPHOMATOSIS |STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|HASHIMOTO'S THYROIDITIS |STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|STRUMA LYMPHOMATOSIS|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|HASHIMOTO'S STRUMA|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|AUTOIMMUNE THYROIDITIS|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|LYMPHOCYTIC THYROIDITIS|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|AUTOIMMUNE LYMPHOCYTIC CHRONIC THYROIDITIS|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|HASHIMOTO THYROIDITIS |STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|HASHIMOTO; THYROIDITIS|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|HASHIMOTO|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|CHRONIC; THYROIDITIS, LYMPHADENOID|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|LYMPHOCYTIC; THYROIDITIS|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|LYMPHOID; THYROIDITIS|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|LYMPHOMATOSA; GOITER|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|LYMPHOMATOUS; THYROIDITIS|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|STRUMA; LYMPHOMATOSA|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|THYROIDITIS; HASHIMOTO|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|THYROIDITIS; CHRONIC, LYMPHADENOID|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|THYROIDITIS; LYMPHOCYTIC|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|THYROIDITIS; LYMPHOID|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|THYROIDITIS; LYMPHOMATOUS|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|DISEASE, HASHIMOTO|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|HASHIMOTOS DISEASE|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|DISEASE, HASHIMOTO'S|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|CHRONIC LYMPHOCYTIC THYROIDITIDES|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|HASHIMOTO THYROIDITIDES|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|LYMPHOCYTIC THYROIDITIDES, CHRONIC|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|LYMPHOCYTIC THYROIDITIS, CHRONIC|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|THYROIDITIDES, CHRONIC LYMPHOCYTIC|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|THYROIDITIDES, HASHIMOTO|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|THYROIDITIS, CHRONIC LYMPHOCYTIC|STRUMA LYMPHOMATOSIS (DISORDER)
C0677607|T047|237537002|SNOMEDCT_US|THYROIDITIS, HASHIMOTO|STRUMA LYMPHOMATOSIS (DISORDER)
C4022660|T047||SNOMEDCT_US|AUTOIMMUNE ANTIBODY POSITIVITY
C0242584|T047|142969008|SNOMEDCT_US|AUTOIMMUNE THROMBOCYTOPENIA|THROMBOCYTOPENIA (& [AUTO-IMMUNE]) (FINDING)
C0242584|T047|142969008|SNOMEDCT_US|AUTO-IMMUNE THROMBOCYTOPENIA|THROMBOCYTOPENIA (& [AUTO-IMMUNE]) (FINDING)
C0242584|T047|142969008|SNOMEDCT_US|THROMBOCYTOPENIA, AUTOIMMUNE|THROMBOCYTOPENIA (& [AUTO-IMMUNE]) (FINDING)
C0242584|T047|142969008|SNOMEDCT_US|THROMBOCYTOPENIA (& [AUTO-IMMUNE])|THROMBOCYTOPENIA (& [AUTO-IMMUNE]) (FINDING)
C0242584|T047|142969008|SNOMEDCT_US|AUTOIMMUNE THROMBOCYTOPENIA |THROMBOCYTOPENIA (& [AUTO-IMMUNE]) (FINDING)
C0242584|T047|142969008|SNOMEDCT_US|THROMBOCYTOPENIA (& [AUTO-IMMUNE]) |THROMBOCYTOPENIA (& [AUTO-IMMUNE]) (FINDING)
C0242584|T047|142969008|SNOMEDCT_US|THROMBOCYTOPENIA (& [AUTO-IMMUNE]) |THROMBOCYTOPENIA (& [AUTO-IMMUNE]) (FINDING)
C0242584|T047|142969008|SNOMEDCT_US|IMMUNE THROMBOCYTOPENIA|THROMBOCYTOPENIA (& [AUTO-IMMUNE]) (FINDING)
C0342410|T047|237706000|SNOMEDCT_US|AUTOIMMUNE HYPOPHYSITIS|AUTOIMMUNE HYPOPHYSITIS (DISORDER)
C0342410|T047|237706000|SNOMEDCT_US|HYPOPHYSITIDES, AUTOIMMUNE|AUTOIMMUNE HYPOPHYSITIS (DISORDER)
C0342410|T047|237706000|SNOMEDCT_US|LYMPHOID HYPOPHYSITIDES|AUTOIMMUNE HYPOPHYSITIS (DISORDER)
C0342410|T047|237706000|SNOMEDCT_US|HYPOPHYSITIS, LYMPHOID|AUTOIMMUNE HYPOPHYSITIS (DISORDER)
C0342410|T047|237706000|SNOMEDCT_US|LYMPHOCYTIC HYPOPHYSITIDES|AUTOIMMUNE HYPOPHYSITIS (DISORDER)
C0342410|T047|237706000|SNOMEDCT_US|HYPOPHYSITIDES, LYMPHOID|AUTOIMMUNE HYPOPHYSITIS (DISORDER)
C0342410|T047|237706000|SNOMEDCT_US|HYPOPHYSITIDES, LYMPHOCYTIC|AUTOIMMUNE HYPOPHYSITIS (DISORDER)
C0342410|T047|237706000|SNOMEDCT_US|AUTOIMMUNE HYPOPHYSITIDES|AUTOIMMUNE HYPOPHYSITIS (DISORDER)
C0342410|T047|237706000|SNOMEDCT_US|AUTOIMMUNE HYPOPHYSITIS [DISEASE/FINDING]|AUTOIMMUNE HYPOPHYSITIS (DISORDER)
C0342410|T047|237706000|SNOMEDCT_US|HYPOPHYSITIS, LYMPHOCYTIC|AUTOIMMUNE HYPOPHYSITIS (DISORDER)
C0342410|T047|237706000|SNOMEDCT_US|HYPOPHYSITIS, AUTOIMMUNE|AUTOIMMUNE HYPOPHYSITIS (DISORDER)
C0342410|T047|237706000|SNOMEDCT_US|LYMPHOCYTIC HYPOPHYSITIS|AUTOIMMUNE HYPOPHYSITIS (DISORDER)
C0342410|T047|237706000|SNOMEDCT_US|LYMPHOID HYPOPHYSITIS|AUTOIMMUNE HYPOPHYSITIS (DISORDER)
C0342410|T047|237706000|SNOMEDCT_US|AUTOIMMUNE HYPOPHYSITIS |AUTOIMMUNE HYPOPHYSITIS (DISORDER)
C0393639|T047|95643007|SNOMEDCT_US|HASHIMOTO'S ENCEPHALOPATHY|AUTOIMMUNE ENCEPHALITIS (DISORDER)
C0393639|T047|95643007|SNOMEDCT_US|HASHIMOTO'S ENCEPHALITIS|AUTOIMMUNE ENCEPHALITIS (DISORDER)
C0393639|T047|95643007|SNOMEDCT_US|STEROID-RESPONSIVE ENCEPHALOPATHY ASSOCIATED WITH AUTOIMMUNE THYROIDITIS|AUTOIMMUNE ENCEPHALITIS (DISORDER)
C0393639|T047|95643007|SNOMEDCT_US|AUTOIMMUNE ENCEPHALITIS|AUTOIMMUNE ENCEPHALITIS (DISORDER)
C0393639|T047|95643007|SNOMEDCT_US|ENCEPHALITIS AUTOIMMUNE|AUTOIMMUNE ENCEPHALITIS (DISORDER)
C0393639|T047|95643007|SNOMEDCT_US|AUTOIMMUNE ENCEPHALOPATHY|AUTOIMMUNE ENCEPHALITIS (DISORDER)
C0393639|T047|95643007|SNOMEDCT_US|ENCEPHALITIS ALLERGIC (AUTOIMMUNE)|AUTOIMMUNE ENCEPHALITIS (DISORDER)
C0393639|T047|95643007|SNOMEDCT_US|AUTOIMMUNE ENCEPHALITIS |AUTOIMMUNE ENCEPHALITIS (DISORDER)
C0393639|T047|95643007|SNOMEDCT_US|AUTOIMMUNE ENCEPHALITIS, NOS|AUTOIMMUNE ENCEPHALITIS (DISORDER)
C4075851|T047|713654004|SNOMEDCT_US|AUTOIMMUNE CHOLANGITIS |AUTOIMMUNE CHOLANGITIS (DISORDER)
C4075851|T047|713654004|SNOMEDCT_US|AUTOIMMUNE CHOLANGITIS|AUTOIMMUNE CHOLANGITIS (DISORDER)
C0271893|T047|183005|SNOMEDCT_US|AUTOIMMUNE PANCYTOPENIA|AUTOIMMUNE PANCYTOPENIA (DISORDER)
C0271893|T047|183005|SNOMEDCT_US|PANCYTOPENIA AUTOIMMUNE|AUTOIMMUNE PANCYTOPENIA (DISORDER)
C0271893|T047|183005|SNOMEDCT_US|PANCYTOPENIA AUTOIMMUNE |AUTOIMMUNE PANCYTOPENIA (DISORDER)
C0271893|T047|183005|SNOMEDCT_US|AUTOIMMUNE PANCYTOPENIA |AUTOIMMUNE PANCYTOPENIA (DISORDER)
C0543694|T047|123777002|SNOMEDCT_US|AUTOIMMUNE LEUKOPENIA|AUTOIMMUNE LEUKOPENIA (DISORDER)
C0543694|T047|123777002|SNOMEDCT_US|AUTOIMMUNE LEUCOPENIA|AUTOIMMUNE LEUKOPENIA (DISORDER)
C0543694|T047|123777002|SNOMEDCT_US|AUTOIMMUNE LEUKOPENIA |AUTOIMMUNE LEUKOPENIA (DISORDER)
C0395947|T047|232308006|SNOMEDCT_US|AUTOIMMUNE DISORDER OF INNER EAR|AUTOIMMUNE DISORDER OF INNER EAR (DISORDER)
C0395947|T047|232308006|SNOMEDCT_US|AUTOIMMUNE LABYRINTHITIS|AUTOIMMUNE DISORDER OF INNER EAR (DISORDER)
C0395947|T047|232308006|SNOMEDCT_US|AUTOIMMUNE DISORDER OF INNER EAR |AUTOIMMUNE DISORDER OF INNER EAR (DISORDER)
C0406632|T047|95329006|SNOMEDCT_US|AUTOIMMUNE DISEASES AFFECTING SKIN|AUTOIMMUNE SKIN DISEASE (DISORDER)
C0406632|T047|95329006|SNOMEDCT_US|AUTOIMMUNE SKIN DISEASE |AUTOIMMUNE SKIN DISEASE (DISORDER)
C0406632|T047|95329006|SNOMEDCT_US|AUTOIMMUNE SKIN DISEASE|AUTOIMMUNE SKIN DISEASE (DISORDER)
C0406632|T047|95329006|SNOMEDCT_US|AUTOIMMUNE SKIN DISEASE, NOS|AUTOIMMUNE SKIN DISEASE (DISORDER)
C0086981|T047|267875002|SNOMEDCT_US|SICCA SYNDROME|SICCA SYNDROME (DISORDER)
C0086981|T047|267875002|SNOMEDCT_US|SYNDROME, SICCA|SICCA SYNDROME (DISORDER)
C0086981|T047|267875002|SNOMEDCT_US|XERODERMOSTEOSIS|SICCA SYNDROME (DISORDER)
C0086981|T047|267875002|SNOMEDCT_US|SICCA SYNDROME |SICCA SYNDROME (DISORDER)
C0086981|T047|267875002|SNOMEDCT_US|SICCA|SICCA SYNDROME (DISORDER)
C0086981|T047|267875002|SNOMEDCT_US|SICCA SYNDROME, UNSPECIFIED|SICCA SYNDROME (DISORDER)
C0086981|T047|267875002|SNOMEDCT_US|SICCA SYNDROME |SICCA SYNDROME (DISORDER)
C0086981|T047|267875002|SNOMEDCT_US|SYNDROME SICCA|SICCA SYNDROME (DISORDER)
C0086981|T047|267875002|SNOMEDCT_US|SICCA; SYNDROME|SICCA SYNDROME (DISORDER)
C0086981|T047|267875002|SNOMEDCT_US|SYNDROME; SICCA|SICCA SYNDROME (DISORDER)
C1328835|T047||SNOMEDCT_US|AUTOIMMUNE DERMATOLOGIC DISORDER
C1328836|T047||SNOMEDCT_US|AUTOIMMUNE GASTROINTESTINAL AND LIVER DISORDER
C1328837|T047||SNOMEDCT_US|AUTOIMMUNE GENITOURINARY DISORDER
C1328837|T047||SNOMEDCT_US|AUTOIMMUNE UROGENITAL DISORDER
C1328837|T047||SNOMEDCT_US|UROGENITAL AUTOIMMUNE DISORDER
C1328841|T047||SNOMEDCT_US|AUTOIMMUNE RESPIRATORY DISORDER
C1328842|T047||SNOMEDCT_US|AUTOIMMUNE RHEUMATOLOGIC DISEASE
C0175816|T047|234382005|SNOMEDCT_US|COLD TYPE HAEMOLYTIC ANAEMIA|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|COLD AGGLUTININ DIS|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|COLD HEMAGGLUTININ DISEASE|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|COLD ANTIBODY HEMOLYTIC ANEMIA|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|HEMOLYTIC ANEMIA DUE TO COLD AGGLUTININ DISEASE |COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|HEMOLYTIC ANEMIA DUE TO COLD AGGLUTININ DISEASE|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|COLD AGGLUTININ DISEASE|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|DISEASES, COLD ANTIBODY|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|DISEASE, COLD ANTIBODY|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|COLD ANTIBODY DISEASES|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|HAEMOLYTIC ANAEMIA DUE TO COLD ANTIBODY|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|CRYOPATHIC HEMOLYTIC ANEMIA|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|COLD HAEMAGGLUTININ DISEASE|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|AIHA - COLD AUTOIMMUNE HEMOLYTIC ANEMIA|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|HEMOLYTIC ANEMIA DUE TO COLD ANTIBODY|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|COLD AUTOIMMUNE HEMOLYTIC ANEMIA |COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|COLD AUTOIMMUNE HAEMOLYTIC ANAEMIA|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|CHAD - COLD HEMAGGLUTININ DISEASE|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|COLD AUTOIMMUNE HEMOLYTIC ANEMIA|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|AIHA - COLD AUTOIMMUNE HAEMOLYTIC ANAEMIA|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|COLD TYPE HEMOLYTIC ANEMIA|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|COLD HEMOLYTIC DISEASE|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|COLD ANTIBODY HAEMOLYTIC ANAEMIA|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|CRYOPATHIC HAEMOLYTIC ANAEMIA|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|COLD HAEMOLYTIC DISEASE|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|COLD HAEMAGGLUTININ DISEASE |COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|CHAD - COLD HAEMAGGLUTININ DISEASE|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|ANEMIA, HEMOLYTIC, COLD ANTIBODY|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|COLD ANTIBODY DISEASE|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|HEMOLYTIC ANEMIA DUE TO COLD ANTIBODY, NOS|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|AGGLUTININ DISEASE, COLD|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|AGGLUTININ DISEASES, COLD|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|COLD AGGLUTININ DISEASES|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|DISEASE, COLD AGGLUTININ|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0175816|T047|234382005|SNOMEDCT_US|DISEASES, COLD AGGLUTININ|COLD HAEMAGGLUTININ DISEASE (DISORDER)
C0011644|T047|287005009|SNOMEDCT_US|SCLERODERMA|SCLERODERMA NOS (DISORDER)
C0011644|T047|287005009|SNOMEDCT_US|DERMATOSCLEROSIS|SCLERODERMA NOS (DISORDER)
C0011644|T047|287005009|SNOMEDCT_US|SCLERODERMA |SCLERODERMA NOS (DISORDER)
C0011644|T047|287005009|SNOMEDCT_US|SCLERODERMA |SCLERODERMA NOS (DISORDER)
C0011644|T047|287005009|SNOMEDCT_US|SCLERODERMA NOS|SCLERODERMA NOS (DISORDER)
C0011644|T047|287005009|SNOMEDCT_US|SCLERODERMA NOS |SCLERODERMA NOS (DISORDER)
C0011644|T047|287005009|SNOMEDCT_US|SCLERODERMA |SCLERODERMA NOS (DISORDER)
C0011644|T047|287005009|SNOMEDCT_US|PROGRESSIVE SYSTEMIC SCLERODERMA|SCLERODERMA NOS (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|DERMATOMYOSITIDES|[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|DERMATOMYOSITIS|[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|DERMATOPOLYMYOSITIS|[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|DERMATOPOLYMYOSITIS, UNSPECIFIED|[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|POLYMYOSITIS DERMATOMYOSITIS|[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|POLYMYOSITIS-DERMATOMYOSITIDES|[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|DERMATOPOLYMYOSITIDES|[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|DERMATOPOLYMYOSITIS, UNSPECIFIED, ORGAN INVOLVEMENT UNSPECIFIED|[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|POLYMYOSITIS-DERMATOMYOSITIS|[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|DERMATOMYOSITIS [DISEASE/FINDING]|[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|DERMATOPOLYMYOSITIS, UNSP, ORGAN INVOLVEMENT UNSPECIFIED|[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|[X]DERMATOPOLYMYOSITIS, UNSPECIFIED|[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|POLYMYOSITIS WITH SKIN INVOLVEMENT|[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|DM - DERMATOMYOSITIS|[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|DERMATOMYOSITIS |[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|[X]DERMATOPOLYMYOSITIS, UNSPECIFIED |[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|WAGNER-UNVERRICHT SYNDROME|[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|DERMATOPOLYMYOSITIS |[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|POLYMYOSITIS/DERMATOMYOSITIS|[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|DERMATOMYOSITIS |[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|POLYMYOSITIS; WITH INVOLVEMENT OF SKIN|[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0011633|T047|201448000|SNOMEDCT_US|DERMATOMUCOSOMYOSITIS|[X]DERMATOPOLYMYOSITIS, UNSPECIFIED (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|DISEASE, SCHAUMANN|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SARCOID, BOECK'S|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SARCOIDOSES|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SARCOIDOSIS|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BESNIER BOECK DISEASE|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BOECK SARCOID|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BOECKS SARCOID|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SARCOIDOSIS, UNSPECIFIED|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BOECK'S SARCOIDOSIS|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BOECKS SARCOIDOSIS|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SCHAUMANN DIS|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BESNIER BOECK DIS|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|LYMPHOGRANULOMATOSIS (BENIGN)|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SARCOIDOSIS |SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BENIGN LYMPHOGRANULOMATOSIS|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BOECK'S SARCOID|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BENIGN LYMPHOGRANULOMATOSIS |SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BENIGN LYMPHOGRANULOMATOSIS OF SCHAUMANN|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SYNDROME, BESNIER-BOECK-SCHAUMANN|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SYNDROME, SCHAUMANN|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SCHAUMANN'S SYNDROMES|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BESNIER BOECK SCHAUMANN SYNDROME|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BOECKS DISEASE|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SYNDROME, SCHAUMANN'S|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SCHAUMANN DISEASE|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SARCOIDOSIS [DISEASE/FINDING]|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BESNIER-BOECK DISEASE|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BOECK DISEASE|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SCHAUMANN SYNDROME|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BESNIER-BOECK-SCHAUMANN SYNDROME|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SCHAUMANN'S SYNDROME|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BOECK'S DISEASE|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|LYMPHOGRANULOMATOSIS|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SARCOIDOSIS |SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SARCOID|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SCHAUMANN'S DISEASE|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BESNIER-BOECK-SCHAUMANN'S DISEASE|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SARCOIDOSIS NOS|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|DARIER-ROUSSY SARCOID|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|LUPUS PERNIO OF BESNIER|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|MILIARY LUPOID OF BOECK|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BENIGN; LYMPHOGRANULOMATOSIS|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|HUTCHINSON-BOECK|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SCHAUMANN; BENIGN LYMPHOGRANULOMATOSIS|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SCHAUMANN; DISEASE OR SYNDROME|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BESNIER-BOECK|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BESNIER; LUPUS PERNIO|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BOECK; DISEASE|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BOECK; SARCOID|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|LYMPHOGRANULOMATOSIS; BENIGN|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SARCOID; BOECK|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SARCOID; DARIER-ROUSSY|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SYNDROME; SCHAUMANN|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|DARIER-ROUSSY; SARCOID|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SARCOIDOSIS, NOS|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BESNIER-BOECK-SCHAUMANN DISEASE|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BOECK SARCOID, ANY SITE|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|BENIGN LYMPHOGRANULOMATOSIS, SCHAUMANN'S|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|LUPUS PERNIO, BESNIER|SARCOIDOSIS (DISORDER)
C0036202|T047|31541009|SNOMEDCT_US|SARCOID NOS|SARCOIDOSIS (DISORDER)
C0272126|T047|75331009|SNOMEDCT_US|EVANS SYNDROME|EVANS SYNDROME (DISORDER)
C0272126|T047|75331009|SNOMEDCT_US|EVANS' SYNDROME |EVANS SYNDROME (DISORDER)
C0272126|T047|75331009|SNOMEDCT_US|EVANS' SYNDROME|EVANS SYNDROME (DISORDER)
C0272126|T047|75331009|SNOMEDCT_US|AUTOIMMUNE HEMOLYTIC ANEMIA AND AUTOIMMUNE THROMBOCYTOPENIA|EVANS SYNDROME (DISORDER)
C0272126|T047|75331009|SNOMEDCT_US|EVAN'S SYNDROME|EVANS SYNDROME (DISORDER)
C0272126|T047|75331009|SNOMEDCT_US|EVANS SYNDROME |EVANS SYNDROME (DISORDER)
C0272126|T047|75331009|SNOMEDCT_US|EVANS|EVANS SYNDROME (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|DISEASE, PERIODIC|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|FAMILIAL MEDITERRANEAN FEVER|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|BENIGN PAROXYSMAL PERITONITIS|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|RECURRENT POLYSEROSITIS|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|FMF|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|WOLFFS PERIODIC DIS|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|WOLFF PERIODIC DIS|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PERIODIC DIS WOLFFS|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PERIODIC DIS|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|FAMILIAL MEDITERRANEAN FEVER |FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|FAMILIAL MEDITERRANEAN FEVER WITH RECURRENT POLYSEROSITIS|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|FAMILIAL MEDITERRANEAN FEVER WITH RECURRENT POLYSEROSITIS |FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|DISEASE, WOLFF PERIODIC|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|DISEASE, WOLFF'S PERIODIC|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PERIODIC DISEASE, WOLFF|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|WOLFFS PERIODIC DISEASE|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|FAM MEDITERRANEAN FEVER|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|DISEASES, PERIODIC|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PERIODIC DISEASE, WOLFFS|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PERIODIC DISEASES|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|WOLFF PERIODIC DISEASE|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PERIODIC DISEASE, WOLFF'S|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|FAMILIAL MEDITERRANEAN FEVER [DISEASE/FINDING]|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|WOLFF'S PERIODIC DISEASE|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|MEDITERRANEAN FEVER, FAMILIAL|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PERIODIC DISEASE|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PERITONITIS, PERIODIC|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PERITONITIDES, BENIGN PAROXYSMAL|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PERITONITIS, BENIGN PAROXYSMAL|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|FAMILIAL PAROXYSMAL POLYSEROSITIDES|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PERIODIC PERITONITIDES|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PERITONITIDES, PERIODIC|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PAROXYSMAL POLYSEROSITIS, FAMILIAL|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PAROXYSMAL PERITONITIDES, BENIGN|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PAROXYSMAL POLYSEROSITIDES, FAMILIAL|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|BENIGN PAROXYSMAL PERITONITIDES|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PAROXYSMAL PERITONITIS, BENIGN|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|POLYSEROSITIDES, FAMILIAL PAROXYSMAL|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|POLYSEROSITIDES, RECURRENT|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|RECURRENT POLYSEROSITIDES|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PERIODIC PERITONITIS|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|FAMILIAL PAROXYSMAL POLYSEROSITIS|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|POLYSEROSITIS, RECURRENT|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|POLYSEROSITIS, FAMILIAL PAROXYSMAL|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|FAMILIAL MEDITERRANEAN FEVER, AUTOSOMAL RECESSIVE|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|FAMILIAL MEDITERRANEAN FEVER AUTOSOMAL RECESSIVE|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|FMF AUTOSOMAL RECESSIVE|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|FAMILIAL MEDITERRANEAN FEVER AUTOSOMAL RECESSIVE |FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|FAMILIAL RECURRENT POLYSEROSITIS|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PAROXYSMAL POLYSEROSITIS|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|FMF - FAMILIAL MEDITERRANEAN FEVER|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PERIODIC FAMILIAL PERITONITIS|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PERIODIC POLYSEROSITIS|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|MEF - FAMILIAL MEDITERRANEAN FEVER|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|FAMILIAL MEDITERRANEAN FEVER |FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|FEVER; MEDITERRANEAN, FAMILIAL|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|MEDITERRANEAN; FEVER, FAMILIAL|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PERIODIC; PERITONITIS|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PERIODIC; POLYSEROSITIS|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PERITONITIS; PERIODIC|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|POLYSEROSITIS; PERIODIC|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
C0031069|T047|12579009|SNOMEDCT_US|PERIODIC FEVER|FAMILIAL MEDITERRANEAN FEVER (DISORDER)
