C1305855|T034|9300|MEDCIN|BODY MASS INDEX|BODY MASS INDEX (PHYSICAL FINDING)
C0005893|T034||MEDCIN|BODY MASS INDEX PROCEDURE
C4229017|T034||MEDCIN|NORMAL BMI
C0424671|T034||MEDCIN|BODY MASS INDEX 30+ OBESITY
C1561729|T034||MEDCIN|BODY MASS INDEX (BMI) 40 OR GREATER, ADULT
C2724372|T034||MEDCIN|BODY MASS INDEX (BMI), DOCUMENTED (PV)
C2240399|T034||MEDCIN|ENCOUNTER FOR BODY MASS INDEX [BMI]
C0578022|T034||MEDCIN|FINDING OF BODY MASS INDEX
C1305855|T034|9300|MEDCIN|QUETELET INDEX|BODY MASS INDEX (PHYSICAL FINDING)
C1305855|T034|9300|MEDCIN|BODY MASS INDEX|BODY MASS INDEX (PHYSICAL FINDING)
C1305855|T034|9300|MEDCIN|BMI|BODY MASS INDEX (PHYSICAL FINDING)
C1305855|T034|9300|MEDCIN|BODY MASS INDEX (PHYSICAL FINDING)|BODY MASS INDEX (PHYSICAL FINDING)
C1305855|T034|9300|MEDCIN|QUETELET INDEX (OBSERVABLE ENTITY)|BODY MASS INDEX (PHYSICAL FINDING)
C1305855|T034|9300|MEDCIN|BODY MASS INDEX - OBSERVATION|BODY MASS INDEX (PHYSICAL FINDING)
C1305855|T034|9300|MEDCIN|BODY MASS INDEX (OBSERVABLE ENTITY)|BODY MASS INDEX (PHYSICAL FINDING)
C1305855|T034|9300|MEDCIN|BMI - BODY MASS INDEX|BODY MASS INDEX (PHYSICAL FINDING)
C1305855|T034|9300|MEDCIN|BODY MASS INDEX, NOS|BODY MASS INDEX (PHYSICAL FINDING)
C1305855|T034|9300|MEDCIN|BODY MASS INDEX [DUP] (OBSERVABLE ENTITY)|BODY MASS INDEX (PHYSICAL FINDING)
C2227318|T034|268430|MEDCIN|BMI ___ PERCENTILE|BODY MASS INDEX PERCENTILE (PHYSICAL FINDING)
C2227318|T034|268430|MEDCIN|BODY MASS INDEX PERCENTILE (PHYSICAL FINDING)|BODY MASS INDEX PERCENTILE (PHYSICAL FINDING)
C2227318|T034|268430|MEDCIN|BODY MASS INDEX PERCENTILE|BODY MASS INDEX PERCENTILE (PHYSICAL FINDING)
C0578022|T034||MEDCIN|OBSERVATION OF BODY MASS INDEX
C0578022|T034||MEDCIN|FINDING OF BODY MASS INDEX 
C0578022|T034||MEDCIN|FINDING OF BODY MASS INDEX
C3695134|T034|297651|MEDCIN|BODY MASS INDEX SCREENING SCORE (PHYSICAL FINDING)|BODY MASS INDEX SCREENING SCORE (PHYSICAL FINDING)
C3695134|T034|297651|MEDCIN|BODY MASS INDEX SCREENING SCORE|BODY MASS INDEX SCREENING SCORE (PHYSICAL FINDING)
C0231255|T034|297796|MEDCIN|BODY MASS INDEX DECREASED|BODY MASS INDEX LOW (PHYSICAL FINDING)
C0231255|T034|297796|MEDCIN|BODY MASS INDEX DECREASED (PHYSICAL FINDING)|BODY MASS INDEX LOW (PHYSICAL FINDING)
C0231255|T034|297796|MEDCIN|BODY MASS INDEX LOW (PHYSICAL FINDING)|BODY MASS INDEX LOW (PHYSICAL FINDING)
C0231255|T034|297796|MEDCIN|BODY MASS INDEX LOW|BODY MASS INDEX LOW (PHYSICAL FINDING)
C0231255|T034|297796|MEDCIN|DECREASED BODY MASS INDEX|BODY MASS INDEX LOW (PHYSICAL FINDING)
C0231255|T034|297796|MEDCIN|LOW BODY MASS INDEX|BODY MASS INDEX LOW (PHYSICAL FINDING)
C0231255|T034|297796|MEDCIN|DECREASED BODY MASS INDEX |BODY MASS INDEX LOW (PHYSICAL FINDING)
C0231253|T034|297751|MEDCIN|BODY MASS INDEX NORMAL|NORMAL BODY MASS INDEX (PHYSICAL FINDING)
C0231253|T034|297751|MEDCIN|NORMAL BODY MASS INDEX (PHYSICAL FINDING)|NORMAL BODY MASS INDEX (PHYSICAL FINDING)
C0231253|T034|297751|MEDCIN|NORMAL BODY MASS INDEX|NORMAL BODY MASS INDEX (PHYSICAL FINDING)
C0231253|T034|297751|MEDCIN|NORMAL BODY MASS INDEX |NORMAL BODY MASS INDEX (PHYSICAL FINDING)
C0231254|T034|297795|MEDCIN|BODY MASS INDEX INCREASED|BODY MASS INDEX HIGH (PHYSICAL FINDING)
C0231254|T034|297795|MEDCIN|INCREASED BODY MASS INDEX|BODY MASS INDEX HIGH (PHYSICAL FINDING)
C0231254|T034|297795|MEDCIN|BODY MASS INDEX INCREASED (PHYSICAL FINDING)|BODY MASS INDEX HIGH (PHYSICAL FINDING)
C0231254|T034|297795|MEDCIN|BODY MASS INDEX HIGH|BODY MASS INDEX HIGH (PHYSICAL FINDING)
C0231254|T034|297795|MEDCIN|BODY MASS INDEX HIGH (PHYSICAL FINDING)|BODY MASS INDEX HIGH (PHYSICAL FINDING)
C0231254|T034|297795|MEDCIN|INCREASE IN BODY MASS INDEX|BODY MASS INDEX HIGH (PHYSICAL FINDING)
C0231254|T034|297795|MEDCIN|INCREASED BODY MASS INDEX |BODY MASS INDEX HIGH (PHYSICAL FINDING)
C2911062|T034|298297|MEDCIN|BODY MASS INDEX, PEDIATRIC|BMI, PEDIATRIC
C2911062|T034|298297|MEDCIN|BODY MASS INDEX (BMI) PEDIATRIC|BMI, PEDIATRIC
C2911062|T034|298297|MEDCIN|BODY MASS INDEX PEDIATRIC|BMI, PEDIATRIC
C2911062|T034|298297|MEDCIN|BODY MASS INDEX, PEDIATRIC (PHYSICAL FINDING)|BMI, PEDIATRIC
C0005893|T034||MEDCIN|BODY MASS INDEX
C0005893|T034||MEDCIN|INDEX, BODY MASS
C0005893|T034||MEDCIN|QUETELETS INDEX
C0005893|T034||MEDCIN|QUETELET'S INDEX
C0005893|T034||MEDCIN|QUETELET INDEX
C0005893|T034||MEDCIN|BODY MASS INDEX PROCEDURE
C0005893|T034||MEDCIN|INDEX, QUETELET
C0424671|T034||MEDCIN|BODY MASS INDEX 30+ - OBESITY
C0424671|T034||MEDCIN|OBESITY (BMI>30)
C0424671|T034||MEDCIN|BODY MASS INDEX 30+ - OBESITY 
C0424671|T034||MEDCIN|BMI 30+ - OBESITY
C2921312|T034||MEDCIN|BMI 40.0-44.9, ADULT
C2921312|T034||MEDCIN|BODY MASS INDEX 40.0-44.9, ADULT
C2921313|T034||MEDCIN|BODY MASS INDEX 45.0-49.9, ADULT
C2921313|T034||MEDCIN|BMI 45.0-49.9, ADULT
C2921314|T034||MEDCIN|BMI 50.0-59.9, ADULT
C2921314|T034||MEDCIN|BODY MASS INDEX 50.0-59.9, ADULT
C2921315|T034||MEDCIN|BODY MASS INDEX 60.0-69.9, ADULT
C2921315|T034||MEDCIN|BMI 60.0-69.9, ADULT
C2921316|T034||MEDCIN|BMI 70 AND OVER, ADULT
C2921316|T034||MEDCIN|BODY MASS INDEX 70 AND OVER, ADULT
C2977643|T034||MEDCIN|BODY MASS INDEX (BMI) 40.0-44.9, ADULT
C2977644|T034||MEDCIN|BODY MASS INDEX (BMI) 45.0-49.9, ADULT
C2977645|T034||MEDCIN|BODY MASS INDEX (BMI) 50-59.9 , ADULT
C2977646|T034||MEDCIN|BODY MASS INDEX (BMI) 60.0-69.9, ADULT
C2977647|T034||MEDCIN|BODY MASS INDEX (BMI) 70 OR GREATER, ADULT
C2724372|T034||MEDCIN|BODY MASS INDEX DOCD
C2724372|T034||MEDCIN|BODY MASS INDEX (BMI), DOCUMENTED (PV)
C2724372|T034||MEDCIN|BODY MASS INDEX DOCUMENTED
C2911038|T034||MEDCIN|BODY MASS INDEX (BMI) 19 OR LESS, ADULT
C2911039|T034||MEDCIN|BODY MASS INDEX (BMI) 20-29, ADULT
C2911050|T034||MEDCIN|BODY MASS INDEX (BMI) 30-39, ADULT
C1561729|T034||MEDCIN|BODY MASS INDEX 40 AND OVER, ADULT
C1561729|T034||MEDCIN|BODY MASS INDEX (BMI) 40 OR GREATER, ADULT
C2240399|T034||MEDCIN|BODY MASS INDEX
C2240399|T034||MEDCIN|BODY MASS INDEX [BMI]
C2240399|T034||MEDCIN|ENCOUNTER FOR BODY MASS INDEX [BMI]
C2240399|T034||MEDCIN|BODY MASS INDEX [BMI] (Z68)
C1561711|T034||MEDCIN|BMI BETWEEN 19-24,ADULT
C1561711|T034||MEDCIN|BODY MASS INDEX BETWEEN 19-24, ADULT
C1561717|T034||MEDCIN|BODY MASS INDEX BETWEEN 25-29, ADULT
C1561728|T034||MEDCIN|BODY MASS INDEX BETWEEN 30-39, ADULT
C1561710|T034||MEDCIN|BMI LESS THAN 19,ADULT
C1561710|T034||MEDCIN|BODY MASS INDEX LESS THAN 19, ADULT
C1319441|T034||MEDCIN|BODY MASS INDEX 40+ - MORBIDLY OBESE
C1319441|T034||MEDCIN|OBESE CLASS III
C1319441|T034||MEDCIN|BODY MASS INDEX 40+ - SEVERELY OBESE 
C1319441|T034||MEDCIN|BODY MASS INDEX 40+ - SEVERELY OBESE
C0587773|T034||MEDCIN|BODY MASS INDEX LESS THAN 20 
C0587773|T034||MEDCIN|BODY MASS INDEX LESS THAN 20
C0587773|T034||MEDCIN|BMI LESS THAN 20
C0424672|T034||MEDCIN|BODY MASS INDEX 25-29 - OVERWEIGHT 
C0424672|T034||MEDCIN|BODY MASS INDEX INDEX 25-29 - OVERWEIGHT
C0424672|T034||MEDCIN|BODY MASS INDEX 25-29 - OVERWEIGHT
C0424672|T034||MEDCIN|BODY MASS INDEX INDEX 25-29 - OVERWEIGHT 
C0424672|T034||MEDCIN|BMI 25-29 - OVERWEIGHT
C1445936|T034||MEDCIN|BODY MASS INDEX 20-24 - NORMAL 
C1445936|T034||MEDCIN|BODY MASS INDEX 20-24 - NORMAL
C0424674|T034||MEDCIN|BODY MASS INDEX HIGH K/M2
C0424674|T034||MEDCIN|BODY MASS INDEX HIGH K/M2 
C0424673|T034||MEDCIN|BODY MASS INDEX LOW K/M2
C0424673|T034||MEDCIN|BODY MASS INDEX LOW K/M2 
C0424675|T034||MEDCIN|BODY MASS INDEX NORMAL K/M2 
C0424675|T034||MEDCIN|BODY MASS INDEX NORMAL K/M2
