C0014544|T047|267698007|SNOMEDCT_US|EPILEPSY|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0751495|T047|3485007|SNOMEDCT_US|PARTIAL SEIZURE|LOCAL CONVULSION (DISORDER)
C0751495|T047|3485007|SNOMEDCT_US|FOCAL SEIZURE|LOCAL CONVULSION (DISORDER)
C0751495|T047|3485007|SNOMEDCT_US|SEIZURES, PARTIAL, AFEBRILE|LOCAL CONVULSION (DISORDER)
C0751495|T047|3485007|SNOMEDCT_US|PARTIAL SEIZURE (PHYSICAL FINDING)|LOCAL CONVULSION (DISORDER)
C0751495|T047|3485007|SNOMEDCT_US|SEIZURE PARTIAL (FOCAL)|LOCAL CONVULSION (DISORDER)
C0751495|T047|3485007|SNOMEDCT_US|CONVULSIONS LOCAL|LOCAL CONVULSION (DISORDER)
C0751495|T047|3485007|SNOMEDCT_US|PARTIAL SEIZURES, NOS|LOCAL CONVULSION (DISORDER)
C0751495|T047|3485007|SNOMEDCT_US|FOCAL SEIZURES|LOCAL CONVULSION (DISORDER)
C0751495|T047|3485007|SNOMEDCT_US|SEIZURE, FOCAL|LOCAL CONVULSION (DISORDER)
C0751495|T047|3485007|SNOMEDCT_US|SEIZURES, PARTIAL|LOCAL CONVULSION (DISORDER)
C0751495|T047|3485007|SNOMEDCT_US|PARTIAL SEIZURES|LOCAL CONVULSION (DISORDER)
C0751495|T047|3485007|SNOMEDCT_US|LOCAL CONVULSION|LOCAL CONVULSION (DISORDER)
C0751495|T047|3485007|SNOMEDCT_US|PARTIAL SEIZURE |LOCAL CONVULSION (DISORDER)
C0751495|T047|3485007|SNOMEDCT_US|LOCAL CONVULSION |LOCAL CONVULSION (DISORDER)
C0751495|T047|3485007|SNOMEDCT_US|SEIZURES, FOCAL|LOCAL CONVULSION (DISORDER)
C0751495|T047|3485007|SNOMEDCT_US|PARTIAL SEIZURES NOS|LOCAL CONVULSION (DISORDER)
C0751495|T047|3485007|SNOMEDCT_US|FOCAL FITS|LOCAL CONVULSION (DISORDER)
C0751495|T047|3485007|SNOMEDCT_US|LOCAL SEIZURE|LOCAL CONVULSION (DISORDER)
C0751495|T047|3485007|SNOMEDCT_US|PARTIAL SEIZURE |LOCAL CONVULSION (DISORDER)
C0751495|T047|3485007|SNOMEDCT_US|FOCAL SEIZURE, NOS|LOCAL CONVULSION (DISORDER)
C0234533|T047|246545002|SNOMEDCT_US|GENERALIZED SEIZURE|GENERALIZED SEIZURE (FINDING)
C0234533|T047|246545002|SNOMEDCT_US|GENERALIZED SEIZURES|GENERALIZED SEIZURE (FINDING)
C0234533|T047|246545002|SNOMEDCT_US|GENERALIZED CONVULSIONS |GENERALIZED SEIZURE (FINDING)
C0234533|T047|246545002|SNOMEDCT_US|GENERALIZED CONVULSIONS|GENERALIZED SEIZURE (FINDING)
C0234533|T047|246545002|SNOMEDCT_US|GENERALIZED SEIZURE (PHYSICAL FINDING)|GENERALIZED SEIZURE (FINDING)
C0234533|T047|246545002|SNOMEDCT_US|SEIZURE GENERALIZED|GENERALIZED SEIZURE (FINDING)
C0234533|T047|246545002|SNOMEDCT_US|SEIZURE, GENERALIZED|GENERALIZED SEIZURE (FINDING)
C0234533|T047|246545002|SNOMEDCT_US|SEIZURES, GENERALIZED|GENERALIZED SEIZURE (FINDING)
C0234533|T047|246545002|SNOMEDCT_US|GENERALIZED CONVULSION|GENERALIZED SEIZURE (FINDING)
C0234533|T047|246545002|SNOMEDCT_US|GENERALISED CONVULSION|GENERALIZED SEIZURE (FINDING)
C0234533|T047|246545002|SNOMEDCT_US|GENERALIZED CONVULSION |GENERALIZED SEIZURE (FINDING)
C0234533|T047|246545002|SNOMEDCT_US|CONVULSIONS GENERALIZED|GENERALIZED SEIZURE (FINDING)
C0234533|T047|246545002|SNOMEDCT_US|CONVULSIONS GENERALISED|GENERALIZED SEIZURE (FINDING)
C0234533|T047|246545002|SNOMEDCT_US|GENERALISED SEIZURE|GENERALIZED SEIZURE (FINDING)
C0234533|T047|246545002|SNOMEDCT_US|GENERALISED FIT|GENERALIZED SEIZURE (FINDING)
C0234533|T047|246545002|SNOMEDCT_US|GENERALIZED FIT|GENERALIZED SEIZURE (FINDING)
C0234533|T047|246545002|SNOMEDCT_US|GENERALIZED SEIZURE |GENERALIZED SEIZURE (FINDING)
C0234533|T047|246545002|SNOMEDCT_US|CONVULSIONS; GENERALIZED|GENERALIZED SEIZURE (FINDING)
C0234533|T047|246545002|SNOMEDCT_US|GENERALIZED; CONVULSIONS|GENERALIZED SEIZURE (FINDING)
C0234533|T047|246545002|SNOMEDCT_US|GENERALIZED CONVULSION, NOS|GENERALIZED SEIZURE (FINDING)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPSIES|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPSY|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPSY, UNSPECIFIED|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPTIC SEIZURE|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|SEIZURE, EPILEPTIC|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|SEIZURE DISORDER NOS|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|SEIZURE DISORDER|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|SEIZURE DIS|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPSIA|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPSY |(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|SEIZURE DISORDER |(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|SEIZURE DISORDERS|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPTIC CONVULSIONS NOS|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPTIC FITS NOS|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPSY NOS|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPTIC SEIZURES NOS|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPSY [DISEASE/FINDING]|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPTIC SEIZURES|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|SEIZURES, EPILEPTIC|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|SEIZURE;EPILEPTIC|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPTIC ATTACK|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPSY NOS |(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|(EPILEPSY) OR (EPILEPTIC ATTACK) |(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|(EPILEPSY) OR |(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|ATTACK - EPILEPTIC|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPTIC FIT|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EF - EPILEPTIC FIT|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EP - EPILEPSY|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPTIC|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPSY |(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPTIC CONVULSIONS|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPTIC DISORDER|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPTIC FITS|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPTIC SEIZURE |(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|SEIZURE DISORDER |(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|CADUCUS; MORBUS|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|CEREBRAL; EPILEPTIC|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|CONVULSIONS; EPILEPTIC|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPSY; CEREBRAL|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPSY; CORTICAL|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPSY; FIT|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPSY; SEIZURE|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPTIC; CONVULSIONS|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPTIC; SYNDROME|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|FIT; EPILEPTIC|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|MORBUS; CADUCUS|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|SEIZURE; EPILEPTIC|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|SYNDROME; EPILEPTIC|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILECTIC ATTACK, NOS|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPSY, NOS|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPTIC CONVULSIONS, NOS|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPTIC DISORDER, NOS|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPTIC FITS, NOS|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPTIC SEIZURES, NOS|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0014544|T047|267698007|SNOMEDCT_US|EPILEPTIC ATTACK, NOS|(EPILEPSY) OR (EPILEPTIC ATTACK) (DISORDER)
C0270850|T047|36803009|SNOMEDCT_US|GENERALIZED IDIOPATHIC EPILEPSY AND EPILEPTIC SYNDROMES|IDIOPATHIC GENERALIZED EPILEPSY (DISORDER)
C0270850|T047|36803009|SNOMEDCT_US|EPILEPSY, IDIOPATHIC GENERALIZED|IDIOPATHIC GENERALIZED EPILEPSY (DISORDER)
C0270850|T047|36803009|SNOMEDCT_US|IDIOPATHIC GENERALIZED EPILEPSY|IDIOPATHIC GENERALIZED EPILEPSY (DISORDER)
C0270850|T047|36803009|SNOMEDCT_US|GENERALIZED IDIOPATHIC EPILEPSY AND EPILEPTIC SYNDROMES NOS|IDIOPATHIC GENERALIZED EPILEPSY (DISORDER)
C0270850|T047|36803009|SNOMEDCT_US|IDIOPATHIC GENERALISED EPILEPSY|IDIOPATHIC GENERALIZED EPILEPSY (DISORDER)
C0270850|T047|36803009|SNOMEDCT_US|EPILEPSY GENERALIZED IDIOPATHIC|IDIOPATHIC GENERALIZED EPILEPSY (DISORDER)
C0270850|T047|36803009|SNOMEDCT_US|EPILEPSY GENERALIZED IDIOPATHIC |IDIOPATHIC GENERALIZED EPILEPSY (DISORDER)
C0270850|T047|36803009|SNOMEDCT_US|PRIMARY GENERALISED EPILEPSY|IDIOPATHIC GENERALIZED EPILEPSY (DISORDER)
C0270850|T047|36803009|SNOMEDCT_US|PRIMARY GENERALIZED EPILEPSY|IDIOPATHIC GENERALIZED EPILEPSY (DISORDER)
C0270850|T047|36803009|SNOMEDCT_US|IDIOPATHIC GENERALIZED EPILEPSY |IDIOPATHIC GENERALIZED EPILEPSY (DISORDER)
C0270850|T047|36803009|SNOMEDCT_US|EPILEPSY; GENERALIZED, IDIOPATHIC|IDIOPATHIC GENERALIZED EPILEPSY (DISORDER)
C0270850|T047|36803009|SNOMEDCT_US|EPILEPSY; IDIOPATHIC, GENERALIZED|IDIOPATHIC GENERALIZED EPILEPSY (DISORDER)
C0270850|T047|36803009|SNOMEDCT_US|EPILEPSY; SYNDROME, GENERALIZED, IDIOPATHIC|IDIOPATHIC GENERALIZED EPILEPSY (DISORDER)
C0270850|T047|36803009|SNOMEDCT_US|GENERALIZED; EPILEPTIC, IDIOPATHIC|IDIOPATHIC GENERALIZED EPILEPSY (DISORDER)
C0270850|T047|36803009|SNOMEDCT_US|SYNDROME; EPILEPTIC, GENERALIZED, IDIOPATHIC|IDIOPATHIC GENERALIZED EPILEPSY (DISORDER)
C0270850|T047|36803009|SNOMEDCT_US|IDIOPATHIC GENERALIZED EPILEPSY, NOS|IDIOPATHIC GENERALIZED EPILEPSY (DISORDER)
C0494475|T047|65155005|SNOMEDCT_US|GRAND MAL SEIZURES, UNSPECIFIED (WITH OR WITHOUT PETIT MAL)|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|GENERALIZED TONIC-CLONIC SEIZURE|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|GRAND MAL SEIZURE|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|GRAND MAL|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|GRAND-MAL SEIZURE|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|GENERALIZED TONIC CLONIC SEIZURES|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|GENERALIZED TONIC-CLONIC SEIZURES|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|SEIZURES, GENERALIZED TONIC-CLONIC|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|GENERALIZED CLONIC-TONIC SEIZURES|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|SEIZURES, TONIC-CLONIC|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|GENERALIZED TONIC-CLONIC SEIZURES (GTCS)|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|GENERALISED TONIC-CLONIC SEIZURES|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|SEIZURE, TONIC-CLONIC|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|SEIZURES, TONIC CLONIC|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|TONIC-CLONIC SEIZURE|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|TONIC-CLONIC SEIZURES|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|SEIZURES, CLONIC-TONIC|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|SEIZURE;TONIC-CLONIC|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|GRAND MAL SEIZURES|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|GRAND MAL SEIZURE NOS|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|SEIZURES, GENERALIZED TONIC-CLONIC (GTCS)|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|GRAND MAL SEIZURE |GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|GRAND MAL CONVULSION|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|GRAND MAL SEIZURE |GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|GENERALISED TONIC-CLONIC SEIZURE|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|SEIZURES, GRAND-MAL|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|GRAND-MAL SEIZURES|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|SEIZURES, GENERALIZED, TONIC-CLONIC|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|GRAND MAL EPILEPTIC FIT|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|GRAND MAL FIT|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|SEIZURE GRAND MAL|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|TONIC-CLONIC SEIZURE (PHYSICAL FINDING)|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|SEIZURE GENERALIZED TONIC-CLONIC|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|TONIC-CLONIC CONVULSION|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|TONIC-CLONIC CONVULSIONS|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|TONIC-CLONIC SEIZURE |GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|TONIC - CLONIC SEIZURES|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|GRAND MAL; SEIZURE|GRAND MAL SEIZURE (FINDING)
C0494475|T047|65155005|SNOMEDCT_US|SEIZURE; GRAND MAL|GRAND MAL SEIZURE (FINDING)
C0475521|T047|193022009|SNOMEDCT_US|LOCALIZATION-RELATED (FOCAL) (PARTIAL) IDIOPATHIC EPILEPSY AND EPILEPTIC SYNDROMES WITH SEIZURES OF LOCALIZED ONSET|LOCALIZATION-RELATED(FOCAL)(PARTIAL)IDIOPATHIC EPILEPSY AND EPILEPTIC SYNDROMES WITH SEIZURES OF LOCALIZED ONSET (DISORDER)
C0475521|T047|193022009|SNOMEDCT_US|LOCALIZATION-RELATED (FOCAL) (PARTIAL) IDIOPATHIC EPILEPSY AND EPILEPTIC SYNDROMES WITH SEIZURES OF LOCALIZED ONSET NOS|LOCALIZATION-RELATED(FOCAL)(PARTIAL)IDIOPATHIC EPILEPSY AND EPILEPTIC SYNDROMES WITH SEIZURES OF LOCALIZED ONSET (DISORDER)
C0475521|T047|193022009|SNOMEDCT_US|LOCALIZATION-RELATED(FOCAL)(PARTIAL)IDIOPATHIC EPILEPSY AND EPILEPTIC SYNDROMES WITH SEIZURES OF LOCALISED ONSET|LOCALIZATION-RELATED(FOCAL)(PARTIAL)IDIOPATHIC EPILEPSY AND EPILEPTIC SYNDROMES WITH SEIZURES OF LOCALIZED ONSET (DISORDER)
C0475521|T047|193022009|SNOMEDCT_US|LOCALIZATION-RELATED(FOCAL)(PARTIAL)IDIOPATHIC EPILEPSY AND EPILEPTIC SYNDROMES WITH SEIZURES OF LOCALIZED ONSET|LOCALIZATION-RELATED(FOCAL)(PARTIAL)IDIOPATHIC EPILEPSY AND EPILEPTIC SYNDROMES WITH SEIZURES OF LOCALIZED ONSET (DISORDER)
C0475521|T047|193022009|SNOMEDCT_US|LOCALIZATION-RELATED(FOCAL)(PARTIAL)IDIOPATHIC EPILEPSY AND EPILEPTIC SYNDROMES WITH SEIZURES OF LOCALIZED ONSET |LOCALIZATION-RELATED(FOCAL)(PARTIAL)IDIOPATHIC EPILEPSY AND EPILEPTIC SYNDROMES WITH SEIZURES OF LOCALIZED ONSET (DISORDER)
C0494472|T047||SNOMEDCT_US|LOCALIZATION-RELATED (FOCAL) (PARTIAL) SYMPTOMATIC EPILEPSY AND EPILEPTIC SYNDROMES WITH COMPLEX PARTIAL SEIZURES
C0494472|T047||SNOMEDCT_US|LOCALIZATION-RELATED (FOCAL) (PARTIAL) SYMPTOMATIC EPILEPSY AND EPILEPTIC SYNDROMES WITH COMPLEX PARTIAL SEIZURES NOS
C0494471|T047||SNOMEDCT_US|LOCALIZATION-RELATED (FOCAL) (PARTIAL) SYMPTOMATIC EPILEPSY AND EPILEPTIC SYNDROMES WITH SIMPLE PARTIAL SEIZURES
C0494471|T047||SNOMEDCT_US|LOCALIZATION-RELATED (FOCAL) (PARTIAL) SYMPTOMATIC EPILEPSY AND EPILEPTIC SYNDROMES WITH SIMPLE PARTIAL SEIZURES NOS
C0477371|T047|194491006|SNOMEDCT_US|OTHER FORMS OF EPILEPSY|[X]OTHER EPILEPSY (DISORDER)
C0477371|T047|194491006|SNOMEDCT_US|OTHER EPILEPSY|[X]OTHER EPILEPSY (DISORDER)
C0477371|T047|194491006|SNOMEDCT_US|OTHER EPILEPSY NOS|[X]OTHER EPILEPSY (DISORDER)
C0477371|T047|194491006|SNOMEDCT_US|OTHER FORMS OF EPILEPSY NOS |[X]OTHER EPILEPSY (DISORDER)
C0477371|T047|194491006|SNOMEDCT_US|OTHER FORMS OF EPILEPSY |[X]OTHER EPILEPSY (DISORDER)
C0477371|T047|194491006|SNOMEDCT_US|OTHER FORMS OF EPILEPSY NOS|[X]OTHER EPILEPSY (DISORDER)
C0477371|T047|194491006|SNOMEDCT_US|[X]OTHER EPILEPSY|[X]OTHER EPILEPSY (DISORDER)
C0477371|T047|194491006|SNOMEDCT_US|[X]OTHER EPILEPSY |[X]OTHER EPILEPSY (DISORDER)
C0477370|T047|194490007|SNOMEDCT_US|OTHER GENERALIZED EPILEPSY AND EPILEPTIC SYNDROMES|[X]OTHER GENERALIZED EPILEPSY AND EPILEPTIC SYNDROMES (DISORDER)
C0477370|T047|194490007|SNOMEDCT_US|OTHER GENERALIZED EPILEPSY AND EPILEPTIC SYNDROMES NOS|[X]OTHER GENERALIZED EPILEPSY AND EPILEPTIC SYNDROMES (DISORDER)
C0477370|T047|194490007|SNOMEDCT_US|[X]OTHER GENERALIZED EPILEPSY AND EPILEPTIC SYNDROMES |[X]OTHER GENERALIZED EPILEPSY AND EPILEPTIC SYNDROMES (DISORDER)
C0477370|T047|194490007|SNOMEDCT_US|[X]OTHER GENERALIZED EPILEPSY AND EPILEPTIC SYNDROMES|[X]OTHER GENERALIZED EPILEPSY AND EPILEPTIC SYNDROMES (DISORDER)
C0477370|T047|194490007|SNOMEDCT_US|[X]OTHER GENERALISED EPILEPSY AND EPILEPTIC SYNDROMES|[X]OTHER GENERALIZED EPILEPSY AND EPILEPTIC SYNDROMES (DISORDER)
C0477370|T047|194490007|SNOMEDCT_US|SYNDROME; EPILEPTIC, GENERALIZED|[X]OTHER GENERALIZED EPILEPSY AND EPILEPTIC SYNDROMES (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|ABSENCE EPILEPSY|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|EPILEPSY, ABSENCE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|PETIT MAL EPILEPSIES|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|PYKNOLEPSIES|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|SEIZURE, ABSENCE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|ABSENCE SEIZURE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|ABSENCE SEIZURES|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|PETIT MAL, UNSPECIFIED, WITHOUT GRAND MAL SEIZURES|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|PETIT MAL SEIZURE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|PETIT MAL|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|PETIT-MAL SEIZURE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|SEIZURES, ABSENCE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|ABSENCE SEIZURE DIS|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|SEIZURE DIS ABSENCE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|PYKNOLEPSY|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|EPILEPSY GENERALIZED NONCONVULSIVE PYKNO-EPILEPSY |PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|EPILEPSY GENERALIZED NONCONVULSIVE PYKNO-EPILEPSY|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|GENERALIZED NONCONVULSIVE PETIT MAL SEIZURE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|PETIT MAL SEIZURE |PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|PYKNO-EPILEPSY|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|PETIT MAL EPILEPSY|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|ABSENCE SEIZURE DISORDERS|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|SEIZURE DISORDERS, ABSENCE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|CONVULSION, PETIT MAL|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|MINOR EPILEPSIES|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|MINOR EPILEPSY|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|PYKNO EPILEPSY|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|PYKNO-EPILEPSIES|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|CHILDHOOD ABSENCE SEIZURES|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|EPILEPSY, MINOR|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|EPILEPSY, ABSENCE [DISEASE/FINDING]|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|JUVENILE ABSENCE EPILEPSY|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|CHILDHOOD ABSENCE EPILEPSY|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|ABSENCE SEIZURE DISORDER|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|EPILEPSY, PETIT MAL|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|PETIT MAL CONVULSION|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|SEIZURE DISORDER, ABSENCE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|SEIZURE;ABSENCE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|TYPICAL ABSENCE SEIZURE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|TYPICAL ABSENCE SEIZURE |PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|EPILEPSY JUVENILE ABSENCES|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|JUVENILE ABSENCES, EPILEPSY|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|JUVENILE ABSENCE, EPILEPSY|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|JUVENILE ABSENCE EPILEPSY |PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|ABSENCE SEIZURE |PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|CHILDHOOD ABSENCE EPILEPSY |PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|PETIT MAL |PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|EPILEPSY JUVENILE ABSENCE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|PETIT-MAL SEIZURES|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|SEIZURES, PETIT-MAL|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|PETIT MAL SEIZURES|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|TYPICAL ABSENCE SEIZURES|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|CONVULSION PETIT MAL|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|EPILEPSY PETIT MAL|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|SEIZURE GENERALIZED ABSENCE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|ABSENCE SEIZURE (PHYSICAL FINDING)|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|CHILDHOOD ABSENCE SEIZURE |PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|JUVENILE ABSENCE SEIZURE |PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|JUVENILE ABSENCE SEIZURE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|CHILDHOOD ABSENCE SEIZURE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|CHILDHOOD - JUVENILE - ABSENCE EPILEPSY|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|PETIT-MAL EPILEPSY|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|ABSENCE SEIZURE |PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|EPILEPSY; ABSENCE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|EPILEPSY; MINOR|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|EPILEPSY; PETIT MAL|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|ABSENCE; EPILEPTIC|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|ABSENCES; EPILEPTIC|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|PETIT MAL; EPILEPSY|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|ABSENCE EPILEPSIES, CHILDHOOD|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|ABSENCE EPILEPSY, CHILDHOOD|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|CHILDHOOD ABSENCE EPILEPSIES|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|EPILEPSIES, CHILDHOOD ABSENCE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|EPILEPSY, CHILDHOOD ABSENCE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|ABSENCE EPILEPSIES, JUVENILE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|ABSENCE EPILEPSY, JUVENILE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|EPILEPSIES, JUVENILE ABSENCE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|EPILEPSY, JUVENILE ABSENCE|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|JUVENILE ABSENCE EPILEPSIES|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|ABSENCES, TYPICAL|PETIT MAL (DISORDER)
C0014553|T047|16757004|SNOMEDCT_US|ABSENCE OF SEIZURE|PETIT MAL (DISORDER)
C0494474|T047||SNOMEDCT_US|SPECIAL EPILEPTIC SYNDROMES
C0494474|T047||SNOMEDCT_US|EPILEPSY; SYNDROME, SPECIAL
C0494474|T047||SNOMEDCT_US|EPILEPTIC; SYNDROME, SPECIAL
C0494474|T047||SNOMEDCT_US|SYNDROME; EPILEPTIC, SPECIAL
C0014547|T047|67139004|SNOMEDCT_US|EPILEPSIES, FOCAL|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|EPILEPSIES, LOCALIZATION-RELATED|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|EPILEPSIES, PARTIAL|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|FOCAL EPILEPSIES|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|FOCAL EPILEPSY|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|LOCALIZATION-RELATED EPILEPSIES|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|LOCALIZATION-RELATED EPILEPSY|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|PARTIAL EPILEPSIES|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|FOCAL SEIZURE DIS|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|PARTIAL SEIZURE DIS|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|SEIZURE DIS PARTIAL|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|EPILEPSY LOCALIZATION RELAT|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|SEIZURE DIS FOCAL|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|LOCALIZATION-RELATED EPILEPSY -RETIRED-|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|LOCALISATION-RELATED EPILEPSY -RETIRED-|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|DISORDERS, FOCAL SEIZURE|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|FOCAL SEIZURE DISORDERS|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|SEIZURE DISORDERS, FOCAL|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|DISORDERS, PARTIAL SEIZURE|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|PARTIAL SEIZURE DISORDERS|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|SEIZURE DISORDERS, PARTIAL|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|EPILEPSIES, PARTIAL [DISEASE/FINDING]|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|EPILEPSY, PARTIAL|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|FOCAL SEIZURE DISORDER|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|SEIZURE DISORDER, FOCAL|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|EPILEPSY, FOCAL|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|EPILEPSY, LOCALIZATION-RELATED|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|SEIZURE DISORDER, PARTIAL|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|PARTIAL EPILEPSY|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|PARTIAL SEIZURE DISORDER|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|LOCALISATION-RELATED EPILEPSY|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|LOCALISATION-RELATED EPILEPSY |LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|LOCALIZATION-RELATED EPILEPSY |LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|LOCALISATION RELATED EPILEPSY|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|LOCALIZATION RELATED EPILEPSY|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|LOCAL EPILEPSY|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|EPILEPSY; FOCAL|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|EPILEPSY; LOCALIZATION-RELATED|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|EPILEPSY; PARTIAL|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|FOCAL; EPILEPTIC|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|PARTIAL; EPILEPTIC|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|FOCAL EPILEPSY, NOS|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|LOCALIZATION-RELATED EPILEPSY, NOS|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|EPILEPSY, FOCAL NOS|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014547|T047|67139004|SNOMEDCT_US|EPILEPSY, PARTIAL NOS|LOCALIZATION-RELATED EPILEPSY -RETIRED-
C0014548|T047|19598007|SNOMEDCT_US|EPILEPSIES, GENERALIZED|GENERALIZED EPILEPSY (DISORDER)
C0014548|T047|19598007|SNOMEDCT_US|EPILEPSY, GENERALIZED|GENERALIZED EPILEPSY (DISORDER)
C0014548|T047|19598007|SNOMEDCT_US|GENERALIZED EPILEPSIES|GENERALIZED EPILEPSY (DISORDER)
C0014548|T047|19598007|SNOMEDCT_US|GENERALIZED EPILEPSY|GENERALIZED EPILEPSY (DISORDER)
C0014548|T047|19598007|SNOMEDCT_US|SEIZURE DIS GENERALIZED|GENERALIZED EPILEPSY (DISORDER)
C0014548|T047|19598007|SNOMEDCT_US|GENERALIZED SEIZURE DISORDER|GENERALIZED EPILEPSY (DISORDER)
C0014548|T047|19598007|SNOMEDCT_US|GENERALIZED SEIZURE DISORDERS|GENERALIZED EPILEPSY (DISORDER)
C0014548|T047|19598007|SNOMEDCT_US|SEIZURE DISORDERS, GENERALIZED|GENERALIZED EPILEPSY (DISORDER)
C0014548|T047|19598007|SNOMEDCT_US|EPILEPSY, GENERALIZED [DISEASE/FINDING]|GENERALIZED EPILEPSY (DISORDER)
C0014548|T047|19598007|SNOMEDCT_US|SEIZURE DISORDER, GENERALIZED|GENERALIZED EPILEPSY (DISORDER)
C0014548|T047|19598007|SNOMEDCT_US|EPILEPSY GENERALIZED|GENERALIZED EPILEPSY (DISORDER)
C0014548|T047|19598007|SNOMEDCT_US|GENERALIZED EPILEPSY |GENERALIZED EPILEPSY (DISORDER)
C0014548|T047|19598007|SNOMEDCT_US|GENERALISED EPILEPSY |GENERALIZED EPILEPSY (DISORDER)
C0014548|T047|19598007|SNOMEDCT_US|GENERALISED EPILEPSY|GENERALIZED EPILEPSY (DISORDER)
C0014548|T047|19598007|SNOMEDCT_US|GENERALIZED EPILEPSY |GENERALIZED EPILEPSY (DISORDER)
C0014548|T047|19598007|SNOMEDCT_US|EPILEPSY; GENERALIZED|GENERALIZED EPILEPSY (DISORDER)
C0014548|T047|19598007|SNOMEDCT_US|EPILEPSY; SYNDROME, GENERALIZED|GENERALIZED EPILEPSY (DISORDER)
C0014548|T047|19598007|SNOMEDCT_US|GENERALIZED; EPILEPTIC|GENERALIZED EPILEPSY (DISORDER)
C0014548|T047|19598007|SNOMEDCT_US|GENERALIZED EPILEPSY, NOS|GENERALIZED EPILEPSY (DISORDER)
C0014548|T047|19598007|SNOMEDCT_US|GENERALISED EPILEPSY [AMBIGUOUS]|GENERALIZED EPILEPSY (DISORDER)
C0014550|T047||SNOMEDCT_US|EPILEPSIES, MYOCLONIC
C0014550|T047||SNOMEDCT_US|EPILEPSY, MYOCLONIC
C0014550|T047||SNOMEDCT_US|MYOCLONIC EPILEPSIES
C0014550|T047||SNOMEDCT_US|MYOCLONUS EPILEPSIES
C0014550|T047||SNOMEDCT_US|MYOCLONUS EPILEPSY
C0014550|T047||SNOMEDCT_US|SEIZURES, MYOCLONIC
C0014550|T047||SNOMEDCT_US|MYOCLONIC SEIZURES
C0014550|T047||SNOMEDCT_US|MYOCLONIC EPILEPSY
C0014550|T047||SNOMEDCT_US|MYOCLONIC SEIZURE DIS
C0014550|T047||SNOMEDCT_US|MYOCLONIA EPILEPTICA
C0014550|T047||SNOMEDCT_US|MYOCLONIC SEIZURE
C0014550|T047||SNOMEDCT_US|MYOCLONIC SEIZURE DISORDER
C0014550|T047||SNOMEDCT_US|MYOCLONIC EPILEPSY 
C0014550|T047||SNOMEDCT_US|GENERALIZED CONVULSIVE MYOCLONIC SEIZURE
C0014550|T047||SNOMEDCT_US|DISORDER, MYOCLONIC SEIZURE
C0014550|T047||SNOMEDCT_US|DISORDERS, MYOCLONIC SEIZURE
C0014550|T047||SNOMEDCT_US|MYOCLONIC SEIZURE DISORDERS
C0014550|T047||SNOMEDCT_US|SEIZURE DISORDER, MYOCLONIC
C0014550|T047||SNOMEDCT_US|SEIZURE DISORDERS, MYOCLONIC
C0014550|T047||SNOMEDCT_US|EPILEPSIES, MYOCLONIC [DISEASE/FINDING]
C0014550|T047||SNOMEDCT_US|EPILEPSY, MYOCLONUS
C0014550|T047||SNOMEDCT_US|SEIZURE;MYOCLONIC
C0014550|T047||SNOMEDCT_US|MYOCLONIC SEIZURE NOS
C0014550|T047||SNOMEDCT_US|SEIZURE GENERALIZED MYOCLONIC
C0014550|T047||SNOMEDCT_US|MYOCLONIC SEIZURE (PHYSICAL FINDING)
C0014550|T047||SNOMEDCT_US|EPILEPTIC SEIZURES - MYOCLONIC
C0014550|T047||SNOMEDCT_US|EPILEPTIC SEIZURES - MYOCLONIC 
C0014550|T047||SNOMEDCT_US|MYOCLONIC SEIZURE 
C0014550|T047||SNOMEDCT_US|EPILEPSY; MYOCLONUS
C0014550|T047||SNOMEDCT_US|EPILEPTICA; MYOCLONUS
C0014550|T047||SNOMEDCT_US|EPILEPTIC SEIZURES, MYOCLONIC
C0014557|T047|157437008|SNOMEDCT_US|EPILEPSIES, POST-TRAUMATIC|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|EPILEPSIES, TRAUMATIC|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|EPILEPSY, POST TRAUMATIC|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|EPILEPSY, POST-TRAUMATIC|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|POST-TRAUMATIC EPILEPSIES|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|POST-TRAUMATIC EPILEPSY|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|TRAUMATIC EPILEPSIES|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|TRAUMATIC EPILEPSY|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|SEIZURE DIS POST TRAUMATIC|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|POST TRAUMATIC SEIZURE DIS|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|DISORDER, POST-TRAUMATIC SEIZURE|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|DISORDERS, POST-TRAUMATIC SEIZURE|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|POST TRAUMATIC SEIZURE DISORDER|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|POST-TRAUMATIC SEIZURE DISORDERS|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|SEIZURE DISORDER, POST TRAUMATIC|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|SEIZURE DISORDERS, POST-TRAUMATIC|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|EPILEPSY, POST-TRAUMATIC [DISEASE/FINDING]|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|POST-TRAUMATIC SEIZURE DISORDER|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|EPILEPSY, TRAUMATIC|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|SEIZURE DISORDER, POST-TRAUMATIC|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|TRAUMATIC EPILEPSY |TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|PTE - POST-TRAUMATIC EPILEPSY|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|POST-TRAUMATIC EPILEPSY |TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|EPILEPSY; TRAUMATIC|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T047|157437008|SNOMEDCT_US|TRAUMATIC; EPILEPTIC|TRAUMATIC EPILEPSY (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|SEIZURE|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|CONVULSIONS|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|SEIZURES|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|CONVULSION|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|[D]CONVULSION NOS (CONTEXT-DEPENDENT CATEGORY)|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|[D]CONVULSIONS (CONTEXT-DEPENDENT CATEGORY)|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|[D]FIT (CONTEXT-DEPENDENT CATEGORY)|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|SEIZURE NOS|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|SEIZURE (PHYSICAL FINDING)|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|CONVULSIONS |FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|FIT, NOS|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|SEIZURE, NOS|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|CONVULSION, NOS|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|UNSPECIFIED CONVULSIONS|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|FIT NOS|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|SEIZURES [DISEASE/FINDING]|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|FIT(S)|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|FITS - CONVULSIONS|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|[D]CONVULSIONS|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|[D]CONVULSIONS |FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|[D]FIT |FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|[D]FIT|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|[D]CONVULSION NOS|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|FITS - CONVULSIONS |FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|[D]CONVULSION NOS |FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|[D]SEIZURE NOS|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|FIT - CONVULSION |FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|FIT|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|FIT - CONVULSION|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|CONVULSION |FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|FITTING|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|CONVULSION (NOS)|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|FITS NOS|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|CONVULSIONS NOS|FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|SEIZURE |FITS - CONVULSIONS (DISORDER)
C0036572|T047|313290005|SNOMEDCT_US|FITS|FITS - CONVULSIONS (DISORDER)
C0038220|T047|230456007|SNOMEDCT_US|STATUS EPILEPTICUS|STATUS EPILEPTICUS (DISORDER)
C0038220|T047|230456007|SNOMEDCT_US|STATUS EPILEPTICUS, UNSPECIFIED|STATUS EPILEPTICUS (DISORDER)
C0038220|T047|230456007|SNOMEDCT_US|GENERALIZED STATUS EPILEPTICUS|STATUS EPILEPTICUS (DISORDER)
C0038220|T047|230456007|SNOMEDCT_US|STATUS EPILEPTICUS [DISEASE/FINDING]|STATUS EPILEPTICUS (DISORDER)
C0038220|T047|230456007|SNOMEDCT_US|STATUS EPILEPTICUS, GENERALIZED|STATUS EPILEPTICUS (DISORDER)
C0038220|T047|230456007|SNOMEDCT_US|[X]STATUS EPILEPTICUS, UNSPECIFIED |STATUS EPILEPTICUS (DISORDER)
C0038220|T047|230456007|SNOMEDCT_US|[X]STATUS EPILEPTICUS, UNSPECIFIED|STATUS EPILEPTICUS (DISORDER)
C0038220|T047|230456007|SNOMEDCT_US|STATUS EPILEPTICUS |STATUS EPILEPTICUS (DISORDER)
C0038220|T047|230456007|SNOMEDCT_US|EPILEPSY; STATUS|STATUS EPILEPTICUS (DISORDER)
C0038220|T047|230456007|SNOMEDCT_US|EPILEPTICUS; STATUS|STATUS EPILEPTICUS (DISORDER)
C0038220|T047|230456007|SNOMEDCT_US|STATUS; EPILEPTICUS|STATUS EPILEPTICUS (DISORDER)
C0038220|T047|230456007|SNOMEDCT_US|STATUS; EPILEPTIC|STATUS EPILEPTICUS (DISORDER)
C0038220|T047|230456007|SNOMEDCT_US|STATUS EPILEPTICUS NOS|STATUS EPILEPTICUS (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|ACQUIRED EPILEPTIC APHASIA|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|ACQUIRED EPILEPTIC APHASIAS|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|EPILEPTIC APHASIA, ACQUIRED|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|EPILEPTIC APHASIAS, ACQUIRED|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|LANDAU KLEFFNER SYNDROME|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|LANDAU-KLEFFNER SYNDROME|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|SYNDROME, LANDAU-KLEFFNER|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|ACQUIRED APHASIA WITH EPILEPSY [LANDAU-KLEFFNER]|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|ACQUIRED CHILDHOOD APHASIA WITH CONVULSIVE DIS|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|ACQUIRED CHILDHOOOD APHASIA WITH CONVULSIVE DISORDER|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|APHASIA, EPILEPTIC, ACQUIRED|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|LANDAU-KLEFFNER ACQUIRED EPILEPTIFORM APHASIA|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|APHASIA, ACQUIRED EPILEPTIC|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|LANDAU-KLEFFNER SYNDROME [DISEASE/FINDING]|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|ACQUIRED EPILEPTIFORM APHASIAS|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|EPILEPTIFORM APHASIAS, ACQUIRED|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|EPILEPTIFORM APHASIA, ACQUIRED|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|ACQUIRED APHASIA WITH CONVULSIVE DISORDER|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|ACQUIRED EPILEPTIFORM APHASIA|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|LANDAU KLEFFNER ACQUIRED EPILEPTIFORM APHASIA|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|APHASIA, ACQUIRED, WITH CONVULSIVE DISORDER|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|ACQUIRED APHASIA WITH EPILEPSY|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|ACQUIRED EPILEPTIC APHASIA |ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|ACQUIRED EPILEPTIC APHASIA |ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0282512|T047|230438007|SNOMEDCT_US|DEVELOPMENTAL DISORDER - SPEECH ACQUIRED EPILEPTIC APHASIA|ACQUIRED EPILEPTIC APHASIA (DISORDER)
C0270857|T047|79745005|SNOMEDCT_US|EPILEPSIES, REFLEX|REFLEX EPILEPSY (DISORDER)
C0270857|T047|79745005|SNOMEDCT_US|EPILEPSY, REFLEX|REFLEX EPILEPSY (DISORDER)
C0270857|T047|79745005|SNOMEDCT_US|REFLEX EPILEPSIES|REFLEX EPILEPSY (DISORDER)
C0270857|T047|79745005|SNOMEDCT_US|REFLEX EPILEPSY|REFLEX EPILEPSY (DISORDER)
C0270857|T047|79745005|SNOMEDCT_US|EPILEPSY, REFLEX [DISEASE/FINDING]|REFLEX EPILEPSY (DISORDER)
C0270857|T047|79745005|SNOMEDCT_US|EPILEPSY ASSOCIATED WITH SPECIFIC STIMULI|REFLEX EPILEPSY (DISORDER)
C0270857|T047|79745005|SNOMEDCT_US|SENSORY-INDUCED EPILEPSY|REFLEX EPILEPSY (DISORDER)
C0270857|T047|79745005|SNOMEDCT_US|REFLEX EPILEPSY |REFLEX EPILEPSY (DISORDER)
C0270857|T047|79745005|SNOMEDCT_US|EPILEPSY; REFLEX|REFLEX EPILEPSY (DISORDER)
C0270857|T047|79745005|SNOMEDCT_US|EPILEPSY, SENSORY-INDUCED|REFLEX EPILEPSY (DISORDER)
C0270851|T047|276724002|SNOMEDCT_US|BENIGN NEONATAL CONVULSION|BENIGN NEONATAL SEIZURES (DISORDER)
C0270851|T047|276724002|SNOMEDCT_US|CONVULSION, BENIGN NEONATAL|BENIGN NEONATAL SEIZURES (DISORDER)
C0270851|T047|276724002|SNOMEDCT_US|CONVULSIONS, BENIGN NEONATAL|BENIGN NEONATAL SEIZURES (DISORDER)
C0270851|T047|276724002|SNOMEDCT_US|NEONATAL CONVULSION, BENIGN|BENIGN NEONATAL SEIZURES (DISORDER)
C0270851|T047|276724002|SNOMEDCT_US|BENIGN NEONATAL EPILEPSIES|BENIGN NEONATAL SEIZURES (DISORDER)
C0270851|T047|276724002|SNOMEDCT_US|EPILEPSIES, BENIGN NEONATAL|BENIGN NEONATAL SEIZURES (DISORDER)
C0270851|T047|276724002|SNOMEDCT_US|EPILEPSY, BENIGN NEONATAL|BENIGN NEONATAL SEIZURES (DISORDER)
C0270851|T047|276724002|SNOMEDCT_US|NEONATAL EPILEPSIES, BENIGN|BENIGN NEONATAL SEIZURES (DISORDER)
C0270851|T047|276724002|SNOMEDCT_US|NEONATAL EPILEPSY, BENIGN|BENIGN NEONATAL SEIZURES (DISORDER)
C0270851|T047|276724002|SNOMEDCT_US|BENIGN NEONATAL EPILEPSY|BENIGN NEONATAL SEIZURES (DISORDER)
C0270851|T047|276724002|SNOMEDCT_US|NEONATAL CONVULSIONS, BENIGN|BENIGN NEONATAL SEIZURES (DISORDER)
C0270851|T047|276724002|SNOMEDCT_US|BENIGN NEONATAL CONVULSIONS|BENIGN NEONATAL SEIZURES (DISORDER)
C0270851|T047|276724002|SNOMEDCT_US|EPILEPSY, BENIGN NEONATAL [DISEASE/FINDING]|BENIGN NEONATAL SEIZURES (DISORDER)
C0270851|T047|276724002|SNOMEDCT_US|BENIGN NEONATAL SEIZURES|BENIGN NEONATAL SEIZURES (DISORDER)
C0270851|T047|276724002|SNOMEDCT_US|BENIGN NEONATAL SEIZURES |BENIGN NEONATAL SEIZURES (DISORDER)
C0270851|T047|276724002|SNOMEDCT_US|BENIGN NEONATAL CONVULSIONS |BENIGN NEONATAL SEIZURES (DISORDER)
C0270851|T047|276724002|SNOMEDCT_US|BENIGN NEONATAL SEIZURES [AMBIGUOUS]|BENIGN NEONATAL SEIZURES (DISORDER)
C1856931|T047||SNOMEDCT_US|EPILEPSY, PHOTOGENIC, WITH SPASTIC DIPLEGIA AND MENTAL RETARDATION
C1856930|T047||SNOMEDCT_US|EPILEPSY WITH BILATERAL OCCIPITAL CALCIFICATIONS
C1856930|T047||SNOMEDCT_US|EPILEPSY OCCIPITAL CALCIFICATIONS
C1856930|T047||SNOMEDCT_US|BILATERAL OCCIPITAL CALCIFICATIONS WITH EPILEPSY
C1856930|T047||SNOMEDCT_US|FAMILIAL UNILATERAL AND BILATERAL OCCIPITAL CALCIFICATIONS AND EPILEPSY
C2584947|T047|438156004|SNOMEDCT_US|ANOXIC EPILEPTIC SEIZURE|ANOXIC EPILEPTIC SEIZURE (FINDING)
C2584947|T047|438156004|SNOMEDCT_US|ANOXIC EPILEPTIC SEIZURE |ANOXIC EPILEPTIC SEIZURE (FINDING)
C0270853|T047|6204001|SNOMEDCT_US|JUVENILE MYOCLONIC EPILEPSY|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|GENERALIZED CONVULSIVE MYOCLONIC SEIZURE, JUVENILE|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|JUVENILE MYOCLONIC EPILEPSY |JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|ADOLESCENT MYOCLONIC EPILEPSIES|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|EPILEPSIES, ADOLESCENT MYOCLONIC|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|EPILEPSY, ADOLESCENT MYOCLONIC|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|MYOCLONIC EPILEPSIES, ADOLESCENT|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|EPILEPSIES, JUVENILE MYOCLONIC|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|EPILEPSY, JUVENILE MYOCLONIC|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|JUVENILE MYOCLONIC EPILEPSIES|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|MYOCLONIC EPILEPSIES, JUVENILE|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|MYOCLONIC EPILEPSY, JUVENILE|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|SYNDROME, JANZ|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|MUCH MORE COMMONLY USED ABBREV.|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|EPILEPSY, MYOCLONIC JUVENILE|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|ADOLESCENT MYOCLONIC EPILEPSY|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|JANZ JUVENILE MYOCLONIC EPILEPSY|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|EPILEPSY, MYOCLONIC, JUVENILE|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|MYOCLONIC EPILEPSY, JUVENILE [DISEASE/FINDING]|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|IMPULSIVE PETIT MAL, JANZ|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|JANZ SYNDROME|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|MYOCLONIC EPILEPSY, ADOLESCENT|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|PETIT MAL, IMPULSIVE, JANZ|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|JUVENILE MYOCLONIC EPILEPSY OF JANZ|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|IMPULSIVE PETIT MAL EPILEPSY|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|JME (JUVENILE MYOCLONIC EPILEPSY)|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|JANZ IMPULSIVE PETIT MAL|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|PETIT MALS, IMPULSIVE|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|MYOCLONIC EPILEPSY, JUVENILE, 1|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|PETIT MAL, IMPULSIVE|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|JMES (JUVENILE MYOCLONIC EPILEPSY)|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|IMPULSIVE PETIT MAL OF JANZ|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|IMPULSIVE PETIT-MAL EPILEPSY|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|MYOCLONIC EPILEPSY OF ADOLESCENCE|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|JME - JUVENILE MYOCLONIC EPILEPSY|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|JUVENILE MYOCLONIC EPILEPSY |JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|IMPULSIVE; PETIT MAL|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C0270853|T047|6204001|SNOMEDCT_US|MYOCLONIC; EPILEPTIC, JUVENILE|JUVENILE MYOCLONIC EPILEPSY (DISORDER)
C1848137|T047||SNOMEDCT_US|EFMR
C1848137|T047||SNOMEDCT_US|EPILEPSY, FEMALE-RESTRICTED, WITH MENTAL RETARDATION 
C1848137|T047||SNOMEDCT_US|EPILEPTIC ENCEPHALOPATHY, EARLY INFANTILE, 9
C1848137|T047||SNOMEDCT_US|EIEE9
C1848137|T047||SNOMEDCT_US|CONVULSIVE DISORDER AND MENTAL RETARDATION
C1848137|T047||SNOMEDCT_US|EPILEPSY, FEMALE-RESTRICTED, WITH MENTAL RETARDATION
C1848137|T047||SNOMEDCT_US|JUBERG-HELLMAN SYNDROME
C2875138|T047||SNOMEDCT_US|EPILEPSY, UNSPECIFIED, NOT INTRACTABLE
C2875141|T047||SNOMEDCT_US|EPILEPSY, UNSPECIFIED, INTRACTABLE
C2919602|T047|445095002|SNOMEDCT_US|EPILEPTIC SEIZURE WITNESSED BY PROVIDER OF HISTORY OTHER THAN SUBJECT|EPILEPTIC SEIZURE WITNESSED BY PROVIDER OF HISTORY OTHER THAN SUBJECT (FINDING)
C2919602|T047|445095002|SNOMEDCT_US|WITNESSED EPILEPTIC SEIZURE|EPILEPTIC SEIZURE WITNESSED BY PROVIDER OF HISTORY OTHER THAN SUBJECT (FINDING)
C2919602|T047|445095002|SNOMEDCT_US|EPILEPTIC SEIZURE WITNESSED BY PROVIDER OF HISTORY OTHER THAN SUBJECT |EPILEPTIC SEIZURE WITNESSED BY PROVIDER OF HISTORY OTHER THAN SUBJECT (FINDING)
C1096063|T047|445355009|SNOMEDCT_US|INTRACTABLE EPILEPSY|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|REFRACTORY EPILEPSY |REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|REFRACTORY EPILEPSY|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|EPILEPSY INTRACTABLE|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|EPILEPSY INTRACTABLE |REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|EPILEPSIES, DRUG RESISTANT|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|INTRACTABLE EPILEPSIES|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|EPILEPSIES, DRUG REFRACTORY|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|RESISTANT EPILEPSY, DRUG|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|MEDICATION RESISTANT EPILEPSIES|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|RESISTANT EPILEPSIES, MEDICATION|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|EPILEPSY, MEDICATION RESISTANT|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|REFRACTORY EPILEPSY, DRUG|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|DRUG RESISTANT EPILEPSY|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|EPILEPSIES, INTRACTABLE|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|DRUG RESISTANT EPILEPSIES|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|RESISTANT EPILEPSIES, DRUG|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|EPILEPSIES, MEDICATION RESISTANT|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|DRUG REFRACTORY EPILEPSIES|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|RESISTANT EPILEPSY, MEDICATION|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|REFRACTORY EPILEPSIES, DRUG|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|EPILEPSY, DRUG REFRACTORY|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|EPILEPSY, DRUG RESISTANT|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|EPILEPSY, INTRACTABLE|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|DRUG REFRACTORY EPILEPSY|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|MEDICATION RESISTANT EPILEPSY|REFRACTORY EPILEPSY (DISORDER)
C1096063|T047|445355009|SNOMEDCT_US|DRUG RESISTANT EPILEPSY [DISEASE/FINDING]|REFRACTORY EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|GENERALIZED NONCONVULSIVE EPILEPSY|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|GENERALIZED SEIZURE DIS NONCONVULSIVE|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|NONCONVULSIVE SEIZURE DIS GENERALIZED|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|SEIZURE DIS NONCONVULSIVE GENERALIZED|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|GENERALIZED NONCONVULSIVE SEIZURE DIS|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|NONCONVULSIVE GENERALIZED SEIZURE DIS|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|SEIZURE DIS GENERALIZED NONCONVULSIVE|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|GENERALIZED NONCONVULSIVE SEIZURE |GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|GENERALIZED NONCONVULSIVE SEIZURE|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|GENERALISED NON-CONVULSIVE EPILEPSY|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|EPILEPSY, GENERALIZED NONCONVULSIVE|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|NONCONVULSIVE EPILEPSY, GENERALIZED|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|GENERALIZED NONCONVULSIVE EPILEPSY |GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|GENERALISED NON-CONVULSIVE EPILEPSY NOS|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|GENERALIZED NON-CONVULSIVE EPILEPSY NOS|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|GENERALIZED NON-CONVULSIVE EPILEPSY NOS |GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|GENERALISED NONCONVULSIVE EPILEPSY|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|GENERALIZED NON-CONVULSIVE EPILEPSY|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|SEIZURE DISORDER, NONCONVULSIVE GENERALIZED|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|SEIZURE DISORDER, GENERALIZED NONCONVULSIVE|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|GENERALIZED SEIZURE DISORDER, NONCONVULSIVE|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|NONCONVULSIVE GENERALIZED SEIZURE DISORDER|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|NONCONVULSIVE SEIZURE DISORDER, GENERALIZED|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|GENERALIZED NON-CONVULSIVE EPILEPSY |GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|EPILEPSY; GENERALIZED, NONCONVULSIVE|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|GENERALIZED; EPILEPTIC, NONCONVULSIVE|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|GENERALIZED NONCONVULSIVE EPILEPSY, NOS|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0017332|T047|35796005|SNOMEDCT_US|GENERALIZED NONCONVULSIVE SEIZURE DISORDER|GENERALIZED NONCONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|CONVULSIVE GENERALIZED SEIZURE DIS|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|CONVULSIVE SEIZURE DIS GENERALIZED|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|SEIZURE DIS GENERALIZED ONSET|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|SEIZURE DIS CONVULSIVE GENERALIZED|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|SEIZURE DIS GENERALIZED CONVULSIVE|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|GENERALIZED SEIZURE DIS CONVULSIVE|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|GENERALIZED ONSET SEIZURE DIS|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|CONVULSIVE EPILEPSIES, GENERALIZED|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|CONVULSIVE EPILEPSY, GENERALIZED|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|EPILEPSIES, GENERALIZED CONVULSIVE|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|EPILEPSY, GENERALIZED CONVULSIVE|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|GENERALIZED CONVULSIVE EPILEPSIES|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|GENERALIZED CONVULSIVE EPILEPSY |GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|GENERALIZED CONVULSIVE EPILEPSY NOS|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|GENERALISED CONVULSIVE EPILEPSY|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|GENERALISED CONVULSIVE EPILEPSY NOS|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|GENERALIZED CONVULSIVE EPILEPSY|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|GENERALIZED CONVULSIVE EPILEPSY NOS |GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|GENERALIZED CONVULSIVE SEIZURE |GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|GENERALIZED CONVULSIVE SEIZURE|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|EPILEPSY GENERALIZED CONVULSIVE|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|CONVULSIVE SEIZURE DISORDER, GENERALIZED|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|SEIZURE DISORDER, GENERALIZED ONSET|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|SEIZURE DISORDER, GENERALIZED, CONVULSIVE|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|SEIZURE DISORDER, CONVULSIVE, GENERALIZED|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|GENERALIZED SEIZURE DISORDER, CONVULSIVE|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|GENERALIZED ONSET SEIZURE DISORDER|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|GENERALISED-ONSET SEIZURES|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|GENERALIZED-ONSET SEIZURES |GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|GENERALIZED-ONSET SEIZURES|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|EPILEPSY; GENERALIZED, CONVULSIVE|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|GENERALIZED; EPILEPTIC, CONVULSIVE|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|GENERALIZED CONVULSIVE EPILEPSY, NOS|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|GENERALIZED-ONSET SEIZURES, NOS|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|GENERALIZED CONVULSIVE EPILEPSY [DUP] |GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0311334|T047|65120008|SNOMEDCT_US|CONVULSIVE GENERALIZED SEIZURE DISORDER|GENERALIZED CONVULSIVE EPILEPSY (DISORDER)
C0149958|T047|393577005|SNOMEDCT_US|COMPLEX PARTIAL SEIZURES|PARTIAL COMPLEX SEIZURE (DISORDER)
C0149958|T047|393577005|SNOMEDCT_US|SEIZURE PARTIAL (FOCAL) COMPLEX|PARTIAL COMPLEX SEIZURE (DISORDER)
C0149958|T047|393577005|SNOMEDCT_US|COMPLEX PARTIAL SEIZURE|PARTIAL COMPLEX SEIZURE (DISORDER)
C0149958|T047|393577005|SNOMEDCT_US|COMPLEX PARTIAL SEIZURE (PHYSICAL FINDING)|PARTIAL COMPLEX SEIZURE (DISORDER)
C0149958|T047|393577005|SNOMEDCT_US|PARTIAL COMPLEX SEIZURE |PARTIAL COMPLEX SEIZURE (DISORDER)
C0149958|T047|393577005|SNOMEDCT_US|PARTIAL COMPLEX SEIZURE|PARTIAL COMPLEX SEIZURE (DISORDER)
C0149958|T047|393577005|SNOMEDCT_US|PARTIAL COMPLEX SEIZURES|PARTIAL COMPLEX SEIZURE (DISORDER)
C0149958|T047|393577005|SNOMEDCT_US|SEIZURES, COMPLEX PARTIAL|PARTIAL COMPLEX SEIZURE (DISORDER)
C0149958|T047|393577005|SNOMEDCT_US|PARTIAL COMPLEX SEIZURE |PARTIAL COMPLEX SEIZURE (DISORDER)
C0149958|T047|393577005|SNOMEDCT_US|PARTIAL SEIZURES, COMPLEX|PARTIAL COMPLEX SEIZURE (DISORDER)
C0149958|T047|393577005|SNOMEDCT_US|PSYCHOMOTOR FIT|PARTIAL COMPLEX SEIZURE (DISORDER)
C0234972|T047||SNOMEDCT_US|CONVULSIVE DISORDER
C0234972|T047||SNOMEDCT_US|CONVULSIVE DISORDER 
C0234972|T047||SNOMEDCT_US|CONVULSION DISORDER
C0234972|T047||SNOMEDCT_US|DISORDER CONVULSIVE
C0234972|T047||SNOMEDCT_US|CONVULSIVE DISORDER NOS
C0238111|T047|230418006|SNOMEDCT_US|LENNOX-GASTAUT SYNDROME|LENNOX-GASTAUT SYNDROME (DISORDER)
C0238111|T047|230418006|SNOMEDCT_US|LENNOX-GASTAT SYNDROME|LENNOX-GASTAUT SYNDROME (DISORDER)
C0238111|T047|230418006|SNOMEDCT_US|LENNOX GASTAUT SYNDROME|LENNOX-GASTAUT SYNDROME (DISORDER)
C0238111|T047|230418006|SNOMEDCT_US|GASTAUT SYNDROME|LENNOX-GASTAUT SYNDROME (DISORDER)
C0238111|T047|230418006|SNOMEDCT_US|LENNOX-GASTANT SYNDROME|LENNOX-GASTAUT SYNDROME (DISORDER)
C0238111|T047|230418006|SNOMEDCT_US|LENNOX-GASTANT SYNDROME |LENNOX-GASTAUT SYNDROME (DISORDER)
C0238111|T047|230418006|SNOMEDCT_US|LENNOX-GASTAUT SYNDROME |LENNOX-GASTAUT SYNDROME (DISORDER)
C0238111|T047|230418006|SNOMEDCT_US|SYNDROME, LENNOX GASTAUT|LENNOX-GASTAUT SYNDROME (DISORDER)
C0238111|T047|230418006|SNOMEDCT_US|GASTAUT SYNDROME, LENNOX|LENNOX-GASTAUT SYNDROME (DISORDER)
C0238111|T047|230418006|SNOMEDCT_US|LENNOX GASTAUT SYNDROMES|LENNOX-GASTAUT SYNDROME (DISORDER)
C0238111|T047|230418006|SNOMEDCT_US|GASTAUT SYNDROMES, LENNOX|LENNOX-GASTAUT SYNDROME (DISORDER)
C0238111|T047|230418006|SNOMEDCT_US|SYNDROMES, LENNOX GASTAUT|LENNOX-GASTAUT SYNDROME (DISORDER)
C0238111|T047|230418006|SNOMEDCT_US|LENNOX GASTAUT SYNDROME [DISEASE/FINDING]|LENNOX-GASTAUT SYNDROME (DISORDER)
C0238111|T047|230418006|SNOMEDCT_US|LGS|LENNOX-GASTAUT SYNDROME (DISORDER)
C0238111|T047|230418006|SNOMEDCT_US|LENNOX-GASTAUT|LENNOX-GASTAUT SYNDROME (DISORDER)
C0238111|T047|230418006|SNOMEDCT_US|LENNOX-GASTAUT SYNDROME  [AMBIGUOUS]|LENNOX-GASTAUT SYNDROME (DISORDER)
C2236802|T047||SNOMEDCT_US|NONEPILEPTIC SEIZURES 
C2236802|T047||SNOMEDCT_US|NONEPILEPTIC SEIZURES
C2080645|T047||SNOMEDCT_US|PHOTOSENSITIVE SEIZURES 
C2080645|T047||SNOMEDCT_US|PHOTOSENSITIVE SEIZURES
C2349436|T047||SNOMEDCT_US|MIGRAINE TRIGGERED SEIZURES
C2349436|T047||SNOMEDCT_US|MIGRAINE TRIGGERED SEIZURES 
C2349436|T047||SNOMEDCT_US|MIGRAINE-TRIGGERED SEIZURE
C0234974|T047|79348005|SNOMEDCT_US|EPILEPSY, PARTIAL NOS, WITHOUT IMPAIRMENT OF CONSCIOUSNESS|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|EPILEPSY, PARTIAL, WITHOUT IMPAIRMENT OF CONSCIOUSNESS|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|SIMPLE PARTIAL SEIZURES|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|SIMPLE PARTIAL SEIZURES WITH CONSCIOUSNESS PRESERVED|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|SEIZURE PARTIAL (FOCAL) SIMPLE|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|SIMPLE PARTIAL SEIZURE|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|SIMPLE PARTIAL SEIZURE (PHYSICAL FINDING)|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|PARTIAL SIMPLE SEIZURE |SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|PARTIAL SIMPLE SEIZURE WITHOUT IMPAIRMENT OF CONSCIOUSNESS |SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|PARTIAL SIMPLE SEIZURE|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|PARTIAL SIMPLE SEIZURE WITHOUT IMPAIRMENT OF CONSCIOUSNESS|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|PARTIAL SEIZURES, SIMPLE|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|SEIZURES, SIMPLE PARTIAL|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|SEIZURE;FOCAL;SIMPLE PARTIAL|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|PARTIAL EPILEPSY WITHOUT MENTION OF IMPAIRMENT OF CONSCIOUSNESS|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|PARTIAL EPILEPSY WITHOUT MENTION OF IMPAIRMENT OF CONSCIOUSNESS |SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|SIMPLE PARTIAL SEIZURE |SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|PARTIAL EPILEPSY WITHOUT MENTION OF IMPAIRMENT OF CONSCIOUSNESS NOS |SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|PARTIAL EPILEPSY WITHOUT MENTION OF IMPAIRMENT OF CONSCIOUSNESS NOS|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|FOCAL SEIZURES WITHOUT IMPAIRMENT OF CONSCIOUSNESS OR AWARENESS|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|PARTIAL SEIZURES, SIMPLE, CONSCIOUSNESS PRESERVED|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED |SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|SEIZURE; EPILEPTIC, SIMPLE, PARTIAL|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|SIMPLE PARTIAL SEIZURES; EPILEPTIC|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED |SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|SIMPLE PARTIAL FOCAL SEIZURE|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0234974|T047|79348005|SNOMEDCT_US|PARTIAL EPILEPSY, WITHOUT MENTION OF IMPAIRMENT OF CONSCIOUSNESS|SIMPLE PARTIAL SEIZURE, CONSCIOUSNESS NOT IMPAIRED (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|STATUS, PETIT MAL|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|PETIT MAL STATUS|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|PETIT MAL STATUS EPILEPTICUS|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|PETIT MAL EPILEPSY STATUS|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|PETIT MAL EPILEPSY STATUS |PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|STATUS, ABSENCE|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|STATUS EPILEPTICUS;PETIT MAL|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|PETIT MAL STATUS, EPILEPTIC|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|STATUS EPILEPTICUS PETIT MAL|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|ABSENCE STATUS|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|EPILEPTIC ABSENCE STATUS|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|EPILEPSIA MINORIS CONTINUA|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|PETIT-MAL STATUS|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|PROLONGED EPILEPTIC TWILIGHT STATE|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|STATUS PYKNOLEPTICUS|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|NON-CONVULSIVE STATUS EPILEPTICUS WITH IMPAIRED CONSCIOUSNESS|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|SPIKE WAVE STUPOR|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|PETIT MAL STATUS |PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|CONFUSIONAL; STATE, EPILEPTIC|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|EPILEPSY; STATUS, ABSENCE|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|EPILEPSY; STATUS, PETIT MAL|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|EPILEPTICUS; STATUS, PETIT MAL|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|ABSENCE; STATUS|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|PETIT MAL; STATUS|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|STATE; CONFUSIONAL, EPILEPTIC|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|STATUS; ABSENCES|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|STATUS; ABSENCE|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|STATUS; EPILEPTIC, ABSENCE|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|STATUS; EPILEPTIC, PETIT MAL|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|STATUS; EPILEPTICUS, PETIT MAL|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|STATUS; PETIT MAL|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|TWILIGHT STATE; EPILEPTIC|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|EPILEPTIC CONFUSIONAL STATE|PETIT MAL STATUS (DISORDER)
C0270823|T047|7033004|SNOMEDCT_US|EPILEPTIC TWILIGHT STATE|PETIT MAL STATUS (DISORDER)
C0311335|T047|13973009|SNOMEDCT_US|GRAND MAL STATUS EPILEPTICUS|GRAND MAL STATUS (DISORDER)
C0311335|T047|13973009|SNOMEDCT_US|GRAND MAL EPILEPSY STATUS|GRAND MAL STATUS (DISORDER)
C0311335|T047|13973009|SNOMEDCT_US|GRAND MAL EPILEPSY STATUS |GRAND MAL STATUS (DISORDER)
C0311335|T047|13973009|SNOMEDCT_US|GRAND MAL STATUS|GRAND MAL STATUS (DISORDER)
C0311335|T047|13973009|SNOMEDCT_US|STATUS EPILEPTICUS;GRAND MAL|GRAND MAL STATUS (DISORDER)
C0311335|T047|13973009|SNOMEDCT_US|GRAND MAL STATUS, EPILEPTIC|GRAND MAL STATUS (DISORDER)
C0311335|T047|13973009|SNOMEDCT_US|CONVULSIVE STATUS EPILEPTICUS|GRAND MAL STATUS (DISORDER)
C0311335|T047|13973009|SNOMEDCT_US|STATUS EPILEPTICUS GRAND MAL|GRAND MAL STATUS (DISORDER)
C0311335|T047|13973009|SNOMEDCT_US|STATUS EPILEPTICUS, GRAND MAL|GRAND MAL STATUS (DISORDER)
C0311335|T047|13973009|SNOMEDCT_US|GENERALIZED CONVULSIVE STATUS EPILEPTICUS|GRAND MAL STATUS (DISORDER)
C0311335|T047|13973009|SNOMEDCT_US|STATUS EPILEPTICUS, GENERALIZED CONVULSIVE|GRAND MAL STATUS (DISORDER)
C0311335|T047|13973009|SNOMEDCT_US|GRAND MAL STATUS |GRAND MAL STATUS (DISORDER)
C0311335|T047|13973009|SNOMEDCT_US|EPILEPSY; STATUS, GRAND MAL|GRAND MAL STATUS (DISORDER)
C0311335|T047|13973009|SNOMEDCT_US|EPILEPTICUS; STATUS, GRAND MAL|GRAND MAL STATUS (DISORDER)
C0311335|T047|13973009|SNOMEDCT_US|GRAND MAL; STATUS|GRAND MAL STATUS (DISORDER)
C0311335|T047|13973009|SNOMEDCT_US|STATUS; EPILEPTIC, GRAND MAL|GRAND MAL STATUS (DISORDER)
C0311335|T047|13973009|SNOMEDCT_US|STATUS; EPILEPTICUS, GRAND MAL|GRAND MAL STATUS (DISORDER)
C0311335|T047|13973009|SNOMEDCT_US|STATUS; GRAND MAL|GRAND MAL STATUS (DISORDER)
C0751777|T047||SNOMEDCT_US|PROGRESSIVE FAMILIAL MYOCLONIC EPILEPSY
C0751777|T047||SNOMEDCT_US|PROGRESSIVE FAMILIAL MYOCLONIC EPILEPSY 
C0751777|T047||SNOMEDCT_US|FAMILIAL PROGRESSIVE MYOCLONIC EPILEPSY
C0751777|T047||SNOMEDCT_US|MYOCLONIC; EPILEPTIC, PROGRESSIVE (FAMILIAL)
C0751783|T047|230425004|SNOMEDCT_US|DISEASE, LAFORA|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|LAFORA DISEASE|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|LAFORA'S DISEASE|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|MYOCLONIC EPILEPSY OF LAFORA|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|EPM2A|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|LAFORA DIS|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|LAFORA BODY DIS|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|LAFORA BODY DISEASE |LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|LAFORA BODY DISEASE|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|DISEASE, LAFORA BODY|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|LAFORA TYPE PROGRESSIVE MYOCLONIC EPILEPSY|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|EPILEPSY, PROGRESSIVE MYOCLONIC, LAFORA|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|PROGRESSIVE MYOCLONIC EPILEPSY, LAFORA TYPE|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|LAFORA DISEASE [DISEASE/FINDING]|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|PROGRESSIVE MYOCLONIC EPILEPSY, LAFORA|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|LAFORA PROGRESSIVE MYOCLONIC EPILEPSY|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|DISORDER, LAFORA BODY|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|LAFORA MYOCLONIC EPILEPSY|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|LAFORA BODY DISORDER|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|EPILEPSY PROGRESSIVE MYOCLONIC 2|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|LAFORA'S MYOCLONIC EPILEPSY|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|LAFORA PROGRESSIVE MYOCLONUS EPILEPSY|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|PROGRESSIVE MYOCLONUS EPILEPSY, LAFORA TYPE|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|PROGRESSIVE MYOCLONIC EPILEPSY TYPE 2|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|EPILEPSY, PROGRESSIVE MYOCLONIC 2A|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|EPILEPSY, PROGRESSIVE MYOCLONIC, 2A|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|MELF|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|EPM2|LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|LAFORA DISEASE |LAFORA DISEASE (DISORDER)
C0751783|T047|230425004|SNOMEDCT_US|LAFORA|LAFORA DISEASE (DISORDER)
C0037769|T047|288197007|SNOMEDCT_US|INFANTILE SPASMS|WEST SYNDROME (FINDING)
C0037769|T047|288197007|SNOMEDCT_US|INFANTILE SPASM|WEST SYNDROME (FINDING)
C0037769|T047|288197007|SNOMEDCT_US|SPASMS, INFANTILE|WEST SYNDROME (FINDING)
C0037769|T047|288197007|SNOMEDCT_US|SYNDROME, WEST|WEST SYNDROME (FINDING)
C0037769|T047|288197007|SNOMEDCT_US|INFANTILE SPASMS |WEST SYNDROME (FINDING)
C0037769|T047|288197007|SNOMEDCT_US|WEST SYNDROME|WEST SYNDROME (FINDING)
C0037769|T047|288197007|SNOMEDCT_US|SPASMS, INFANTILE [DISEASE/FINDING]|WEST SYNDROME (FINDING)
C0037769|T047|288197007|SNOMEDCT_US|SEIZURE;INFANT SPASMS|WEST SYNDROME (FINDING)
C0037769|T047|288197007|SNOMEDCT_US|WEST'S SYNDROME|WEST SYNDROME (FINDING)
C0037769|T047|288197007|SNOMEDCT_US|WEST SYNDROME |WEST SYNDROME (FINDING)
C0037769|T047|288197007|SNOMEDCT_US|INFANTILE SPASMS NOS|WEST SYNDROME (FINDING)
C0037769|T047|288197007|SNOMEDCT_US|WEST SYNDROME |WEST SYNDROME (FINDING)
C0037769|T047|288197007|SNOMEDCT_US|INFANTILE SPASMS NOS |WEST SYNDROME (FINDING)
C0037769|T047|288197007|SNOMEDCT_US|INFANTILE SPASMS - HYPSARRYTHMIA|WEST SYNDROME (FINDING)
C0037769|T047|288197007|SNOMEDCT_US|INFANTILE SPASMS - HYPSARRHYTHMIA|WEST SYNDROME (FINDING)
C0037769|T047|288197007|SNOMEDCT_US|LIGHTNING SPASMS|WEST SYNDROME (FINDING)
C0037769|T047|288197007|SNOMEDCT_US|INFANTILE; SPASM|WEST SYNDROME (FINDING)
C0037769|T047|288197007|SNOMEDCT_US|LIGHTNING; SPASM|WEST SYNDROME (FINDING)
C0037769|T047|288197007|SNOMEDCT_US|SPASM; INFANTILE|WEST SYNDROME (FINDING)
C0037769|T047|288197007|SNOMEDCT_US|SPASM; LIGHTNING|WEST SYNDROME (FINDING)
C0270819|T047|71427006|SNOMEDCT_US|CURSIVE EPILEPSY|CURSIVE SEIZURE (DISORDER)
C0270819|T047|71427006|SNOMEDCT_US|CURSIVE SEIZURE |CURSIVE SEIZURE (DISORDER)
C0270819|T047|71427006|SNOMEDCT_US|CURSIVE SEIZURE|CURSIVE SEIZURE (DISORDER)
C0270819|T047|71427006|SNOMEDCT_US|EPILEPSIES, CURSIVE|CURSIVE SEIZURE (DISORDER)
C0270819|T047|71427006|SNOMEDCT_US|EPILEPSY, CURSIVE|CURSIVE SEIZURE (DISORDER)
C0270819|T047|71427006|SNOMEDCT_US|REFLEX EPILEPSIES, CURSIVE (RUNNING)|CURSIVE SEIZURE (DISORDER)
C0270819|T047|71427006|SNOMEDCT_US|CURSIVE REFLEX EPILEPSIES (RUNNING)|CURSIVE SEIZURE (DISORDER)
C0270819|T047|71427006|SNOMEDCT_US|CURSIVE REFLEX EPILEPSY (RUNNING)|CURSIVE SEIZURE (DISORDER)
C0270819|T047|71427006|SNOMEDCT_US|EPILEPSY, CURSIVE REFLEX (RUNNING)|CURSIVE SEIZURE (DISORDER)
C0270819|T047|71427006|SNOMEDCT_US|RUNNING EPILEPSY|CURSIVE SEIZURE (DISORDER)
C0270819|T047|71427006|SNOMEDCT_US|CURSIVE (RUNNING) EPILEPSY|CURSIVE SEIZURE (DISORDER)
C0270819|T047|71427006|SNOMEDCT_US|CURSIVE (RUNNING) EPILEPSY |CURSIVE SEIZURE (DISORDER)
C0270819|T047|71427006|SNOMEDCT_US|CURSIVE SEIZURE |CURSIVE SEIZURE (DISORDER)
C0270819|T047|71427006|SNOMEDCT_US|REFLEX EPILEPSY, CURSIVE (RUNNING)|CURSIVE SEIZURE (DISORDER)
C0270819|T047|71427006|SNOMEDCT_US|EPILEPSY, RUNNING|CURSIVE SEIZURE (DISORDER)
C0270820|T047|89525009|SNOMEDCT_US|GELASTIC EPILEPSY|GELASTIC SEIZURE (DISORDER)
C0270820|T047|89525009|SNOMEDCT_US|GELASTIC SEIZURE|GELASTIC SEIZURE (DISORDER)
C0270820|T047|89525009|SNOMEDCT_US|GELASTIC SEIZURE |GELASTIC SEIZURE (DISORDER)
C0270820|T047|89525009|SNOMEDCT_US|EPILEPSIES, GELASTIC|GELASTIC SEIZURE (DISORDER)
C0270820|T047|89525009|SNOMEDCT_US|GELASTIC EPILEPSIES|GELASTIC SEIZURE (DISORDER)
C0270820|T047|89525009|SNOMEDCT_US|GELASTIC SEIZURES|GELASTIC SEIZURE (DISORDER)
C0270820|T047|89525009|SNOMEDCT_US|GELASTIC SEIZURE |GELASTIC SEIZURE (DISORDER)
C0270820|T047|89525009|SNOMEDCT_US|EPILEPSY, GELASTIC|GELASTIC SEIZURE (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|EPILEPSIA PARTIALIS CONTINUA|KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|SYNDROME, KOJEWNIKOW'S|KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|SYNDROME, KOZHEVNIKOV'S|KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|EPILEPSY, KOJEVNIKOV'S|KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|EPILEPSIA PARTIALIS CONTINUA |KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|KOJEVNIKOV EPILEPSY|KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|EPILEPSY, KOJEWNIKOV'S|KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|KOJEWNIKOV EPILEPSY|KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|SYNDROME, KOJEWNIKOW|KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|SYNDROME, KOZHEVNIKOV|KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|KOJEVNIKOV'S EPILEPSY|KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|KOJEWNIKOW SYNDROME|KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|KOJEWNIKOW'S SYNDROME|KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|KOZHEVNIKOV'S SYNDROME|KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|KOJEWNIKOV'S EPILEPSY|KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|EPILEPSIA PARTIALIS CONTINUA [DISEASE/FINDING]|KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|KOZHEVNIKOV SYNDROME|KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|KOJEVNIKOV'S EPILEPSIES|KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|EPILEPSIES, KOJEVNIKOV'S|KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|KOJEVNIKOV'S EPILEPSY |KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|FOCAL STATUS EPILEPTICUS|KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|MOTOR SIMPLE PARTIAL STATUS|KOJEVNIKOV'S EPILEPSY (DISORDER)
C0085543|T047|193017009|SNOMEDCT_US|EPILEPSIA PARTIALIS CONTINUA |KOJEVNIKOV'S EPILEPSY (DISORDER)
C0796133|T047||SNOMEDCT_US|RAMON SYNDROME
C0796133|T047||SNOMEDCT_US|GINGIVAL FIBROMATOSIS COMBINED WITH CHERUBISM
C0796133|T047||SNOMEDCT_US|CHERUBISM, GINGIVAL FIBROMATOSIS, EPILEPSY, MENTAL DEFICIENCY, HYPERTRICHOSIS, AND STUNTED GROWTH
C1856929|T047||SNOMEDCT_US|EPILEPSY-TELANGIECTASIA
C1856929|T047||SNOMEDCT_US|EPILEPSY TELANGIECTASIA
C0270709|T047|2355008|SNOMEDCT_US|RUD SYNDROME|RUD'S SYNDROME (DISORDER)
C0270709|T047|2355008|SNOMEDCT_US|RUDS|RUD'S SYNDROME (DISORDER)
C0270709|T047|2355008|SNOMEDCT_US|ICHTHYOSIS HYPOGONADISM MENTAL RETARDATION EPILEPSY SYNDROME|RUD'S SYNDROME (DISORDER)
C0270709|T047|2355008|SNOMEDCT_US|ICHTHYOSIS MENTAL RETARDATION-EPILEPSY HYPOGONADISM SYNDROME|RUD'S SYNDROME (DISORDER)
C0270709|T047|2355008|SNOMEDCT_US|RUD'S SYNDROME|RUD'S SYNDROME (DISORDER)
C0270709|T047|2355008|SNOMEDCT_US|NEUROICHTHYOSIS HYPOGONADISM SYNDROME|RUD'S SYNDROME (DISORDER)
C0270709|T047|2355008|SNOMEDCT_US|DWARFISM ICHTHYOSIFORM ERYTHRODERMA MENTAL DEFICIENCY SYNDROME|RUD'S SYNDROME (DISORDER)
C0270709|T047|2355008|SNOMEDCT_US|ICHTHYOSIS OLIGOPHRENIA EPILEPSY SYNDROME|RUD'S SYNDROME (DISORDER)
C0270709|T047|2355008|SNOMEDCT_US|ICHTHYOSIS MALE HYPOGONADISM SYNDROME|RUD'S SYNDROME (DISORDER)
C0270709|T047|2355008|SNOMEDCT_US|DWARFISM-ICHTHYOSIFORM ERYTHRODERMA-MENTAL DEFICIENCY SYNDROME|RUD'S SYNDROME (DISORDER)
C0270709|T047|2355008|SNOMEDCT_US|RUD'S SYNDROME |RUD'S SYNDROME (DISORDER)
C1849508|T047|734434007|SNOMEDCT_US|EPILEPSY, PYRIDOXINE-DEPENDENT|PYRIDOXINE-DEPENDENT EPILEPSY (DISORDER)
C1849508|T047|734434007|SNOMEDCT_US|PYRIDOXINE DEPENDENCY WITH SEIZURES|PYRIDOXINE-DEPENDENT EPILEPSY (DISORDER)
C1849508|T047|734434007|SNOMEDCT_US|PYRIDOXINE-DEPENDENT EPILEPSY|PYRIDOXINE-DEPENDENT EPILEPSY (DISORDER)
C1849508|T047|734434007|SNOMEDCT_US|PYRIDOXINE DEPENDENCY|PYRIDOXINE-DEPENDENT EPILEPSY (DISORDER)
C1849508|T047|734434007|SNOMEDCT_US|AASA DEHYDROGENASE DEFICIENCY|PYRIDOXINE-DEPENDENT EPILEPSY (DISORDER)
C1849508|T047|734434007|SNOMEDCT_US|PYRIDOXINE-DEPENDENT SEIZURES|PYRIDOXINE-DEPENDENT EPILEPSY (DISORDER)
C1849508|T047|734434007|SNOMEDCT_US|VITAMIN B6-DEPENDENT SEIZURES|PYRIDOXINE-DEPENDENT EPILEPSY (DISORDER)
C0795900|T047||SNOMEDCT_US|DWARFISM, LEAN SPASTIC TYPE
C0795900|T047||SNOMEDCT_US|COFFIN SYNDROME 1
C0795900|T047||SNOMEDCT_US|LEAN SPASTIC DWARFISM
C0265339|T047|21634003|SNOMEDCT_US|BFLS|BORJESON-FORSSMAN-LEHMANN SYNDROME (DISORDER)
C0265339|T047|21634003|SNOMEDCT_US|BORJESON-FORSSMAN-LEHMANN SYNDROME|BORJESON-FORSSMAN-LEHMANN SYNDROME (DISORDER)
C0265339|T047|21634003|SNOMEDCT_US|BORJESON SYNDROME|BORJESON-FORSSMAN-LEHMANN SYNDROME (DISORDER)
C0265339|T047|21634003|SNOMEDCT_US|MENTAL DEFICIENCY, EPILEPSY AND ENDOCRINE DISORDERS|BORJESON-FORSSMAN-LEHMANN SYNDROME (DISORDER)
C0265339|T047|21634003|SNOMEDCT_US|MRXSBFL|BORJESON-FORSSMAN-LEHMANN SYNDROME (DISORDER)
C0265339|T047|21634003|SNOMEDCT_US|MENTAL DEFICIENCY, EPILEPSY, AND ENDOCRINE DISORDERS|BORJESON-FORSSMAN-LEHMANN SYNDROME (DISORDER)
C0265339|T047|21634003|SNOMEDCT_US|BORJESON-FORSSMAN-LEHMANN SYNDROME |BORJESON-FORSSMAN-LEHMANN SYNDROME (DISORDER)
C0265339|T047|21634003|SNOMEDCT_US|MENTAL RETARDATION, EPILEPSY, AND ENDOCRINE DISORDERS|BORJESON-FORSSMAN-LEHMANN SYNDROME (DISORDER)
C0265339|T047|21634003|SNOMEDCT_US|MENTAL RETARDATION, X-LINKED, SYNDROMIC, BORJESON-FORSSMAN-LEHMANN TYPE|BORJESON-FORSSMAN-LEHMANN SYNDROME (DISORDER)
C0265339|T047|21634003|SNOMEDCT_US|BORJESON-FORSSMAN-LEHMANN SYNDROME |BORJESON-FORSSMAN-LEHMANN SYNDROME (DISORDER)
C0796202|T047||SNOMEDCT_US|WITTWER SYNDROME
C0265328|T047|45167004|SNOMEDCT_US|ALOPECIA-EPILEPSY-OLIGOPHRENIA SYNDROME OF MOYNAHAN|MOYNAHAN'S SYNDROME (DISORDER)
C0265328|T047|45167004|SNOMEDCT_US|MOYNAHAN'S SYNDROME |MOYNAHAN'S SYNDROME (DISORDER)
C0265328|T047|45167004|SNOMEDCT_US|MOYNAHAN'S SYNDROME|MOYNAHAN'S SYNDROME (DISORDER)
C0265328|T047|45167004|SNOMEDCT_US|MOYNAHAN SYNDROME|MOYNAHAN'S SYNDROME (DISORDER)
C0265328|T047|45167004|SNOMEDCT_US|ALOPECIA EPILEPSY OLIGOPHRENIA SYNDROME OF MOYNAHAN|MOYNAHAN'S SYNDROME (DISORDER)
C0265328|T047|45167004|SNOMEDCT_US|MOYNAHAN ALOPECIA SYNDROME|MOYNAHAN'S SYNDROME (DISORDER)
C0265328|T047|45167004|SNOMEDCT_US|PROGRESSIVE CARDIOMYOPATHIC LENTIGINOSIS|MOYNAHAN'S SYNDROME (DISORDER)
C0265328|T047|45167004|SNOMEDCT_US|MOYNAHAN'S SYNDROME |MOYNAHAN'S SYNDROME (DISORDER)
C1863090|T047|720980004|SNOMEDCT_US|ALOPECIA, PSYCHOMOTOR EPILEPSY, PYORRHEA, AND MENTAL SUBNORMALITY|SHOKEIR SYNDROME
C1863090|T047|720980004|SNOMEDCT_US|CONGENITAL UNIVERSAL ALOPECIA, EPILEPSY, MENTAL SUBNORMALITY AND PYORRHEA|SHOKEIR SYNDROME
C1863090|T047|720980004|SNOMEDCT_US|ALOPECIA, EPILEPSY, PYORRHEA, MENTAL SUBNORMALITY|SHOKEIR SYNDROME
C1863090|T047|720980004|SNOMEDCT_US|SHOKEIR SYNDROME|SHOKEIR SYNDROME
C0406740|T047|109478007|SNOMEDCT_US|KOHLSCHUTTER-TONZ SYNDROME|KOHLSCHUTTER'S SYNDROME (DISORDER)
C0406740|T047|109478007|SNOMEDCT_US|EPILEPSY DEMENTIA AMELOGENESIS IMPERFECTA|KOHLSCHUTTER'S SYNDROME (DISORDER)
C0406740|T047|109478007|SNOMEDCT_US|EPILEPSY AND YELLOW TEETH|KOHLSCHUTTER'S SYNDROME (DISORDER)
C0406740|T047|109478007|SNOMEDCT_US|KOHLSCHUTTER SYNDROME|KOHLSCHUTTER'S SYNDROME (DISORDER)
C0406740|T047|109478007|SNOMEDCT_US|KOHLSCHUTTER TONZ SYNDROME|KOHLSCHUTTER'S SYNDROME (DISORDER)
C0406740|T047|109478007|SNOMEDCT_US|EPILEPSY, DEMENTIA, AND AMELOGENESIS IMPERFECTA|KOHLSCHUTTER'S SYNDROME (DISORDER)
C0406740|T047|109478007|SNOMEDCT_US|KTZS|KOHLSCHUTTER'S SYNDROME (DISORDER)
C0406740|T047|109478007|SNOMEDCT_US|KOHLSCHUTTER'S SYNDROME|KOHLSCHUTTER'S SYNDROME (DISORDER)
C0406740|T047|109478007|SNOMEDCT_US|DISORDERS OF CENTRAL NERVOUS SYSTEM KOHLSCHUTTER'S SYNDROME|KOHLSCHUTTER'S SYNDROME (DISORDER)
C0406740|T047|109478007|SNOMEDCT_US|KOHLSCHUTTER'S SYNDROME |KOHLSCHUTTER'S SYNDROME (DISORDER)
C0406740|T047|109478007|SNOMEDCT_US|AMELOCEREBROHYPOHIDROTIC SYNDROME|KOHLSCHUTTER'S SYNDROME (DISORDER)
C0406740|T047|109478007|SNOMEDCT_US|EPILEPSY, DEMENTIA AND AMELOGENESIS IMPERFECTA|KOHLSCHUTTER'S SYNDROME (DISORDER)
C0406740|T047|109478007|SNOMEDCT_US|EPILEPSY, MENTAL DETERIORATION AND YELLOW TEETH|KOHLSCHUTTER'S SYNDROME (DISORDER)
C0406740|T047|109478007|SNOMEDCT_US|KOHLSCHUTTER'S SYNDROME |KOHLSCHUTTER'S SYNDROME (DISORDER)
C2931451|T047||SNOMEDCT_US|SANDHAUS BEN-AMI SYNDROME
C2931451|T047||SNOMEDCT_US|PATELLA HYPOPLASIA SKELETAL MALFORMATIONS
C2931495|T047||SNOMEDCT_US|ARTHROGRYPOSIS MULTIPLEX CONGENITA WITH EPILEPTIC SEIZURES AND MIGRATIONAL BRAIN DISORDER
C2931495|T047||SNOMEDCT_US|ARTHROGRYPOSIS EPILEPTIC SEIZURES MIGRATIONAL BRAIN DISORDER
C1846278|T047|722037004|SNOMEDCT_US|MENTAL RETARDATION, EPILEPTIC SEIZURES, HYPOGONADISM AND HYPOGENITALISM, MICROCEPHALY, AND OBESITY|MEHMO (MENTAL RETARDATION, EPILEPTIC SEIZURES, HYPOGONADISM AND HYPOGENITALISM, MICROCEPHALY, OBESITY) SYNDROME
C1846278|T047|722037004|SNOMEDCT_US|MEHMO|MEHMO (MENTAL RETARDATION, EPILEPTIC SEIZURES, HYPOGONADISM AND HYPOGENITALISM, MICROCEPHALY, OBESITY) SYNDROME
C1846278|T047|722037004|SNOMEDCT_US|MENTAL RETARDATION, EPILEPTIC SEIZURES, HYPOGONADISM AND HYPOGENITALISM, MICROCEPHALY, AND OBESITY |MEHMO (MENTAL RETARDATION, EPILEPTIC SEIZURES, HYPOGONADISM AND HYPOGENITALISM, MICROCEPHALY, OBESITY) SYNDROME
C1846278|T047|722037004|SNOMEDCT_US|MEHMO SYNDROME|MEHMO (MENTAL RETARDATION, EPILEPTIC SEIZURES, HYPOGONADISM AND HYPOGENITALISM, MICROCEPHALY, OBESITY) SYNDROME
C1846278|T047|722037004|SNOMEDCT_US|X-LINKED MEHMO SYNDROME|MEHMO (MENTAL RETARDATION, EPILEPTIC SEIZURES, HYPOGONADISM AND HYPOGENITALISM, MICROCEPHALY, OBESITY) SYNDROME
C1846278|T047|722037004|SNOMEDCT_US|MRXS20|MEHMO (MENTAL RETARDATION, EPILEPTIC SEIZURES, HYPOGONADISM AND HYPOGENITALISM, MICROCEPHALY, OBESITY) SYNDROME
C1846278|T047|722037004|SNOMEDCT_US|MRXS25|MEHMO (MENTAL RETARDATION, EPILEPTIC SEIZURES, HYPOGONADISM AND HYPOGENITALISM, MICROCEPHALY, OBESITY) SYNDROME
C1846278|T047|722037004|SNOMEDCT_US|MENTAL RETARDATION, X-LINKED, SYNDROMIC 25|MEHMO (MENTAL RETARDATION, EPILEPTIC SEIZURES, HYPOGONADISM AND HYPOGENITALISM, MICROCEPHALY, OBESITY) SYNDROME
C1846278|T047|722037004|SNOMEDCT_US|MENTAL RETARDATION, X-LINKED, SYNDROMIC 20|MEHMO (MENTAL RETARDATION, EPILEPTIC SEIZURES, HYPOGONADISM AND HYPOGENITALISM, MICROCEPHALY, OBESITY) SYNDROME
C0796046|T047|715428003|SNOMEDCT_US|GURRIERI SYNDROME|SKELETAL DYSPLASIA WITH EPILEPSY AND SHORT STATURE SYNDROME (DISORDER)
C0796046|T047|715428003|SNOMEDCT_US|SKELETAL DYSPLASIA EPILEPSY SHORT STATURE|SKELETAL DYSPLASIA WITH EPILEPSY AND SHORT STATURE SYNDROME (DISORDER)
C0796046|T047|715428003|SNOMEDCT_US|GURRIERI SAMMITO BELLUSSI SYNDROME|SKELETAL DYSPLASIA WITH EPILEPSY AND SHORT STATURE SYNDROME (DISORDER)
C2931579|T047|733031004|SNOMEDCT_US|BATTAGLIA NERI SYNDROME|EPILEPSY, MICROCEPHALY, SKELETAL DYSPLASIA SYNDROME (DISORDER)
C0796010|T047||SNOMEDCT_US|KIFAFA SEIZURE DISORDER
C0796010|T047||SNOMEDCT_US|COMPLEX FAMILIAL SEIZURE DISORDER
C0796010|T047||SNOMEDCT_US|VITSALA
C2931668|T047||SNOMEDCT_US|BOUDHINA YEDES KHIARI SYNDROME
C1838491|T047||SNOMEDCT_US|PACHYGYRIA, MENTAL RETARDATION AND EPILEPSY
C1838491|T047||SNOMEDCT_US|PACHYGYRIA WITH MENTAL RETARDATION AND SEIZURES
C1838491|T047||SNOMEDCT_US|KUZNIECKY SYNDROME
C1838491|T047||SNOMEDCT_US|PACHYGYRIA WITH MENTAL RETARDATION, SEIZURES, AND ARACHNOID CYSTS
C3472688|T047|981000119108|SNOMEDCT_US|SINGLE EPILEPTIC SEIZURE |SINGLE EPILEPTIC SEIZURE (FINDING)
C3472688|T047|981000119108|SNOMEDCT_US|SINGLE EPILEPTIC SEIZURE|SINGLE EPILEPTIC SEIZURE (FINDING)
C0751111|T047||SNOMEDCT_US|EPILEPSY, AWAKENING
C0751111|T047||SNOMEDCT_US|AWAKENING EPILEPSY
C0751110|T047|703150000|SNOMEDCT_US|SEIZURE, SINGLE|SINGLE SEIZURE (FINDING)
C0751110|T047|703150000|SNOMEDCT_US|SEIZURES, SINGLE|SINGLE SEIZURE (FINDING)
C0751110|T047|703150000|SNOMEDCT_US|SINGLE SEIZURES|SINGLE SEIZURE (FINDING)
C0751110|T047|703150000|SNOMEDCT_US|SINGLE SEIZURE|SINGLE SEIZURE (FINDING)
C0751110|T047|703150000|SNOMEDCT_US|SINGLE SEIZURE |SINGLE SEIZURE (FINDING)
C0086237|T047||SNOMEDCT_US|CRYPTOGENIC EPILEPSIES
C0086237|T047||SNOMEDCT_US|CRYPTOGENIC EPILEPSY
C0086237|T047||SNOMEDCT_US|EPILEPSIES, CRYPTOGENIC
C0086237|T047||SNOMEDCT_US|EPILEPSY, CRYPTOGENIC
C0553754|T047|309847002|SNOMEDCT_US|FIT (IN KNOWN EPILEPTIC) NOS|FIT (IN KNOWN EPILEPTIC) NOS (DISORDER)
C0553754|T047|309847002|SNOMEDCT_US|FIT (IN KNOWN EPILEPTIC) NOS |FIT (IN KNOWN EPILEPTIC) NOS (DISORDER)
C0553754|T047|309847002|SNOMEDCT_US|FIT (IN KNOWN EPILEPTIC)|FIT (IN KNOWN EPILEPTIC) NOS (DISORDER)
C1827389|T047|422513000|SNOMEDCT_US|EPILEPSY, NOT REFRACTORY |EPILEPSY, NOT INTRACTABLE
C1827389|T047|422513000|SNOMEDCT_US|EPILEPSY, NOT REFRACTORY|EPILEPSY, NOT INTRACTABLE
C1827389|T047|422513000|SNOMEDCT_US|EPILEPSY, NOT INTRACTABLE|EPILEPSY, NOT INTRACTABLE
C1827389|T047|422513000|SNOMEDCT_US|EPILEPSY NOT INTRACTABLE|EPILEPSY, NOT INTRACTABLE
C1827389|T047|422513000|SNOMEDCT_US|EPILEPSY, NOT INTRACTABLE |EPILEPSY, NOT INTRACTABLE
C3649195|T047||SNOMEDCT_US|EPILEPSY, NOT INTRACTABLE, WITH STATUS EPILEPTICUS
C3649195|T047||SNOMEDCT_US|EPILEPSY NOT INTRACTABLE WITH STATUS EPILEPTICUS
C3649195|T047||SNOMEDCT_US|EPILEPSY, NOT INTRACTABLE, WITH STATUS EPILEPTICUS 
C3646244|T047||SNOMEDCT_US|SEIZURES RELATED TO EXTERNAL CAUSES 
C3646244|T047||SNOMEDCT_US|SEIZURES RELATED TO EXTERNAL CAUSES
C0472349|T047|230390002|SNOMEDCT_US|LOCALIZATION-RELATED SYMPTOMATIC EPILEPSY|LOCALIZATION-RELATED SYMPTOMATIC EPILEPSY (DISORDER)
C0472349|T047|230390002|SNOMEDCT_US|EPILEPSY LOCALIZATION-RELATED SYMPTOMATIC|LOCALIZATION-RELATED SYMPTOMATIC EPILEPSY (DISORDER)
C0472349|T047|230390002|SNOMEDCT_US|LOCALIZATION-RELATED SYMPTOMATIC EPILEPSY |LOCALIZATION-RELATED SYMPTOMATIC EPILEPSY (DISORDER)
C0472349|T047|230390002|SNOMEDCT_US|LOCALISATION-RELATED SYMPTOMATIC EPILEPSY|LOCALIZATION-RELATED SYMPTOMATIC EPILEPSY (DISORDER)
C0472349|T047|230390002|SNOMEDCT_US|LOCALIZATION-RELATED SYMPTOMATIC EPILEPSY |LOCALIZATION-RELATED SYMPTOMATIC EPILEPSY (DISORDER)
C0472349|T047|230390002|SNOMEDCT_US|EPILEPSY; LOCALIZATION-RELATED, SYMPTOMATIC|LOCALIZATION-RELATED SYMPTOMATIC EPILEPSY (DISORDER)
C0472348|T047|278510009|SNOMEDCT_US|EPILEPSY LOCALIZATION-RELATED IDIOPATHIC |LOCALIZATION-RELATED IDIOPATHIC EPILEPSY (DISORDER)
C0472348|T047|278510009|SNOMEDCT_US|EPILEPSY LOCALIZATION-RELATED IDIOPATHIC|LOCALIZATION-RELATED IDIOPATHIC EPILEPSY (DISORDER)
C0472348|T047|278510009|SNOMEDCT_US|LOCALISATION-RELATED IDIOPATHIC EPILEPSY|LOCALIZATION-RELATED IDIOPATHIC EPILEPSY (DISORDER)
C0472348|T047|278510009|SNOMEDCT_US|LOCALIZATION-RELATED IDIOPATHIC EPILEPSY|LOCALIZATION-RELATED IDIOPATHIC EPILEPSY (DISORDER)
C0472348|T047|278510009|SNOMEDCT_US|LOCALIZATION-RELATED IDIOPATHIC EPILEPSY |LOCALIZATION-RELATED IDIOPATHIC EPILEPSY (DISORDER)
C0472348|T047|278510009|SNOMEDCT_US|EPILEPSY; IDIOPATHIC, LOCALIZATION-RELATED|LOCALIZATION-RELATED IDIOPATHIC EPILEPSY (DISORDER)
C0472348|T047|278510009|SNOMEDCT_US|EPILEPSY; LOCALIZATION-RELATED, IDIOPATHIC|LOCALIZATION-RELATED IDIOPATHIC EPILEPSY (DISORDER)
C3662042|T047|137991000119103|SNOMEDCT_US|SEIZURE DISORDER AS SEQUELA OF STROKE|SEIZURE DISORDER AS SEQUELA OF STROKE (DISORDER)
C3662042|T047|137991000119103|SNOMEDCT_US|SEIZURE DISORDER AS SEQUELA OF STROKE |SEIZURE DISORDER AS SEQUELA OF STROKE (DISORDER)
C0751124|T047|187931000119106|SNOMEDCT_US|ATYPICAL ABSENCE EPILEPSY|ATYPICAL ABSENCE EPILEPSY (DISORDER)
C0751124|T047|187931000119106|SNOMEDCT_US|ATYPICAL ABSENCE EPILEPSY |ATYPICAL ABSENCE EPILEPSY (DISORDER)
C0751124|T047|187931000119106|SNOMEDCT_US|EPILEPSY, ABSENCE, ATYPICAL|ATYPICAL ABSENCE EPILEPSY (DISORDER)
C0086236|T047|192981006|SNOMEDCT_US|ATONIC EPILEPSIES|EPILEPTIC SEIZURES - ATONIC (FINDING)
C0086236|T047|192981006|SNOMEDCT_US|ATONIC EPILEPSY|EPILEPTIC SEIZURES - ATONIC (FINDING)
C0086236|T047|192981006|SNOMEDCT_US|EPILEPSIES, ATONIC|EPILEPTIC SEIZURES - ATONIC (FINDING)
C0086236|T047|192981006|SNOMEDCT_US|ATONIC EPILEPSY |EPILEPTIC SEIZURES - ATONIC (FINDING)
C0086236|T047|192981006|SNOMEDCT_US|EPILEPSY, ATONIC|EPILEPTIC SEIZURES - ATONIC (FINDING)
C0086236|T047|192981006|SNOMEDCT_US|EPILEPTIC SEIZURES - ATONIC|EPILEPTIC SEIZURES - ATONIC (FINDING)
C0086236|T047|192981006|SNOMEDCT_US|EPILEPTIC SEIZURES - ATONIC |EPILEPTIC SEIZURES - ATONIC (FINDING)
C3697594|T047|698767004|SNOMEDCT_US|POST-CEREBROVASCULAR ACCIDENT EPILEPSY |POST-CEREBROVASCULAR ACCIDENT EPILEPSY (DISORDER)
C3697594|T047|698767004|SNOMEDCT_US|POST-CEREBROVASCULAR ACCIDENT EPILEPSY|POST-CEREBROVASCULAR ACCIDENT EPILEPSY (DISORDER)
C1837530|T047||SNOMEDCT_US|AICAR TRANSFORMYLASE/IMP CYCLOHYDROLASE DEFICIENCY
C1837530|T047||SNOMEDCT_US|AICA RIBOSURIA DUE TO ATIC DEFICIENCY
C1837530|T047||SNOMEDCT_US|AICAR TRANSFORMYLASE INOSINE MONOPHOSPHATE CYCLOHYDROLASE DEFICIENCY
C1837530|T047||SNOMEDCT_US|ATIC DEFICIENCY
C1837530|T047||SNOMEDCT_US|AICA-RIBOSURIA DUE TO ATIC DEFICIENCY
C1845343|T047||SNOMEDCT_US|EPILEPSY, X-LINKED, WITH VARIABLE LEARNING DISABILITIES AND BEHAVIOR DISORDERS
C1849416|T047||SNOMEDCT_US|RETINAL DEGENERATION AND EPILEPSY
C1845102|T047||SNOMEDCT_US|EPILEPTIC ENCEPHALOPATHY, EARLY INFANTILE, 8
C1845102|T047||SNOMEDCT_US|EIEE8
C1845102|T047||SNOMEDCT_US|HYPEREKPLEXIA AND EPILEPSY
C2751195|T047||SNOMEDCT_US|EPILEPSY, BENIGN NEONATAL, 1, AND/OR MYOKYMIA
C2751195|T047||SNOMEDCT_US|EPILEPSY, BENIGN NEONATAL, 1, AND-OR MYOKYMIA
C1845543|T047||SNOMEDCT_US|MRXSH
C1845543|T047||SNOMEDCT_US|MRXE
C1845543|T047||SNOMEDCT_US|MENTAL RETARDATION, X-LINKED, SYNDROMIC, HEDERA TYPE
C1845543|T047||SNOMEDCT_US|MENTAL RETARDATION, X-LINKED, WITH EPILEPSY
C1836824|T047|722762005|SNOMEDCT_US|AMISH INFANTILE EPILEPSY SYNDROME|GM3 SYNTHASE DEFICIENCY
C1836824|T047|722762005|SNOMEDCT_US|GM3 SYNTHASE DEFICIENCY|GM3 SYNTHASE DEFICIENCY
C1836824|T047|722762005|SNOMEDCT_US|EPILEPSY SYNDROME, INFANTILE-ONSET SYMPTOMATIC|GM3 SYNTHASE DEFICIENCY
C1836824|T047|722762005|SNOMEDCT_US|SALT AND PEPPER MENTAL RETARDATION SYNDROME|GM3 SYNTHASE DEFICIENCY
C1843852|T047|699328003|SNOMEDCT_US|SPINOCEREBELLAR ATAXIA WITH EPILEPSY|MYOCLONIC EPILEPSY MYOPATHY SENSORY ATAXIA (DISORDER)
C1843852|T047|699328003|SNOMEDCT_US|MYOCLONIC EPILEPSY MYOPATHY SENSORY ATAXIA|MYOCLONIC EPILEPSY MYOPATHY SENSORY ATAXIA (DISORDER)
C1843852|T047|699328003|SNOMEDCT_US|MYOCLONIC EPILEPSY MYOPATHY SENSORY ATAXIA |MYOCLONIC EPILEPSY MYOPATHY SENSORY ATAXIA (DISORDER)
C1843852|T047|699328003|SNOMEDCT_US|MEMSA - MYOCLONIC EPILEPSY MYOPATHY SENSORY ATAXIA|MYOCLONIC EPILEPSY MYOPATHY SENSORY ATAXIA (DISORDER)
C1970203|T047||SNOMEDCT_US|POLYHYDRAMNIOS, MEGALENCEPHALY, AND SYMPTOMATIC EPILEPSY
C1970203|T047||SNOMEDCT_US|PMSE SYNDROME
C1832437|T047||SNOMEDCT_US|MENTAL RETARDATION, MICROCEPHALY, EPILEPSY, AND COARSE FACE
C1853564|T047||SNOMEDCT_US|DEND
C1853564|T047||SNOMEDCT_US|DEVELOPMENTAL DELAY, EPILEPSY, AND NEONATAL DIABETES
C1853623|T047||SNOMEDCT_US|FRYNS-AFTIMOS SYNDROME
C1853623|T047||SNOMEDCT_US|CEREBROOCULOFACIAL LYMPHATIC SYNDROME
C1853623|T047||SNOMEDCT_US|PACHYGYRIA, MENTAL RETARDATION, EPILEPSY, AND CHARACTERISTIC FACIES
C1853623|T047||SNOMEDCT_US|MENTAL RETARDATION WITH EPILEPSY AND CHARACTERISTIC FACIES
C1853623|T047||SNOMEDCT_US|COFL SYNDROME
C2678194|T047|702354007|SNOMEDCT_US|MENTAL RETARDATION, X-LINKED, SYNDROMIC, CHRISTIANSON TYPE|X-LINKED MENTAL RETARDATION SYNDROME, CHRISTIANSON TYPE
C2678194|T047|702354007|SNOMEDCT_US|MRXSCH|X-LINKED MENTAL RETARDATION SYNDROME, CHRISTIANSON TYPE
C2678194|T047|702354007|SNOMEDCT_US|MENTAL RETARDATION, MICROCEPHALY, EPILEPSY, AND ATAXIA SYNDROME|X-LINKED MENTAL RETARDATION SYNDROME, CHRISTIANSON TYPE
C2678194|T047|702354007|SNOMEDCT_US|ANGELMAN-LIKE SYNDROME, X-LINKED|X-LINKED MENTAL RETARDATION SYNDROME, CHRISTIANSON TYPE
C2678194|T047|702354007|SNOMEDCT_US|CHRISTIANSON SYNDROME |X-LINKED MENTAL RETARDATION SYNDROME, CHRISTIANSON TYPE
C2678194|T047|702354007|SNOMEDCT_US|CHRISTIANSON SYNDROME|X-LINKED MENTAL RETARDATION SYNDROME, CHRISTIANSON TYPE
C2678194|T047|702354007|SNOMEDCT_US|INTELLECTUAL DEFICIT, X-LINKED, SOUTH AFRICAN TYPE|X-LINKED MENTAL RETARDATION SYNDROME, CHRISTIANSON TYPE
C2678194|T047|702354007|SNOMEDCT_US|X-LINKED MENTAL RETARDATION SYNDROME, CHRISTIANSON TYPE |X-LINKED MENTAL RETARDATION SYNDROME, CHRISTIANSON TYPE
C2678194|T047|702354007|SNOMEDCT_US|X-LINKED INTELLECTUAL DEFICIT, SOUTH AFRICAN TYPE|X-LINKED MENTAL RETARDATION SYNDROME, CHRISTIANSON TYPE
C2678194|T047|702354007|SNOMEDCT_US|X-LINKED MENTAL RETARDATION SYNDROME, CHRISTIANSON TYPE|X-LINKED MENTAL RETARDATION SYNDROME, CHRISTIANSON TYPE
C3837709|T047||SNOMEDCT_US|EPILEPSY, NOT INTRACTABLE, WITHOUT STATUS EPILEPTICUS
C3837709|T047||SNOMEDCT_US|EPILEPSY NOT INTRACTABLE WITHOUT STATUS EPILEPTICUS
C3837709|T047||SNOMEDCT_US|EPILEPSY, NOT INTRACTABLE, WITHOUT STATUS EPILEPTICUS 
C3826393|T047|100941000119100|SNOMEDCT_US|EPILEPSY IN PREGNANCY|EPILEPSY IN MOTHER COMPLICATING PREGNANCY (DISORDER)
C3826393|T047|100941000119100|SNOMEDCT_US|EPILEPSY IN MOTHER COMPLICATING PREGNANCY |EPILEPSY IN MOTHER COMPLICATING PREGNANCY (DISORDER)
C3826393|T047|100941000119100|SNOMEDCT_US|EPILEPSY IN MOTHER COMPLICATING PREGNANCY|EPILEPSY IN MOTHER COMPLICATING PREGNANCY (DISORDER)
C3840267|T047|10750951000119106|SNOMEDCT_US|EPILEPSY IN CHILDBIRTH|EPILEPSY IN CHILDBIRTH
C3840267|T047|10750951000119106|SNOMEDCT_US|EPILEPSY IN MOTHER COMPLICATING CHILDBIRTH|EPILEPSY IN CHILDBIRTH
C3840267|T047|10750951000119106|SNOMEDCT_US|EPILEPSY IN MOTHER COMPLICATING CHILDBIRTH |EPILEPSY IN CHILDBIRTH
C0751122|T047|230437002|SNOMEDCT_US|SMEI|SEVERE MYOCLONIC EPILEPSY IN INFANCY (DISORDER)
C0751122|T047|230437002|SNOMEDCT_US|INFANTILE SEVERE MYOCLONIC EPILEPSY|SEVERE MYOCLONIC EPILEPSY IN INFANCY (DISORDER)
C0751122|T047|230437002|SNOMEDCT_US|EIEE6|SEVERE MYOCLONIC EPILEPSY IN INFANCY (DISORDER)
C0751122|T047|230437002|SNOMEDCT_US|SYNDROMES, DRAVET|SEVERE MYOCLONIC EPILEPSY IN INFANCY (DISORDER)
C0751122|T047|230437002|SNOMEDCT_US|DRAVET SYNDROMES|SEVERE MYOCLONIC EPILEPSY IN INFANCY (DISORDER)
C0751122|T047|230437002|SNOMEDCT_US|SYNDROME, DRAVET|SEVERE MYOCLONIC EPILEPSY IN INFANCY (DISORDER)
C0751122|T047|230437002|SNOMEDCT_US|DRAVET SYNDROME|SEVERE MYOCLONIC EPILEPSY IN INFANCY (DISORDER)
C0751122|T047|230437002|SNOMEDCT_US|SEVERE MYOCLONIC EPILEPSY OF INFANCY|SEVERE MYOCLONIC EPILEPSY IN INFANCY (DISORDER)
C0751122|T047|230437002|SNOMEDCT_US|EPILEPTIC ENCEPHALOPATHY, EARLY INFANTILE, 6|SEVERE MYOCLONIC EPILEPSY IN INFANCY (DISORDER)
C0751122|T047|230437002|SNOMEDCT_US|SEVERE INFANTILE MYOCLONIC EPILEPSY|SEVERE MYOCLONIC EPILEPSY IN INFANCY (DISORDER)
C0751122|T047|230437002|SNOMEDCT_US|SEVERE MYOCLONIC EPILEPSY, INFANTILE|SEVERE MYOCLONIC EPILEPSY IN INFANCY (DISORDER)
C0751122|T047|230437002|SNOMEDCT_US|EPILEPSY, MYOCLONIC, INFANTILE, SEVERE|SEVERE MYOCLONIC EPILEPSY IN INFANCY (DISORDER)
C0751122|T047|230437002|SNOMEDCT_US|MYOCLONIC EPILEPSY, INFANTILE, SEVERE|SEVERE MYOCLONIC EPILEPSY IN INFANCY (DISORDER)
C0751122|T047|230437002|SNOMEDCT_US|MYOCLONIC EPILEPSY, SEVERE, OF INFANCY|SEVERE MYOCLONIC EPILEPSY IN INFANCY (DISORDER)
C0751122|T047|230437002|SNOMEDCT_US|MYOCLONIC EPILEPSY, SEVERE INFANTILE|SEVERE MYOCLONIC EPILEPSY IN INFANCY (DISORDER)
C0751122|T047|230437002|SNOMEDCT_US|SEVERE MYOCLONIC EPILEPSY IN INFANCY|SEVERE MYOCLONIC EPILEPSY IN INFANCY (DISORDER)
C0751122|T047|230437002|SNOMEDCT_US|SEVERE MYOCLONIC EPILEPSY IN INFANCY |SEVERE MYOCLONIC EPILEPSY IN INFANCY (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|BECTS|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|CENTRALOPATHIC EPILEPSY|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|BENIGN ROLANDIC EPILEPSY|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|EPILEPSIES, CENTROTEMPORAL|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|EPILEPSY, CENTRALOPATHIC|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|ROLANDIC EPILEPSY, BENIGN|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|EPILEPSY, BENIGN ROLANDIC|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|EPILEPSIES, CENTRALOPATHIC|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|CENTROTEMPORAL EPILEPSIES|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|CENTRALOPATHIC EPILEPSIES|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|BENIGN CHILDHOOD EPILEPSY WITH CENTRO TEMPORAL SPIKES|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE |BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|BENIGN EPILEPSY OF CHILDHOOD WITH CENTROTEMPORAL SPIKES|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKES|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|BRE|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|TEMPORAL-CENTRAL FOCAL EPILEPSY|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|CENTROTEMPORAL EPILEPSY|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|BCECTS|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|BENIGN ROLANDIC EPILEPSY OF CHILDHOOD|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|EPILEPSY, CENTROTEMPORAL|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|BENIGN CHILDHOOD EPILEPSY WITH CENTRO-TEMPORAL SPIKES|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|BENIGN EPILEPSY WITH CENTROTEMPORAL SPIKES|BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C2363129|T047|193024005|SNOMEDCT_US|BENIGN ROLANDIC EPILEPSY |BENIGN CHILDHOOD EPILEPSY WITH CENTROTEMPORAL SPIKE (DISORDER)
C3889476|T047||SNOMEDCT_US|BENIGN FAMILIAL NEONATAL SEIZURES
C3889476|T047||SNOMEDCT_US|BENIGN FAMILIAL CONVULSIONS
C3889476|T047||SNOMEDCT_US|BENIGN FAMILAL NEONATAL SEIZURES
C3889476|T047||SNOMEDCT_US|BENIGN FAMILIAL CONVULSION
C1846385|T047||SNOMEDCT_US|FOCAL CORTICAL DYSPLASIA OF TAYLOR
C1846385|T047||SNOMEDCT_US|FCDT
C1846385|T047||SNOMEDCT_US|CORTICAL DYSPLASIA OF TAYLOR
C1846385|T047||SNOMEDCT_US|FOCAL CORTICAL DYSPLASIA, TYPE 2
C1846385|T047||SNOMEDCT_US|FOCAL CORTICAL DYSPLASIA, TYPE II
C4064621|T047||SNOMEDCT_US|MIGRAINE TRIGGERED SEIZURES WITHOUT INTRACTABLE MIGRAINE W/O STATUS MIGRAINOSUS
C4064621|T047||SNOMEDCT_US|MIGRAINE TRIGGERED SEIZURES WITHOUT INTRACTABLE MIGRAINE WITHOUT STATUS MIGRAINOSUS
C4064621|T047||SNOMEDCT_US|MIGRAINE TRIGGERED SEIZURES WITHOUT INTRACTABLE MIGRAINE WITHOUT STATUS MIGRAINOSUS 
C4064624|T047||SNOMEDCT_US|MIGRAINE TRIGGERED SEIZURES WITH INTRACTABLE MIGRAINE WITHOUT STATUS MIGRAINOSUS
C4064624|T047||SNOMEDCT_US|MIGRAINE TRIGGERED SEIZURES WITH INTRACTABLE MIGRAINE WITHOUT STATUS MIGRAINOSUS 
C4064623|T047||SNOMEDCT_US|MIGRAINE TRIGGERED SEIZURES WITHOUT INTRACTABLE MIGRAINE 
C4064623|T047||SNOMEDCT_US|MIGRAINE TRIGGERED SEIZURES WITHOUT INTRACTABLE MIGRAINE
C4064622|T047||SNOMEDCT_US|MIGRAINE TRIGGERED SEIZURES WITHOUT INTRACTABLE MIGRAINE WITH STATUS MIGRAINOSUS 
C4064622|T047||SNOMEDCT_US|MIGRAINE TRIGGERED SEIZURES WITHOUT INTRACTABLE MIGRAINE WITH STATUS MIGRAINOSUS
C0270825|T047|2198002|SNOMEDCT_US|VISCERAL EPILEPSY|VISCERAL EPILEPSY (DISORDER)
C0270825|T047|2198002|SNOMEDCT_US|VISCERAL EPILEPSY |VISCERAL EPILEPSY (DISORDER)
C0270825|T047|2198002|SNOMEDCT_US|EPILEPSY; VISCERAL|VISCERAL EPILEPSY (DISORDER)
C0270825|T047|2198002|SNOMEDCT_US|VISCERAL; EPILEPTIC|VISCERAL EPILEPSY (DISORDER)
C0270825|T047|2198002|SNOMEDCT_US|EPILEPSY, VISCERAL|VISCERAL EPILEPSY (DISORDER)
C0270824|T047|39194005|SNOMEDCT_US|VISUAL PARTIAL SIMPLE SEIZURE |VISUAL EPILEPSY (DISORDER)
C0270824|T047|39194005|SNOMEDCT_US|VISUAL PARTIAL SIMPLE SEIZURE|VISUAL EPILEPSY (DISORDER)
C0270824|T047|39194005|SNOMEDCT_US|SEIZURE, VISUAL|VISUAL EPILEPSY (DISORDER)
C0270824|T047|39194005|SNOMEDCT_US|VISUAL SEIZURE|VISUAL EPILEPSY (DISORDER)
C0270824|T047|39194005|SNOMEDCT_US|VISUAL SEIZURES|VISUAL EPILEPSY (DISORDER)
C0270824|T047|39194005|SNOMEDCT_US|SEIZURES, VISUAL|VISUAL EPILEPSY (DISORDER)
C0270824|T047|39194005|SNOMEDCT_US|VISUAL EPILEPSY|VISUAL EPILEPSY (DISORDER)
C0270824|T047|39194005|SNOMEDCT_US|VISUAL EPILEPSY |VISUAL EPILEPSY (DISORDER)
C0270824|T047|39194005|SNOMEDCT_US|EPILEPSY; VISUAL|VISUAL EPILEPSY (DISORDER)
C0270824|T047|39194005|SNOMEDCT_US|VISUAL; EPILEPTIC|VISUAL EPILEPSY (DISORDER)
C0270824|T047|39194005|SNOMEDCT_US|EPILEPSY, VISUAL|VISUAL EPILEPSY (DISORDER)
C0347873|T047|193002005|SNOMEDCT_US|PSYCHOSENSORY EPILEPSY|PSYCHOSENSORY EPILEPSY (DISORDER)
C0347873|T047|193002005|SNOMEDCT_US|PSYCHOSENSORY EPILEPSY |PSYCHOSENSORY EPILEPSY (DISORDER)
C0347873|T047|193002005|SNOMEDCT_US|EPILEPSY; PSYCHOSENSORY|PSYCHOSENSORY EPILEPSY (DISORDER)
C0347873|T047|193002005|SNOMEDCT_US|PSYCHOSENSORY; EPILEPTIC|PSYCHOSENSORY EPILEPSY (DISORDER)
C0347873|T047|193002005|SNOMEDCT_US|EPILEPSY, PSYCHOSENSORY|PSYCHOSENSORY EPILEPSY (DISORDER)
C0347874|T047|193008009|SNOMEDCT_US|SOMATOSENSORY EPILEPSY|SOMATOSENSORY EPILEPSY (DISORDER)
C0347874|T047|193008009|SNOMEDCT_US|SOMATOSENSORY EPILEPSY |SOMATOSENSORY EPILEPSY (DISORDER)
C0347874|T047|193008009|SNOMEDCT_US|EPILEPSY; SOMATOSENSORY|SOMATOSENSORY EPILEPSY (DISORDER)
C0347874|T047|193008009|SNOMEDCT_US|SOMATOSENSORY; EPILEPTIC|SOMATOSENSORY EPILEPSY (DISORDER)
C0347874|T047|193008009|SNOMEDCT_US|EPILEPSY, SOMATOSENSORY|SOMATOSENSORY EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|EPILEPSIES, TONIC-CLONIC|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|EPILEPSY, TONIC CLONIC|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|EPILEPSY, TONIC-CLONIC|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|GRAND MAL EPILEPSY|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC-CLONIC EPILEPSIES|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC-CLONIC EPILEPSY|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC CLONIC CONVULSION DIS|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|MAJOR MOTOR SEIZURE DIS|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|SEIZURE DIS TONIC CLONIC|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC CLONIC SEIZURE DIS|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|GRAND MAL SEIZURE DIS|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|SEIZURE DIS GRAND MAL|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|SEIZURE DIS MAJOR MOTOR|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|GENERALIZED CONVULSIVE TONIC-CLONIC SEIZURE|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|GENERALIZED CONVULSIVE GRAND MAL SEIZURE|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC-CLONIC EPILEPSY |TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|CONVULSION DISORDER, TONIC-CLONIC|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|CONVULSION DISORDERS, TONIC-CLONIC|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|DISORDER, TONIC-CLONIC CONVULSION|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|DISORDERS, TONIC-CLONIC CONVULSION|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC CLONIC CONVULSION DISORDER|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC-CLONIC CONVULSION DISORDERS|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|CONVULSION SYNDROME, TONIC-CLONIC|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|CONVULSION SYNDROMES, TONIC-CLONIC|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|SYNDROME, TONIC-CLONIC CONVULSION|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|SYNDROMES, TONIC-CLONIC CONVULSION|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC CLONIC CONVULSION SYNDROME|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC-CLONIC CONVULSION SYNDROMES|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|CONVULSION, TONIC CLONIC|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|CONVULSIONS, TONIC CLONIC|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC CLONIC CONVULSION|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|DISORDER, TONIC-CLONIC SEIZURE|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|DISORDERS, TONIC-CLONIC SEIZURE|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|SEIZURE DISORDER, TONIC-CLONIC|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|SEIZURE DISORDERS, TONIC-CLONIC|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC CLONIC SEIZURE DISORDER|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC-CLONIC SEIZURE DISORDERS|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|SEIZURE SYNDROME, TONIC-CLONIC|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|SEIZURE SYNDROMES, TONIC-CLONIC|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|SYNDROME, TONIC-CLONIC SEIZURE|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|SYNDROMES, TONIC-CLONIC SEIZURE|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC CLONIC SEIZURE SYNDROME|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC-CLONIC SEIZURE SYNDROMES|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|CONVULSION, GRAND MAL|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|GRAND MAL CONVULSION|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|GRAND MAL CONVULSIONS|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|MAJOR EPILEPSIES|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|MAJOR EPILEPSY|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|MAJOR MOTOR SEIZURE DISORDER|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC-CLONIC CONVULSION SYNDROME|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|EPILEPSY, TONIC-CLONIC [DISEASE/FINDING]|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC CLONIC CONVULSIONS|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|EPILEPSY, MAJOR|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC-CLONIC CONVULSION DISORDER|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|SEIZURE DISORDER, GRAND MAL|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC-CLONIC SEIZURE SYNDROME|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|EPILEPSY, GRAND MAL|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|GRAND MAL SEIZURE DISORDER|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|SEIZURE DISORDER, MAJOR MOTOR|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|CONVULSIONS, GRAND MAL|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|SEIZURE DISORDER, TONIC CLONIC|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC-CLONIC SEIZURE DISORDER|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|EPILEPSY;GRAND MAL|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC-CLONIC CONVULSION|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|CLONIC-TONIC CONVULSIONS|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|GRAND MAL|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|CONVULSION GRAND MAL|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|MAJOR CONVULSION|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|CONVULSIONS GRAND MAL|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|EPILEPSY GRAND MAL|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC/ CLONIC CONVULSIONS|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|GRAND MAL SEIZURE|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|GRAND MAL SEIZURE |TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|TONIC-CLONIC EPILEPSY |TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|EPILEPSY; GRAND MAL|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|EPILEPSY; MAJOR|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|GRAND MAL; EPILEPSY|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|MAJOR; EPILEPTIC|TONIC-CLONIC EPILEPSY (DISORDER)
C0014549|T047|352818000|SNOMEDCT_US|EPILEPTIC SEIZURES, TONIC-CLONIC|TONIC-CLONIC EPILEPSY (DISORDER)
C0472355|T047|230435005|SNOMEDCT_US|EPILEPSY UNDETERMINED WHETHER FOCAL OR GENERALISED|EPILEPSY UNDETERMINED WHETHER FOCAL OR GENERALIZED (DISORDER)
C0472355|T047|230435005|SNOMEDCT_US|EPILEPSY UNDETERMINED WHETHER FOCAL OR GENERALIZED|EPILEPSY UNDETERMINED WHETHER FOCAL OR GENERALIZED (DISORDER)
C0472355|T047|230435005|SNOMEDCT_US|EPILEPSY UNDETERMINED WHETHER FOCAL OR GENERALIZED |EPILEPSY UNDETERMINED WHETHER FOCAL OR GENERALIZED (DISORDER)
C0438419|T047|193011005|SNOMEDCT_US|UNILATERAL EPILEPSY |UNILATERAL EPILEPSY (SITUATION)
C0438419|T047|193011005|SNOMEDCT_US|UNILATERAL EPILEPSY |UNILATERAL EPILEPSY (SITUATION)
C0438419|T047|193011005|SNOMEDCT_US|UNILATERAL EPILEPSY|UNILATERAL EPILEPSY (SITUATION)
C0477372|T047|194492004|SNOMEDCT_US|OTHER STATUS EPILEPTICUS|[X]OTHER STATUS EPILEPTICUS (DISORDER)
C0477372|T047|194492004|SNOMEDCT_US|[X]OTHER STATUS EPILEPTICUS|[X]OTHER STATUS EPILEPTICUS (DISORDER)
C0477372|T047|194492004|SNOMEDCT_US|[X]OTHER STATUS EPILEPTICUS |[X]OTHER STATUS EPILEPTICUS (DISORDER)
C0270822|T047|49776008|SNOMEDCT_US|CENTERNCEPHALIC EPILEPSY|CENTRENCEPHALIC EPILEPSY (DISORDER)
C0270822|T047|49776008|SNOMEDCT_US|CENTRENCEPHALIC EPILEPSY |CENTRENCEPHALIC EPILEPSY (DISORDER)
C0270822|T047|49776008|SNOMEDCT_US|CENTRENCEPHALIC EPILEPSY|CENTRENCEPHALIC EPILEPSY (DISORDER)
C0270822|T047|49776008|SNOMEDCT_US|CENTRENCEPHALIC ABSENCE|CENTRENCEPHALIC EPILEPSY (DISORDER)
C0270822|T047|49776008|SNOMEDCT_US|CENTERNCEPHALIC ABSENCE|CENTRENCEPHALIC EPILEPSY (DISORDER)
C0347869|T047|192982004|SNOMEDCT_US|AKINETIC EPILEPSY|EPILEPTIC SEIZURES - AKINETIC (FINDING)
C0347869|T047|192982004|SNOMEDCT_US|AKINETIC EPILEPSIES|EPILEPTIC SEIZURES - AKINETIC (FINDING)
C0347869|T047|192982004|SNOMEDCT_US|EPILEPSIES, AKINETIC|EPILEPTIC SEIZURES - AKINETIC (FINDING)
C0347869|T047|192982004|SNOMEDCT_US|AKINETIC SEIZURES|EPILEPTIC SEIZURES - AKINETIC (FINDING)
C0347869|T047|192982004|SNOMEDCT_US|EPILEPSY, AKINETIC|EPILEPTIC SEIZURES - AKINETIC (FINDING)
C0347869|T047|192982004|SNOMEDCT_US|EPILEPTIC SEIZURES - AKINETIC|EPILEPTIC SEIZURES - AKINETIC (FINDING)
C0347869|T047|192982004|SNOMEDCT_US|EPILEPTIC SEIZURES - AKINETIC |EPILEPTIC SEIZURES - AKINETIC (FINDING)
C0347869|T047|192982004|SNOMEDCT_US|EPILEPSY; AKINETIC|EPILEPTIC SEIZURES - AKINETIC (FINDING)
C0347869|T047|192982004|SNOMEDCT_US|AKINETIC; EPILEPTIC|EPILEPTIC SEIZURES - AKINETIC (FINDING)
C0347869|T047|192982004|SNOMEDCT_US|AKINETIC; SEIZURES|EPILEPTIC SEIZURES - AKINETIC (FINDING)
C0347869|T047|192982004|SNOMEDCT_US|SEIZURE; AKINETIC|EPILEPTIC SEIZURES - AKINETIC (FINDING)
C0347869|T047|192982004|SNOMEDCT_US|SEIZURES, AKINETIC|EPILEPTIC SEIZURES - AKINETIC (FINDING)
C0347870|T047|192991000|SNOMEDCT_US|EPILEPTIC SEIZURES - CLONIC|EPILEPTIC SEIZURES - CLONIC (FINDING)
C0347870|T047|192991000|SNOMEDCT_US|EPILEPTIC SEIZURES - CLONIC |EPILEPTIC SEIZURES - CLONIC (FINDING)
C0347870|T047|192991000|SNOMEDCT_US|EPILEPTIC SEIZURES, CLONIC|EPILEPTIC SEIZURES - CLONIC (FINDING)
C0086241|T047|192993002|SNOMEDCT_US|EPILEPSIES, TONIC|EPILEPTIC SEIZURES - TONIC (FINDING)
C0086241|T047|192993002|SNOMEDCT_US|TONIC EPILEPSIES|EPILEPTIC SEIZURES - TONIC (FINDING)
C0086241|T047|192993002|SNOMEDCT_US|TONIC EPILEPSY|EPILEPTIC SEIZURES - TONIC (FINDING)
C0086241|T047|192993002|SNOMEDCT_US|EPILEPTIC SEIZURES - TONIC|EPILEPTIC SEIZURES - TONIC (FINDING)
C0086241|T047|192993002|SNOMEDCT_US|EPILEPTIC SEIZURES - TONIC |EPILEPTIC SEIZURES - TONIC (FINDING)
C0086241|T047|192993002|SNOMEDCT_US|EPILEPSY; TONIC|EPILEPTIC SEIZURES - TONIC (FINDING)
C0086241|T047|192993002|SNOMEDCT_US|TONIC; EPILEPTIC|EPILEPTIC SEIZURES - TONIC (FINDING)
C0086241|T047|192993002|SNOMEDCT_US|EPILEPSY, TONIC|EPILEPTIC SEIZURES - TONIC (FINDING)
C0086241|T047|192993002|SNOMEDCT_US|EPILEPTIC SEIZURES, TONIC|EPILEPTIC SEIZURES - TONIC (FINDING)
C0422855|T047|10800005|SNOMEDCT_US|SEIZURE, VERTIGINOUS|VERTIGINOUS SEIZURE (DISORDER)
C0422855|T047|10800005|SNOMEDCT_US|VERTIGINOUS SEIZURE|VERTIGINOUS SEIZURE (DISORDER)
C0422855|T047|10800005|SNOMEDCT_US|VERTIGINOUS SEIZURES|VERTIGINOUS SEIZURE (DISORDER)
C0422855|T047|10800005|SNOMEDCT_US|SEIZURE, VESTIBULAR|VERTIGINOUS SEIZURE (DISORDER)
C0422855|T047|10800005|SNOMEDCT_US|VESTIBULAR SEIZURE|VERTIGINOUS SEIZURE (DISORDER)
C0422855|T047|10800005|SNOMEDCT_US|VESTIBULAR SEIZURES|VERTIGINOUS SEIZURE (DISORDER)
C0422855|T047|10800005|SNOMEDCT_US|VERTIGINOUS SEIZURE |VERTIGINOUS SEIZURE (DISORDER)
C0422855|T047|10800005|SNOMEDCT_US|SEIZURES, VERTIGINOUS|VERTIGINOUS SEIZURE (DISORDER)
C0422855|T047|10800005|SNOMEDCT_US|SEIZURES, VESTIBULAR|VERTIGINOUS SEIZURE (DISORDER)
C0422855|T047|10800005|SNOMEDCT_US|EPILEPTIC VERTIGO|VERTIGINOUS SEIZURE (DISORDER)
C0422855|T047|10800005|SNOMEDCT_US|VERTIGINOUS EPILEPSY|VERTIGINOUS SEIZURE (DISORDER)
C0422855|T047|10800005|SNOMEDCT_US|EPILEPTIC VERTIGO |VERTIGINOUS SEIZURE (DISORDER)
C0422855|T047|10800005|SNOMEDCT_US|EPILEPTIC; VERTIGO|VERTIGINOUS SEIZURE (DISORDER)
C0422855|T047|10800005|SNOMEDCT_US|VERTIGO; EPILEPTIC|VERTIGINOUS SEIZURE (DISORDER)
C0422855|T047|10800005|SNOMEDCT_US|VERTIGINOUS SEIZURE |VERTIGINOUS SEIZURE (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|CONVULSIONS OF NEWBORN|CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|CONVULSIONS IN NEWBORN |CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|CONVULSIONS IN NEWBORN|CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|CONVULSION NEONATAL|CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|CONVULSIONS IN NEWBORN |CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|NEONATAL SEIZURE|CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|NEONATAL CONVULSION|CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|NEONATAL FIT|CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|NEONATAL SEIZURES|CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|CONVULSIONS NEONATAL|CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|CONVULSIONS IN THE NEWBORN|CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|FITS IN THE NEWBORN|CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|SEIZURES IN THE NEWBORN|CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|FITS IN NEWBORN|CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|NEONATAL CONVULSIONS|CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|SEIZURES IN NEWBORN|CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|CONVULSIONS IN THE NEWBORN |CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|CONVULSIONS; NEONATAL|CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|CONVULSIONS; NEWBORN|CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|FIT; NEWBORN|CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|NEONATAL; CONVULSIONS|CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|NEWBORN; CONVULSIONS|CONVULSIONS IN THE NEWBORN (DISORDER)
C0159020|T047|87476004|SNOMEDCT_US|NEWBORN; FIT|CONVULSIONS IN THE NEWBORN (DISORDER)
C0270826|T047|77450009|SNOMEDCT_US|UNCLASSIFIED EPILEPTIC SEIZURES|UNCLASSIFIED EPILEPTIC SEIZURES (DISORDER)
C0270826|T047|77450009|SNOMEDCT_US|UNCLASSIFIED EPILEPTIC SEIZURES |UNCLASSIFIED EPILEPTIC SEIZURES (DISORDER)
C0393707|T047|230431001|SNOMEDCT_US|SITUATION-RELATED SEIZURES|SITUATION-RELATED SEIZURES (DISORDER)
C0393707|T047|230431001|SNOMEDCT_US|SITUATION-RELATED SEIZURES |SITUATION-RELATED SEIZURES (DISORDER)
C1299598|T047|371022006|SNOMEDCT_US|SEIZURES DUE TO METABOLIC DISORDER |SEIZURES DUE TO METABOLIC DISORDER (DISORDER)
C1299598|T047|371022006|SNOMEDCT_US|SEIZURES DUE TO METABOLIC DISORDER|SEIZURES DUE TO METABOLIC DISORDER (DISORDER)
C0857345|T047||SNOMEDCT_US|LATE ONSET EPILEPSY
C1328935|T047||SNOMEDCT_US|NOCTURNAL FOCAL LOBE EPILEPSY
C0553587|T047|192999003|SNOMEDCT_US|EPILEPSY, PARTIAL, WITH IMPAIRMENT OF CONSCIOUSNESS|PARTIAL EPILEPSY WITH IMPAIRMENT OF CONSCIOUSNESS (DISORDER)
C0553587|T047|192999003|SNOMEDCT_US|PARTIAL EPILEPSY WITH IMPAIRMENT OF CONSCIOUSNESS NOS|PARTIAL EPILEPSY WITH IMPAIRMENT OF CONSCIOUSNESS (DISORDER)
C0553587|T047|192999003|SNOMEDCT_US|PARTIAL EPILEPSY WITH IMPAIRMENT OF CONSCIOUSNESS NOS |PARTIAL EPILEPSY WITH IMPAIRMENT OF CONSCIOUSNESS (DISORDER)
C0553587|T047|192999003|SNOMEDCT_US|PARTIAL EPILEPSY, WITH IMPAIRMENT OF CONSCIOUSNESS|PARTIAL EPILEPSY WITH IMPAIRMENT OF CONSCIOUSNESS (DISORDER)
C0553587|T047|192999003|SNOMEDCT_US|PARTIAL EPILEPSY WITH IMPAIRMENT OF CONSCIOUSNESS|PARTIAL EPILEPSY WITH IMPAIRMENT OF CONSCIOUSNESS (DISORDER)
C0553587|T047|192999003|SNOMEDCT_US|PARTIAL EPILEPSY WITH IMPAIRMENT OF CONSCIOUSNESS |PARTIAL EPILEPSY WITH IMPAIRMENT OF CONSCIOUSNESS (DISORDER)
C0544645|T047||SNOMEDCT_US|FOCAL SENSORY SEIZURES
C0544645|T047||SNOMEDCT_US|SEIZURE, FOCAL SENSORY
C0544645|T047||SNOMEDCT_US|SEIZURES, FOCAL SENSORY
C0544645|T047||SNOMEDCT_US|SENSORY SEIZURE, FOCAL
C0544645|T047||SNOMEDCT_US|SENSORY SEIZURES, FOCAL
C0544645|T047||SNOMEDCT_US|PARTIAL SENSORY SEIZURES
C0544645|T047||SNOMEDCT_US|SEIZURE, PARTIAL SENSORY
C0544645|T047||SNOMEDCT_US|SEIZURES, PARTIAL SENSORY
C0544645|T047||SNOMEDCT_US|SENSORY SEIZURE, PARTIAL
C0544645|T047||SNOMEDCT_US|SENSORY SEIZURES, PARTIAL
C0544645|T047||SNOMEDCT_US|PARTIAL SENSORY SEIZURE
C0544645|T047||SNOMEDCT_US|FOCAL SENSORY SEIZURE
C0270854|T047|71831005|SNOMEDCT_US|EPILEPSY, SYMPTOMATIC GENERALIZED|SYMPTOMATIC GENERALIZED EPILEPSY (DISORDER)
C0270854|T047|71831005|SNOMEDCT_US|GENERALIZED EPILEPSY, SYMPTOMATIC|SYMPTOMATIC GENERALIZED EPILEPSY (DISORDER)
C0270854|T047|71831005|SNOMEDCT_US|SYMPTOMATIC GENERALIZED EPILEPSY|SYMPTOMATIC GENERALIZED EPILEPSY (DISORDER)
C0270854|T047|71831005|SNOMEDCT_US|SYMPTOMATIC GENERALISED EPILEPSY|SYMPTOMATIC GENERALIZED EPILEPSY (DISORDER)
C0270854|T047|71831005|SNOMEDCT_US|SYMPTOMATIC GENERALIZED EPILEPSY |SYMPTOMATIC GENERALIZED EPILEPSY (DISORDER)
C0270854|T047|71831005|SNOMEDCT_US|SYMPTOMATIC GENERALIZED EPILEPSY, NOS|SYMPTOMATIC GENERALIZED EPILEPSY (DISORDER)
C0154721|T047||SNOMEDCT_US|EPILEPSY, UNSPECIFIED, WITHOUT MENTION OF INTRACTABLE EPILEPSY
C0154721|T047||SNOMEDCT_US|EPILEP NOS W/O INTR EPIL
C0154722|T047||SNOMEDCT_US|EPILEPSY, UNSPECIFIED, WITH INTRACTABLE EPILEPSY
C0154722|T047||SNOMEDCT_US|EPILEPSY NOS W INTR EPIL
C1395129|T047||SNOMEDCT_US|DEMENTIA; EPILEPSY (ETIOLOGY)
C1395129|T047||SNOMEDCT_US|DEMENTIA; EPILEPSY (MANIFESTATION)
C1395129|T047||SNOMEDCT_US|EPILEPSY; DEMENTIA (ETIOLOGY)
C1395129|T047||SNOMEDCT_US|EPILEPSY; DEMENTIA (MANIFESTATION)
C1387228|T047||SNOMEDCT_US|POSTICTAL IN EPILEPSY; AMNESIA
C1387228|T047||SNOMEDCT_US|AMNESIA; POSTICTAL IN EPILEPSY
C1392243|T047||SNOMEDCT_US|CEREBRAL; DYSRHYTHMIA
C1394140|T047||SNOMEDCT_US|CORTICAL; DYSRHYTHMIA
C1395970|T047||SNOMEDCT_US|DYSRHYTHMIA; CEREBRAL OR CORTICAL
C0391957|T047||SNOMEDCT_US|EPILEPSY; IDIOPATHIC
C0391957|T047||SNOMEDCT_US|IDIOPATHIC; EPILEPTIC
C1397835|T047||SNOMEDCT_US|FUGUE; POSTICTAL IN EPILEPSY
C1397835|T047||SNOMEDCT_US|POSTICTAL IN EPILEPSY; FUGUE
C0751778|T047|267581004|SNOMEDCT_US|EPILEPSIES, PROGRESSIVE MYOCLONIC|PROGRESSIVE MYOCLONIC EPILEPSY (DISORDER)
C0751778|T047|267581004|SNOMEDCT_US|MYOCLONIC EPILEPSIES, PROGRESSIVE|PROGRESSIVE MYOCLONIC EPILEPSY (DISORDER)
C0751778|T047|267581004|SNOMEDCT_US|PROGRESSIVE MYOCLONIC EPILEPSIES|PROGRESSIVE MYOCLONIC EPILEPSY (DISORDER)
C0751778|T047|267581004|SNOMEDCT_US|EPILEPSY, PROGRESSIVE MYOCLONIC|PROGRESSIVE MYOCLONIC EPILEPSY (DISORDER)
C0751778|T047|267581004|SNOMEDCT_US|MYOCLONIC EPILEPSY, PROGRESSIVE|PROGRESSIVE MYOCLONIC EPILEPSY (DISORDER)
C0751778|T047|267581004|SNOMEDCT_US|EPILEPSIES, PROGRESSIVE MYOCLONUS|PROGRESSIVE MYOCLONIC EPILEPSY (DISORDER)
C0751778|T047|267581004|SNOMEDCT_US|EPILEPSY, PROGRESSIVE MYOCLONUS|PROGRESSIVE MYOCLONIC EPILEPSY (DISORDER)
C0751778|T047|267581004|SNOMEDCT_US|MYOCLONUS EPILEPSIES, PROGRESSIVE|PROGRESSIVE MYOCLONIC EPILEPSY (DISORDER)
C0751778|T047|267581004|SNOMEDCT_US|PROGRESSIVE MYOCLONUS EPILEPSY|PROGRESSIVE MYOCLONIC EPILEPSY (DISORDER)
C0751778|T047|267581004|SNOMEDCT_US|PROGRESSIVE MYOCLONIC EPILEPSY|PROGRESSIVE MYOCLONIC EPILEPSY (DISORDER)
C0751778|T047|267581004|SNOMEDCT_US|MYOCLONIC EPILEPSIES, PROGRESSIVE [DISEASE/FINDING]|PROGRESSIVE MYOCLONIC EPILEPSY (DISORDER)
C0751778|T047|267581004|SNOMEDCT_US|PROGRESSIVE MYOCLONUS EPILEPSIES|PROGRESSIVE MYOCLONIC EPILEPSY (DISORDER)
C0751778|T047|267581004|SNOMEDCT_US|PROGRESSIVE MYOCLONIC EPILEPSY |PROGRESSIVE MYOCLONIC EPILEPSY (DISORDER)
C0751778|T047|267581004|SNOMEDCT_US|PROGRESSIVE MYOCLONIC EPILEPSY  [AMBIGUOUS]|PROGRESSIVE MYOCLONIC EPILEPSY (DISORDER)
C0852977|T047||SNOMEDCT_US|EPILEPSY AGGRAVATED
C0852977|T047||SNOMEDCT_US|AGGRAVATED EPILEPSY
C0854109|T047||SNOMEDCT_US|EPILEPSY CONGENITAL
C0854109|T047||SNOMEDCT_US|CONGENITAL EPILEPSY
C0270849|T047|111498005|SNOMEDCT_US|EXTRATEMPORAL EPILEPSY|EXTRATEMPORAL EPILEPSY (DISORDER)
C0270849|T047|111498005|SNOMEDCT_US|EXTRATEMPORAL EPILEPSY |EXTRATEMPORAL EPILEPSY (DISORDER)
C1332300|T047||SNOMEDCT_US|ANOSOGNOSTIC EPILEPSY
C1857575|T047||SNOMEDCT_US|CONVULSIVE DISORDER, FAMILIAL, WITH PRENATAL OR EARLY ONSET
