C0193388|T060||CPT|BIOPSY OF LIVER 
C3174660|T060||CPT|PATHOLOGY BIOPSY REPORT:FIND:PT:LIVER:NAR
C1524299|T060||CPT|GUIDANCE FOR BIOPSY:FIND:PT:ABDOMEN>LIVER:DOC:RF
C1628488|T060||CPT|CT AND BIOPSY OF LIVER
C1635159|T060||CPT|US SCAN AND BIOPSY OF LIVER
C1955790|T060||CPT|TRANSJUGULAR BIOPSY OF LIVER
C1955791|T060||CPT|TRANSVENOUS LIVER BIOPSY
C2021366|T060||CPT|LIVER BIOPSY IRON (UG/100 MG OF DRY WEIGHT)
C3836930|T060||CPT|LIVER BIOPSY WITH FLUOROSCOPIC GUIDANCE
C3863012|T060||CPT|LIVER BIOPSY, TRANSJUGULAR APPROACH
C3880782|T060||CPT|LIVER BIOPSY PROCEDURE KIT
C0193388|T060||CPT|BIOPSY OF LIVER 
C0193388|T060||CPT|BIOPSY OF LIVER
C0193388|T060||CPT|LIVER BIOPSY
C0193390|T060|47100|CPT|WEDGE BIOPSY OF LIVER|WEDGE BIOPSY OF LIVER
C0521264|T060||CPT|LAPAROSCOPIC BIOPSY OF LIVER
C0558534|T060||CPT|PERCUTANEOUS LIVER BIOPSY
C0581276|T060|47001|CPT|NEEDLE BIOPSY OF LIVER|NEEDLE BIOPSY OF LIVER
C0842769|T060||CPT|PERCUTANEOUS [CLOSED] LIVER BIOPSY
C0860886|T060||CPT|ULTRASOUND GUIDED LIVER BIOPSY
C1261294|T060|47000|CPT|PERCUTANEOUS NEEDLE BIOPSY LIVER|NEEDLE BIOPSY OF LIVER, ACCESSED THROUGH THE SKIN
C1548877|T060||CPT|CONSENT TYPE - LIVER BIOPSY
C1955790|T060||CPT|TRANSJUGULAR BIOPSY OF LIVER
C1955791|T060||CPT|TRANSVENOUS LIVER BIOPSY
C3522275|T060|47700|CPT|EXPLORATION FOR CONGENITAL ATRESIA OF BILE DUCT WITH LIVER BIOPSY|EXPLORATION FOR CONGENITAL ATRESIA OF BILE DUCT WITH LIVER BIOPSY
C3550399|T060||CPT|INCREASED IRON DEPOSITION SEEN ON LIVER BIOPSY
C0860886|T060||CPT|ULTRASOUND GUIDED LIVER BIOPSY
C0372191|T060|47001|CPT|BIOPSY OF LIVER, NEEDLE; WHEN DONE FOR INDICATED PURPOSE AT TIME OF OTHER MAJOR PROCEDURE (LIST SEPARATELY IN ADDITION TO CODE FOR PRIMARY PROCEDURE)|BX LVR NDL DONE PURPOSE TM OTH MAJOR PX
C0372191|T060|47001|CPT|NEEDLE BIOPSY LIVER ADD-ON|BX LVR NDL DONE PURPOSE TM OTH MAJOR PX
C0372191|T060|47001|CPT|BX LVR NDL DONE PURPOSE TM OTH MAJOR PX|BX LVR NDL DONE PURPOSE TM OTH MAJOR PX
C0176879|T060||CPT|CLOSED LIVER BIOPSY
C0176879|T060||CPT|CLOSED (PERCUTANEOUS) [NEEDLE] BIOPSY OF LIVER
C1955790|T060||CPT|TRANSJUGULAR LIVER BIOPSY
C1955790|T060||CPT|TRANSJUGULAR BIOPSY OF LIVER 
C1955790|T060||CPT|TRANSJUGULAR BIOPSY OF LIVER
C1955790|T060||CPT|TRANSJUGULAR LIVER BX
C2314979|T060||CPT|TRANSJUGULAR BIOPSY OF LIVER USING FLUOROSCOPIC GUIDANCE
C2314979|T060||CPT|TRANSJUGULAR BIOPSY OF LIVER USING FLUOROSCOPIC GUIDANCE 
C0193388|T060||CPT|BIOPSY OF LIVER
C0193388|T060||CPT|LIVER BIOPSY
C0193388|T060||CPT|LIVER BIOPSY 
C0193388|T060||CPT|BIOPSY LIVER
C0193388|T060||CPT|BIOPSY OF LIVER 
C0193388|T060||CPT|BIOPSY OF LIVER, NOS
C2121176|T060||CPT|A LIVER BIOPSY WHEN DONE FOR INDICATED PURPOSE AT TIME OF OTHER MAJOR PROCEDURE
C2121176|T060||CPT|LIVER BIOPSY WHEN DONE FOR INDICATED PURPOSE AT TIME OF OTHER MAJOR PROCEDURE
C2121176|T060||CPT|LIVER BIOPSY WHEN DONE FOR INDICATED PURPOSE AT TIME OF OTHER MAJOR PROCEDURE 
C2021366|T060||CPT|LIVER BIOPSY IRON (UG/100 MG OF DRY WEIGHT) 
C2021366|T060||CPT|LIVER BIOPSY IRON (UG/100 MG OF DRY WEIGHT)
C2021366|T060||CPT|LIVER BIOPSY IRON
C1261294|T060|47000|CPT|BIOPSY OF LIVER, NEEDLE; PERCUTANEOUS|NEEDLE BIOPSY OF LIVER, ACCESSED THROUGH THE SKIN
C1261294|T060|47000|CPT|PERCUTANEOUS NEEDLE BIOPSY LIVER|NEEDLE BIOPSY OF LIVER, ACCESSED THROUGH THE SKIN
C1261294|T060|47000|CPT|PERCUTANEOUS NEEDLE BIOPSY OF LIVER|NEEDLE BIOPSY OF LIVER, ACCESSED THROUGH THE SKIN
C1261294|T060|47000|CPT|PERCUTANEOUS NEEDLE BIOPSY LIVER |NEEDLE BIOPSY OF LIVER, ACCESSED THROUGH THE SKIN
C1261294|T060|47000|CPT|PERCUTANEOUS NEEDLE BIOPSY OF LIVER |NEEDLE BIOPSY OF LIVER, ACCESSED THROUGH THE SKIN
C1261294|T060|47000|CPT|PERCUTANEOUS NEEDLE LIVER BIOPSY |NEEDLE BIOPSY OF LIVER, ACCESSED THROUGH THE SKIN
C1261294|T060|47000|CPT|PERCUTANEOUS NEEDLE LIVER BIOPSY|NEEDLE BIOPSY OF LIVER, ACCESSED THROUGH THE SKIN
C1261294|T060|47000|CPT|BIOPSY LIVER NEEDLE PERCUTANEOUS|NEEDLE BIOPSY OF LIVER, ACCESSED THROUGH THE SKIN
C1261294|T060|47000|CPT|NEEDLE BIOPSY OF LIVER, ACCESSED THROUGH THE SKIN|NEEDLE BIOPSY OF LIVER, ACCESSED THROUGH THE SKIN
C1261294|T060|47000|CPT|NEEDLE BIOPSY OF LIVER|NEEDLE BIOPSY OF LIVER, ACCESSED THROUGH THE SKIN
C0193390|T060|47100|CPT|BIOPSY OF LIVER, WEDGE|WEDGE BIOPSY OF LIVER
C0193390|T060|47100|CPT|WEDGE BIOPSY OF LIVER|WEDGE BIOPSY OF LIVER
C0193390|T060|47100|CPT|WEDGE LIVER BIOPSY|WEDGE BIOPSY OF LIVER
C0193390|T060|47100|CPT|WEDGE LIVER BIOPSY |WEDGE BIOPSY OF LIVER
C0193390|T060|47100|CPT|BIOPSY LIVER WEDGE|WEDGE BIOPSY OF LIVER
C0193390|T060|47100|CPT|WEDGE BIOPSY OF LIVER |WEDGE BIOPSY OF LIVER
C0193393|T060||CPT|PERCUTANEOUS CORE NEEDLE BIOPSY OF LIVER
C0193393|T060||CPT|PERCUTANEOUS CORE NEEDLE BIOPSY OF LIVER 
C0193389|T060||CPT|OPEN LIVER BIOPSY
C0193389|T060||CPT|OPEN BIOPSY OF LIVER
C0193389|T060||CPT|OPEN BIOPSY OF LIVER 
C0193394|T060||CPT|PERCUTANEOUS FINE NEEDLE BIOPSY OF LIVER
C0193394|T060||CPT|PERCUTANEOUS FINE NEEDLE ASPIRATION BIOPSY OF LIVER
C0193394|T060||CPT|PERCUTANEOUS FINE NEEDLE BIOPSY OF LIVER 
C0581276|T060|47001|CPT|NEEDLE BIOPSY OF LIVER|NEEDLE BIOPSY OF LIVER
C0581276|T060|47001|CPT|BIOPSY OF LIVER, NEEDLE|NEEDLE BIOPSY OF LIVER
C0581276|T060|47001|CPT|NEEDLE BIOPSY OF LIVER |NEEDLE BIOPSY OF LIVER
C0521264|T060||CPT|LAPAROSCOPIC LIVER BIOPSY
C0521264|T060||CPT|LAPAROSCOPIC LIVER BX
C0521264|T060||CPT|LAPAROSCOPIC BIOPSY OF LIVER 
C0521264|T060||CPT|LAPAROSCOPIC BIOPSY OF LIVER
C0521264|T060||CPT|LAPAROSCOPIC BIOPSY OF LIVER, NOS
C0400397|T060||CPT|DIAGNOSTIC ENDOSCOPIC EXAMINATION OF LIVER AND BIOPSY OF LESION OF LIVER USING LAPAROSCOPE
C0400397|T060||CPT|DIAGNOSTIC ENDOSCOPIC EXAMINATION OF LIVER AND BIOPSY OF LESION OF LIVER USING LAPAROSCOPE 
C0400418|T060||CPT|BIOPSY OF LIVER NEC 
C0400418|T060||CPT|BIOPSY OF LIVER NEC
C3836930|T060||CPT|LIVER BIOPSY WITH FLUOROSCOPIC GUIDANCE
C3836930|T060||CPT|LIVER BIOPSY WITH FLUOROSCOPIC GUIDANCE 
C3863012|T060||CPT|LIVER BIOPSY, TRANSJUGULAR APPROACH
C3863012|T060||CPT|LIVER BIOPSY TRANSJUGULAR APPROACH
C3863012|T060||CPT|LIVER BIOPSY, TRANSJUGULAR APPROACH 
C4031824|T060||CPT|BIOPSY LIVER LOCATION 
C4031824|T060||CPT|BIOPSY LIVER LOCATION
C4031823|T060||CPT|BIOPSY LIVER SPECIMEN NO. ______
C4031823|T060||CPT|BIOPSY LIVER SPECIMEN NO. ______ 
C4030893|T060||CPT|BIOPSY OF LIVER MALIGNANT NEOPLASM 
C4030893|T060||CPT|BIOPSY OF LIVER MALIGNANT NEOPLASM
C4030863|T060||CPT|BIOPSY OF LIVER SHOWED CARCINOMA IN SITU
C4030863|T060||CPT|BIOPSY OF LIVER SHOWED CARCINOMA IN SITU 
C4030863|T060||CPT|BX LIVER SHOWED CARCINOMA IN SITU
C4030881|T060||CPT|BIOPSY OF LIVER SHOWED BENIGN NEOPLASM
C4030881|T060||CPT|BIOPSY OF LIVER SHOWED BENIGN NEOPLASM 
C0400419|T060||CPT|BIOPSY OF LIVER LESION
C0400419|T060||CPT|BIOPSY OF LIVER LESION 
C0558534|T060||CPT|PERCUTANEOUS LIVER BIOPSY
C0558534|T060||CPT|PERCUTANEOUS LIVER BIOPSY 
C0558560|T060||CPT|SURGICAL BIOPSY OF LIVER 
C0558560|T060||CPT|SURGICAL BIOPSY OF LIVER
C0558560|T060||CPT|LIVER: SURGICAL BIOPSY 
C0558560|T060||CPT|LIVER: SURGICAL BIOPSY
C1628488|T060||CPT|CT AND BIOPSY OF LIVER
C1628488|T060||CPT|COMPUTED TOMOGRAPHY AND BIOPSY OF LIVER 
C1628488|T060||CPT|COMPUTED TOMOGRAPHY AND BIOPSY OF LIVER
C1635159|T060||CPT|US SCAN AND BIOPSY OF LIVER
C1635159|T060||CPT|ULTRASOUND SCAN AND BIOPSY OF LIVER 
C1635159|T060||CPT|ULTRASOUND SCAN AND BIOPSY OF LIVER
C0193392|T060||CPT|OPEN FINE NEEDLE BIOPSY OF LIVER 
C0193392|T060||CPT|OPEN FINE NEEDLE BIOPSY OF LIVER
C0193392|T060||CPT|OPEN FINE NEEDLE ASPIRATION BIOPSY OF LIVER
C0193392|T060||CPT|OPEN FINE NEEDLE ASPIRATION BIOPSY OF LIVER 
C0193392|T060||CPT|OPEN FINE NEEDLE BIOPSY OF LIVER  [AMBIGUOUS]
C3174660|T060||CPT|PATHOLOGY BIOPSY REPORT:FIND:PT:LIVER:NAR
C3174660|T060||CPT|LIVER PATH BX REPORT
C3174660|T060||CPT|PATHOLOGY BIOPSY REPORT:FINDING:POINT IN TIME:LIVER:NARRATIVE
C3174660|T060||CPT|LIVER PATHOLOGY BIOPSY REPORT
C1524299|T060||CPT|FLUOROSCOPY GUIDANCE FOR BIOPSY OF LIVER
C1524299|T060||CPT|LIVER FLR BX GUID
C1524299|T060||CPT|GUIDANCE FOR BIOPSY:FINDING:POINT IN TIME:LIVER:DOCUMENT:XR.FLUOR
C1524299|T060||CPT|GUIDANCE FOR BIOPSY:FIND:PT:LIVER:DOC:XR.FLUOR
C2585711|T060||CPT|BIOPSY OF LIVER USING ULTRASOUND GUIDANCE 
C2585711|T060||CPT|BIOPSY OF LIVER USING ULTRASOUND GUIDANCE
C1960013|T060||CPT|ENDOSCOPIC ULTRASOUND EXAMINATION OF LIVER AND BIOPSY OF LESION OF LIVER 
C1960013|T060||CPT|ENDOSCOPIC ULTRASOUND EXAMINATION OF LIVER AND BIOPSY OF LESION OF LIVER
C3863011|T060||CPT|LIVER BIOPSY TRANSJUGULAR APPROACH WITH FLUOROSCOPIC GUIDANCE
C3863011|T060||CPT|LIVER BIOPSY, TRANSJUGULAR APPROACH WITH FLUOROSCOPIC GUIDANCE 
C3863011|T060||CPT|LIVER BIOPSY, TRANSJUGULAR APPROACH WITH FLUOROSCOPIC GUIDANCE
C0400423|T060||CPT|OPEN WEDGE BIOPSY OF LESION OF LIVER
C0400423|T060||CPT|OPEN WEDGE BIOPSY OF LESION OF LIVER 
C0585492|T060||CPT|LAPAROSCOPIC BIOPSY OF LIVER LESION
C0585492|T060||CPT|LAPAROSCOPIC BIOPSY OF LIVER LESION 
C2315061|T060||CPT|PERCUTANEOUS TRANSJUGULAR BIOPSY OF LIVER USING FLUOROSCOPIC GUIDANCE 
C2315061|T060||CPT|PERCUTANEOUS TRANSJUGULAR BIOPSY OF LIVER USING FLUOROSCOPIC GUIDANCE
C2733386|T060||CPT|PERCUTANEOUS BIOPSY OF LIVER USING ULTRASOUND GUIDANCE 
C2733386|T060||CPT|PERCUTANEOUS BIOPSY OF LIVER USING ULTRASOUND GUIDANCE
C0400422|T060||CPT|PERCUTANEOUS TRANSVASCULAR BIOPSY OF LESION OF LIVER
C0400422|T060||CPT|PERCUTANEOUS TRANSVASCULAR BIOPSY OF LESION OF LIVER 
C2317400|T060||CPT|FINE NEEDLE ASPIRATION BIOPSY OF LIVER
C2317400|T060||CPT|FINE NEEDLE ASPIRATON BIOPSY OF LIVER
C2317400|T060||CPT|FINE NEEDLE ASPIRATION BIOPSY OF LIVER 
C2317400|T060||CPT|FINE NEEDLE ASPIRATON BIOPSY OF LIVER 
C0554070|T060||CPT|NEEDLE BIOPSY OF LIVER NEC
C0554070|T060||CPT|NEEDLE BIOPSY OF LIVER NEC 
C0193391|T060||CPT|OPEN CORE NEEDLE BIOPSY OF LIVER
C0193391|T060||CPT|OPEN CORE NEEDLE BIOPSY OF LIVER 
C0554069|T060||CPT|MENGHINI NEEDLE BIOPSY OF LIVER
C0554069|T060||CPT|MENGHINI NEEDLE BIOPSY OF LIVER 
C0554071|T060||CPT|SHEEBA NEEDLE BIOPSY OF LIVER
C0554071|T060||CPT|SHEEBA NEEDLE BIOPSY OF LIVER 
C2732498|T060||CPT|PERCUTANEOUS NEEDLE BIOPSY OF LIVER USING FLUOROSCOPIC GUIDANCE 
C2732498|T060||CPT|PERCUTANEOUS NEEDLE BIOPSY OF LIVER USING FLUOROSCOPIC GUIDANCE
C3836502|T060||CPT|PERCUTANEOUS NEEDLE LIVER BIOPSY WITH FLUOROSCOPIC GUIDANCE
C3836502|T060||CPT|PERCUTANEOUS NEEDLE LIVER BIOPSY WITH FLUOROSCOPIC GUIDANCE 
C3862599|T060||CPT|PERCUTANEOUS NEEDLE LIVER BIOPSY FINE NEEDLE ASPIRATION 
C3862599|T060||CPT|PERCUTANEOUS NEEDLE LIVER BIOPSY FINE NEEDLE ASPIRATION
