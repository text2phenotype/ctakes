// CUI|TUI|CODE|VOCAB|TXT|PREF TEXT
C000001|T109|1|CUSTOM|Aspirin|Aspirin