C3494624|T053|428061000124105|SNOMEDCT_US|CURRENT HEAVY TOBACCO SMOKER (SNOMED:428071000124103)|LIGHT TOBACCO SMOKER (FINDING)
C3494624|T053|428061000124105|SNOMEDCT_US|CURRENT LIGHT TOBACCO SMOKER (SNOMED:428061000124105)|LIGHT TOBACCO SMOKER (FINDING)
C1880200|T053|428041000124106|SNOMEDCT_US|CURRENT SOME DAY SMOKER	 (SNOMED:428041000124106)|OCCASIONAL TOBACCO SMOKER (FINDING)
C0337671|T053|8517006|SNOMEDCT_US|EX-SMOKER 	FORMER SMOKER(SNOMED:8517006)|EX-SMOKER (LIFE STYLE)
C0425293|T053|266919005|SNOMEDCT_US|NEVER SMOKED TOBACCO 	NEVER SMOKER (SNOMED:266919005)|NEVER SMOKED TOBACCO (LIFE STYLE)
C0337664|T053|77176002|SNOMEDCT_US|SMOKER 	SMOKER, CURRENT STATUS UNKNOWN (SNOMED:77176002)|SMOKER (LIFE STYLE)
C3266136|T053|449868002|SNOMEDCT_US|SMOKES TOBACCO DAILY 	CURRENT EVERY DAY SMOKER (SNOMED:449868002)|CURRENT EVERY DAY SMOKER
C0425306|T053|266927001|SNOMEDCT_US|TOBACCO SMOKING CONSUMPTION UNKNOWN 	UNKNOWN IF EVER SMOKED (SNOMED:266927001)|TOBACCO SMOKING CONSUMPTION UNKNOWN (FINDING)
C3494624|T053|428061000124105|SNOMEDCT_US|LIGHT TOBACCO SMOKER |LIGHT TOBACCO SMOKER (FINDING)
C3494624|T053|428061000124105|SNOMEDCT_US|LIGHT TOBACCO SMOKER|LIGHT TOBACCO SMOKER (FINDING)
C3494624|T053|428061000124105|SNOMEDCT_US|CURRENT LIGHT TOBACCO SMOKER|LIGHT TOBACCO SMOKER (FINDING)
C3494624|T053|428061000124105|SNOMEDCT_US|CURRENT LIGHT TOBACCO SMOKER |LIGHT TOBACCO SMOKER (FINDING)
C1880200|T053|428041000124106|SNOMEDCT_US|SOME DAY SMOKER|OCCASIONAL TOBACCO SMOKER (FINDING)
C1880200|T053|428041000124106|SNOMEDCT_US|NON-DAILY SMOKER|OCCASIONAL TOBACCO SMOKER (FINDING)
C1880200|T053|428041000124106|SNOMEDCT_US|OCCASIONAL SMOKER|OCCASIONAL TOBACCO SMOKER (FINDING)
C1880200|T053|428041000124106|SNOMEDCT_US|CURRENT SOME DAY SMOKER|OCCASIONAL TOBACCO SMOKER (FINDING)
C1880200|T053|428041000124106|SNOMEDCT_US|CURRENT SOME DAY SMOKER |OCCASIONAL TOBACCO SMOKER (FINDING)
C1880200|T053|428041000124106|SNOMEDCT_US|OCCASIONAL TOBACCO SMOKER|OCCASIONAL TOBACCO SMOKER (FINDING)
C1880200|T053|428041000124106|SNOMEDCT_US|OCCASIONAL TOBACCO SMOKER |OCCASIONAL TOBACCO SMOKER (FINDING)
C1880200|T053|428041000124106|SNOMEDCT_US|SOME-DAY SMOKER|OCCASIONAL TOBACCO SMOKER (FINDING)
C3649460|T053||SNOMEDCT_US|CURRENT OCCASIONAL TOBACCO SMOKER
C3649460|T053||SNOMEDCT_US|CURRENT OCCASIONAL TOBACCO SMOKER 
C2114448|T053||SNOMEDCT_US|PREVIOUS HISTORY OF SMOKING
C2114448|T053||SNOMEDCT_US|PREVIOUS HISTORY OF SMOKING 
C3468596|T053||SNOMEDCT_US|FORMER CIGARETTE CHAIN SMOKER
C3468596|T053||SNOMEDCT_US|FORMER CIGARETTE CHAIN SMOKER 
C0337671|T053|8517006|SNOMEDCT_US|FORMER SMOKER|EX-SMOKER (LIFE STYLE)
C0337671|T053|8517006|SNOMEDCT_US|PRIOR SMOKER|EX-SMOKER (LIFE STYLE)
C0337671|T053|8517006|SNOMEDCT_US|PAST TOBACCO SMOKER|EX-SMOKER (LIFE STYLE)
C0337671|T053|8517006|SNOMEDCT_US|EX-SMOKER|EX-SMOKER (LIFE STYLE)
C0337671|T053|8517006|SNOMEDCT_US|EX-SMOKER |EX-SMOKER (LIFE STYLE)
C0337671|T053|8517006|SNOMEDCT_US|PREVIOUS TOBACCO USE|EX-SMOKER (LIFE STYLE)
C0337671|T053|8517006|SNOMEDCT_US|RECOVERED SMOKER|EX-SMOKER (LIFE STYLE)
C0337671|T053|8517006|SNOMEDCT_US|CESSATION OF SMOKING|EX-SMOKER (LIFE STYLE)
C0337671|T053|8517006|SNOMEDCT_US|EX-SMOKER |EX-SMOKER (LIFE STYLE)
C3494626|T053|428081000124100|SNOMEDCT_US|FORMER HEAVY TOBACCO SMOKER |FORMER HEAVY TOBACCO SMOKER (FINDING)
C3494626|T053|428081000124100|SNOMEDCT_US|EX-HEAVY TOBACCO SMOKER|FORMER HEAVY TOBACCO SMOKER (FINDING)
C3494626|T053|428081000124100|SNOMEDCT_US|FORMER HEAVY TOBACCO SMOKER|FORMER HEAVY TOBACCO SMOKER (FINDING)
C3494626|T053|428081000124100|SNOMEDCT_US|FORMER HEAVY TOBACCO SMOKER |FORMER HEAVY TOBACCO SMOKER (FINDING)
C3494627|T053|428091000124102|SNOMEDCT_US|EX-LIGHT TOBACCO SMOKER|FORMER LIGHT TOBACCO SMOKER (FINDING)
C3494627|T053|428091000124102|SNOMEDCT_US|FORMER LIGHT TOBACCO SMOKER|FORMER LIGHT TOBACCO SMOKER (FINDING)
C3494627|T053|428091000124102|SNOMEDCT_US|FORMER LIGHT TOBACCO SMOKER |FORMER LIGHT TOBACCO SMOKER (FINDING)
C3494627|T053|428091000124102|SNOMEDCT_US|FORMER LIGHT TOBACCO SMOKER |FORMER LIGHT TOBACCO SMOKER (FINDING)
C3693442|T053||SNOMEDCT_US|STOPPED SMOKING ___ YEARS AGO
C3693442|T053||SNOMEDCT_US|STOPPED SMOKING ___ YEARS AGO 
C4041321|T053|48031000119106|SNOMEDCT_US|EX-SMOKER FOR MORE THAN 1 YEAR |EX-SMOKER FOR MORE THAN 1 YEAR (FINDING)
C4041321|T053|48031000119106|SNOMEDCT_US|EX-SMOKER FOR MORE THAN 1 YEAR|EX-SMOKER FOR MORE THAN 1 YEAR (FINDING)
C0521323|T053|65909009|SNOMEDCT_US|AGGRESSIVE EX-SMOKER |AGGRESSIVE EX-SMOKER (LIFE STYLE)
C0521323|T053|65909009|SNOMEDCT_US|AGGRESSIVE EX-SMOKER|AGGRESSIVE EX-SMOKER (LIFE STYLE)
C0521323|T053|65909009|SNOMEDCT_US|AGGRESSIVE EX-SMOKER |AGGRESSIVE EX-SMOKER (LIFE STYLE)
C0521323|T053|65909009|SNOMEDCT_US|AGGRESSIVE EX-SMOKER  [AMBIGUOUS]|AGGRESSIVE EX-SMOKER (LIFE STYLE)
C0425314|T053|160621008|SNOMEDCT_US|EX-CIGAR SMOKER|EX-CIGAR SMOKER (LIFE STYLE)
C0425314|T053|160621008|SNOMEDCT_US|EX-CIGAR SMOKER |EX-CIGAR SMOKER (LIFE STYLE)
C0425314|T053|160621008|SNOMEDCT_US|FORMER CIGAR SMOKER |EX-CIGAR SMOKER (LIFE STYLE)
C0425314|T053|160621008|SNOMEDCT_US|FORMER CIGAR SMOKER|EX-CIGAR SMOKER (LIFE STYLE)
C0425314|T053|160621008|SNOMEDCT_US|EX-CIGAR SMOKER |EX-CIGAR SMOKER (LIFE STYLE)
C0459838|T053|281018007|SNOMEDCT_US|EX-CIGARETTE SMOKER|EX-CIGARETTE SMOKER (LIFE STYLE)
C0459838|T053|281018007|SNOMEDCT_US|EX-CIGARETTE SMOKER |EX-CIGARETTE SMOKER (LIFE STYLE)
C0459838|T053|281018007|SNOMEDCT_US|EX-CIGARETTE SMOKER |EX-CIGARETTE SMOKER (LIFE STYLE)
C0425313|T053|160620009|SNOMEDCT_US|EX-PIPE SMOKER|EX-PIPE SMOKER (LIFE STYLE)
C0425313|T053|160620009|SNOMEDCT_US|EX-PIPE SMOKER |EX-PIPE SMOKER (LIFE STYLE)
C0425313|T053|160620009|SNOMEDCT_US|FORMER PIPE SMOKER|EX-PIPE SMOKER (LIFE STYLE)
C0425313|T053|160620009|SNOMEDCT_US|FORMER PIPE SMOKER |EX-PIPE SMOKER (LIFE STYLE)
C0425313|T053|160620009|SNOMEDCT_US|EX-PIPE SMOKER |EX-PIPE SMOKER (LIFE STYLE)
C1261257|T053|360890004|SNOMEDCT_US|INTOLERANT EX-SMOKER|INTOLERANT EX-SMOKER (LIFE STYLE)
C1261257|T053|360890004|SNOMEDCT_US|INTOLERANT EX-SMOKER |INTOLERANT EX-SMOKER (LIFE STYLE)
C1261257|T053|360890004|SNOMEDCT_US|INTOLERANT EX-SMOKER |INTOLERANT EX-SMOKER (LIFE STYLE)
C0425310|T053|160617001|SNOMEDCT_US|STOPPED SMOKING|STOPPED SMOKING (LIFE STYLE)
C0425310|T053|160617001|SNOMEDCT_US|STOPPED SMOKING |STOPPED SMOKING (LIFE STYLE)
C0425310|T053|160617001|SNOMEDCT_US|STOPPED SMOKING |STOPPED SMOKING (LIFE STYLE)
C0521322|T053|53896009|SNOMEDCT_US|TOLERANT EX-SMOKER|TOLERANT EX-SMOKER (LIFE STYLE)
C0521322|T053|53896009|SNOMEDCT_US|TOLERANT EX-SMOKER |TOLERANT EX-SMOKER (LIFE STYLE)
C0521322|T053|53896009|SNOMEDCT_US|TOLERANT EX-SMOKER |TOLERANT EX-SMOKER (LIFE STYLE)
C0558928|T053|160608001|SNOMEDCT_US|EX-LIGHT SMOKER (1-9/DAY) |EX-LIGHT SMOKER (1-9/DAY) (LIFE STYLE)
C0558928|T053|160608001|SNOMEDCT_US|EX-LIGHT SMOKER (1-9/DAY)|EX-LIGHT SMOKER (1-9/DAY) (LIFE STYLE)
C0558928|T053|160608001|SNOMEDCT_US|EX-LIGHT SMOKER (1-9/DAY) |EX-LIGHT SMOKER (1-9/DAY) (LIFE STYLE)
C0558927|T053|160607006|SNOMEDCT_US|EX-TRIVIAL SMOKER (<1/DAY)|EX-TRIVIAL SMOKER (<1/DAY) (LIFE STYLE)
C0558927|T053|160607006|SNOMEDCT_US|EX-TRIVIAL SMOKER (<1/DAY) |EX-TRIVIAL SMOKER (<1/DAY) (LIFE STYLE)
C0558927|T053|160607006|SNOMEDCT_US|EX-TRIVIAL SMOKER (<1/DAY) |EX-TRIVIAL SMOKER (<1/DAY) (LIFE STYLE)
C0558929|T053|160609009|SNOMEDCT_US|EX-MODERATE SMOKER (10-19/DAY)|EX-MODERATE SMOKER (10-19/DAY) (LIFE STYLE)
C0558929|T053|160609009|SNOMEDCT_US|EX-MODERATE SMOKER (10-19/DAY) |EX-MODERATE SMOKER (10-19/DAY) (LIFE STYLE)
C0558929|T053|160609009|SNOMEDCT_US|EX-MODERATE SMOKER (10-19/DAY) |EX-MODERATE SMOKER (10-19/DAY) (LIFE STYLE)
C0558930|T053|160610004|SNOMEDCT_US|EX-HEAVY SMOKER (20-39/DAY)|EX-HEAVY SMOKER (20-39/DAY) (LIFE STYLE)
C0558930|T053|160610004|SNOMEDCT_US|EX-HEAVY SMOKER (20-39/DAY) |EX-HEAVY SMOKER (20-39/DAY) (LIFE STYLE)
C0558930|T053|160610004|SNOMEDCT_US|EX-HEAVY SMOKER (20-39/DAY) |EX-HEAVY SMOKER (20-39/DAY) (LIFE STYLE)
C0558931|T053|160611000|SNOMEDCT_US|EX-VERY HEAVY SMOKER (40+/DAY) |EX-VERY HEAVY SMOKER (40+/DAY) (LIFE STYLE)
C0558931|T053|160611000|SNOMEDCT_US|EX-VERY HEAVY SMOKER (40+/DAY)|EX-VERY HEAVY SMOKER (40+/DAY) (LIFE STYLE)
C0558931|T053|160611000|SNOMEDCT_US|EX-VERY HEAVY SMOKER (40+/DAY) |EX-VERY HEAVY SMOKER (40+/DAY) (LIFE STYLE)
C0558932|T053|160615009|SNOMEDCT_US|EX-SMOKER - AMOUNT UNKNOWN|EX-SMOKER - AMOUNT UNKNOWN (LIFE STYLE)
C0558932|T053|160615009|SNOMEDCT_US|EX-SMOKER - AMOUNT UNKNOWN |EX-SMOKER - AMOUNT UNKNOWN (LIFE STYLE)
C0558932|T053|160615009|SNOMEDCT_US|EX-SMOKER - AMOUNT UNKNOWN |EX-SMOKER - AMOUNT UNKNOWN (LIFE STYLE)
C3469008|T053||SNOMEDCT_US|NEVER A SMOKER - TOLERANT
C3469008|T053||SNOMEDCT_US|NEVER A SMOKER - TOLERANT 
C3469007|T053||SNOMEDCT_US|NEVER A SMOKER - INTOLERANT
C3469007|T053||SNOMEDCT_US|NEVER A SMOKER - INTOLERANT 
C3469006|T053||SNOMEDCT_US|NEVER A SMOKER - AGGRESSIVE 
C3469006|T053||SNOMEDCT_US|NEVER A SMOKER - AGGRESSIVE
C3472670|T053|221000119102|SNOMEDCT_US|NEVER SMOKED ANY SUBSTANCE|NEVER SMOKED ANY SUBSTANCE (FINDING)
C3472670|T053|221000119102|SNOMEDCT_US|NEVER SMOKED ANY SUBSTANCE |NEVER SMOKED ANY SUBSTANCE (FINDING)
C0425293|T053|266919005|SNOMEDCT_US|NEVER SMOKED|NEVER SMOKED TOBACCO (LIFE STYLE)
C0425293|T053|266919005|SNOMEDCT_US|NEVER SMOKER|NEVER SMOKED TOBACCO (LIFE STYLE)
C0425293|T053|266919005|SNOMEDCT_US|NEVER SMOKED |NEVER SMOKED TOBACCO (LIFE STYLE)
C0425293|T053|266919005|SNOMEDCT_US|NON-SMOKER|NEVER SMOKED TOBACCO (LIFE STYLE)
C0425293|T053|266919005|SNOMEDCT_US|NEVER SMOKED TOBACCO|NEVER SMOKED TOBACCO (LIFE STYLE)
C0425293|T053|266919005|SNOMEDCT_US|NEVER SMOKED TOBACCO |NEVER SMOKED TOBACCO (LIFE STYLE)
C0425293|T053|266919005|SNOMEDCT_US|NEVER SMOKED TOBACCO |NEVER SMOKED TOBACCO (LIFE STYLE)
C3241966|T053||SNOMEDCT_US|CURRENT SMOKER
C3241966|T053||SNOMEDCT_US|CURRENT SMOKER 
C0337664|T053|77176002|SNOMEDCT_US|SMOKER|SMOKER (LIFE STYLE)
C0337664|T053|77176002|SNOMEDCT_US|SMOKER, NOS|SMOKER (LIFE STYLE)
C0337664|T053|77176002|SNOMEDCT_US|SMOKER |SMOKER (LIFE STYLE)
C0337664|T053|77176002|SNOMEDCT_US|SMOKER |SMOKER (LIFE STYLE)
C3494625|T053|428071000124103|SNOMEDCT_US|CURRENT HEAVY TOBACCO SMOKER|HEAVY TOBACCO SMOKER (FINDING)
C3494625|T053|428071000124103|SNOMEDCT_US|HEAVY TOBACCO SMOKER |HEAVY TOBACCO SMOKER (FINDING)
C3494625|T053|428071000124103|SNOMEDCT_US|HEAVY TOBACCO SMOKER|HEAVY TOBACCO SMOKER (FINDING)
C3494625|T053|428071000124103|SNOMEDCT_US|CURRENT HEAVY TOBACCO SMOKER |HEAVY TOBACCO SMOKER (FINDING)
C1883049|T053||SNOMEDCT_US|SMOKER, CURRENT STATUS UNKNOWN
C1883049|T053||SNOMEDCT_US|SMOKER, CURRENT STATUS UNKNOWN 
C3694955|T053||SNOMEDCT_US|CURRENT SMOKER DURATION (___ YEARS) 
C3694955|T053||SNOMEDCT_US|CURRENT SMOKER DURATION (___ YEARS)
C0459847|T053|230063004|SNOMEDCT_US|HEAVY CIGARETTE SMOKER|HEAVY CIGARETTE SMOKER (LIFE STYLE)
C0459847|T053|230063004|SNOMEDCT_US|HEAVY CIGARETTE SMOKER |HEAVY CIGARETTE SMOKER (LIFE STYLE)
C0459847|T053|230063004|SNOMEDCT_US|HEAVY CIGARETTE SMOKER |HEAVY CIGARETTE SMOKER (LIFE STYLE)
C0337666|T053|59978006|SNOMEDCT_US|CIGAR SMOKER|CIGAR SMOKER (LIFE STYLE)
C0337666|T053|59978006|SNOMEDCT_US|SMOKING, CIGAR|CIGAR SMOKER (LIFE STYLE)
C0337666|T053|59978006|SNOMEDCT_US|CIGAR SMOKING|CIGAR SMOKER (LIFE STYLE)
C0337666|T053|59978006|SNOMEDCT_US|CIGAR SMOKER |CIGAR SMOKER (LIFE STYLE)
C0337666|T053|59978006|SNOMEDCT_US|CIGAR SMOKER |CIGAR SMOKER (LIFE STYLE)
C0337667|T053|65568007|SNOMEDCT_US|SMOKING CIGARETTES|CIGARETTE SMOKER (LIFE STYLE)
C0337667|T053|65568007|SNOMEDCT_US|CIGARETTE SMOKER|CIGARETTE SMOKER (LIFE STYLE)
C0337667|T053|65568007|SNOMEDCT_US|SMOKING CIGARETTES |CIGARETTE SMOKER (LIFE STYLE)
C0337667|T053|65568007|SNOMEDCT_US|SMOKES CIGARETTES|CIGARETTE SMOKER (LIFE STYLE)
C0337667|T053|65568007|SNOMEDCT_US|CIGARETTE SMOKER |CIGARETTE SMOKER (LIFE STYLE)
C0337667|T053|65568007|SNOMEDCT_US|CIGARETTE SMOKER, NOS|CIGARETTE SMOKER (LIFE STYLE)
C0337667|T053|65568007|SNOMEDCT_US|CIGARETTE SMOKER |CIGARETTE SMOKER (LIFE STYLE)
C0337669|T053|56771006|SNOMEDCT_US|HEAVY SMOKER (OVER 20 PER DAY)|HEAVY SMOKER (OVER 20 PER DAY) (LIFE STYLE)
C0337669|T053|56771006|SNOMEDCT_US|HEAVY SMOKER (OVER 20 PER DAY) |HEAVY SMOKER (OVER 20 PER DAY) (LIFE STYLE)
C0337669|T053|56771006|SNOMEDCT_US|HEAVY SMOKER (OVER 20 PER DAY) |HEAVY SMOKER (OVER 20 PER DAY) (LIFE STYLE)
C0337668|T053|56578002|SNOMEDCT_US|CURRENT MODERATE TOBACCO SMOKER |MODERATE SMOKER (20 OR LESS PER DAY) (LIFE STYLE)
C0337668|T053|56578002|SNOMEDCT_US|CURRENT MODERATE TOBACCO SMOKER|MODERATE SMOKER (20 OR LESS PER DAY) (LIFE STYLE)
C0337668|T053|56578002|SNOMEDCT_US|MODERATE SMOKER (20 OR LESS PER DAY)|MODERATE SMOKER (20 OR LESS PER DAY) (LIFE STYLE)
C0337668|T053|56578002|SNOMEDCT_US|MODERATE SMOKER (20 OR LESS PER DAY) |MODERATE SMOKER (20 OR LESS PER DAY) (LIFE STYLE)
C0337668|T053|56578002|SNOMEDCT_US|MODERATE SMOKER (20 OR LESS PER DAY) |MODERATE SMOKER (20 OR LESS PER DAY) (LIFE STYLE)
C0337665|T053|82302008|SNOMEDCT_US|PIPE SMOKER|PIPE SMOKER (LIFE STYLE)
C0337665|T053|82302008|SNOMEDCT_US|PIPE SMOKER |PIPE SMOKER (LIFE STYLE)
C0337665|T053|82302008|SNOMEDCT_US|PIPE SMOKER |PIPE SMOKER (LIFE STYLE)
C0425315|T053|266929003|SNOMEDCT_US|SMOKING STARTED - FINDING|SMOKING STARTED (LIFE STYLE)
C0425315|T053|266929003|SNOMEDCT_US|SMOKING STARTED|SMOKING STARTED (LIFE STYLE)
C0425315|T053|266929003|SNOMEDCT_US|SMOKING STARTED |SMOKING STARTED (LIFE STYLE)
C0425315|T053|266929003|SNOMEDCT_US|SMOKING STARTED |SMOKING STARTED (LIFE STYLE)
C3266136|T053|449868002|SNOMEDCT_US|DAILY SMOKER|CURRENT EVERY DAY SMOKER
C3266136|T053|449868002|SNOMEDCT_US|CURRENT EVERY DAY SMOKER|CURRENT EVERY DAY SMOKER
C3266136|T053|449868002|SNOMEDCT_US|EVERY DAY SMOKER|CURRENT EVERY DAY SMOKER
C3266136|T053|449868002|SNOMEDCT_US|CURRENT EVERY DAY SMOKER |CURRENT EVERY DAY SMOKER
C3266136|T053|449868002|SNOMEDCT_US|SMOKES TOBACCO DAILY|CURRENT EVERY DAY SMOKER
C3266136|T053|449868002|SNOMEDCT_US|SMOKES TOBACCO DAILY |CURRENT EVERY DAY SMOKER
C3266136|T053|449868002|SNOMEDCT_US|DAILY TOBACCO SMOKER|CURRENT EVERY DAY SMOKER
C3266136|T053|449868002|SNOMEDCT_US|EVERY-DAY SMOKER|CURRENT EVERY DAY SMOKER
C1883465|T053||SNOMEDCT_US|UNKNOWN IF EVER SMOKED
C1883465|T053||SNOMEDCT_US|UNKNOWN IF EVER SMOKED 
