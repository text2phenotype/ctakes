C0421451|T079|152322001|SNOMEDCT_US|PATIENT DATE OF BIRTH|DATE OF BIRTH (FINDING)
C2967445|T079||SNOMEDCT_US|BIRTH DATE PATIENT
C2348576|T079||SNOMEDCT_US|SUBJECT BIRTH DATE
C2919018|T079||SNOMEDCT_US|BIRTH DATE AND TIME
C2348576|T079||SNOMEDCT_US|SUBJECT BIRTH DATE
C2986369|T079||SNOMEDCT_US|BIOLOGIC ENTITY BIRTH DATE
C2986369|T079||SNOMEDCT_US|BIOLOGICENTITY.BIRTHDATE
C0421451|T079|152322001|SNOMEDCT_US|PATIENT DATE OF BIRTH|DATE OF BIRTH (FINDING)
C0421451|T079|152322001|SNOMEDCT_US|DOB|DATE OF BIRTH (FINDING)
C0421451|T079|152322001|SNOMEDCT_US|DATE OF BIRTH|DATE OF BIRTH (FINDING)
C0421451|T079|152322001|SNOMEDCT_US|BIRTH DATE|DATE OF BIRTH (FINDING)
C0421451|T079|152322001|SNOMEDCT_US|DATE OF BIRTH |DATE OF BIRTH (FINDING)
C0421451|T079|152322001|SNOMEDCT_US|BRTHDAT|DATE OF BIRTH (FINDING)
C0421451|T079|152322001|SNOMEDCT_US|BIRTHDATE|DATE OF BIRTH (FINDING)
C0421451|T079|152322001|SNOMEDCT_US|DOB - DATE OF BIRTH|DATE OF BIRTH (FINDING)
C0421451|T079|152322001|SNOMEDCT_US|DATE OF BIRTH (OBSERVABLE ENTITY)|DATE OF BIRTH (FINDING)
C0421451|T079|152322001|SNOMEDCT_US|DATE OF BIRTH OF PERSON CARED FOR|DATE OF BIRTH (FINDING)
C0421451|T079|152322001|SNOMEDCT_US|DATE OF BIRTH OF RECIPIENT OF CARE (OBSERVABLE ENTITY)|DATE OF BIRTH (FINDING)
C0421451|T079|152322001|SNOMEDCT_US|DATE OF BIRTH OF RECIPIENT OF CARE|DATE OF BIRTH (FINDING)
C2967445|T079||SNOMEDCT_US|BIRTH DATE &#X7C; PATIENT
C0803906|T079||SNOMEDCT_US|BIRTH DATE:TIME STAMP -- DATE AND TIME:POINT IN TIME:^PATIENT:QUANTITATIVE
C0803906|T079||SNOMEDCT_US|BIRTH DATE
C0803906|T079||SNOMEDCT_US|BIRTH DATE:TMSTP:PT:^PATIENT:QN
