C2367785|T034||LNC|HEPATITIS C GENOTYPE TESTING DOCUMENTED
C1533728|T034||LNC|HEPATITIS C VIRUS GENOTYPE DETERMINATION
C1148363|T034|MTHU014928|LNC|HEPATITIS C VIRUS GENOTYPE |HEPATITIS C VIRUS GENOTYPE
C4272868|T034||LNC|HEPATITIS C VIRAL GENOTYPE
C3532919|T034|MTHU054600|LNC|HEPATITIS C VIRUS GENOTYPE 1|HEPATITIS C VIRUS GENOTYPE 1
C3532920|T034||LNC|HEPATITIS C VIRUS GENOTYPE 2
C3532921|T034|MTHU054601|LNC|HEPATITIS C VIRUS GENOTYPE 3|HEPATITIS C VIRUS GENOTYPE 3
C3532922|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4
C3532923|T034||LNC|HEPATITIS C VIRUS GENOTYPE 5
C3532924|T034||LNC|HEPATITIS C VIRUS GENOTYPE 6
C3532919|T034|MTHU054600|LNC|HCV GENOTYPE 1|HEPATITIS C VIRUS GENOTYPE 1
C3532920|T034||LNC|HCV GENOTYPE 2
C3532921|T034|MTHU054601|LNC|HCV GENOTYPE 3|HEPATITIS C VIRUS GENOTYPE 3
C3532922|T034||LNC|HCV GENOTYPE 4
C3532923|T034||LNC|HCV GENOTYPE 5
C3532924|T034||LNC|HCV GENOTYPE 6
C3805156|T034||LNC|CHRONIC HEPATITIS C VIRUS GENOTYPE 1
C4049392|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 1
C4049393|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 1A
C4049394|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 1B
C4049395|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 2
C4049396|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 2A
C4049397|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 2B
C4049416|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4I
C4049417|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4J
C4049418|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 5
C4049419|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 5A
C4049420|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 6
C4049421|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 6A
C4049422|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4C
C4049423|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4D
C4049424|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4E
C4049425|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4F
C4049426|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4G
C4049427|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4H
C4049428|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 3D
C4049429|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 3E
C4049430|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 3F
C4049431|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4
C4049432|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4A
C4049433|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 2C
C4049434|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 2D
C4049435|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 3
C4049436|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 3A
C4049437|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 3B
C4049438|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 3C
C4049588|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4B
C3805156|T034||LNC|CHRONIC HCV GENOTYPE 1
C4049392|T034||LNC|CHRONIC HCV GENOTYPE 1
C4049393|T034||LNC|CHRONIC HCV GENOTYPE 1A
C4049394|T034||LNC|CHRONIC HCV GENOTYPE 1B
C4049395|T034||LNC|CHRONIC HCV GENOTYPE 2
C4049396|T034||LNC|CHRONIC HCV GENOTYPE 2A
C4049397|T034||LNC|CHRONIC HCV GENOTYPE 2B
C4049416|T034||LNC|CHRONIC HCV GENOTYPE 4I
C4049417|T034||LNC|CHRONIC HCV GENOTYPE 4J
C4049418|T034||LNC|CHRONIC HCV GENOTYPE 5
C4049419|T034||LNC|CHRONIC HCV GENOTYPE 5A
C4049420|T034||LNC|CHRONIC HCV GENOTYPE 6
C4049421|T034||LNC|CHRONIC HCV GENOTYPE 6A
C4049422|T034||LNC|CHRONIC HCV GENOTYPE 4C
C4049423|T034||LNC|CHRONIC HCV GENOTYPE 4D
C4049424|T034||LNC|CHRONIC HCV GENOTYPE 4E
C4049425|T034||LNC|CHRONIC HCV GENOTYPE 4F
C4049426|T034||LNC|CHRONIC HCV GENOTYPE 4G
C4049427|T034||LNC|CHRONIC HCV GENOTYPE 4H
C4049428|T034||LNC|CHRONIC HCV GENOTYPE 3D
C4049429|T034||LNC|CHRONIC HCV GENOTYPE 3E
C4049430|T034||LNC|CHRONIC HCV GENOTYPE 3F
C4049431|T034||LNC|CHRONIC HCV GENOTYPE 4
C4049432|T034||LNC|CHRONIC HCV GENOTYPE 4A
C4049433|T034||LNC|CHRONIC HCV GENOTYPE 2C
C4049434|T034||LNC|CHRONIC HCV GENOTYPE 2D
C4049435|T034||LNC|CHRONIC HCV GENOTYPE 3
C4049436|T034||LNC|CHRONIC HCV GENOTYPE 3A
C4049437|T034||LNC|CHRONIC HCV GENOTYPE 3B
C4049438|T034||LNC|CHRONIC HCV GENOTYPE 3C
C4049588|T034||LNC|CHRONIC HCV GENOTYPE 4B
C4272862|T034||LNC|HEPATITIS C VIRAL GENOTYPE 6
C4272863|T034||LNC|HEPATITIS C VIRAL GENOTYPE 5
C4272864|T034||LNC|HEPATITIS C VIRAL GENOTYPE 4
C4272865|T034||LNC|HEPATITIS C VIRAL GENOTYPE 3
C4272866|T034||LNC|HEPATITIS C VIRAL GENOTYPE 2
C4272867|T034||LNC|HEPATITIS C VIRAL GENOTYPE 1
C4272862|T034||LNC|HCV VIRAL GENOTYPE 6
C4272863|T034||LNC|HCV VIRAL GENOTYPE 5
C4272864|T034||LNC|HCV VIRAL GENOTYPE 4
C4272865|T034||LNC|HCV VIRAL GENOTYPE 3
C4272866|T034||LNC|HCV VIRAL GENOTYPE 2
C4272867|T034||LNC|HCV VIRAL GENOTYPE 1
C4284773|T034|MTHU054613|LNC|HEPATITIS C VIRUS GENOTYPE PANEL|HEPATITIS C VIRUS GENOTYPE PANEL
C4284909|T034|82525-7|LNC|HEPATITIS C VIRUS GENOTYPE PANEL|HEPATITIS C VIRUS GENOTYPE PANEL:-:POINT IN TIME:ISOLATE+SERUM:-
C0973340|T034||LNC|INFECTIOUS AGENT GENOTYPE ANALYSIS BY NUCLEIC ACID (DNA OR RNA); HEPATITIS C VIRUS
C2030676|T034||LNC|HEPATITIS C VIRUS GENOTYPE ANALYSIS BY NUCLEIC ACID
C4064267|T034||LNC|PROBE AND TARGET AMPLIFICATION FOR HEPATITIS C VIRUS GENOTYPE
C4284773|T034|MTHU054613|LNC|HCV GENOTYPE PANEL|HEPATITIS C VIRUS GENOTYPE PANEL
C4284909|T034|82525-7|LNC|HCV GENOTYPE PANEL|HEPATITIS C VIRUS GENOTYPE PANEL:-:POINT IN TIME:ISOLATE+SERUM:-
C0973340|T034||LNC|INFECTIOUS AGENT HCV GENOTYPE ANALYSIS
C1971440|T034||LNC|HCV GENOTYPE TESTING
C2030676|T034||LNC|HCV GENOTYPE ANALYSIS BY NUCLEIC ACID
C4064267|T034||LNC|HCV PROBE AND TARGET AMPLIFICATION
C1742607|T034||LNC|HCV MOLECULAR ASSAY
C3495939|T034||LNC|HEPATITIS C VIRUS GENOTYPE 1A POSITIVE
C3495940|T034||LNC|HEPATITIS C VIRUS GENOTYPE 1B POSITIVE
C3495941|T034||LNC|HEPATITIS C VIRUS GENOTYPE 3A POSITIVE
C3495942|T034||LNC|HEPATITIS C VIRUS GENOTYPE 3B POSITIVE
C3495943|T034||LNC|HEPATITIS C VIRUS GENOTYPE 1 POSITIVE
C3495944|T034||LNC|HEPATITIS C VIRUS GENOTYPE 3 POSITIVE
C3495939|T034||LNC|HCV GENOTYPE 1A POSITIVE
C3495940|T034||LNC|HCV GENOTYPE 1B POSITIVE
C3495941|T034||LNC|HCV GENOTYPE 3A POSITIVE
C3495942|T034||LNC|HCV GENOTYPE 3B POSITIVE
C3495943|T034||LNC|HCV GENOTYPE 1 POSITIVE
C3495944|T034||LNC|HCV GENOTYPE 3 POSITIVE
C3854557|T034||LNC|HEPATITIS C VIRUS GENOTYPE 2B POSITIVE
C3854558|T034||LNC|HEPATITIS C VIRUS GENOTYPE 2 POSITIVE
C3889043|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4 POSITIVE
C3889044|T034||LNC|HEPATITIS C VIRUS GENOTYPE 5 POSITIVE
C3889045|T034||LNC|HEPATITIS C VIRUS GENOTYPE 6 POSITIVE
C4049398|T034||LNC|HEPATITIS C VIRUS GENOTYPE 6A POSITIVE
C4049399|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4F POSITIVE
C4049400|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4G POSITIVE
C4049401|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4H POSITIVE
C4049402|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4I POSITIVE
C4049403|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4J POSITIVE
C4049404|T034||LNC|HEPATITIS C VIRUS GENOTYPE 5A POSITIVE
C4049405|T034||LNC|HEPATITIS C VIRUS GENOTYPE 3F POSITIVE
C4049406|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4A POSITIVE
C4049407|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4B POSITIVE
C4049408|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4C POSITIVE
C4049409|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4D POSITIVE
C4049410|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4E POSITIVE
C4049411|T034||LNC|HEPATITIS C VIRUS GENOTYPE 2A POSITIVE
C4049412|T034||LNC|HEPATITIS C VIRUS GENOTYPE 2C POSITIVE
C4049413|T034||LNC|HEPATITIS C VIRUS GENOTYPE 2D POSITIVE
C4049414|T034||LNC|HEPATITIS C VIRUS GENOTYPE 3C POSITIVE
C4049415|T034||LNC|HEPATITIS C VIRUS GENOTYPE 3E POSITIVE
C4049587|T034||LNC|HEPATITIS C VIRUS GENOTYPE 3D POSITIVE
C1954138|T034|48574-8|LNC|HEPATITIS C VIRUS GENOTYPE|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:WHOLE BLOOD:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR
C1977372|T034|49607-5|LNC|HEPATITIS C VIRUS GENOTYPE|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:TISSUE, UNSPECIFIED:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR
C4298651|T034|82513-3|LNC|HEPATITIS C VIRUS GENOTYPE 3|HCV GENTYP 3 SERPL QL NAA+PROBE
C4298652|T034|82512-5|LNC|HEPATITIS C VIRUS GENOTYPE 1|HEPATITIS C VIRUS GENOTYPE 1 [TYPE] IN SERUM OR PLASMA BY NAA WITH PROBE DETECTION
C4064283|T034||LNC|PROBE WITH TARGET AMPLIFICATION FOR HEPATITIS C VIRUS GENOTYPE IN SERUM OR PLASMA
C1147970|T034|32286-7|LNC|HEPATITIS C VIRUS GENOTYPE|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:SERUM/PLASMA:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR
C1954139|T034|48575-5|LNC|HEPATITIS C VIRUS GENOTYPE|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:TO BE SPECIFIED IN ANOTHER PART OF THE MESSAGE:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR
C4300371|T034|LP220401-6|LNC|HEPATITIS C VIRUS GENOTYPE 3 NS5A GENE|HEPATITIS C VIRUS GENOTYPE 3 NS5A GENE
C4300372|T034|LP220303-4|LNC|HEPATITIS C VIRUS GENOTYPE 1 NS5B GENE|HEPATITIS C VIRUS GENOTYPE 1 NS5B GENE
C4300373|T034|LP220405-7|LNC|HEPATITIS C VIRUS GENOTYPE 1 NS5A GENE|HEPATITIS C VIRUS GENOTYPE 1 NS5A GENE
C3654330|T034|73655-3|LNC|HEPATITIS C VIRUS NS5 GENE MUTATIONS DETECTED|HEPATITIS C VIRUS NS5 GENE MUTATIONS DETECTED:PRESENCE OR IDENTITY:POINT IN TIME:ISOLATE:NOMINAL:GENOTYPING
C3654331|T034|73654-6|LNC|HEPATITIS C VIRUS NS3 GENE MUTATIONS DETECTED|HCV NS3 MUT DET ISLT GENOTYP
C4285206|T034|82381-5|LNC|HEPATITIS C VIRUS GENOTYPE 1 NS5B GENE MUTATIONS DETECTED|HEPATITIS C VIRUS GENOTYPE 1 NS5B GENE MUTATIONS DETECTED:PRESENCE OR IDENTITY:POINT IN TIME:ISOLATE:NOMINAL:GENOTYPING
C4285533|T034|82514-1|LNC|HEPATITIS C VIRUS GENOTYPE 3 NS5A GENE MUTATIONS DETECTED|HEPATITIS C VIRUS GENOTYPE 3 NS5A GENE MUTATIONS DETECTED:PRESENCE OR IDENTITY:POINT IN TIME:ISOLATE:NOMINAL:GENOTYPING
C4296735|T034|MTHU054602|LNC|HEPATITIS C VIRUS GENOTYPE 3 NS5A GENE MUTATIONS DETECTED|HEPATITIS C VIRUS GENOTYPE 3 NS5A GENE MUTATIONS DETECTED
C4296782|T034|MTHU054535|LNC|HEPATITIS C VIRUS GENOTYPE 1 NS5B GENE MUTATIONS DETECTED|HEPATITIS C VIRUS GENOTYPE 1 NS5B GENE MUTATIONS DETECTED
C4296783|T034|MTHU054534|LNC|HEPATITIS C VIRUS GENOTYPE 1 NS5A GENE MUTATIONS DETECTED|HEPATITIS C VIRUS GENOTYPE 1 NS5A GENE MUTATIONS DETECTED
C4298748|T034|82380-7|LNC|HEPATITIS C VIRUS GENOTYPE 1 NS5A GENE MUTATIONS DETECTED|HCV GENTYP 1 NS5A MUT DET ISLT
C1269856|T034||LNC|PCR POSITIVE FOR HCV VIRAL RNA (GENOTYPE 1A)
C1148363|T034|MTHU014928|LNC|HEPATITIS C VIRUS GENOTYPE |HEPATITIS C VIRUS GENOTYPE
C1148363|T034|MTHU014928|LNC|HEPATITIS C VIRUS GENOTYPE|HEPATITIS C VIRUS GENOTYPE
C1533728|T034||LNC|HEPATITIS C VIRUS GENOTYPE
C1533728|T034||LNC|HEPATITIS C VIRUS GENOTYPE 
C1533728|T034||LNC|HCV GENOTYPING
C1533728|T034||LNC|HEPATITIS C VIRUS GENOTYPE ASSAY
C1533728|T034||LNC|HCV GENOTYPE ASSAY
C1533728|T034||LNC|HCV GENOTYPE MEASUREMENT
C1533728|T034||LNC|HCV GENOTYPE
C1533728|T034||LNC|HEPATITIS C VIRUS GENOTYPE DETERMINATION 
C1533728|T034||LNC|HEPATITIS C VIRUS GENOTYPE DETERMINATION
C4064267|T034||LNC|PROBE WITH TARGET AMPLIFICATION HEPATITIS C VIRUS GENOTYPE
C4064267|T034||LNC|PROBE WITH TARGET AMPLIFICATION HEPATITIS C VIRUS GENOTYPE 
C4064283|T034||LNC|PROBE WITH TARGET AMPLIFICATION FOR HEPATITIS C VIRUS GENOTYPE IN SERUM OR PLASMA 
C4064283|T034||LNC|PROBE WITH TARGET AMPLIFICATION FOR HEPATITIS C VIRUS GENOTYPE IN SERUM OR PLASMA
C4064283|T034||LNC|PROBE & TARGET AMPLIF HEPATITIS C VIRUS GENOTYPE SERUM / PLASMA
C3494966|T034||LNC|HEPATITIS C VIRUS SUBTYPE 1A 
C3494966|T034||LNC|HEPATITIS C VIRUS SUBTYPE 1A
C3494965|T034||LNC|HEPATITIS C VIRUS SUBTYPE 1B 
C3494965|T034||LNC|HEPATITIS C VIRUS SUBTYPE 1B
C3532925|T034||LNC|HEPATITIS C VIRUS SUBTYPE 1C
C3532925|T034||LNC|HEPATITIS C VIRUS SUBTYPE 1C 
C3494964|T034||LNC|HEPATITIS C VIRUS SUBTYPE 2A
C3494964|T034||LNC|HEPATITIS C VIRUS SUBTYPE 2A 
C3494963|T034||LNC|HEPATITIS C VIRUS SUBTYPE 2B 
C3494963|T034||LNC|HEPATITIS C VIRUS SUBTYPE 2B
C3532926|T034||LNC|HEPATITIS C VIRUS SUBTYPE 2C
C3532926|T034||LNC|HEPATITIS C VIRUS SUBTYPE 2C 
C3494962|T034||LNC|HEPATITIS C VIRUS SUBTYPE 3A
C3494962|T034||LNC|HEPATITIS C VIRUS SUBTYPE 3A 
C3494961|T034||LNC|HEPATITIS C VIRUS SUBTYPE 3B 
C3494961|T034||LNC|HEPATITIS C VIRUS SUBTYPE 3B
C3532918|T034||LNC|HEPATITIS C VIRUS SUBTYPE 4A
C3532918|T034||LNC|HEPATITIS C VIRUS SUBTYPE 4A 
C3532927|T034||LNC|HEPATITIS C VIRUS SUBTYPE 4B
C3532927|T034||LNC|HEPATITIS C VIRUS SUBTYPE 4B 
C3532928|T034||LNC|HEPATITIS C VIRUS SUBTYPE 4C
C3532928|T034||LNC|HEPATITIS C VIRUS SUBTYPE 4C 
C3532929|T034||LNC|HEPATITIS C VIRUS SUBTYPE 4D 
C3532929|T034||LNC|HEPATITIS C VIRUS SUBTYPE 4D
C3494960|T034||LNC|HEPATITIS C VIRUS SUBTYPE 4E 
C3494960|T034||LNC|HEPATITIS C VIRUS SUBTYPE 4E
C3494959|T034||LNC|HEPATITIS C VIRUS SUBTYPE 5A 
C3494959|T034||LNC|HEPATITIS C VIRUS SUBTYPE 5A
C3494958|T034||LNC|HEPATITIS C VIRUS SUBTYPE 6A 
C3494958|T034||LNC|HEPATITIS C VIRUS SUBTYPE 6A
C3805156|T034||LNC|CHRONIC HEPATITIS C VIRUS GENOTYPE 1
C4049392|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 1
C4049393|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 1A
C4049394|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 1B
C4049395|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 2
C4049396|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 2A
C4049397|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 2B
C4049416|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4I
C4049417|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4J
C4049418|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 5
C4049419|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 5A
C4049420|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 6
C4049421|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 6A
C4049422|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4C
C4049423|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4D
C4049424|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4E
C4049425|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4F
C4049426|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4G
C4049427|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4H
C4049428|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 3D
C4049429|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 3E
C4049430|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 3F
C4049431|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4
C4049432|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4A
C4049433|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 2C
C4049434|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 2D
C4049435|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 3
C4049436|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 3A
C4049437|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 3B
C4049438|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 3C
C4049588|T034||LNC|CHRONIC HEPATITIS C GENOTYPE 4B
C0973340|T034||LNC|NFCT AGNT GENOTYP NUCLEIC ACID HEPATITIS C VIRUS
C0973340|T034||LNC|INFECTIOUS AGENT GENOTYPE ANALYSIS BY NUCLEIC ACID (DNA OR RNA); HEPATITIS C VIRUS
C0973340|T034||LNC|GENOTYPE DNA/RNA HEP C
C0973340|T034||LNC|ANALYSIS OF INFECTIOUS AGENT GENOTYPE OF HEPATITIS C VIRUS
C1971440|T034||LNC|HEPC GN TSTNG DOCD B/4TXMNT
C1971440|T034||LNC|HEPATITIS C GENOTYPE PRIOR ANTIVIRAL TREATMENT
C3495939|T034||LNC|HEPATITIS C VIRUS GENOTYPE 1A POSITIVE
C3495940|T034||LNC|HEPATITIS C VIRUS GENOTYPE 1B POSITIVE
C3495941|T034||LNC|HEPATITIS C VIRUS GENOTYPE 3A POSITIVE
C3495942|T034||LNC|HEPATITIS C VIRUS GENOTYPE 3B POSITIVE
C3495943|T034||LNC|HEPATITIS C VIRUS GENOTYPE 1 POSITIVE
C3495944|T034||LNC|HEPATITIS C VIRUS GENOTYPE 3 POSITIVE
C4049415|T034||LNC|HEPATITIS C VIRUS GENOTYPE 3E POSITIVE
C3854557|T034||LNC|HEPATITIS C VIRUS GENOTYPE 2B POSITIVE
C3854558|T034||LNC|HEPATITIS C VIRUS GENOTYPE 2 POSITIVE
C3889043|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4 POSITIVE
C3889044|T034||LNC|HEPATITIS C VIRUS GENOTYPE 5 POSITIVE
C3889045|T034||LNC|HEPATITIS C VIRUS GENOTYPE 6 POSITIVE
C4049398|T034||LNC|HEPATITIS C VIRUS GENOTYPE 6A POSITIVE
C4049399|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4F POSITIVE
C4049400|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4G POSITIVE
C4049401|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4H POSITIVE
C4049402|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4I POSITIVE
C4049403|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4J POSITIVE
C4049404|T034||LNC|HEPATITIS C VIRUS GENOTYPE 5A POSITIVE
C4049405|T034||LNC|HEPATITIS C VIRUS GENOTYPE 3F POSITIVE
C4049406|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4A POSITIVE
C4049407|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4B POSITIVE
C4049408|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4C POSITIVE
C4049409|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4D POSITIVE
C4049410|T034||LNC|HEPATITIS C VIRUS GENOTYPE 4E POSITIVE
C4049411|T034||LNC|HEPATITIS C VIRUS GENOTYPE 2A POSITIVE
C4049412|T034||LNC|HEPATITIS C VIRUS GENOTYPE 2C POSITIVE
C4049413|T034||LNC|HEPATITIS C VIRUS GENOTYPE 2D POSITIVE
C4049414|T034||LNC|HEPATITIS C VIRUS GENOTYPE 3C POSITIVE
C4049587|T034||LNC|HEPATITIS C VIRUS GENOTYPE 3D POSITIVE
C1954138|T034|48574-8|LNC|HEPATITIS C VIRUS GENOTYPE:PRID:PT:BLD:NOM:PROBE.AMP.TAR|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:WHOLE BLOOD:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR
C1954138|T034|48574-8|LNC|HCV GENTYP BLD PCR|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:WHOLE BLOOD:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR
C1954138|T034|48574-8|LNC|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:WHOLE BLOOD:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:WHOLE BLOOD:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR
C1954138|T034|48574-8|LNC|HEPATITIS C VIRUS GENOTYPE [IDENTIFIER] IN BLOOD BY PROBE AND TARGET AMPLIFICATION METHOD|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:WHOLE BLOOD:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR
C1977372|T034|49607-5|LNC|HEPATITIS C VIRUS GENOTYPE:PRID:PT:TISS:NOM:PROBE.AMP.TAR|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:TISSUE, UNSPECIFIED:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR
C1977372|T034|49607-5|LNC|HCV GENTYP TISS PCR|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:TISSUE, UNSPECIFIED:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR
C1977372|T034|49607-5|LNC|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:TISSUE, UNSPECIFIED:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:TISSUE, UNSPECIFIED:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR
C1977372|T034|49607-5|LNC|HEPATITIS C VIRUS GENOTYPE [IDENTIFIER] IN TISSUE BY PROBE AND TARGET AMPLIFICATION METHOD|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:TISSUE, UNSPECIFIED:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR
C1147970|T034|32286-7|LNC|HEPATITIS C VIRUS GENOTYPE:PRID:PT:SER/PLAS:NOM:PROBE.AMP.TAR|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:SERUM/PLASMA:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR
C1147970|T034|32286-7|LNC|HCV GENTYP SERPL PCR|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:SERUM/PLASMA:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR
C1147970|T034|32286-7|LNC|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:SERUM/PLASMA:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:SERUM/PLASMA:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR
C1147970|T034|32286-7|LNC|HEPATITIS C VIRUS GENOTYPE [IDENTIFIER] IN SERUM OR PLASMA BY PROBE AND TARGET AMPLIFICATION METHOD|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:SERUM/PLASMA:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR
C1954139|T034|48575-5|LNC|HEPATITIS C VIRUS GENOTYPE:PRID:PT:XXX:NOM:PROBE.AMP.TAR|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:TO BE SPECIFIED IN ANOTHER PART OF THE MESSAGE:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR
C1954139|T034|48575-5|LNC|HCV GENTYP XXX PCR|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:TO BE SPECIFIED IN ANOTHER PART OF THE MESSAGE:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR
C1954139|T034|48575-5|LNC|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:TO BE SPECIFIED IN ANOTHER PART OF THE MESSAGE:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:TO BE SPECIFIED IN ANOTHER PART OF THE MESSAGE:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR
C1954139|T034|48575-5|LNC|HEPATITIS C VIRUS GENOTYPE [IDENTIFIER] IN UNSPECIFIED SPECIMEN BY PROBE AND TARGET AMPLIFICATION METHOD|HEPATITIS C VIRUS GENOTYPE:PRESENCE OR IDENTITY:POINT IN TIME:TO BE SPECIFIED IN ANOTHER PART OF THE MESSAGE:NOMINAL:DNA NUCLEIC ACID PROBE.AMP.TAR
C3654330|T034|73655-3|LNC|HEPATITIS C VIRUS NS5 GENE MUTATIONS DETECTED:PRID:PT:ISOLATE:NOM:GENOTYPING|HEPATITIS C VIRUS NS5 GENE MUTATIONS DETECTED:PRESENCE OR IDENTITY:POINT IN TIME:ISOLATE:NOMINAL:GENOTYPING
C3654330|T034|73655-3|LNC|HEPATITIS C VIRUS NS5 GENE MUTATIONS DETECTED:PRESENCE OR IDENTITY:POINT IN TIME:ISOLATE:NOMINAL:GENOTYPING|HEPATITIS C VIRUS NS5 GENE MUTATIONS DETECTED:PRESENCE OR IDENTITY:POINT IN TIME:ISOLATE:NOMINAL:GENOTYPING
C3654330|T034|73655-3|LNC|HCV NS5 MUT DET ISLT GENOTYP|HEPATITIS C VIRUS NS5 GENE MUTATIONS DETECTED:PRESENCE OR IDENTITY:POINT IN TIME:ISOLATE:NOMINAL:GENOTYPING
C3654330|T034|73655-3|LNC|HEPATITIS C VIRUS NS5 GENE MUTATIONS DETECTED [IDENTIFIER] BY GENOTYPE METHOD|HEPATITIS C VIRUS NS5 GENE MUTATIONS DETECTED:PRESENCE OR IDENTITY:POINT IN TIME:ISOLATE:NOMINAL:GENOTYPING
C3654331|T034|73654-6|LNC|HCV NS3 MUT DET ISLT GENOTYP|HCV NS3 MUT DET ISLT GENOTYP
C3654331|T034|73654-6|LNC|HEPATITIS C VIRUS NS3 GENE MUTATIONS DETECTED:PRESENCE OR IDENTITY:POINT IN TIME:ISOLATE:NOMINAL:GENOTYPING|HCV NS3 MUT DET ISLT GENOTYP
C3654331|T034|73654-6|LNC|HEPATITIS C VIRUS NS3 GENE MUTATIONS DETECTED:PRID:PT:ISOLATE:NOM:GENOTYPING|HCV NS3 MUT DET ISLT GENOTYP
C3654331|T034|73654-6|LNC|HEPATITIS C VIRUS NS3 GENE MUTATIONS DETECTED [IDENTIFIER] BY GENOTYPE METHOD|HCV NS3 MUT DET ISLT GENOTYP
