C0000731|T033|SY|60728008|SNOMEDCT_CORE|Abdomen distended|Swollen abdomen
C0000731|T033|OAP|41931001|SNOMEDCT_CORE|Abdominal distension|Swollen abdomen
C0000731|T033|OAF|41931001|SNOMEDCT_CORE|Abdominal distension|Swollen abdomen
C0000731|T033|IS|41931001|SNOMEDCT_CORE|Abdominal distention|Swollen abdomen
C0000731|T033|SY|60728008|SNOMEDCT_CORE|Abdominal distention|Swollen abdomen
C0000731|T033|SY|60728008|SNOMEDCT_CORE|Abdominal swelling|Swollen abdomen
C0000731|T033|SY|60728008|SNOMEDCT_CORE|Swelling of abdomen|Swollen abdomen
C0000731|T033|PT|60728008|SNOMEDCT_CORE|Swollen abdomen|Swollen abdomen
C0000731|T033|FN|60728008|SNOMEDCT_CORE|Swollen abdomen|Swollen abdomen
C0000734|T033|SY|271860004|SNOMEDCT_CORE|Abdominal lump|Abdominal mass
C0000734|T033|PT|271860004|SNOMEDCT_CORE|Abdominal mass|Abdominal mass
C0000734|T033|FN|271860004|SNOMEDCT_CORE|Abdominal mass|Abdominal mass
C0000737|T184|PT|21522001|SNOMEDCT_CORE|Abdominal pain|Abdominal pain
C0000737|T184|FN|21522001|SNOMEDCT_CORE|Abdominal pain|Abdominal pain
C0000737|T184|SY|21522001|SNOMEDCT_CORE|AP - Abdominal pain|Abdominal pain
C0000768|T019|SY|276654001|SNOMEDCT_CORE|CM - Congenital malformation|Congenital malformation
C0000768|T019|SY|276654001|SNOMEDCT_CORE|Congenital abnormality|Congenital malformation
C0000768|T019|SY|276654001|SNOMEDCT_CORE|Congenital anomaly|Congenital malformation
C0000768|T019|PT|276654001|SNOMEDCT_CORE|Congenital malformation|Congenital malformation
C0000768|T019|FN|276654001|SNOMEDCT_CORE|Congenital malformation|Congenital malformation
C0000768|T019|SY|276654001|SNOMEDCT_CORE|Fetal developmental abnormality|Congenital malformation
C0000768|T019|SY|276654001|SNOMEDCT_CORE|Fetal malformation|Congenital malformation
C0000768|T019|SYGB|276654001|SNOMEDCT_CORE|Foetal developmental abnormality|Congenital malformation
C0000768|T019|SY|276654001|SNOMEDCT_CORE|Foetal malformation|Congenital malformation
C0000772|T019|IS|67024003|SNOMEDCT_CORE|Multiple anomalies, NOS|Multiple congenital anomalies
C0000772|T019|OP|444406006|SNOMEDCT_CORE|Multiple congenital anomalies|Multiple congenital anomalies
C0000772|T019|OAP|67024003|SNOMEDCT_CORE|Multiple congenital anomalies|Multiple congenital anomalies
C0000772|T019|OAF|67024003|SNOMEDCT_CORE|Multiple congenital anomalies|Multiple congenital anomalies
C0000772|T019|OAF|444406006|SNOMEDCT_CORE|Multiple congenital anomalies|Multiple congenital anomalies
C0000772|T019|IS|67024003|SNOMEDCT_CORE|Multiple congenital anomalies, NOS|Multiple congenital anomalies
C0000772|T019|OAP|444406006|SNOMEDCT_CORE|Multiple congenital malformations|Multiple congenital anomalies
C0000786|T046|PT|17369002|SNOMEDCT_CORE|Miscarriage|Miscarriage
C0000786|T046|FN|17369002|SNOMEDCT_CORE|Miscarriage|Miscarriage
C0000786|T046|IS|17369002|SNOMEDCT_CORE|Miscarriage, NOS|Miscarriage
C0000786|T046|SY|17369002|SNOMEDCT_CORE|Spontaneous abortion|Miscarriage
C0000786|T046|OF|17369002|SNOMEDCT_CORE|Spontaneous abortion|Miscarriage
C0000786|T046|IS|17369002|SNOMEDCT_CORE|Spontaneous abortion, NOS|Miscarriage
C0000786|T046|SY|17369002|SNOMEDCT_CORE|Vaginal expulsion of fetus|Miscarriage
C0000786|T046|SY|17369002|SNOMEDCT_CORE|Vaginal expulsion of foetus|Miscarriage
C0000786|T046|SY|17369002|SNOMEDCT_CORE|Vaginal expulsion of product of conception|Miscarriage
C0000790|T033|OAP|267014009|SNOMEDCT_CORE|H/O: abortion|History of pregnancy with abortive outcome
C0000790|T033|OAS|267014009|SNOMEDCT_CORE|H/O: termination|History of pregnancy with abortive outcome
C0000790|T033|IS|267014009|SNOMEDCT_CORE|History of - abortion|History of pregnancy with abortive outcome
C0000790|T033|OF|267014009|SNOMEDCT_CORE|History of - abortion|History of pregnancy with abortive outcome
C0000790|T033|IS|267014009|SNOMEDCT_CORE|History of - fetal loss|History of pregnancy with abortive outcome
C0000790|T033|IS|267014009|SNOMEDCT_CORE|History of - foetal loss|History of pregnancy with abortive outcome
C0000790|T033|OAS|267014009|SNOMEDCT_CORE|History of abortion|History of pregnancy with abortive outcome
C0000790|T033|OAF|267014009|SNOMEDCT_CORE|History of abortion|History of pregnancy with abortive outcome
C0000790|T033|IS|267014009|SNOMEDCT_CORE|History of fetal loss|History of pregnancy with abortive outcome
C0000790|T033|SY|713651007|SNOMEDCT_CORE|History of fetal loss|History of pregnancy with abortive outcome
C0000790|T033|IS|267014009|SNOMEDCT_CORE|History of foetal loss|History of pregnancy with abortive outcome
C0000790|T033|SYGB|713651007|SNOMEDCT_CORE|History of foetal loss|History of pregnancy with abortive outcome
C0000790|T033|PT|713651007|SNOMEDCT_CORE|History of pregnancy with abortive outcome|History of pregnancy with abortive outcome
C0000790|T033|FN|713651007|SNOMEDCT_CORE|History of pregnancy with abortive outcome|History of pregnancy with abortive outcome
C0000810|T046|OAP|16863000|SNOMEDCT_CORE|Incomplete miscarriage|Incomplete miscarriage
C0000810|T046|PT|156072005|SNOMEDCT_CORE|Incomplete miscarriage|Incomplete miscarriage
C0000810|T046|FN|156072005|SNOMEDCT_CORE|Incomplete miscarriage|Incomplete miscarriage
C0000810|T046|SY|156072005|SNOMEDCT_CORE|Incomplete spontaneous abortion|Incomplete miscarriage
C0000810|T046|OAS|16863000|SNOMEDCT_CORE|Incomplete spontaneous abortion|Incomplete miscarriage
C0000810|T046|PT|275425008|SNOMEDCT_CORE|Retained products after miscarriage|Incomplete miscarriage
C0000810|T046|FN|275425008|SNOMEDCT_CORE|Retained products after miscarriage|Incomplete miscarriage
C0000810|T046|SY|275425008|SNOMEDCT_CORE|Retained products after spontaneous abortion|Incomplete miscarriage
C0000810|T046|OF|275425008|SNOMEDCT_CORE|Retained products after spontaneous abortion|Incomplete miscarriage
C0000810|T046|SY|275425008|SNOMEDCT_CORE|Retained tissue after pregnancy loss|Incomplete miscarriage
C0000814|T047|SY|16607004|SNOMEDCT_CORE|Foetal death before 22 weeks with retention of dead foetus|Missed miscarriage
C0000814|T047|SY|16607004|SNOMEDCT_CORE|MA - Missed abortion|Missed miscarriage
C0000814|T047|SY|16607004|SNOMEDCT_CORE|Missed abortion|Missed miscarriage
C0000814|T047|FN|16607004|SNOMEDCT_CORE|Missed abortion|Missed miscarriage
C0000814|T047|PT|16607004|SNOMEDCT_CORE|Missed miscarriage|Missed miscarriage
C0000814|T047|SY|16607004|SNOMEDCT_CORE|Silent miscarriage|Missed miscarriage
C0000821|T046|SY|54048003|SNOMEDCT_CORE|Threatened abortion|Threatened miscarriage
C0000821|T046|FN|54048003|SNOMEDCT_CORE|Threatened abortion|Threatened miscarriage
C0000821|T046|IS|54048003|SNOMEDCT_CORE|Threatened abortion, NOS|Threatened miscarriage
C0000821|T046|PT|54048003|SNOMEDCT_CORE|Threatened miscarriage|Threatened miscarriage
C0000832|T046|SY|415105001|SNOMEDCT_CORE|Ablatio placentae|Placental abruption
C0000832|T046|SY|415105001|SNOMEDCT_CORE|Abruptio placentae|Placental abruption
C0000832|T046|PT|415105001|SNOMEDCT_CORE|Placental abruption|Placental abruption
C0000832|T046|FN|415105001|SNOMEDCT_CORE|Placental abruption|Placental abruption
C0000832|T046|SY|415105001|SNOMEDCT_CORE|Premature detachment of normally implanted placenta|Placental abruption
C0000832|T046|SY|415105001|SNOMEDCT_CORE|Premature detachment of placenta|Placental abruption
C0000832|T046|SY|415105001|SNOMEDCT_CORE|Premature separation of placenta|Placental abruption
C0000833|T047|PT|128477000|SNOMEDCT_CORE|Abscess|Abscess
C0000833|T047|FN|128477000|SNOMEDCT_CORE|Abscess|Abscess
C0000889|T047|PT|402599005|SNOMEDCT_CORE|Acanthosis nigricans|Acanthosis nigricans
C0000889|T047|FN|402599005|SNOMEDCT_CORE|Acanthosis nigricans|Acanthosis nigricans
C0000921|T037|PT|217082002|SNOMEDCT_CORE|Accidental fall|Accidental fall
C0000921|T037|OF|217082002|SNOMEDCT_CORE|Accidental fall|Accidental fall
C0000921|T037|FN|217082002|SNOMEDCT_CORE|Accidental fall|Accidental fall
C0000921|T037|SY|217082002|SNOMEDCT_CORE|Fall - accidental|Accidental fall
C0001122|T046|PT|51387008|SNOMEDCT_CORE|Acidosis|Acidosis
C0001122|T046|FN|51387008|SNOMEDCT_CORE|Acidosis|Acidosis
C0001122|T046|IS|51387008|SNOMEDCT_CORE|Acidosis, NOS|Acidosis
C0001125|T047|PT|91273001|SNOMEDCT_CORE|Lactic acidosis|Lactic acidosis
C0001125|T047|FN|91273001|SNOMEDCT_CORE|Lactic acidosis|Lactic acidosis
C0001126|T047|PT|1776003|SNOMEDCT_CORE|Renal tubular acidosis|Renal tubular acidosis
C0001126|T047|FN|1776003|SNOMEDCT_CORE|Renal tubular acidosis|Renal tubular acidosis
C0001126|T047|IS|1776003|SNOMEDCT_CORE|Renal tubular acidosis, NOS|Renal tubular acidosis
C0001126|T047|IS|1776003|SNOMEDCT_CORE|RTA|Renal tubular acidosis
C0001126|T047|SY|1776003|SNOMEDCT_CORE|RTA - Renal tubular acidosis|Renal tubular acidosis
C0001126|T047|IS|1776003|SNOMEDCT_CORE|RTA, NOS|Renal tubular acidosis
C0001144|T047|OAP|88616000|SNOMEDCT_CORE|Acne vulgaris|Common acne
C0001144|T047|OAF|88616000|SNOMEDCT_CORE|Acne vulgaris|Common acne
C0001144|T047|OAS|88616000|SNOMEDCT_CORE|Common acne|Common acne
C0001145|T047|PT|238746008|SNOMEDCT_CORE|Acne keloid|Acne keloid
C0001145|T047|FN|238746008|SNOMEDCT_CORE|Acne keloid|Acne keloid
C0001173|T020|PT|416605008|SNOMEDCT_CORE|Acquired obstruction of pylorus|Acquired obstruction of pylorus
C0001173|T020|FN|416605008|SNOMEDCT_CORE|Acquired obstruction of pylorus|Acquired obstruction of pylorus
C0001173|T020|SY|416605008|SNOMEDCT_CORE|Acquired pyloric obstruction|Acquired obstruction of pylorus
C0001175|T047|SY|62479008|SNOMEDCT_CORE|Acquired immune deficiency syndrome|AIDS
C0001175|T047|OF|62479008|SNOMEDCT_CORE|Acquired immune deficiency syndrome|AIDS
C0001175|T047|FN|62479008|SNOMEDCT_CORE|Acquired immune deficiency syndrome|AIDS
C0001175|T047|IS|62479008|SNOMEDCT_CORE|Acquired immune deficiency syndrome, NOS|AIDS
C0001175|T047|SY|62479008|SNOMEDCT_CORE|Acquired immunodeficiency syndrome|AIDS
C0001175|T047|IS|62479008|SNOMEDCT_CORE|Acquired immunodeficiency syndrome, NOS|AIDS
C0001175|T047|PT|62479008|SNOMEDCT_CORE|AIDS|AIDS
C0001175|T047|OF|62479008|SNOMEDCT_CORE|AIDS|AIDS
C0001175|T047|SY|62479008|SNOMEDCT_CORE|AIDS - Acquired immunodeficiency syndrome|AIDS
C0001175|T047|IS|62479008|SNOMEDCT_CORE|AIDS, NOS|AIDS
C0001175|T047|SY|62479008|SNOMEDCT_CORE|Immunodeficiency due to human immunodeficiency virus infection|AIDS
C0001206|T047|SY|74107003|SNOMEDCT_CORE|Acromegalia|Acromegaly
C0001206|T047|PT|74107003|SNOMEDCT_CORE|Acromegaly|Acromegaly
C0001206|T047|FN|74107003|SNOMEDCT_CORE|Acromegaly|Acromegaly
C0001206|T047|SY|74107003|SNOMEDCT_CORE|Anterior pituitary adenoma syndrome|Acromegaly
C0001206|T047|SY|74107003|SNOMEDCT_CORE|Growth hormone hypersecretion syndrome|Acromegaly
C0001206|T047|SY|74107003|SNOMEDCT_CORE|Marie disease|Acromegaly
C0001206|T047|SY|74107003|SNOMEDCT_CORE|STH hypersecretion syndrome|Acromegaly
C0001306|T047|SY|9953008|SNOMEDCT_CORE|Acute alcoholic hepatitis|Acute alcoholic liver disease
C0001306|T047|PT|9953008|SNOMEDCT_CORE|Acute alcoholic liver disease|Acute alcoholic liver disease
C0001306|T047|FN|9953008|SNOMEDCT_CORE|Acute alcoholic liver disease|Acute alcoholic liver disease
C0001308|T047|FN|197268000|SNOMEDCT_CORE|Acute and subacute liver necrosis|Acute and subacute liver necrosis
C0001308|T047|PT|197268000|SNOMEDCT_CORE|Acute and subacute liver necrosis|Acute and subacute liver necrosis
C0001309|T047|SY|67678004|SNOMEDCT_CORE|Acute allergic conjunctivitis|Acute atopic conjunctivitis
C0001309|T047|PT|67678004|SNOMEDCT_CORE|Acute atopic conjunctivitis|Acute atopic conjunctivitis
C0001309|T047|FN|67678004|SNOMEDCT_CORE|Acute atopic conjunctivitis|Acute atopic conjunctivitis
C0001309|T047|SY|67678004|SNOMEDCT_CORE|Angelucci's syndrome|Acute atopic conjunctivitis
C0001309|T047|SY|67678004|SNOMEDCT_CORE|Critical allergic conjunctivitis syndrome|Acute atopic conjunctivitis
C0001311|T047|PT|5505005|SNOMEDCT_CORE|Acute bronchiolitis|Acute bronchiolitis
C0001311|T047|FN|5505005|SNOMEDCT_CORE|Acute bronchiolitis|Acute bronchiolitis
C0001311|T047|IS|5505005|SNOMEDCT_CORE|Acute bronchiolitis, NOS|Acute bronchiolitis
C0001311|T047|SY|5505005|SNOMEDCT_CORE|Acute capillary bronchiolitis|Acute bronchiolitis
C0001311|T047|SY|5505005|SNOMEDCT_CORE|Capillary pneumonia|Acute bronchiolitis
C0001327|T047|PT|6655004|SNOMEDCT_CORE|Acute laryngitis|Acute laryngitis
C0001327|T047|FN|6655004|SNOMEDCT_CORE|Acute laryngitis|Acute laryngitis
C0001339|T047|PT|197456007|SNOMEDCT_CORE|Acute pancreatitis|Acute pancreatitis
C0001339|T047|FN|197456007|SNOMEDCT_CORE|Acute pancreatitis|Acute pancreatitis
C0001339|T047|SY|197456007|SNOMEDCT_CORE|AP - Acute pancreatitis|Acute pancreatitis
C0001342|T047|SY|21638000|SNOMEDCT_CORE|Acute pericementitis|Acute periodontitis
C0001342|T047|PT|21638000|SNOMEDCT_CORE|Acute periodontitis|Acute periodontitis
C0001342|T047|FN|21638000|SNOMEDCT_CORE|Acute periodontitis|Acute periodontitis
C0001342|T047|IS|21638000|SNOMEDCT_CORE|Aggressive periodontitis|Acute periodontitis
C0001344|T047|PT|363746003|SNOMEDCT_CORE|Acute pharyngitis|Acute pharyngitis
C0001344|T047|FN|363746003|SNOMEDCT_CORE|Acute pharyngitis|Acute pharyngitis
C0001361|T047|PT|17741008|SNOMEDCT_CORE|Acute tonsillitis|Acute tonsillitis
C0001361|T047|FN|17741008|SNOMEDCT_CORE|Acute tonsillitis|Acute tonsillitis
C0001361|T047|SY|17741008|SNOMEDCT_CORE|Infective tonsillitis|Acute tonsillitis
C0001365|T047|PT|288723005|SNOMEDCT_CORE|Acute ill-defined cerebrovascular disease|Acute ill-defined cerebrovascular disease
C0001365|T047|FN|288723005|SNOMEDCT_CORE|Acute ill-defined cerebrovascular disease|Acute ill-defined cerebrovascular disease
C0001403|T047|SY|363732003|SNOMEDCT_CORE|Addison disease|Addison's disease
C0001403|T047|PT|363732003|SNOMEDCT_CORE|Addison's disease|Addison's disease
C0001403|T047|FN|363732003|SNOMEDCT_CORE|Addison's disease|Addison's disease
C0001418|T191|SY|443961001|SNOMEDCT_CORE|Adenocarcinoma|Adenocarcinoma
C0001418|T191|PT|35917007|SNOMEDCT_CORE|Adenocarcinoma|Adenocarcinoma
C0001418|T191|FN|35917007|SNOMEDCT_CORE|Adenocarcinoma, no subtype|Adenocarcinoma
C0001418|T191|SY|35917007|SNOMEDCT_CORE|Adenocarcinoma, no subtype|Adenocarcinoma
C0001418|T191|IS|35917007|SNOMEDCT_CORE|Adenocarcinoma, NOS|Adenocarcinoma
C0001418|T191|PT|443961001|SNOMEDCT_CORE|Malignant adenomatous neoplasm|Adenocarcinoma
C0001418|T191|FN|443961001|SNOMEDCT_CORE|Malignant adenomatous neoplasm|Adenocarcinoma
C0001429|T191|PT|422470007|SNOMEDCT_CORE|Adenolymphoma|Adenolymphoma
C0001429|T191|FN|422470007|SNOMEDCT_CORE|Adenolymphoma|Adenolymphoma
C0001429|T191|SY|422470007|SNOMEDCT_CORE|Papillary cystadenoma lymphomatosum|Adenolymphoma
C0001429|T191|SY|422470007|SNOMEDCT_CORE|Warthin's tumor|Adenolymphoma
C0001429|T191|SYGB|422470007|SNOMEDCT_CORE|Warthin's tumour|Adenolymphoma
C0001430|T191|SY|443416007|SNOMEDCT_CORE|Adenoma|Adenoma
C0001430|T191|PT|32048006|SNOMEDCT_CORE|Adenoma|Adenoma
C0001430|T191|FN|32048006|SNOMEDCT_CORE|Adenoma, no subtype|Adenoma
C0001430|T191|SY|32048006|SNOMEDCT_CORE|Adenoma, no subtype|Adenoma
C0001430|T191|IS|32048006|SNOMEDCT_CORE|Adenoma, NOS|Adenoma
C0001430|T191|SY|443416007|SNOMEDCT_CORE|Benign adenoma|Adenoma
C0001430|T191|FN|443416007|SNOMEDCT_CORE|Benign adenomatous neoplasm|Adenoma
C0001430|T191|PT|443416007|SNOMEDCT_CORE|Benign adenomatous neoplasm|Adenoma
C0001486|T047|SY|25225006|SNOMEDCT_CORE|Adenovirus infection|Disease due to Adenovirus
C0001486|T047|IS|25225006|SNOMEDCT_CORE|Adenovirus infection, NOS|Disease due to Adenovirus
C0001486|T047|FN|25225006|SNOMEDCT_CORE|Disease caused by Adenovirus|Disease due to Adenovirus
C0001486|T047|SY|25225006|SNOMEDCT_CORE|Disease caused by Adenovirus|Disease due to Adenovirus
C0001486|T047|PT|25225006|SNOMEDCT_CORE|Disease due to Adenovirus|Disease due to Adenovirus
C0001486|T047|OF|25225006|SNOMEDCT_CORE|Disease due to Adenovirus|Disease due to Adenovirus
C0001486|T047|IS|25225006|SNOMEDCT_CORE|Disease due to Adenovirus, NOS|Disease due to Adenovirus
C0001539|T048|PT|57194009|SNOMEDCT_CORE|Adjustment disorder with depressed mood|Adjustment disorder with depressed mood
C0001539|T048|FN|57194009|SNOMEDCT_CORE|Adjustment disorder with depressed mood|Adjustment disorder with depressed mood
C0001541|T048|PT|66381006|SNOMEDCT_CORE|Adjustment disorder with mixed disturbance of emotions AND conduct|Adjustment disorder with mixed disturbance of emotions AND conduct
C0001541|T048|IS|66381006|SNOMEDCT_CORE|Adjustment disorder with mixed disturbance of emotions and conduct|Adjustment disorder with mixed disturbance of emotions AND conduct
C0001541|T048|FN|66381006|SNOMEDCT_CORE|Adjustment disorder with mixed disturbance of emotions AND conduct|Adjustment disorder with mixed disturbance of emotions AND conduct
C0001541|T048|SY|66381006|SNOMEDCT_CORE|Adjustment reaction with mixed disturbance of emotion and conduct|Adjustment disorder with mixed disturbance of emotions AND conduct
C0001542|T048|PT|55668003|SNOMEDCT_CORE|Adjustment disorder with mixed emotional features|Adjustment disorder with mixed emotional features
C0001542|T048|FN|55668003|SNOMEDCT_CORE|Adjustment disorder with mixed emotional features|Adjustment disorder with mixed emotional features
C0001542|T048|SY|55668003|SNOMEDCT_CORE|Adjustment reaction with mixed disturbance of emotion|Adjustment disorder with mixed emotional features
C0001546|T048|PT|17226007|SNOMEDCT_CORE|Adjustment disorder|Adjustment disorder
C0001546|T048|FN|17226007|SNOMEDCT_CORE|Adjustment disorder|Adjustment disorder
C0001546|T048|IS|17226007|SNOMEDCT_CORE|Adjustment disorder, NOS|Adjustment disorder
C0001546|T048|SY|192041001|SNOMEDCT_CORE|Brief situational non-psychotic disorder|Adjustment disorder
C0001546|T048|IS|17226007|SNOMEDCT_CORE|Brief situational non-psychotic disorder, NOS|Adjustment disorder
C0001548|T048|PT|192046006|SNOMEDCT_CORE|Brief depressive adjustment reaction|Brief depressive adjustment reaction
C0001548|T048|FN|192046006|SNOMEDCT_CORE|Brief depressive adjustment reaction|Brief depressive adjustment reaction
C0001621|T047|SY|30171000|SNOMEDCT_CORE|Adrenal disease|Disorder of adrenal gland
C0001621|T047|SY|30171000|SNOMEDCT_CORE|Adrenal disorder|Disorder of adrenal gland
C0001621|T047|IS|30171000|SNOMEDCT_CORE|Disease of adrenal gland|Disorder of adrenal gland
C0001621|T047|OF|30171000|SNOMEDCT_CORE|Disease of adrenal gland|Disorder of adrenal gland
C0001621|T047|IS|30171000|SNOMEDCT_CORE|Disease of adrenal gland, NOS|Disorder of adrenal gland
C0001621|T047|PT|30171000|SNOMEDCT_CORE|Disorder of adrenal gland|Disorder of adrenal gland
C0001621|T047|FN|30171000|SNOMEDCT_CORE|Disorder of adrenal gland|Disorder of adrenal gland
C0001621|T047|IS|30171000|SNOMEDCT_CORE|Disorder of adrenal gland, NOS|Disorder of adrenal gland
C0001622|T047|SY|47270006|SNOMEDCT_CORE|Hypercorticism|Hypercortisolism
C0001622|T047|PT|47270006|SNOMEDCT_CORE|Hypercortisolism|Hypercortisolism
C0001622|T047|FN|47270006|SNOMEDCT_CORE|Hypercortisolism|Hypercortisolism
C0001622|T047|SY|47270006|SNOMEDCT_CORE|Overproduction of cortisol|Hypercortisolism
C0001623|T047|OAS|111563005|SNOMEDCT_CORE|Adrenal failure|Hypoadrenalism
C0001623|T047|OAP|111563005|SNOMEDCT_CORE|Adrenal hypofunction|Hypoadrenalism
C0001623|T047|SY|237785004|SNOMEDCT_CORE|Adrenal hypofunction|Hypoadrenalism
C0001623|T047|OAF|111563005|SNOMEDCT_CORE|Adrenal hypofunction|Hypoadrenalism
C0001623|T047|PT|237785004|SNOMEDCT_CORE|Hypoadrenalism|Hypoadrenalism
C0001623|T047|FN|237785004|SNOMEDCT_CORE|Hypoadrenalism|Hypoadrenalism
C0001624|T191|SY|127021009|SNOMEDCT_CORE|Adrenal tumor|Neoplasm of adrenal gland
C0001624|T191|SYGB|127021009|SNOMEDCT_CORE|Adrenal tumour|Neoplasm of adrenal gland
C0001624|T191|PT|127021009|SNOMEDCT_CORE|Neoplasm of adrenal gland|Neoplasm of adrenal gland
C0001624|T191|FN|127021009|SNOMEDCT_CORE|Neoplasm of adrenal gland|Neoplasm of adrenal gland
C0001624|T191|SY|127021009|SNOMEDCT_CORE|Tumor of adrenal gland|Neoplasm of adrenal gland
C0001624|T191|SYGB|127021009|SNOMEDCT_CORE|Tumour of adrenal gland|Neoplasm of adrenal gland
C0001723|T048|PT|441704009|SNOMEDCT_CORE|Affective psychosis|Affective psychosis
C0001723|T048|FN|441704009|SNOMEDCT_CORE|Affective psychosis|Affective psychosis
C0001733|T047|PTGB|278504009|SNOMEDCT_CORE|Afibrinogenaemia|Afibrinogenemia
C0001733|T047|PT|278504009|SNOMEDCT_CORE|Afibrinogenemia|Afibrinogenemia
C0001733|T047|FN|278504009|SNOMEDCT_CORE|Afibrinogenemia|Afibrinogenemia
C0001815|T191|SY|52967002|SNOMEDCT_CORE|Agnogenic myeloid metaplasia|Myelosclerosis with myeloid metaplasia
C0001815|T191|SY|307651005|SNOMEDCT_CORE|Myelofibrosis with myeloid metaplasia|Myelosclerosis with myeloid metaplasia
C0001815|T191|PT|307651005|SNOMEDCT_CORE|Myelosclerosis with myeloid metaplasia|Myelosclerosis with myeloid metaplasia
C0001815|T191|FN|307651005|SNOMEDCT_CORE|Myelosclerosis with myeloid metaplasia|Myelosclerosis with myeloid metaplasia
C0001815|T191|SY|307651005|SNOMEDCT_CORE|Primary myelofibrosis|Myelosclerosis with myeloid metaplasia
C0001818|T048|PT|70691001|SNOMEDCT_CORE|Agoraphobia|Agoraphobia
C0001818|T048|FN|70691001|SNOMEDCT_CORE|Agoraphobia|Agoraphobia
C0001818|T048|IS|70691001|SNOMEDCT_CORE|Agoraphobia, NOS|Agoraphobia
C0001818|T048|SY|70691001|SNOMEDCT_CORE|Fear of open places|Agoraphobia
C0001818|T048|SY|70691001|SNOMEDCT_CORE|Phobia of going out|Agoraphobia
C0001824|T047|PT|17182001|SNOMEDCT_CORE|Agranulocytosis|Agranulocytosis
C0001824|T047|FN|17182001|SNOMEDCT_CORE|Agranulocytosis|Agranulocytosis
C0001824|T047|SY|17182001|SNOMEDCT_CORE|Schultz disease|Agranulocytosis
C0001883|T047|IS|79688008|SNOMEDCT_CORE|Airway obstruction|Respiratory obstruction
C0001883|T047|IS|79688008|SNOMEDCT_CORE|Airway obstruction, NOS|Respiratory obstruction
C0001883|T047|IS|68372009|SNOMEDCT_CORE|Airway obstruction, NOS|Respiratory obstruction
C0001883|T047|SY|79688008|SNOMEDCT_CORE|Embarrassed airway|Respiratory obstruction
C0001883|T047|PT|79688008|SNOMEDCT_CORE|Respiratory obstruction|Respiratory obstruction
C0001883|T047|FN|79688008|SNOMEDCT_CORE|Respiratory obstruction|Respiratory obstruction
C0001925|T033|IS|29738008|SNOMEDCT_CORE|Albuminuria|Albuminuria
C0001925|T033|PT|274769005|SNOMEDCT_CORE|Albuminuria|Albuminuria
C0001925|T033|FN|274769005|SNOMEDCT_CORE|Albuminuria|Albuminuria
C0001925|T033|IS|29738008|SNOMEDCT_CORE|Albuminuria, NOS|Albuminuria
C0001957|T047|PT|8635005|SNOMEDCT_CORE|Alcohol withdrawal delirium|Alcohol withdrawal delirium
C0001957|T047|FN|8635005|SNOMEDCT_CORE|Alcohol withdrawal delirium|Alcohol withdrawal delirium
C0001957|T047|SY|8635005|SNOMEDCT_CORE|Delirium tremens|Alcohol withdrawal delirium
C0001957|T047|SY|8635005|SNOMEDCT_CORE|DTs - delirium tremens|Alcohol withdrawal delirium
C0001969|T048|PT|25702006|SNOMEDCT_CORE|Alcohol intoxication|Alcohol intoxication
C0001969|T048|FN|25702006|SNOMEDCT_CORE|Alcohol intoxication|Alcohol intoxication
C0001969|T048|SY|25702006|SNOMEDCT_CORE|Drunk|Alcohol intoxication
C0001969|T048|SY|25702006|SNOMEDCT_CORE|Drunkenness|Alcohol intoxication
C0001973|T048|PT|66590003|SNOMEDCT_CORE|Alcohol dependence|Alcohol dependence
C0001973|T048|FN|66590003|SNOMEDCT_CORE|Alcohol dependence|Alcohol dependence
C0001973|T048|SY|66590003|SNOMEDCT_CORE|Alcohol dependence syndrome|Alcohol dependence
C0001973|T048|SY|7200002|SNOMEDCT_CORE|Alcohol problem drinking|Alcohol dependence
C0001973|T048|PT|7200002|SNOMEDCT_CORE|Alcoholism|Alcohol dependence
C0001973|T048|FN|7200002|SNOMEDCT_CORE|Alcoholism|Alcohol dependence
C0001973|T048|IS|7200002|SNOMEDCT_CORE|Alcoholism, NOS|Alcohol dependence
C0001973|T048|SY|284591009|SNOMEDCT_CORE|Chronic alcohol abuse|Alcohol dependence
C0001973|T048|SY|66590003|SNOMEDCT_CORE|Chronic alcoholism|Alcohol dependence
C0001973|T048|SY|7200002|SNOMEDCT_CORE|Dipsomania|Alcohol dependence
C0001973|T048|PT|284591009|SNOMEDCT_CORE|Persistent alcohol abuse|Alcohol dependence
C0001973|T048|FN|284591009|SNOMEDCT_CORE|Persistent alcohol abuse|Alcohol dependence
C0002170|T047|PT|56317004|SNOMEDCT_CORE|Alopecia|Alopecia
C0002170|T047|FN|56317004|SNOMEDCT_CORE|Alopecia|Alopecia
C0002170|T047|IS|56317004|SNOMEDCT_CORE|Alopecia, NOS|Alopecia
C0002170|T047|SY|56317004|SNOMEDCT_CORE|Bald|Alopecia
C0002170|T047|SY|56317004|SNOMEDCT_CORE|Baldness|Alopecia
C0002170|T047|SY|56317004|SNOMEDCT_CORE|Hair loss disorder|Alopecia
C0002170|T047|IS|56317004|SNOMEDCT_CORE|Loss of hair|Alopecia
C0002171|T047|SY|68225006|SNOMEDCT_CORE|AA - Alopecia areata|Alopecia areata
C0002171|T047|PT|68225006|SNOMEDCT_CORE|Alopecia areata|Alopecia areata
C0002171|T047|FN|68225006|SNOMEDCT_CORE|Alopecia areata|Alopecia areata
C0002171|T047|SY|68225006|SNOMEDCT_CORE|Alopecia circumscripta|Alopecia areata
C0002171|T047|SY|68225006|SNOMEDCT_CORE|Circumscribed alopecia|Alopecia areata
C0002171|T047|SY|68225006|SNOMEDCT_CORE|Patchy loss of hair|Alopecia areata
C0002312|T047|PTGB|68913001|SNOMEDCT_CORE|Alpha thalassaemia|Alpha thalassemia
C0002312|T047|SYGB|68913001|SNOMEDCT_CORE|alpha thalassaemia|Alpha thalassemia
C0002312|T047|OP|68913001|SNOMEDCT_CORE|alpha Thalassaemia|Alpha thalassemia
C0002312|T047|SYGB|68913001|SNOMEDCT_CORE|Alpha thalassaemia syndrome|Alpha thalassemia
C0002312|T047|PT|68913001|SNOMEDCT_CORE|Alpha thalassemia|Alpha thalassemia
C0002312|T047|SY|68913001|SNOMEDCT_CORE|alpha thalassemia|Alpha thalassemia
C0002312|T047|OP|68913001|SNOMEDCT_CORE|alpha Thalassemia|Alpha thalassemia
C0002312|T047|FN|68913001|SNOMEDCT_CORE|Alpha thalassemia|Alpha thalassemia
C0002312|T047|OF|68913001|SNOMEDCT_CORE|alpha Thalassemia|Alpha thalassemia
C0002312|T047|SY|68913001|SNOMEDCT_CORE|Alpha thalassemia syndrome|Alpha thalassemia
C0002312|T047|IS|68913001|SNOMEDCT_CORE|alpha Thalassemia, NOS|Alpha thalassemia
C0002390|T047|SY|37471005|SNOMEDCT_CORE|Allergic alveolitis|Extrinsic allergic alveolitis
C0002390|T047|IS|37471005|SNOMEDCT_CORE|Allergic alveolitis, NOS|Extrinsic allergic alveolitis
C0002390|T047|SY|37471005|SNOMEDCT_CORE|Allergic interstitial pneumonitis|Extrinsic allergic alveolitis
C0002390|T047|IS|37471005|SNOMEDCT_CORE|Allergic interstitial pneumonitis, NOS|Extrinsic allergic alveolitis
C0002390|T047|SY|37471005|SNOMEDCT_CORE|Allergic pneumonitis|Extrinsic allergic alveolitis
C0002390|T047|IS|37471005|SNOMEDCT_CORE|Allergic pneumonitis, NOS|Extrinsic allergic alveolitis
C0002390|T047|SY|37471005|SNOMEDCT_CORE|Bagpipe lung|Extrinsic allergic alveolitis
C0002390|T047|SY|37471005|SNOMEDCT_CORE|EAA - Extrinsic allergic alveolitis|Extrinsic allergic alveolitis
C0002390|T047|PT|37471005|SNOMEDCT_CORE|Extrinsic allergic alveolitis|Extrinsic allergic alveolitis
C0002390|T047|FN|37471005|SNOMEDCT_CORE|Extrinsic allergic alveolitis|Extrinsic allergic alveolitis
C0002390|T047|IS|37471005|SNOMEDCT_CORE|Extrinsic allergic alveolitis, NOS|Extrinsic allergic alveolitis
C0002390|T047|SY|37471005|SNOMEDCT_CORE|Extrinsic allergic bronchiolo-alveolitis|Extrinsic allergic alveolitis
C0002390|T047|IS|37471005|SNOMEDCT_CORE|Extrinsic allergic bronchiolo-alveolitis, NOS|Extrinsic allergic alveolitis
C0002390|T047|SY|37471005|SNOMEDCT_CORE|Hypersensitivity pneumonia|Extrinsic allergic alveolitis
C0002390|T047|IS|37471005|SNOMEDCT_CORE|Hypersensitivity pneumonia, NOS|Extrinsic allergic alveolitis
C0002390|T047|SY|37471005|SNOMEDCT_CORE|Hypersensitivity pneumonitis|Extrinsic allergic alveolitis
C0002390|T047|IS|37471005|SNOMEDCT_CORE|Hypersensitivity pneumonitis, NOS|Extrinsic allergic alveolitis
C0002395|T047|SY|26929004|SNOMEDCT_CORE|AD - Alzheimer's disease|Alzheimer's disease
C0002395|T047|SY|26929004|SNOMEDCT_CORE|Alzheimer dementia|Alzheimer's disease
C0002395|T047|SY|26929004|SNOMEDCT_CORE|Alzheimer disease|Alzheimer's disease
C0002395|T047|PT|26929004|SNOMEDCT_CORE|Alzheimer's disease|Alzheimer's disease
C0002395|T047|FN|26929004|SNOMEDCT_CORE|Alzheimer's disease|Alzheimer's disease
C0002395|T047|IS|26929004|SNOMEDCT_CORE|Alzheimer's disease, NOS|Alzheimer's disease
C0002395|T047|IS|26929004|SNOMEDCT_CORE|Alzheimers disease|Alzheimer's disease
C0002418|T047|PT|387742006|SNOMEDCT_CORE|Amblyopia|Amblyopia
C0002418|T047|FN|387742006|SNOMEDCT_CORE|Amblyopia|Amblyopia
C0002418|T047|SY|387742006|SNOMEDCT_CORE|Amblyopic|Amblyopia
C0002453|T033|SY|14302001|SNOMEDCT_CORE|Absence of menstruation|Amenorrhea
C0002453|T033|IS|14302001|SNOMEDCT_CORE|Absence of menstruation, NOS|Amenorrhea
C0002453|T033|PT|14302001|SNOMEDCT_CORE|Amenorrhea|Amenorrhea
C0002453|T033|FN|14302001|SNOMEDCT_CORE|Amenorrhea|Amenorrhea
C0002453|T033|IS|14302001|SNOMEDCT_CORE|Amenorrhea, NOS|Amenorrhea
C0002453|T033|PTGB|14302001|SNOMEDCT_CORE|Amenorrhoea|Amenorrhea
C0002453|T033|IS|14302001|SNOMEDCT_CORE|Amenorrhoea, NOS|Amenorrhea
C0002622|T048|PT|48167000|SNOMEDCT_CORE|Amnesia|Amnesia
C0002622|T048|FN|48167000|SNOMEDCT_CORE|Amnesia|Amnesia
C0002622|T048|IS|48167000|SNOMEDCT_CORE|Amnesia, NOS|Amnesia
C0002622|T048|IS|48167000|SNOMEDCT_CORE|Dysmnesia|Amnesia
C0002622|T048|SY|386807006|SNOMEDCT_CORE|Dysmnesia|Amnesia
C0002622|T048|SY|48167000|SNOMEDCT_CORE|LOM - Loss of memory|Amnesia
C0002622|T048|SY|48167000|SNOMEDCT_CORE|Loss of memory|Amnesia
C0002622|T048|SY|48167000|SNOMEDCT_CORE|Memory gone|Amnesia
C0002622|T048|SY|48167000|SNOMEDCT_CORE|Memory loss|Amnesia
C0002622|T048|SY|48167000|SNOMEDCT_CORE|Memory loss - amnesia|Amnesia
C0002726|T047|PT|17602002|SNOMEDCT_CORE|Amyloidosis|Amyloidosis
C0002726|T047|FN|17602002|SNOMEDCT_CORE|Amyloidosis|Amyloidosis
C0002726|T047|IS|17602002|SNOMEDCT_CORE|Amyloidosis, NOS|Amyloidosis
C0002736|T047|SY|86044005|SNOMEDCT_CORE|ALS - Amyotrophic lateral sclerosis|Amyotrophic lateral sclerosis
C0002736|T047|PT|86044005|SNOMEDCT_CORE|Amyotrophic lateral sclerosis|Amyotrophic lateral sclerosis
C0002736|T047|FN|86044005|SNOMEDCT_CORE|Amyotrophic lateral sclerosis|Amyotrophic lateral sclerosis
C0002736|T047|SY|86044005|SNOMEDCT_CORE|Bulbar motor neuron disease|Amyotrophic lateral sclerosis
C0002736|T047|SY|86044005|SNOMEDCT_CORE|Lou Gehrig's disease|Amyotrophic lateral sclerosis
C0002753|T020|FN|197210001|SNOMEDCT_CORE|Anal and rectal polyp|Anal and rectal polyp
C0002753|T020|PT|197210001|SNOMEDCT_CORE|Anal and rectal polyp|Anal and rectal polyp
C0002792|T047|IS|39579001|SNOMEDCT_CORE|Allergic shock|Anaphylaxis
C0002792|T047|SY|39579001|SNOMEDCT_CORE|Anaphylactic reaction|Anaphylaxis
C0002792|T047|IS|39579001|SNOMEDCT_CORE|Anaphylactic shock|Anaphylaxis
C0002792|T047|PT|39579001|SNOMEDCT_CORE|Anaphylaxis|Anaphylaxis
C0002792|T047|FN|39579001|SNOMEDCT_CORE|Anaphylaxis|Anaphylaxis
C0002792|T047|SYGB|39579001|SNOMEDCT_CORE|Generalised anaphylaxis|Anaphylaxis
C0002792|T047|SY|39579001|SNOMEDCT_CORE|Generalized anaphylaxis|Anaphylaxis
C0002792|T047|SY|39579001|SNOMEDCT_CORE|Systemic anaphylaxis|Anaphylaxis
C0002871|T047|PTGB|271737000|SNOMEDCT_CORE|Anaemia|Anemia
C0002871|T047|OP|271737000|SNOMEDCT_CORE|Anaemia|Anemia
C0002871|T047|PT|271737000|SNOMEDCT_CORE|Anemia|Anemia
C0002871|T047|FN|271737000|SNOMEDCT_CORE|Anemia|Anemia
C0002871|T047|IS|271737000|SNOMEDCT_CORE|Anemia|Anemia
C0002873|T047|PTGB|234347009|SNOMEDCT_CORE|Anaemia of chronic disease|Anemia of chronic disease
C0002873|T047|SYGB|234347009|SNOMEDCT_CORE|Anaemia of chronic disorder|Anemia of chronic disease
C0002873|T047|SYGB|234347009|SNOMEDCT_CORE|Anaemia of systemic disease|Anemia of chronic disease
C0002873|T047|PT|234347009|SNOMEDCT_CORE|Anemia of chronic disease|Anemia of chronic disease
C0002873|T047|SY|234347009|SNOMEDCT_CORE|Anemia of chronic disorder|Anemia of chronic disease
C0002873|T047|FN|234347009|SNOMEDCT_CORE|Anemia of chronic disorder|Anemia of chronic disease
C0002873|T047|SY|234347009|SNOMEDCT_CORE|Anemia of systemic disease|Anemia of chronic disease
C0002873|T047|SY|234347009|SNOMEDCT_CORE|Secondary anemia|Anemia of chronic disease
C0002874|T047|PTGB|306058006|SNOMEDCT_CORE|Aplastic anaemia|Aplastic anemia
C0002874|T047|PT|306058006|SNOMEDCT_CORE|Aplastic anemia|Aplastic anemia
C0002874|T047|FN|306058006|SNOMEDCT_CORE|Aplastic anemia|Aplastic anemia
C0002874|T047|SY|306058006|SNOMEDCT_CORE|Erythroid aplasia|Aplastic anemia
C0002875|T047|SYGB|26682008|SNOMEDCT_CORE|Beta thalassaemia major|Homozygous beta thalassemia
C0002875|T047|SYGB|26682008|SNOMEDCT_CORE|Cooley's anaemia|Homozygous beta thalassemia
C0002875|T047|SY|26682008|SNOMEDCT_CORE|Cooley's anemia|Homozygous beta thalassemia
C0002875|T047|PTGB|26682008|SNOMEDCT_CORE|Homozygous beta thalassaemia|Homozygous beta thalassemia
C0002875|T047|PT|26682008|SNOMEDCT_CORE|Homozygous beta thalassemia|Homozygous beta thalassemia
C0002875|T047|FN|26682008|SNOMEDCT_CORE|Homozygous beta thalassemia|Homozygous beta thalassemia
C0002875|T047|SY|26682008|SNOMEDCT_CORE|Mediterranean anemia|Homozygous beta thalassemia
C0002878|T047|PTGB|61261009|SNOMEDCT_CORE|Haemolytic anaemia|Hemolytic anemia
C0002878|T047|PT|61261009|SNOMEDCT_CORE|Hemolytic anemia|Hemolytic anemia
C0002878|T047|FN|61261009|SNOMEDCT_CORE|Hemolytic anemia|Hemolytic anemia
C0002878|T047|IS|61261009|SNOMEDCT_CORE|Hemolytic anemia, NOS|Hemolytic anemia
C0002879|T047|PTGB|4854004|SNOMEDCT_CORE|Acquired haemolytic anaemia|Acquired hemolytic anemia
C0002879|T047|PT|4854004|SNOMEDCT_CORE|Acquired hemolytic anemia|Acquired hemolytic anemia
C0002879|T047|FN|4854004|SNOMEDCT_CORE|Acquired hemolytic anemia|Acquired hemolytic anemia
C0002879|T047|IS|4854004|SNOMEDCT_CORE|Acquired hemolytic anemia, NOS|Acquired hemolytic anemia
C0002880|T047|PTGB|413603009|SNOMEDCT_CORE|Autoimmune haemolytic anaemia|Autoimmune hemolytic anemia
C0002880|T047|PT|413603009|SNOMEDCT_CORE|Autoimmune hemolytic anemia|Autoimmune hemolytic anemia
C0002880|T047|FN|413603009|SNOMEDCT_CORE|Autoimmune hemolytic anemia|Autoimmune hemolytic anemia
C0002886|T047|PTGB|83414005|SNOMEDCT_CORE|Macrocytic anaemia|Macrocytic anemia
C0002886|T047|PT|83414005|SNOMEDCT_CORE|Macrocytic anemia|Macrocytic anemia
C0002886|T047|FN|83414005|SNOMEDCT_CORE|Macrocytic anemia|Macrocytic anemia
C0002888|T047|PTGB|53165003|SNOMEDCT_CORE|Megaloblastic anaemia|Megaloblastic anemia
C0002888|T047|PT|53165003|SNOMEDCT_CORE|Megaloblastic anemia|Megaloblastic anemia
C0002888|T047|FN|53165003|SNOMEDCT_CORE|Megaloblastic anemia|Megaloblastic anemia
C0002888|T047|IS|53165003|SNOMEDCT_CORE|Megaloblastic anemia, NOS|Megaloblastic anemia
C0002892|T047|SY|84027009|SNOMEDCT_CORE|Addison's anemia|Pernicious anemia
C0002892|T047|SYGB|84027009|SNOMEDCT_CORE|Addisonian pernicious anaemia|Pernicious anemia
C0002892|T047|SY|84027009|SNOMEDCT_CORE|Addisonian pernicious anemia|Pernicious anemia
C0002892|T047|SYGB|84027009|SNOMEDCT_CORE|Biermer's anaemia|Pernicious anemia
C0002892|T047|SY|84027009|SNOMEDCT_CORE|Biermer's anemia|Pernicious anemia
C0002892|T047|SYGB|84027009|SNOMEDCT_CORE|Megaloblastic anaemia due to impaired absorption of cobalamin|Pernicious anemia
C0002892|T047|SY|84027009|SNOMEDCT_CORE|Megaloblastic anemia due to impaired absorption of cobalamin|Pernicious anemia
C0002892|T047|SYGB|84027009|SNOMEDCT_CORE|PA - Pernicious anaemia|Pernicious anemia
C0002892|T047|PTGB|84027009|SNOMEDCT_CORE|Pernicious anaemia|Pernicious anemia
C0002892|T047|PT|84027009|SNOMEDCT_CORE|Pernicious anemia|Pernicious anemia
C0002892|T047|FN|84027009|SNOMEDCT_CORE|Pernicious anemia|Pernicious anemia
C0002892|T047|IS|84027009|SNOMEDCT_CORE|Pernicious anemia, NOS|Pernicious anemia
C0002893|T047|PTGB|128845005|SNOMEDCT_CORE|Refractory anaemia|Refractory anemia
C0002893|T047|PT|128845005|SNOMEDCT_CORE|Refractory anemia|Refractory anemia
C0002893|T047|FN|128845005|SNOMEDCT_CORE|Refractory anemia|Refractory anemia
C0002895|T047|SY|417357006|SNOMEDCT_CORE|Sickle cell disease|Sickling disorder due to hemoglobin S
C0002895|T047|SY|417357006|SNOMEDCT_CORE|Sickle cell syndrome|Sickling disorder due to hemoglobin S
C0002895|T047|PTGB|417357006|SNOMEDCT_CORE|Sickling disorder due to haemoglobin S|Sickling disorder due to hemoglobin S
C0002895|T047|FN|417357006|SNOMEDCT_CORE|Sickling disorder due to hemoglobin S|Sickling disorder due to hemoglobin S
C0002895|T047|PT|417357006|SNOMEDCT_CORE|Sickling disorder due to hemoglobin S|Sickling disorder due to hemoglobin S
C0002940|T046|PT|432119003|SNOMEDCT_CORE|Aneurysm|Aneurysm
C0002940|T046|FN|432119003|SNOMEDCT_CORE|Aneurysm|Aneurysm
C0002962|T184|SY|194828000|SNOMEDCT_CORE|Angina|Angina pectoris
C0002962|T184|FN|194828000|SNOMEDCT_CORE|Angina|Angina pectoris
C0002962|T184|PT|194828000|SNOMEDCT_CORE|Angina pectoris|Angina pectoris
C0002962|T184|SY|194828000|SNOMEDCT_CORE|Anginal syndrome|Angina pectoris
C0002962|T184|SY|194828000|SNOMEDCT_CORE|AP - Angina pectoris|Angina pectoris
C0002962|T184|SY|194828000|SNOMEDCT_CORE|Cardiac angina|Angina pectoris
C0002962|T184|SYGB|194828000|SNOMEDCT_CORE|Ischaemic heart disease - angina|Angina pectoris
C0002962|T184|SY|194828000|SNOMEDCT_CORE|Ischemic heart disease - angina|Angina pectoris
C0002962|T184|SY|194828000|SNOMEDCT_CORE|Stenocardia|Angina pectoris
C0002963|T047|SY|87343002|SNOMEDCT_CORE|Coronary artery spasm angina|Prinzmetal angina
C0002963|T047|IS|87343002|SNOMEDCT_CORE|Prinzmental angina|Prinzmetal angina
C0002963|T047|PT|87343002|SNOMEDCT_CORE|Prinzmetal angina|Prinzmetal angina
C0002963|T047|FN|87343002|SNOMEDCT_CORE|Prinzmetal angina|Prinzmetal angina
C0002963|T047|SY|87343002|SNOMEDCT_CORE|Prinzmetal's angina|Prinzmetal angina
C0002963|T047|SY|87343002|SNOMEDCT_CORE|Variant angina|Prinzmetal angina
C0002963|T047|SY|87343002|SNOMEDCT_CORE|Variant angina pectoris|Prinzmetal angina
C0002965|T047|SY|4557003|SNOMEDCT_CORE|Crescendo angina|Intermediate coronary syndrome
C0002965|T047|IS|4557003|SNOMEDCT_CORE|Impending infarction|Intermediate coronary syndrome
C0002965|T047|SY|4557003|SNOMEDCT_CORE|Intermediate coronary syndrome|Intermediate coronary syndrome
C0002965|T047|OAP|64333001|SNOMEDCT_CORE|Preinfarction angina|Intermediate coronary syndrome
C0002965|T047|OAF|64333001|SNOMEDCT_CORE|Preinfarction angina|Intermediate coronary syndrome
C0002965|T047|SY|4557003|SNOMEDCT_CORE|Unstable angina|Intermediate coronary syndrome
C0002965|T047|SY|4557003|SNOMEDCT_CORE|Worsening angina|Intermediate coronary syndrome
C0002991|T191|SY|254750001|SNOMEDCT_CORE|Benign fibrous histiocytoma of skin|Fibrous histiocytoma of skin
C0002991|T191|PT|254750001|SNOMEDCT_CORE|Fibrous histiocytoma of skin|Fibrous histiocytoma of skin
C0002991|T191|FN|254750001|SNOMEDCT_CORE|Fibrous histiocytoma of skin|Fibrous histiocytoma of skin
C0002991|T191|SY|254750001|SNOMEDCT_CORE|Fibrous xanthoma of skin|Fibrous histiocytoma of skin
C0002994|T046|PTGB|41291007|SNOMEDCT_CORE|Angio-oedema|Angioedema
C0002994|T046|SYGB|41291007|SNOMEDCT_CORE|Angio-oedema-urticaria|Angioedema
C0002994|T046|PT|41291007|SNOMEDCT_CORE|Angioedema|Angioedema
C0002994|T046|FN|41291007|SNOMEDCT_CORE|Angioedema|Angioedema
C0002994|T046|SY|41291007|SNOMEDCT_CORE|Angioedema-urticaria|Angioedema
C0002994|T046|IS|41291007|SNOMEDCT_CORE|Angioedema, NOS|Angioedema
C0002994|T046|SY|41291007|SNOMEDCT_CORE|Angioneurotic edema|Angioedema
C0002994|T046|IS|41291007|SNOMEDCT_CORE|Angioneurotic edema, NOS|Angioedema
C0002994|T046|SYGB|41291007|SNOMEDCT_CORE|Angioneurotic oedema|Angioedema
C0002994|T046|IS|41291007|SNOMEDCT_CORE|Giant urticaria|Angioedema
C0002994|T046|SY|41291007|SNOMEDCT_CORE|Quincke's disease|Angioedema
C0002994|T046|SY|41291007|SNOMEDCT_CORE|Quincke's edema|Angioedema
C0002994|T046|SYGB|41291007|SNOMEDCT_CORE|Quincke's oedema|Angioedema
C0002994|T046|SYGB|41291007|SNOMEDCT_CORE|Urticaria-angio-oedema|Angioedema
C0002994|T046|SY|41291007|SNOMEDCT_CORE|Urticaria-angioedema|Angioedema
C0003079|T033|PT|13045009|SNOMEDCT_CORE|Anisocoria|Anisocoria
C0003079|T033|FN|13045009|SNOMEDCT_CORE|Anisocoria|Anisocoria
C0003079|T033|SY|13045009|SNOMEDCT_CORE|Anisocoria - unequal pupil diameter|Anisocoria
C0003079|T033|SY|13045009|SNOMEDCT_CORE|Unequal pupil diameter|Anisocoria
C0003079|T033|SY|13045009|SNOMEDCT_CORE|Unequal pupils|Anisocoria
C0003081|T047|PT|3289004|SNOMEDCT_CORE|Anisometropia|Anisometropia
C0003081|T047|FN|3289004|SNOMEDCT_CORE|Anisometropia|Anisometropia
C0003090|T046|PT|111227009|SNOMEDCT_CORE|Ankylosis of joint|Ankylosis of joint
C0003090|T046|FN|111227009|SNOMEDCT_CORE|Ankylosis of joint|Ankylosis of joint
C0003119|T019|IS|7183006|SNOMEDCT_CORE|Agenesis of eye|Anophthalmos
C0003119|T019|SY|7183006|SNOMEDCT_CORE|Agenesis of eyes|Anophthalmos
C0003119|T019|SY|7183006|SNOMEDCT_CORE|Anophthalmia|Anophthalmos
C0003119|T019|PT|7183006|SNOMEDCT_CORE|Anophthalmos|Anophthalmos
C0003119|T019|FN|7183006|SNOMEDCT_CORE|Anophthalmos|Anophthalmos
C0003119|T019|IS|7183006|SNOMEDCT_CORE|Anophthalmos, NOS|Anophthalmos
C0003119|T019|SY|7183006|SNOMEDCT_CORE|Clinical anophthalmos|Anophthalmos
C0003119|T019|IS|7183006|SNOMEDCT_CORE|Clinical anophthalmos, NOS|Anophthalmos
C0003119|T019|SY|7183006|SNOMEDCT_CORE|Congenital absence of eye|Anophthalmos
C0003119|T019|SY|7183006|SNOMEDCT_CORE|Congenital absence of eyes|Anophthalmos
C0003125|T048|SY|56882008|SNOMEDCT_CORE|AN - Anorexia nervosa|Anorexia nervosa
C0003125|T048|PT|56882008|SNOMEDCT_CORE|Anorexia nervosa|Anorexia nervosa
C0003125|T048|FN|56882008|SNOMEDCT_CORE|Anorexia nervosa|Anorexia nervosa
C0003126|T033|IS|44169009|SNOMEDCT_CORE|Absent sense of smell|Loss of sense of smell
C0003126|T033|SY|44169009|SNOMEDCT_CORE|Absent smell|Loss of sense of smell
C0003126|T033|SY|44169009|SNOMEDCT_CORE|Anosmia|Loss of sense of smell
C0003126|T033|PT|44169009|SNOMEDCT_CORE|Loss of sense of smell|Loss of sense of smell
C0003126|T033|FN|44169009|SNOMEDCT_CORE|Loss of sense of smell|Loss of sense of smell
C0003126|T033|SY|44169009|SNOMEDCT_CORE|Loss of the sense of smell|Loss of sense of smell
C0003126|T033|SY|44169009|SNOMEDCT_CORE|No sense of smell|Loss of sense of smell
C0003126|T033|SY|44169009|SNOMEDCT_CORE|Sense of smell absent|Loss of sense of smell
C0003126|T033|SY|44169009|SNOMEDCT_CORE|Sense of smell lost|Loss of sense of smell
C0003128|T047|PT|34571000|SNOMEDCT_CORE|Anovulation|Anovulation
C0003128|T047|FN|34571000|SNOMEDCT_CORE|Anovulation|Anovulation
C0003128|T047|SY|34571000|SNOMEDCT_CORE|Ovulation absent|Anovulation
C0003132|T046|SY|389098007|SNOMEDCT_CORE|Anoxic brain damage|Anoxic encephalopathy
C0003132|T046|SY|389098007|SNOMEDCT_CORE|Anoxic brain injury|Anoxic encephalopathy
C0003132|T046|PT|389098007|SNOMEDCT_CORE|Anoxic encephalopathy|Anoxic encephalopathy
C0003132|T046|FN|389098007|SNOMEDCT_CORE|Anoxic encephalopathy|Anoxic encephalopathy
C0003431|T048|PT|26665006|SNOMEDCT_CORE|Antisocial personality disorder|Antisocial personality disorder
C0003431|T048|FN|26665006|SNOMEDCT_CORE|Antisocial personality disorder|Antisocial personality disorder
C0003431|T048|SY|26665006|SNOMEDCT_CORE|Dissocial personality disorder|Antisocial personality disorder
C0003431|T048|SY|26665006|SNOMEDCT_CORE|Psychopathic personality disorder|Antisocial personality disorder
C0003431|T048|SY|26665006|SNOMEDCT_CORE|Sociopathic personality disorder|Antisocial personality disorder
C0003467|T048|PT|48694002|SNOMEDCT_CORE|Anxiety|Anxiety
C0003467|T048|FN|48694002|SNOMEDCT_CORE|Anxiety|Anxiety
C0003467|T048|SY|48694002|SNOMEDCT_CORE|Anxiety reaction|Anxiety
C0003467|T048|SY|48694002|SNOMEDCT_CORE|Anxiousness|Anxiety
C0003467|T048|SY|48694002|SNOMEDCT_CORE|Feeling anxious|Anxiety
C0003469|T048|PT|197480006|SNOMEDCT_CORE|Anxiety disorder|Anxiety disorder
C0003469|T048|FN|197480006|SNOMEDCT_CORE|Anxiety disorder|Anxiety disorder
C0003477|T048|FN|126943008|SNOMEDCT_CORE|Separation anxiety|Separation anxiety
C0003477|T048|PT|126943008|SNOMEDCT_CORE|Separation anxiety|Separation anxiety
C0003486|T047|SY|67362008|SNOMEDCT_CORE|AA - Aortic aneurysm|Aortic aneurysm
C0003486|T047|SY|67362008|SNOMEDCT_CORE|Aneurysm of aorta|Aortic aneurysm
C0003486|T047|IS|67362008|SNOMEDCT_CORE|Aneurysm of aorta, NOS|Aortic aneurysm
C0003486|T047|PT|67362008|SNOMEDCT_CORE|Aortic aneurysm|Aortic aneurysm
C0003486|T047|FN|67362008|SNOMEDCT_CORE|Aortic aneurysm|Aortic aneurysm
C0003486|T047|IS|67362008|SNOMEDCT_CORE|Aortic aneurysm, NOS|Aortic aneurysm
C0003490|T047|SY|359789008|SNOMEDCT_CORE|Aortic arch syndrome|Aortic arch syndrome
C0003492|T019|SY|7305005|SNOMEDCT_CORE|Aortic coarctation|Coarctation of aorta
C0003492|T019|SY|7305005|SNOMEDCT_CORE|Coarctation|Coarctation of aorta
C0003492|T019|PT|7305005|SNOMEDCT_CORE|Coarctation of aorta|Coarctation of aorta
C0003492|T019|FN|7305005|SNOMEDCT_CORE|Coarctation of aorta|Coarctation of aorta
C0003504|T047|SY|60234000|SNOMEDCT_CORE|AI - Aortic incompetence|Aortic valve regurgitation
C0003504|T047|SY|60234000|SNOMEDCT_CORE|Aortic incompetence|Aortic valve regurgitation
C0003504|T047|SY|60234000|SNOMEDCT_CORE|Aortic insufficiency|Aortic valve regurgitation
C0003504|T047|SY|60234000|SNOMEDCT_CORE|Aortic regurgitation|Aortic valve regurgitation
C0003504|T047|IS|60234000|SNOMEDCT_CORE|Aortic regurgitation, NOS|Aortic valve regurgitation
C0003504|T047|SY|60234000|SNOMEDCT_CORE|Aortic valve incompetence|Aortic valve regurgitation
C0003504|T047|IS|60234000|SNOMEDCT_CORE|Aortic valve incompetence, NOS|Aortic valve regurgitation
C0003504|T047|SY|60234000|SNOMEDCT_CORE|Aortic valve insufficiency|Aortic valve regurgitation
C0003504|T047|IS|60234000|SNOMEDCT_CORE|Aortic valve insufficiency, NOS|Aortic valve regurgitation
C0003504|T047|PT|60234000|SNOMEDCT_CORE|Aortic valve regurgitation|Aortic valve regurgitation
C0003504|T047|FN|60234000|SNOMEDCT_CORE|Aortic valve regurgitation|Aortic valve regurgitation
C0003504|T047|IS|60234000|SNOMEDCT_CORE|Aortic valve regurgitation, NOS|Aortic valve regurgitation
C0003504|T047|SY|60234000|SNOMEDCT_CORE|AR - Aortic regurgitation|Aortic valve regurgitation
C0003507|T047|IS|60573004|SNOMEDCT_CORE|Aortic stenosis|Aortic valve stenosis
C0003507|T047|PT|60573004|SNOMEDCT_CORE|Aortic valve stenosis|Aortic valve stenosis
C0003507|T047|FN|60573004|SNOMEDCT_CORE|Aortic valve stenosis|Aortic valve stenosis
C0003507|T047|IS|60573004|SNOMEDCT_CORE|Aortic valve stenosis, NOS|Aortic valve stenosis
C0003507|T047|IS|60573004|SNOMEDCT_CORE|AS - Aortic stenosis|Aortic valve stenosis
C0003507|T047|SY|60573004|SNOMEDCT_CORE|Stenosed aortic valve|Aortic valve stenosis
C0003510|T047|SY|359789008|SNOMEDCT_CORE|Aortitis syndrome|Aortitis syndrome
C0003534|T190|SY|24010005|SNOMEDCT_CORE|Absence of lens|Aphakia
C0003534|T190|PT|24010005|SNOMEDCT_CORE|Aphakia|Aphakia
C0003534|T190|FN|24010005|SNOMEDCT_CORE|Aphakia|Aphakia
C0003537|T048|PT|87486003|SNOMEDCT_CORE|Aphasia|Aphasia
C0003537|T048|FN|87486003|SNOMEDCT_CORE|Aphasia|Aphasia
C0003537|T048|IS|87486003|SNOMEDCT_CORE|Aphasia, NOS|Aphasia
C0003537|T048|SY|87486003|SNOMEDCT_CORE|Aphasic disturbance|Aphasia
C0003537|T048|IS|87486003|SNOMEDCT_CORE|Aphasic disturbance, NOS|Aphasia
C0003537|T048|SY|87486003|SNOMEDCT_CORE|Loss of power of expression or comprehension|Aphasia
C0003564|T184|SY|44564008|SNOMEDCT_CORE|Absence of voice|Loss of voice
C0003564|T184|IS|44564008|SNOMEDCT_CORE|Aphonia|Loss of voice
C0003564|T184|SY|44564008|SNOMEDCT_CORE|Does not phonate|Loss of voice
C0003564|T184|SY|44564008|SNOMEDCT_CORE|Does not produce voice|Loss of voice
C0003564|T184|SYGB|44564008|SNOMEDCT_CORE|Does not vocalise|Loss of voice
C0003564|T184|SY|44564008|SNOMEDCT_CORE|Does not vocalize|Loss of voice
C0003564|T184|PT|44564008|SNOMEDCT_CORE|Loss of voice|Loss of voice
C0003564|T184|FN|44564008|SNOMEDCT_CORE|Loss of voice|Loss of voice
C0003578|T184|PT|1023001|SNOMEDCT_CORE|Apnea|Apnea
C0003578|T184|FN|1023001|SNOMEDCT_CORE|Apnea|Apnea
C0003578|T184|IS|1023001|SNOMEDCT_CORE|Apnea, NOS|Apnea
C0003578|T184|SY|1023001|SNOMEDCT_CORE|Apneic|Apnea
C0003578|T184|PTGB|1023001|SNOMEDCT_CORE|Apnoea|Apnea
C0003578|T184|IS|1023001|SNOMEDCT_CORE|Apnoea, NOS|Apnea
C0003578|T184|SYGB|1023001|SNOMEDCT_CORE|Apnoeic|Apnea
C0003578|T184|SY|1023001|SNOMEDCT_CORE|Has stopped breathing|Apnea
C0003578|T184|SY|1023001|SNOMEDCT_CORE|Not breathing|Apnea
C0003615|T047|PT|74400008|SNOMEDCT_CORE|Appendicitis|Appendicitis
C0003615|T047|FN|74400008|SNOMEDCT_CORE|Appendicitis|Appendicitis
C0003615|T047|IS|74400008|SNOMEDCT_CORE|Appendicitis, NOS|Appendicitis
C0003635|T048|PT|68345001|SNOMEDCT_CORE|Apraxia|Apraxia
C0003635|T048|FN|68345001|SNOMEDCT_CORE|Apraxia|Apraxia
C0003635|T048|IS|68345001|SNOMEDCT_CORE|Apraxia, NOS|Apraxia
C0003708|T047|PT|8217007|SNOMEDCT_CORE|Arachnoiditis|Arachnoiditis
C0003708|T047|FN|8217007|SNOMEDCT_CORE|Arachnoiditis|Arachnoiditis
C0003708|T047|IS|8217007|SNOMEDCT_CORE|Arachnoiditis, NOS|Arachnoiditis
C0003794|T037|SY|127278005|SNOMEDCT_CORE|Arm injury|Injury of upper extremity
C0003794|T037|PT|127278005|SNOMEDCT_CORE|Injury of upper extremity|Injury of upper extremity
C0003794|T037|FN|127278005|SNOMEDCT_CORE|Injury of upper extremity|Injury of upper extremity
C0003794|T037|SY|127278005|SNOMEDCT_CORE|Injury of upper limb|Injury of upper extremity
C0003803|T019|SY|253184003|SNOMEDCT_CORE|Arnold-Chiari syndrome|Chiari malformation
C0003803|T019|PT|253184003|SNOMEDCT_CORE|Chiari malformation|Chiari malformation
C0003803|T019|FN|253184003|SNOMEDCT_CORE|Chiari malformation|Chiari malformation
C0003811|T047|IS|44808001|SNOMEDCT_CORE|Arrhythmia|Arrhythmia
C0003811|T047|IS|44808001|SNOMEDCT_CORE|Cardiac arrhythmia|Arrhythmia
C0003811|T047|IS|44808001|SNOMEDCT_CORE|Cardiac arrhythmias|Arrhythmia
C0003811|T047|IS|44808001|SNOMEDCT_CORE|Cardiac dysrhythmia|Arrhythmia
C0003811|T047|IS|44808001|SNOMEDCT_CORE|Cardiac dysrhythmias|Arrhythmia
C0003811|T047|IS|44808001|SNOMEDCT_CORE|Disorder of heart rhythm|Arrhythmia
C0003813|T033|SY|71792006|SNOMEDCT_CORE|Sinus arrhythmia|Sinus arrhythmia
C0003838|T047|SY|2929001|SNOMEDCT_CORE|Arterial occlusive disease|Arterial occlusive disease
C0003850|T047|PT|72092001|SNOMEDCT_CORE|Arteriosclerotic vascular disease|Arteriosclerotic vascular disease
C0003850|T047|FN|72092001|SNOMEDCT_CORE|Arteriosclerotic vascular disease|Arteriosclerotic vascular disease
C0003850|T047|IS|72092001|SNOMEDCT_CORE|Arteriosclerotic vascular disease, NOS|Arteriosclerotic vascular disease
C0003851|T047|PT|361133006|SNOMEDCT_CORE|Arteriosclerosis obliterans|Arteriosclerosis obliterans
C0003851|T047|FN|361133006|SNOMEDCT_CORE|Arteriosclerosis obliterans|Arteriosclerosis obliterans
C0003855|T190|PT|439470001|SNOMEDCT_CORE|Arteriovenous fistula|Arteriovenous fistula
C0003855|T190|FN|439470001|SNOMEDCT_CORE|Arteriovenous fistula|Arteriovenous fistula
C0003857|T019|IS|234141001|SNOMEDCT_CORE|Arteriovenous malformation|Congenital arteriovenous malformation
C0003857|T019|SY|234141001|SNOMEDCT_CORE|AV - Congenital arteriovenous anomaly|Congenital arteriovenous malformation
C0003857|T019|SY|234141001|SNOMEDCT_CORE|AV - Congenital arteriovenous malformation|Congenital arteriovenous malformation
C0003857|T019|SY|234141001|SNOMEDCT_CORE|AVM - Congenital arteriovenous malformation|Congenital arteriovenous malformation
C0003857|T019|PT|234141001|SNOMEDCT_CORE|Congenital arteriovenous malformation|Congenital arteriovenous malformation
C0003857|T019|FN|234141001|SNOMEDCT_CORE|Congenital arteriovenous malformation|Congenital arteriovenous malformation
C0003860|T046|PT|52089001|SNOMEDCT_CORE|Arteritis|Arteritis
C0003860|T046|FN|52089001|SNOMEDCT_CORE|Arteritis|Arteritis
C0003860|T046|IS|52089001|SNOMEDCT_CORE|Arteritis, NOS|Arteritis
C0003860|T046|SY|52089001|SNOMEDCT_CORE|Inflammation of artery|Arteritis
C0003862|T184|SY|57676002|SNOMEDCT_CORE|Arthralgia|Joint pain
C0003862|T184|SY|57676002|SNOMEDCT_CORE|Articular pain|Joint pain
C0003862|T184|PT|57676002|SNOMEDCT_CORE|Joint pain|Joint pain
C0003862|T184|FN|57676002|SNOMEDCT_CORE|Joint pain|Joint pain
C0003862|T184|SY|57676002|SNOMEDCT_CORE|Painful joint|Joint pain
C0003864|T047|PT|3723001|SNOMEDCT_CORE|Arthritis|Arthritis
C0003864|T047|FN|3723001|SNOMEDCT_CORE|Arthritis|Arthritis
C0003864|T047|IS|3723001|SNOMEDCT_CORE|Arthritis, NOS|Arthritis
C0003864|T047|SY|3723001|SNOMEDCT_CORE|Inflammatory arthritis|Arthritis
C0003864|T047|SY|3723001|SNOMEDCT_CORE|Joint inflammation|Arthritis
C0003868|T047|PT|190828008|SNOMEDCT_CORE|Gouty arthropathy|Gouty arthropathy
C0003868|T047|FN|190828008|SNOMEDCT_CORE|Gouty arthropathy|Gouty arthropathy
C0003869|T047|SY|396234004|SNOMEDCT_CORE|Infection-associated arthritis|Infective arthritis
C0003869|T047|PT|396234004|SNOMEDCT_CORE|Infective arthritis|Infective arthritis
C0003869|T047|FN|396234004|SNOMEDCT_CORE|Infective arthritis|Infective arthritis
C0003872|T047|IS|33339001|SNOMEDCT_CORE|PA - Psoriatic arthritis|Psoriasis with arthropathy
C0003872|T047|IS|33339001|SNOMEDCT_CORE|PsA - Psoriatic arthritis|Psoriasis with arthropathy
C0003872|T047|PT|33339001|SNOMEDCT_CORE|Psoriasis with arthropathy|Psoriasis with arthropathy
C0003872|T047|FN|33339001|SNOMEDCT_CORE|Psoriasis with arthropathy|Psoriasis with arthropathy
C0003872|T047|IS|33339001|SNOMEDCT_CORE|Psoriatic arthritis|Psoriasis with arthropathy
C0003872|T047|SY|33339001|SNOMEDCT_CORE|Psoriatic arthropathy|Psoriasis with arthropathy
C0003873|T047|SY|69896004|SNOMEDCT_CORE|Atrophic arthritis|Rheumatoid arthritis
C0003873|T047|SY|69896004|SNOMEDCT_CORE|Chronic rheumatic arthritis|Rheumatoid arthritis
C0003873|T047|SY|69896004|SNOMEDCT_CORE|RA - Rheumatoid arthritis|Rheumatoid arthritis
C0003873|T047|SY|69896004|SNOMEDCT_CORE|RhA - Rheumatoid arthritis|Rheumatoid arthritis
C0003873|T047|SY|69896004|SNOMEDCT_CORE|Rheumatic gout|Rheumatoid arthritis
C0003873|T047|PT|69896004|SNOMEDCT_CORE|Rheumatoid arthritis|Rheumatoid arthritis
C0003873|T047|FN|69896004|SNOMEDCT_CORE|Rheumatoid arthritis|Rheumatoid arthritis
C0003873|T047|SY|69896004|SNOMEDCT_CORE|Rheumatoid disease|Rheumatoid arthritis
C0003892|T047|PT|67536000|SNOMEDCT_CORE|Arthropathy associated with a neurological disorder|Arthropathy associated with a neurological disorder
C0003892|T047|FN|67536000|SNOMEDCT_CORE|Arthropathy associated with a neurological disorder|Arthropathy associated with a neurological disorder
C0003892|T047|SY|67536000|SNOMEDCT_CORE|Neuropathic arthropathy|Arthropathy associated with a neurological disorder
C0003910|T048|SY|386701004|SNOMEDCT_CORE|Articulation disorder|Articulation impairment
C0003910|T048|SY|386701004|SNOMEDCT_CORE|Articulation impairment|Articulation impairment
C0003949|T047|SY|22607003|SNOMEDCT_CORE|Amianthosis|Asbestosis
C0003949|T047|SY|22607003|SNOMEDCT_CORE|Asbestos pneumoconiosis|Asbestosis
C0003949|T047|PT|22607003|SNOMEDCT_CORE|Asbestosis|Asbestosis
C0003949|T047|FN|22607003|SNOMEDCT_CORE|Asbestosis|Asbestosis
C0003949|T047|SY|22607003|SNOMEDCT_CORE|Pulmonary asbestosis|Asbestosis
C0003962|T047|IS|389026000|SNOMEDCT_CORE|Abdominal dropsy|Ascites
C0003962|T047|PT|389026000|SNOMEDCT_CORE|Ascites|Ascites
C0003962|T047|FN|389026000|SNOMEDCT_CORE|Ascites|Ascites
C0003962|T047|SY|389026000|SNOMEDCT_CORE|Hydroperitoneum|Ascites
C0003962|T047|SY|389026000|SNOMEDCT_CORE|Hydroperitonia|Ascites
C0003962|T047|SY|389026000|SNOMEDCT_CORE|Hydrops abdominis|Ascites
C0003962|T047|IS|389026000|SNOMEDCT_CORE|Peritoneal dropsy|Ascites
C0003977|T047|IS|29281007|SNOMEDCT_CORE|Aseptic necrosis of head and neck of femur|Aseptic necrosis of head AND/OR neck of femur
C0003977|T047|PT|29281007|SNOMEDCT_CORE|Aseptic necrosis of head AND/OR neck of femur|Aseptic necrosis of head AND/OR neck of femur
C0003977|T047|FN|29281007|SNOMEDCT_CORE|Aseptic necrosis of head AND/OR neck of femur|Aseptic necrosis of head AND/OR neck of femur
C0004030|T047|PT|65553006|SNOMEDCT_CORE|Aspergillosis|Aspergillosis
C0004030|T047|FN|65553006|SNOMEDCT_CORE|Aspergillosis|Aspergillosis
C0004030|T047|IS|65553006|SNOMEDCT_CORE|Aspergillosis, NOS|Aspergillosis
C0004030|T047|SY|65553006|SNOMEDCT_CORE|Infection due to Aspergillus|Aspergillosis
C0004063|T037|PT|52684005|SNOMEDCT_CORE|Assault|Assault
C0004063|T037|IS|52684005|SNOMEDCT_CORE|Assault|Assault
C0004063|T037|OF|52684005|SNOMEDCT_CORE|Assault|Assault
C0004063|T037|FN|52684005|SNOMEDCT_CORE|Assault|Assault
C0004063|T037|IS|52684005|SNOMEDCT_CORE|Attacked|Assault
C0004063|T037|IS|52684005|SNOMEDCT_CORE|Mugged|Assault
C0004093|T184|PT|13791008|SNOMEDCT_CORE|Asthenia|Asthenia
C0004093|T184|FN|13791008|SNOMEDCT_CORE|Asthenia|Asthenia
C0004096|T047|SY|195967001|SNOMEDCT_CORE|Airway hyperreactivity|Asthma
C0004096|T047|PT|195967001|SNOMEDCT_CORE|Asthma|Asthma
C0004096|T047|FN|195967001|SNOMEDCT_CORE|Asthma|Asthma
C0004096|T047|SY|195967001|SNOMEDCT_CORE|Asthmatic|Asthma
C0004096|T047|SY|195967001|SNOMEDCT_CORE|Bronchial asthma|Asthma
C0004099|T047|SY|31387002|SNOMEDCT_CORE|EIA - Exercise-induced asthma|Exercise-induced asthma
C0004099|T047|SY|31387002|SNOMEDCT_CORE|Exercise induced asthma|Exercise-induced asthma
C0004099|T047|PT|31387002|SNOMEDCT_CORE|Exercise-induced asthma|Exercise-induced asthma
C0004099|T047|FN|31387002|SNOMEDCT_CORE|Exercise-induced asthma|Exercise-induced asthma
C0004106|T047|PT|82649003|SNOMEDCT_CORE|Astigmatism|Astigmatism
C0004106|T047|FN|82649003|SNOMEDCT_CORE|Astigmatism|Astigmatism
C0004106|T047|IS|82649003|SNOMEDCT_CORE|Astigmatism, NOS|Astigmatism
C0004134|T184|PT|20262006|SNOMEDCT_CORE|Ataxia|Ataxia
C0004134|T184|FN|20262006|SNOMEDCT_CORE|Ataxia|Ataxia
C0004134|T184|IS|20262006|SNOMEDCT_CORE|Ataxia, NOS|Ataxia
C0004144|T046|PT|46621007|SNOMEDCT_CORE|Atelectasis|Atelectasis
C0004144|T046|FN|46621007|SNOMEDCT_CORE|Atelectasis|Atelectasis
C0004144|T046|IS|46621007|SNOMEDCT_CORE|Atelectasis, NOS|Atelectasis
C0004144|T046|SY|46621007|SNOMEDCT_CORE|Collapse of lung|Atelectasis
C0004144|T046|SY|46621007|SNOMEDCT_CORE|Pulmonary atelectasis|Atelectasis
C0004144|T046|SY|46621007|SNOMEDCT_CORE|Pulmonary collapse|Atelectasis
C0004144|T046|SY|46621007|SNOMEDCT_CORE|Pulmonary collapse with atelectasis|Atelectasis
C0004153|T047|SY|38716007|SNOMEDCT_CORE|Atheromatosis|Atherosclerosis
C0004153|T047|IS|38716007|SNOMEDCT_CORE|Atheromatosis, NOS|Atherosclerosis
C0004153|T047|PT|38716007|SNOMEDCT_CORE|Atherosclerosis|Atherosclerosis
C0004153|T047|FN|38716007|SNOMEDCT_CORE|Atherosclerosis|Atherosclerosis
C0004153|T047|IS|38716007|SNOMEDCT_CORE|Atherosclerosis, NOS|Atherosclerosis
C0004161|T037|OAP|23294000|SNOMEDCT_CORE|Sports injury|Sports injury
C0004161|T037|OAF|23294000|SNOMEDCT_CORE|Sports injury|Sports injury
C0004161|T037|IS|23294000|SNOMEDCT_CORE|Sports injury, NOS|Sports injury, NOS
C0004238|T047|SY|49436004|SNOMEDCT_CORE|AF - Atrial fibrillation|Atrial fibrillation
C0004238|T047|PT|49436004|SNOMEDCT_CORE|Atrial fibrillation|Atrial fibrillation
C0004238|T047|FN|49436004|SNOMEDCT_CORE|Atrial fibrillation|Atrial fibrillation
C0004239|T046|PT|5370000|SNOMEDCT_CORE|Atrial flutter|Atrial flutter
C0004239|T046|FN|5370000|SNOMEDCT_CORE|Atrial flutter|Atrial flutter
C0004245|T047|PT|233917008|SNOMEDCT_CORE|Atrioventricular block|Atrioventricular block
C0004245|T047|FN|233917008|SNOMEDCT_CORE|Atrioventricular block|Atrioventricular block
C0004245|T047|SY|233917008|SNOMEDCT_CORE|AV block|Atrioventricular block
C0004245|T047|SY|233917008|SNOMEDCT_CORE|AVB - Atrioventricular block|Atrioventricular block
C0004269|T047|PT|192127007|SNOMEDCT_CORE|Child attention deficit disorder|Child attention deficit disorder
C0004269|T047|FN|192127007|SNOMEDCT_CORE|Child attention deficit disorder|Child attention deficit disorder
C0004352|T048|SY|408856003|SNOMEDCT_CORE|Autism|Autistic disorder
C0004352|T048|SY|408856003|SNOMEDCT_CORE|Autism disorder|Autistic disorder
C0004352|T048|PT|408856003|SNOMEDCT_CORE|Autistic disorder|Autistic disorder
C0004352|T048|FN|408856003|SNOMEDCT_CORE|Autistic disorder|Autistic disorder
C0004352|T048|SY|408856003|SNOMEDCT_CORE|Kanner's syndrome|Autistic disorder
C0004364|T047|PT|85828009|SNOMEDCT_CORE|Autoimmune disease|Autoimmune disease
C0004364|T047|FN|85828009|SNOMEDCT_CORE|Autoimmune disease|Autoimmune disease
C0004364|T047|IS|85828009|SNOMEDCT_CORE|Autoimmune disease, NOS|Autoimmune disease
C0004364|T047|SY|85828009|SNOMEDCT_CORE|Autoimmune disorder|Autoimmune disease
C0004364|T047|IS|85828009|SNOMEDCT_CORE|Autoimmune disorder, NOS|Autoimmune disease
C0004444|T048|PT|37746008|SNOMEDCT_CORE|Avoidant personality disorder|Avoidant personality disorder
C0004444|T048|FN|37746008|SNOMEDCT_CORE|Avoidant personality disorder|Avoidant personality disorder
C0004601|T037|OAS|81102000|SNOMEDCT_CORE|Back injury|Traumatic and/or non-traumatic injury of back
C0004601|T037|OAP|81102000|SNOMEDCT_CORE|Injury of back|Traumatic and/or non-traumatic injury of back
C0004601|T037|OAF|81102000|SNOMEDCT_CORE|Injury of back|Traumatic and/or non-traumatic injury of back
C0004601|T037|PT|712893003|SNOMEDCT_CORE|Traumatic and/or non-traumatic injury of back|Traumatic and/or non-traumatic injury of back
C0004601|T037|FN|712893003|SNOMEDCT_CORE|Traumatic and/or non-traumatic injury of back|Traumatic and/or non-traumatic injury of back
C0004604|T184|SY|161891005|SNOMEDCT_CORE|Back ache|Backache
C0004604|T184|SY|161891005|SNOMEDCT_CORE|Back pain|Backache
C0004604|T184|OF|161891005|SNOMEDCT_CORE|Backache|Backache
C0004604|T184|PT|161891005|SNOMEDCT_CORE|Backache|Backache
C0004604|T184|FN|161891005|SNOMEDCT_CORE|Backache|Backache
C0004604|T184|SY|161891005|SNOMEDCT_CORE|Pain in back|Backache
C0004606|T047|SY|390834004|SNOMEDCT_CORE|Background diabetic retinopathy|Nonproliferative retinopathy due to diabetes mellitus
C0004606|T047|SY|390834004|SNOMEDCT_CORE|BDR - Background diabetic retinopathy|Nonproliferative retinopathy due to diabetes mellitus
C0004606|T047|SY|390834004|SNOMEDCT_CORE|Non proliferative diabetic retinopathy|Nonproliferative retinopathy due to diabetes mellitus
C0004606|T047|OF|390834004|SNOMEDCT_CORE|Non proliferative diabetic retinopathy|Nonproliferative retinopathy due to diabetes mellitus
C0004606|T047|SY|390834004|SNOMEDCT_CORE|Nonproliferative diabetic retinopathy|Nonproliferative retinopathy due to diabetes mellitus
C0004606|T047|OF|390834004|SNOMEDCT_CORE|Nonproliferative diabetic retinopathy|Nonproliferative retinopathy due to diabetes mellitus
C0004606|T047|IS|390834004|SNOMEDCT_CORE|Nonproliferative retinopathy co-occurrent and due to diabetes mellitus|Nonproliferative retinopathy due to diabetes mellitus
C0004606|T047|OF|390834004|SNOMEDCT_CORE|Nonproliferative retinopathy co-occurrent and due to diabetes mellitus|Nonproliferative retinopathy due to diabetes mellitus
C0004606|T047|PT|390834004|SNOMEDCT_CORE|Nonproliferative retinopathy due to diabetes mellitus|Nonproliferative retinopathy due to diabetes mellitus
C0004606|T047|FN|390834004|SNOMEDCT_CORE|Nonproliferative retinopathy due to diabetes mellitus|Nonproliferative retinopathy due to diabetes mellitus
C0004606|T047|SY|390834004|SNOMEDCT_CORE|NPDR - Non proliferative diabetic retinopathy|Nonproliferative retinopathy due to diabetes mellitus
C0004610|T047|PTGB|5758002|SNOMEDCT_CORE|Bacteraemia|Bacteremia
C0004610|T047|PT|5758002|SNOMEDCT_CORE|Bacteremia|Bacteremia
C0004610|T047|OF|5758002|SNOMEDCT_CORE|Bacteremia|Bacteremia
C0004610|T047|FN|5758002|SNOMEDCT_CORE|Bacteremia|Bacteremia
C0004610|T047|IS|5758002|SNOMEDCT_CORE|Bacteremia, NOS|Bacteremia
C0004623|T047|SY|87628006|SNOMEDCT_CORE|Bacterial disease|Bacterial infectious disease
C0004623|T047|SY|87628006|SNOMEDCT_CORE|Bacterial infection|Bacterial infectious disease
C0004623|T047|IS|87628006|SNOMEDCT_CORE|Bacterial infection, NOS|Bacterial infectious disease
C0004623|T047|PT|87628006|SNOMEDCT_CORE|Bacterial infectious disease|Bacterial infectious disease
C0004623|T047|FN|87628006|SNOMEDCT_CORE|Bacterial infectious disease|Bacterial infectious disease
C0004623|T047|IS|87628006|SNOMEDCT_CORE|Bacterial infectious disease, NOS|Bacterial infectious disease
C0004623|T047|SY|87628006|SNOMEDCT_CORE|Disease caused by bacteria|Bacterial infectious disease
C0004623|T047|IS|87628006|SNOMEDCT_CORE|Disease caused by bacteria, NOS|Bacterial infectious disease
C0004626|T047|PT|53084003|SNOMEDCT_CORE|Bacterial pneumonia|Bacterial pneumonia
C0004626|T047|FN|53084003|SNOMEDCT_CORE|Bacterial pneumonia|Bacterial pneumonia
C0004626|T047|IS|53084003|SNOMEDCT_CORE|Bacterial pneumonia, NOS|Bacterial pneumonia
C0004690|T047|PT|44882003|SNOMEDCT_CORE|Balanitis|Balanitis
C0004690|T047|FN|44882003|SNOMEDCT_CORE|Balanitis|Balanitis
C0004763|T047|SY|302914006|SNOMEDCT_CORE|Barrett esophagus|Barrett's esophagus
C0004763|T047|PT|302914006|SNOMEDCT_CORE|Barrett's esophagus|Barrett's esophagus
C0004763|T047|FN|302914006|SNOMEDCT_CORE|Barrett's esophagus|Barrett's esophagus
C0004763|T047|PTGB|302914006|SNOMEDCT_CORE|Barrett's oesophagus|Barrett's esophagus
C0004763|T047|SY|302914006|SNOMEDCT_CORE|Barrett's syndrome|Barrett's esophagus
C0004763|T047|SY|302914006|SNOMEDCT_CORE|Barretts esophagus|Barrett's esophagus
C0004763|T047|IS|302914006|SNOMEDCT_CORE|BO - Barrett's esophagus|Barrett's esophagus
C0004763|T047|SYGB|302914006|SNOMEDCT_CORE|BO - Barrett's oesophagus|Barrett's esophagus
C0004763|T047|SY|302914006|SNOMEDCT_CORE|CELLO - Columnar epithelial-lined lower esophagus|Barrett's esophagus
C0004763|T047|SYGB|302914006|SNOMEDCT_CORE|CELLO - Columnar epithelial-lined lower oesophagus|Barrett's esophagus
C0004763|T047|SY|302914006|SNOMEDCT_CORE|CLE - Columnar-lined esophagus|Barrett's esophagus
C0004763|T047|SYGB|302914006|SNOMEDCT_CORE|CLE - Columnar-lined oesophagus|Barrett's esophagus
C0004763|T047|SY|302914006|SNOMEDCT_CORE|Columnar epithelial-lined lower esophagus|Barrett's esophagus
C0004763|T047|SYGB|302914006|SNOMEDCT_CORE|Columnar epithelial-lined lower oesophagus|Barrett's esophagus
C0004763|T047|SY|302914006|SNOMEDCT_CORE|Columnar-lined esophagus|Barrett's esophagus
C0004763|T047|SYGB|302914006|SNOMEDCT_CORE|Columnar-lined oesophagus|Barrett's esophagus
C0004763|T047|SY|302914006|SNOMEDCT_CORE|Gastric metaplasia of esophagus|Barrett's esophagus
C0004763|T047|SYGB|302914006|SNOMEDCT_CORE|Gastric metaplasia of oesophagus|Barrett's esophagus
C0004766|T046|SY|67624004|SNOMEDCT_CORE|Abscess of Bartholin gland|Abscess of Bartholin's gland
C0004766|T046|PT|67624004|SNOMEDCT_CORE|Abscess of Bartholin's gland|Abscess of Bartholin's gland
C0004766|T046|FN|67624004|SNOMEDCT_CORE|Abscess of Bartholin's gland|Abscess of Bartholin's gland
C0004766|T046|SY|67624004|SNOMEDCT_CORE|Bartholin's abscess|Abscess of Bartholin's gland
C0004766|T046|SY|67624004|SNOMEDCT_CORE|Vulvovaginal gland abscess|Abscess of Bartholin's gland
C0004767|T047|SY|57044006|SNOMEDCT_CORE|Bartholin's cyst|Cyst of Bartholin's gland duct
C0004767|T047|IS|57044006|SNOMEDCT_CORE|Bartholin's duct cyst|Cyst of Bartholin's gland duct
C0004767|T047|SY|57044006|SNOMEDCT_CORE|Bartholin's gland cyst|Cyst of Bartholin's gland duct
C0004767|T047|SY|57044006|SNOMEDCT_CORE|Bartholin's gland duct cyst|Cyst of Bartholin's gland duct
C0004767|T047|SY|57044006|SNOMEDCT_CORE|Cyst of Bartholin gland duct|Cyst of Bartholin's gland duct
C0004767|T047|IS|57044006|SNOMEDCT_CORE|Cyst of Bartholin's duct|Cyst of Bartholin's gland duct
C0004767|T047|SY|57044006|SNOMEDCT_CORE|Cyst of Bartholin's gland|Cyst of Bartholin's gland duct
C0004767|T047|PT|57044006|SNOMEDCT_CORE|Cyst of Bartholin's gland duct|Cyst of Bartholin's gland duct
C0004767|T047|FN|57044006|SNOMEDCT_CORE|Cyst of Bartholin's gland duct|Cyst of Bartholin's gland duct
C0004812|T047|PT|64009001|SNOMEDCT_CORE|Basilar artery syndrome|Basilar artery syndrome
C0004812|T047|FN|64009001|SNOMEDCT_CORE|Basilar artery syndrome|Basilar artery syndrome
C0004812|T047|SY|64009001|SNOMEDCT_CORE|Insufficiency - basilar artery|Basilar artery syndrome
C0004936|T048|SY|74732009|SNOMEDCT_CORE|Mental disease|Mental disorder
C0004936|T048|PT|74732009|SNOMEDCT_CORE|Mental disorder|Mental disorder
C0004936|T048|FN|74732009|SNOMEDCT_CORE|Mental disorder|Mental disorder
C0004936|T048|IS|74732009|SNOMEDCT_CORE|Mental disorder, NOS|Mental disorder
C0004936|T048|SY|74732009|SNOMEDCT_CORE|Mental health disorder|Mental disorder
C0004936|T048|SY|74732009|SNOMEDCT_CORE|Mental illness|Mental disorder
C0004936|T048|SY|74732009|SNOMEDCT_CORE|Psychiatric disorder|Mental disorder
C0004936|T048|SY|74732009|SNOMEDCT_CORE|Psychiatric illness|Mental disorder
C0004943|T047|SY|310701003|SNOMEDCT_CORE|Adamantiades-Behcet disease|Behcet's syndrome
C0004943|T047|OF|310701003|SNOMEDCT_CORE|Beh?et's syndrome|Behcet's syndrome
C0004943|T047|IS|310701003|SNOMEDCT_CORE|Beh?et's syndrome|Behcet's syndrome
C0004943|T047|SY|310701003|SNOMEDCT_CORE|Behcet syndrome|Behcet's syndrome
C0004943|T047|SY|310701003|SNOMEDCT_CORE|Behcet's disease|Behcet's syndrome
C0004943|T047|PT|310701003|SNOMEDCT_CORE|Behcet's syndrome|Behcet's syndrome
C0004943|T047|FN|310701003|SNOMEDCT_CORE|Behcet's syndrome|Behcet's syndrome
C0004991|T191|PT|92065004|SNOMEDCT_CORE|Benign neoplasm of colon|Benign neoplasm of colon
C0004991|T191|FN|92065004|SNOMEDCT_CORE|Benign neoplasm of colon|Benign neoplasm of colon
C0004991|T191|IS|92065004|SNOMEDCT_CORE|Benign neoplasm of colon, NOS|Benign neoplasm of colon
C0004991|T191|SY|92065004|SNOMEDCT_CORE|Benign tumor of colon|Benign neoplasm of colon
C0004991|T191|SYGB|92065004|SNOMEDCT_CORE|Benign tumour of colon|Benign neoplasm of colon
C0004992|T191|PT|92071005|SNOMEDCT_CORE|Benign neoplasm of cranial nerve|Benign neoplasm of cranial nerve
C0004992|T191|FN|92071005|SNOMEDCT_CORE|Benign neoplasm of cranial nerve|Benign neoplasm of cranial nerve
C0004992|T191|IS|92071005|SNOMEDCT_CORE|Benign neoplasm of cranial nerve, NOS|Benign neoplasm of cranial nerve
C0004997|T191|PT|92260003|SNOMEDCT_CORE|Benign neoplasm of ovary|Benign neoplasm of ovary
C0004997|T191|FN|92260003|SNOMEDCT_CORE|Benign neoplasm of ovary|Benign neoplasm of ovary
C0004997|T191|SY|92260003|SNOMEDCT_CORE|Benign ovarian tumor|Benign neoplasm of ovary
C0004997|T191|SYGB|92260003|SNOMEDCT_CORE|Benign ovarian tumour|Benign neoplasm of ovary
C0004998|T191|PT|92384009|SNOMEDCT_CORE|Benign neoplasm of skin|Benign neoplasm of skin
C0004998|T191|FN|92384009|SNOMEDCT_CORE|Benign neoplasm of skin|Benign neoplasm of skin
C0004998|T191|IS|92384009|SNOMEDCT_CORE|Benign neoplasm of skin, NOS|Benign neoplasm of skin
C0004998|T191|SY|92384009|SNOMEDCT_CORE|Benign tumor of skin|Benign neoplasm of skin
C0004998|T191|SYGB|92384009|SNOMEDCT_CORE|Benign tumour of skin|Benign neoplasm of skin
C0005001|T046|SY|266569009|SNOMEDCT_CORE|Benign enlargement of prostate|Benign prostatic hypertrophy
C0005001|T046|SY|266569009|SNOMEDCT_CORE|Benign prostatic hypertrophy|Benign prostatic hypertrophy
C0005001|T046|SY|266569009|SNOMEDCT_CORE|BEP - Benign enlargement of prostate|Benign prostatic hypertrophy
C0005001|T046|IS|266569009|SNOMEDCT_CORE|BPH|Benign prostatic hypertrophy
C0005001|T046|IS|266569009|SNOMEDCT_CORE|BPH - Benign prostatic hypertrophy|Benign prostatic hypertrophy
C0005136|T046|PT|277196008|SNOMEDCT_CORE|Berry aneurysm|Berry aneurysm
C0005136|T046|FN|277196008|SNOMEDCT_CORE|Berry aneurysm|Berry aneurysm
C0005136|T046|IS|277196008|SNOMEDCT_CORE|Berry aneurysm - disorder|Berry aneurysm
C0005136|T046|SY|277196008|SNOMEDCT_CORE|Berry aneurysm disorder|Berry aneurysm
C0005136|T046|SY|277196008|SNOMEDCT_CORE|Saccular aneurysm|Berry aneurysm
C0005283|T047|PTGB|65959000|SNOMEDCT_CORE|Beta thalassaemia|Beta thalassemia
C0005283|T047|SYGB|65959000|SNOMEDCT_CORE|beta thalassaemia|Beta thalassemia
C0005283|T047|OP|65959000|SNOMEDCT_CORE|beta Thalassaemia|Beta thalassemia
C0005283|T047|SYGB|65959000|SNOMEDCT_CORE|Beta thalassaemia syndrome|Beta thalassemia
C0005283|T047|OP|65959000|SNOMEDCT_CORE|beta Thalassemia|Beta thalassemia
C0005283|T047|PT|65959000|SNOMEDCT_CORE|Beta thalassemia|Beta thalassemia
C0005283|T047|SY|65959000|SNOMEDCT_CORE|beta thalassemia|Beta thalassemia
C0005283|T047|FN|65959000|SNOMEDCT_CORE|Beta thalassemia|Beta thalassemia
C0005283|T047|OF|65959000|SNOMEDCT_CORE|beta Thalassemia|Beta thalassemia
C0005283|T047|SY|65959000|SNOMEDCT_CORE|Beta thalassemia syndrome|Beta thalassemia
C0005283|T047|IS|65959000|SNOMEDCT_CORE|beta Thalassemia, NOS|Beta thalassemia
C0005411|T019|SY|77480004|SNOMEDCT_CORE|Atresia of bile ducts|Congenital biliary atresia
C0005411|T019|SY|77480004|SNOMEDCT_CORE|BA - Biliary atresia|Congenital biliary atresia
C0005411|T019|SY|77480004|SNOMEDCT_CORE|Biliary atresia|Congenital biliary atresia
C0005411|T019|PT|77480004|SNOMEDCT_CORE|Congenital biliary atresia|Congenital biliary atresia
C0005411|T019|FN|77480004|SNOMEDCT_CORE|Congenital biliary atresia|Congenital biliary atresia
C0005416|T047|PT|197432008|SNOMEDCT_CORE|Biliary dyskinesia|Biliary dyskinesia
C0005416|T047|FN|197432008|SNOMEDCT_CORE|Biliary dyskinesia|Biliary dyskinesia
C0005424|T047|SY|105997008|SNOMEDCT_CORE|Disease of biliary system|Disorder of biliary tract
C0005424|T047|IS|105997008|SNOMEDCT_CORE|Disease of biliary tract|Disorder of biliary tract
C0005424|T047|OF|105997008|SNOMEDCT_CORE|Disease of biliary tract|Disorder of biliary tract
C0005424|T047|PT|105997008|SNOMEDCT_CORE|Disorder of biliary tract|Disorder of biliary tract
C0005424|T047|FN|105997008|SNOMEDCT_CORE|Disorder of biliary tract|Disorder of biliary tract
C0005586|T048|SY|13746004|SNOMEDCT_CORE|Bipolar affective disorder|Bipolar disorder
C0005586|T048|PT|13746004|SNOMEDCT_CORE|Bipolar disorder|Bipolar disorder
C0005586|T048|FN|13746004|SNOMEDCT_CORE|Bipolar disorder|Bipolar disorder
C0005586|T048|IS|13746004|SNOMEDCT_CORE|Bipolar disorder, NOS|Bipolar disorder
C0005586|T048|SY|13746004|SNOMEDCT_CORE|Manic-depressive illness|Bipolar disorder
C0005586|T048|SY|13746004|SNOMEDCT_CORE|Manic-depressive psychosis|Bipolar disorder
C0005586|T048|SY|13746004|SNOMEDCT_CORE|MDI - Manic-depressive illness|Bipolar disorder
C0005587|T048|PT|191627008|SNOMEDCT_CORE|Bipolar affective disorder, current episode depression|Bipolar affective disorder, current episode depression
C0005587|T048|FN|191627008|SNOMEDCT_CORE|Bipolar affective disorder, current episode depression|Bipolar affective disorder, current episode depression
C0005587|T048|SY|191627008|SNOMEDCT_CORE|Manic-depressive - now depressed|Bipolar affective disorder, current episode depression
C0005683|T047|SY|70650003|SNOMEDCT_CORE|Bladder calculus|Urinary bladder stone
C0005683|T047|SY|70650003|SNOMEDCT_CORE|Bladder stone|Urinary bladder stone
C0005683|T047|SY|70650003|SNOMEDCT_CORE|Calculus of bladder|Urinary bladder stone
C0005683|T047|PT|70650003|SNOMEDCT_CORE|Urinary bladder stone|Urinary bladder stone
C0005683|T047|FN|70650003|SNOMEDCT_CORE|Urinary bladder stone|Urinary bladder stone
C0005683|T047|SY|70650003|SNOMEDCT_CORE|Vesical calculus|Urinary bladder stone
C0005683|T047|SY|70650003|SNOMEDCT_CORE|Vesicolithiasis|Urinary bladder stone
C0005684|T191|SY|399326009|SNOMEDCT_CORE|Bladder cancer|Malignant tumor of urinary bladder
C0005684|T191|SY|399326009|SNOMEDCT_CORE|CA - Bladder cancer|Malignant tumor of urinary bladder
C0005684|T191|SY|399326009|SNOMEDCT_CORE|Malignant neoplasm of urinary bladder|Malignant tumor of urinary bladder
C0005684|T191|PT|399326009|SNOMEDCT_CORE|Malignant tumor of urinary bladder|Malignant tumor of urinary bladder
C0005684|T191|FN|399326009|SNOMEDCT_CORE|Malignant tumor of urinary bladder|Malignant tumor of urinary bladder
C0005684|T191|PTGB|399326009|SNOMEDCT_CORE|Malignant tumour of urinary bladder|Malignant tumor of urinary bladder
C0005686|T047|IS|42643001|SNOMEDCT_CORE|Disease of bladder|Disorder of bladder
C0005686|T047|OF|42643001|SNOMEDCT_CORE|Disease of bladder|Disorder of bladder
C0005686|T047|IS|42643001|SNOMEDCT_CORE|Disease of bladder, NOS|Disorder of bladder
C0005686|T047|PT|42643001|SNOMEDCT_CORE|Disorder of bladder|Disorder of bladder
C0005686|T047|SY|42643001|SNOMEDCT_CORE|Disorder of bladder and bladder neck|Disorder of bladder
C0005686|T047|IS|42643001|SNOMEDCT_CORE|Disorder of bladder, NOS|Disorder of bladder
C0005686|T047|SY|42643001|SNOMEDCT_CORE|Disorder of urinary bladder|Disorder of bladder
C0005686|T047|FN|42643001|SNOMEDCT_CORE|Disorder of urinary bladder|Disorder of bladder
C0005694|T047|PT|399072004|SNOMEDCT_CORE|Bladder neck obstruction|Bladder neck obstruction
C0005694|T047|FN|399072004|SNOMEDCT_CORE|Bladder neck obstruction|Bladder neck obstruction
C0005694|T047|SY|399072004|SNOMEDCT_CORE|BNO - Bladder neck obstruction|Bladder neck obstruction
C0005694|T047|SY|399072004|SNOMEDCT_CORE|Vesicourethral orifice obstruction|Bladder neck obstruction
C0005695|T191|PT|126885006|SNOMEDCT_CORE|Neoplasm of bladder|Neoplasm of bladder
C0005695|T191|FN|126885006|SNOMEDCT_CORE|Neoplasm of bladder|Neoplasm of bladder
C0005695|T191|SY|126885006|SNOMEDCT_CORE|NGB - New growth of bladder|Neoplasm of bladder
C0005695|T191|SY|126885006|SNOMEDCT_CORE|Tumor of urinary bladder|Neoplasm of bladder
C0005695|T191|SYGB|126885006|SNOMEDCT_CORE|Tumour of urinary bladder|Neoplasm of bladder
C0005697|T047|PT|398064005|SNOMEDCT_CORE|Neurogenic bladder|Neurogenic bladder
C0005697|T047|FN|398064005|SNOMEDCT_CORE|Neurogenic bladder|Neurogenic bladder
C0005697|T047|SY|398064005|SNOMEDCT_CORE|Neuropathic bladder|Neurogenic bladder
C0005741|T047|PT|41446000|SNOMEDCT_CORE|Blepharitis|Blepharitis
C0005741|T047|FN|41446000|SNOMEDCT_CORE|Blepharitis|Blepharitis
C0005741|T047|IS|41446000|SNOMEDCT_CORE|Blepharitis, NOS|Blepharitis
C0005741|T047|SY|41446000|SNOMEDCT_CORE|Eyelid inflammation|Blepharitis
C0005741|T047|SY|41446000|SNOMEDCT_CORE|Inflammation of eyelid|Blepharitis
C0005741|T047|IS|41446000|SNOMEDCT_CORE|Inflammation of eyelid, NOS|Blepharitis
C0005745|T047|SY|11934000|SNOMEDCT_CORE|Blepharoptosis|Ptosis of eyelid
C0005745|T047|SY|11934000|SNOMEDCT_CORE|Drooping eyelid|Ptosis of eyelid
C0005745|T047|SY|11934000|SNOMEDCT_CORE|Droopy eyelid|Ptosis of eyelid
C0005745|T047|SY|11934000|SNOMEDCT_CORE|Ptosis|Ptosis of eyelid
C0005745|T047|SY|11934000|SNOMEDCT_CORE|Ptosis eyelid|Ptosis of eyelid
C0005745|T047|PT|11934000|SNOMEDCT_CORE|Ptosis of eyelid|Ptosis of eyelid
C0005745|T047|FN|11934000|SNOMEDCT_CORE|Ptosis of eyelid|Ptosis of eyelid
C0005745|T047|IS|11934000|SNOMEDCT_CORE|Ptosis of eyelid, NOS|Ptosis of eyelid
C0005747|T047|PT|59026006|SNOMEDCT_CORE|Blepharospasm|Blepharospasm
C0005747|T047|SY|59026006|SNOMEDCT_CORE|Blepharospasm|Blepharospasm
C0005747|T047|FN|59026006|SNOMEDCT_CORE|Blepharospasm|Blepharospasm
C0005747|T047|SY|59026006|SNOMEDCT_CORE|Spasm of eyelids|Blepharospasm
C0005750|T047|PT|66379009|SNOMEDCT_CORE|Bacterial overgrowth syndrome|Blind loop syndrome
C0005750|T047|FN|66379009|SNOMEDCT_CORE|Bacterial overgrowth syndrome|Blind loop syndrome
C0005750|T047|PT|77225009|SNOMEDCT_CORE|Blind loop syndrome|Blind loop syndrome
C0005750|T047|FN|77225009|SNOMEDCT_CORE|Blind loop syndrome|Blind loop syndrome
C0005750|T047|IS|77225009|SNOMEDCT_CORE|Blind loop syndrome, NOS|Blind loop syndrome
C0005750|T047|SY|77225009|SNOMEDCT_CORE|Contaminated small bowel syndrome|Blind loop syndrome
C0005750|T047|SY|77225009|SNOMEDCT_CORE|Stagnant loop syndrome|Blind loop syndrome
C0005779|T047|SY|64779008|SNOMEDCT_CORE|Blood clotting disorder|Blood coagulation disorder
C0005779|T047|IS|64779008|SNOMEDCT_CORE|Blood clotting disorder, NOS|Blood coagulation disorder
C0005779|T047|PT|64779008|SNOMEDCT_CORE|Blood coagulation disorder|Blood coagulation disorder
C0005779|T047|FN|64779008|SNOMEDCT_CORE|Blood coagulation disorder|Blood coagulation disorder
C0005779|T047|IS|64779008|SNOMEDCT_CORE|Blood coagulation disorder, NOS|Blood coagulation disorder
C0005779|T047|SY|64779008|SNOMEDCT_CORE|Clotting disorder|Blood coagulation disorder
C0005779|T047|SY|64779008|SNOMEDCT_CORE|Coagulation disorder|Blood coagulation disorder
C0005779|T047|IS|64779008|SNOMEDCT_CORE|Coagulation disorder, NOS|Blood coagulation disorder
C0005779|T047|SY|64779008|SNOMEDCT_CORE|Coagulopathy|Blood coagulation disorder
C0005779|T047|IS|64779008|SNOMEDCT_CORE|Coagulopathy, NOS|Blood coagulation disorder
C0005779|T047|SYGB|64779008|SNOMEDCT_CORE|Disorder of haemostasis|Blood coagulation disorder
C0005779|T047|IS|64779008|SNOMEDCT_CORE|Disorder of haemostasis, NOS|Blood coagulation disorder
C0005779|T047|SY|64779008|SNOMEDCT_CORE|Disorder of hemostasis|Blood coagulation disorder
C0005779|T047|IS|64779008|SNOMEDCT_CORE|Disorder of hemostasis, NOS|Blood coagulation disorder
C0005818|T047|PT|22716005|SNOMEDCT_CORE|Platelet disorder|Platelet disorder
C0005818|T047|FN|22716005|SNOMEDCT_CORE|Platelet disorder|Platelet disorder
C0005818|T047|IS|22716005|SNOMEDCT_CORE|Platelet disorder, NOS|Platelet disorder
C0005818|T047|SY|22716005|SNOMEDCT_CORE|Thrombocytopathy|Platelet disorder
C0005818|T047|IS|22716005|SNOMEDCT_CORE|Thrombocytopathy, NOS|Platelet disorder
C0005826|T033|PT|38936003|SNOMEDCT_CORE|Abnormal blood pressure|Abnormal blood pressure
C0005826|T033|FN|38936003|SNOMEDCT_CORE|Abnormal blood pressure|Abnormal blood pressure
C0005826|T033|IS|38936003|SNOMEDCT_CORE|Abnormal blood pressure, NOS|Abnormal blood pressure
C0005858|T184|OAP|73009009|SNOMEDCT_CORE|Bloodshot eye|Bloodshot eye
C0005858|T184|OAS|246676003|SNOMEDCT_CORE|Bloodshot eye|Bloodshot eye
C0005858|T184|OAF|73009009|SNOMEDCT_CORE|Bloodshot eye|Bloodshot eye
C0005858|T184|IS|73009009|SNOMEDCT_CORE|Bloodshot eyes|Bloodshot eye
C0005858|T184|OAS|73009009|SNOMEDCT_CORE|Red eye|Bloodshot eye
C0005937|T190|PT|203465002|SNOMEDCT_CORE|Bone cyst|Bone cyst
C0005937|T190|FN|203465002|SNOMEDCT_CORE|Bone cyst|Bone cyst
C0005940|T047|SY|76069003|SNOMEDCT_CORE|Bone disease|Disorder of bone
C0005940|T047|IS|76069003|SNOMEDCT_CORE|Bone disease, NOS|Disorder of bone
C0005940|T047|IS|76069003|SNOMEDCT_CORE|Disease of bone|Disorder of bone
C0005940|T047|OF|76069003|SNOMEDCT_CORE|Disease of bone|Disorder of bone
C0005940|T047|IS|76069003|SNOMEDCT_CORE|Disease of bone, NOS|Disorder of bone
C0005940|T047|PT|76069003|SNOMEDCT_CORE|Disorder of bone|Disorder of bone
C0005940|T047|FN|76069003|SNOMEDCT_CORE|Disorder of bone|Disorder of bone
C0005940|T047|SY|76069003|SNOMEDCT_CORE|Osteopathia|Disorder of bone
C0005940|T047|IS|76069003|SNOMEDCT_CORE|Osteopathia, NOS|Disorder of bone
C0006012|T048|PT|20010003|SNOMEDCT_CORE|Borderline personality disorder|Borderline personality disorder
C0006012|T048|FN|20010003|SNOMEDCT_CORE|Borderline personality disorder|Borderline personality disorder
C0006091|T047|SY|3548001|SNOMEDCT_CORE|Brachial plexus lesion|Brachial plexus lesion
C0006091|T047|IS|3548001|SNOMEDCT_CORE|Brachial plexus lesion, NOS|Brachial plexus lesion
C0006105|T047|IS|60404007|SNOMEDCT_CORE|Brain abscess|Brain abscess
C0006107|T037|SY|110030002|SNOMEDCT_CORE|Brain concussion|Concussion injury of brain
C0006107|T037|IS|110030002|SNOMEDCT_CORE|Cerebral concussion|Concussion injury of brain
C0006107|T037|SY|110030002|SNOMEDCT_CORE|Commotio cerebri|Concussion injury of brain
C0006107|T037|IS|110030002|SNOMEDCT_CORE|Concussion|Concussion injury of brain
C0006107|T037|FN|110030002|SNOMEDCT_CORE|Concussion injury of brain|Concussion injury of brain
C0006107|T037|PT|110030002|SNOMEDCT_CORE|Concussion injury of brain|Concussion injury of brain
C0006107|T037|SY|110030002|SNOMEDCT_CORE|Mild traumatic brain injury|Concussion injury of brain
C0006107|T037|SY|110030002|SNOMEDCT_CORE|MTBI - Mild traumatic brain injury|Concussion injury of brain
C0006111|T047|IS|81308009|SNOMEDCT_CORE|Disease of brain|Disorder of brain
C0006111|T047|OF|81308009|SNOMEDCT_CORE|Disease of brain|Disorder of brain
C0006111|T047|IS|81308009|SNOMEDCT_CORE|Disease of brain, NOS|Disorder of brain
C0006111|T047|PT|81308009|SNOMEDCT_CORE|Disorder of brain|Disorder of brain
C0006111|T047|FN|81308009|SNOMEDCT_CORE|Disorder of brain|Disorder of brain
C0006114|T046|PT|2032001|SNOMEDCT_CORE|Cerebral edema|Cerebral edema
C0006114|T046|FN|2032001|SNOMEDCT_CORE|Cerebral edema|Cerebral edema
C0006114|T046|PTGB|2032001|SNOMEDCT_CORE|Cerebral oedema|Cerebral edema
C0006118|T191|PT|126952004|SNOMEDCT_CORE|Neoplasm of brain|Neoplasm of brain
C0006118|T191|FN|126952004|SNOMEDCT_CORE|Neoplasm of brain|Neoplasm of brain
C0006123|T047|PT|50821009|SNOMEDCT_CORE|Arterial retinal branch occlusion|Arterial retinal branch occlusion
C0006123|T047|FN|50821009|SNOMEDCT_CORE|Arterial retinal branch occlusion|Arterial retinal branch occlusion
C0006123|T047|SY|50821009|SNOMEDCT_CORE|Branch retinal artery occlusion|Arterial retinal branch occlusion
C0006123|T047|SY|50821009|SNOMEDCT_CORE|BRAO - Branch retinal artery occlusion|Arterial retinal branch occlusion
C0006142|T191|SY|254837009|SNOMEDCT_CORE|Breast cancer|Malignant tumor of breast
C0006142|T191|SY|254837009|SNOMEDCT_CORE|CA - Breast cancer|Malignant tumor of breast
C0006142|T191|SY|254837009|SNOMEDCT_CORE|Malignant neoplasm of breast|Malignant tumor of breast
C0006142|T191|FN|254837009|SNOMEDCT_CORE|Malignant neoplasm of breast|Malignant tumor of breast
C0006142|T191|PT|254837009|SNOMEDCT_CORE|Malignant tumor of breast|Malignant tumor of breast
C0006142|T191|OF|254837009|SNOMEDCT_CORE|Malignant tumor of breast|Malignant tumor of breast
C0006142|T191|PTGB|254837009|SNOMEDCT_CORE|Malignant tumour of breast|Malignant tumor of breast
C0006144|T020|PT|399294002|SNOMEDCT_CORE|Cyst of breast|Cyst of breast
C0006144|T020|FN|399294002|SNOMEDCT_CORE|Cyst of breast|Cyst of breast
C0006145|T047|SY|79604008|SNOMEDCT_CORE|Breast disease|Disorder of breast
C0006145|T047|IS|79604008|SNOMEDCT_CORE|Disease of breast|Disorder of breast
C0006145|T047|OF|79604008|SNOMEDCT_CORE|Disease of breast|Disorder of breast
C0006145|T047|IS|79604008|SNOMEDCT_CORE|Disease of breast, NOS|Disorder of breast
C0006145|T047|PT|79604008|SNOMEDCT_CORE|Disorder of breast|Disorder of breast
C0006145|T047|FN|79604008|SNOMEDCT_CORE|Disorder of breast|Disorder of breast
C0006145|T047|IS|79604008|SNOMEDCT_CORE|Disorder of breast, NOS|Disorder of breast
C0006157|T046|PT|6096002|SNOMEDCT_CORE|Breech presentation|Breech presentation
C0006157|T046|FN|6096002|SNOMEDCT_CORE|Breech presentation|Breech presentation
C0006266|T047|SY|4386001|SNOMEDCT_CORE|Bronchial spasm|Bronchospasm
C0006266|T047|PT|4386001|SNOMEDCT_CORE|Bronchospasm|Bronchospasm
C0006266|T047|FN|4386001|SNOMEDCT_CORE|Bronchospasm|Bronchospasm
C0006267|T047|PT|12295008|SNOMEDCT_CORE|Bronchiectasis|Bronchiectasis
C0006267|T047|FN|12295008|SNOMEDCT_CORE|Bronchiectasis|Bronchiectasis
C0006267|T047|IS|12295008|SNOMEDCT_CORE|Bronchiectasis, NOS|Bronchiectasis
C0006271|T047|PT|4120002|SNOMEDCT_CORE|Bronchiolitis|Bronchiolitis
C0006271|T047|FN|4120002|SNOMEDCT_CORE|Bronchiolitis|Bronchiolitis
C0006271|T047|IS|4120002|SNOMEDCT_CORE|Bronchiolitis, NOS|Bronchiolitis
C0006272|T047|SY|40100001|SNOMEDCT_CORE|Bronchiolitis fibrosa obliterans|Obliterative bronchiolitis
C0006272|T047|SY|40100001|SNOMEDCT_CORE|Bronchiolitis obliterans|Obliterative bronchiolitis
C0006272|T047|SY|40100001|SNOMEDCT_CORE|OB - Obliterative bronchiolitis|Obliterative bronchiolitis
C0006272|T047|PT|40100001|SNOMEDCT_CORE|Obliterative bronchiolitis|Obliterative bronchiolitis
C0006272|T047|FN|40100001|SNOMEDCT_CORE|Obliterative bronchiolitis|Obliterative bronchiolitis
C0006272|T047|IS|40100001|SNOMEDCT_CORE|Obliterative bronchiolitis, NOS|Obliterative bronchiolitis
C0006277|T047|PT|32398004|SNOMEDCT_CORE|Bronchitis|Bronchitis
C0006277|T047|FN|32398004|SNOMEDCT_CORE|Bronchitis|Bronchitis
C0006277|T047|IS|32398004|SNOMEDCT_CORE|Bronchitis, NOS|Bronchitis
C0006285|T047|SY|396285007|SNOMEDCT_CORE|Bronchial pneumonia|Bronchopneumonia
C0006285|T047|PT|396285007|SNOMEDCT_CORE|Bronchopneumonia|Bronchopneumonia
C0006285|T047|FN|396285007|SNOMEDCT_CORE|Bronchopneumonia|Bronchopneumonia
C0006285|T047|SY|396285007|SNOMEDCT_CORE|Lobular pneumonia|Bronchopneumonia
C0006287|T047|SY|67569000|SNOMEDCT_CORE|BPD - Bronchopulmonary dysplasia|Bronchopulmonary dysplasia of newborn
C0006287|T047|SY|67569000|SNOMEDCT_CORE|Bronchopulmonary dysplasia|Bronchopulmonary dysplasia of newborn
C0006287|T047|PT|67569000|SNOMEDCT_CORE|Bronchopulmonary dysplasia of newborn|Bronchopulmonary dysplasia of newborn
C0006287|T047|FN|67569000|SNOMEDCT_CORE|Bronchopulmonary dysplasia of newborn|Bronchopulmonary dysplasia of newborn
C0006287|T047|SY|67569000|SNOMEDCT_CORE|Chronic lung disease of prematurity|Bronchopulmonary dysplasia of newborn
C0006287|T047|SY|67569000|SNOMEDCT_CORE|Perinatal bronchopulmonary dysplasia|Bronchopulmonary dysplasia of newborn
C0006287|T047|SY|67569000|SNOMEDCT_CORE|Ventilator lung in newborn|Bronchopulmonary dysplasia of newborn
C0006318|T033|PT|70466008|SNOMEDCT_CORE|Bruit|Bruit
C0006318|T033|FN|70466008|SNOMEDCT_CORE|Bruit|Bruit
C0006325|T048|SY|191983006|SNOMEDCT_CORE|Bruxism|Bruxism
C0006325|T048|PT|191983006|SNOMEDCT_CORE|Bruxism|Bruxism
C0006325|T048|FN|191983006|SNOMEDCT_CORE|Bruxism|Bruxism
C0006325|T048|OF|191983006|SNOMEDCT_CORE|Bruxism|Bruxism
C0006370|T048|SY|78004001|SNOMEDCT_CORE|Bulimia|Bulimia
C0006384|T047|SY|6374002|SNOMEDCT_CORE|BBB - Bundle branch block|Bundle branch block
C0006384|T047|PT|6374002|SNOMEDCT_CORE|Bundle branch block|Bundle branch block
C0006384|T047|FN|6374002|SNOMEDCT_CORE|Bundle branch block|Bundle branch block
C0006384|T047|IS|6374002|SNOMEDCT_CORE|Bundle branch block, NOS|Bundle branch block
C0006386|T020|PT|415692008|SNOMEDCT_CORE|Bunion|Bunion
C0006386|T020|SY|415692008|SNOMEDCT_CORE|Bunion of great toe|Bunion
C0006386|T020|FN|415692008|SNOMEDCT_CORE|Swelling of first metatarsophalangeal joint of hallux|Bunion
C0006386|T020|SY|415692008|SNOMEDCT_CORE|Swelling of first metatarsophalangeal joint of hallux|Bunion
C0006430|T047|SY|399165002|SNOMEDCT_CORE|BMS - Burning mouth syndrome|Burning mouth syndrome
C0006430|T047|PT|399165002|SNOMEDCT_CORE|Burning mouth syndrome|Burning mouth syndrome
C0006430|T047|FN|399165002|SNOMEDCT_CORE|Burning mouth syndrome|Burning mouth syndrome
C0006430|T047|SY|399165002|SNOMEDCT_CORE|Orodynia|Burning mouth syndrome
C0006430|T047|SY|399165002|SNOMEDCT_CORE|Stomatopyrosis|Burning mouth syndrome
C0006434|T037|PT|125666000|SNOMEDCT_CORE|Burn|Burn
C0006434|T037|FN|125666000|SNOMEDCT_CORE|Burn|Burn
C0006435|T037|SY|426284001|SNOMEDCT_CORE|Caustic burn|Chemical burn
C0006435|T037|PT|426284001|SNOMEDCT_CORE|Chemical burn|Chemical burn
C0006435|T037|FN|426284001|SNOMEDCT_CORE|Chemical burn|Chemical burn
C0006444|T047|PT|84017003|SNOMEDCT_CORE|Bursitis|Bursitis
C0006444|T047|FN|84017003|SNOMEDCT_CORE|Bursitis|Bursitis
C0006444|T047|IS|84017003|SNOMEDCT_CORE|Bursitis, NOS|Bursitis
C0006444|T047|SY|84017003|SNOMEDCT_CORE|Inflammation of bursa|Bursitis
C0006625|T184|SY|238108007|SNOMEDCT_CORE|Cachectic|Cachexia
C0006625|T184|PT|238108007|SNOMEDCT_CORE|Cachexia|Cachexia
C0006625|T184|FN|238108007|SNOMEDCT_CORE|Cachexia|Cachexia
C0006625|T184|IS|238108007|SNOMEDCT_CORE|General body deterioration|Cachexia
C0006625|T184|SY|285384003|SNOMEDCT_CORE|General body deterioration|Cachexia
C0006826|T191|SY|363346000|SNOMEDCT_CORE|CA - Cancer|Malignant neoplastic disease
C0006826|T191|SY|363346000|SNOMEDCT_CORE|Cancer|Malignant neoplastic disease
C0006826|T191|SY|363346000|SNOMEDCT_CORE|Malignant neoplasm|Malignant neoplastic disease
C0006826|T191|PT|363346000|SNOMEDCT_CORE|Malignant neoplastic disease|Malignant neoplastic disease
C0006826|T191|FN|363346000|SNOMEDCT_CORE|Malignant neoplastic disease|Malignant neoplastic disease
C0006826|T191|SY|363346000|SNOMEDCT_CORE|Malignant tumor|Malignant neoplastic disease
C0006826|T191|OF|363346000|SNOMEDCT_CORE|Malignant tumor|Malignant neoplastic disease
C0006826|T191|SYGB|363346000|SNOMEDCT_CORE|Malignant tumour|Malignant neoplastic disease
C0006840|T047|SY|78048006|SNOMEDCT_CORE|Candida infection|Candidiasis
C0006840|T047|PT|78048006|SNOMEDCT_CORE|Candidiasis|Candidiasis
C0006840|T047|FN|78048006|SNOMEDCT_CORE|Candidiasis|Candidiasis
C0006840|T047|IS|78048006|SNOMEDCT_CORE|Candidiasis, NOS|Candidiasis
C0006840|T047|SY|78048006|SNOMEDCT_CORE|Candidosis|Candidiasis
C0006840|T047|IS|78048006|SNOMEDCT_CORE|Candidosis, NOS|Candidiasis
C0006840|T047|SY|78048006|SNOMEDCT_CORE|Infection by Candida species|Candidiasis
C0006840|T047|SY|78048006|SNOMEDCT_CORE|Monilia infection|Candidiasis
C0006840|T047|SY|78048006|SNOMEDCT_CORE|Moniliasis|Candidiasis
C0006840|T047|IS|78048006|SNOMEDCT_CORE|Moniliasis, NOS|Candidiasis
C0006846|T047|SY|49883006|SNOMEDCT_CORE|Candida of skin|Candidiasis of skin
C0006846|T047|PT|49883006|SNOMEDCT_CORE|Candidiasis of skin|Candidiasis of skin
C0006846|T047|FN|49883006|SNOMEDCT_CORE|Candidiasis of skin|Candidiasis of skin
C0006846|T047|SY|49883006|SNOMEDCT_CORE|Candidosis of skin|Candidiasis of skin
C0006849|T047|SY|79740000|SNOMEDCT_CORE|Candida infection of mouth|Candidiasis of mouth
C0006849|T047|SY|79740000|SNOMEDCT_CORE|Candida of mouth|Candidiasis of mouth
C0006849|T047|PT|79740000|SNOMEDCT_CORE|Candidiasis of mouth|Candidiasis of mouth
C0006849|T047|FN|79740000|SNOMEDCT_CORE|Candidiasis of mouth|Candidiasis of mouth
C0006849|T047|SY|79740000|SNOMEDCT_CORE|Candidosis of mouth|Candidiasis of mouth
C0006849|T047|SY|79740000|SNOMEDCT_CORE|Moniliasis of mouth|Candidiasis of mouth
C0006849|T047|SY|79740000|SNOMEDCT_CORE|Mycotic stomatitis|Candidiasis of mouth
C0006849|T047|SY|79740000|SNOMEDCT_CORE|Oral candidiasis|Candidiasis of mouth
C0006849|T047|SY|79740000|SNOMEDCT_CORE|Oral candidosis|Candidiasis of mouth
C0006849|T047|SY|79740000|SNOMEDCT_CORE|Oral moniliasis|Candidiasis of mouth
C0006849|T047|SY|79740000|SNOMEDCT_CORE|Oral thrush|Candidiasis of mouth
C0006849|T047|IS|79740000|SNOMEDCT_CORE|Thrush|Candidiasis of mouth
C0006849|T047|SY|78048006|SNOMEDCT_CORE|Thrush|Candidiasis of mouth
C0006852|T047|SY|72934000|SNOMEDCT_CORE|Candida of vagina|Candidiasis of vagina
C0006852|T047|PT|72934000|SNOMEDCT_CORE|Candidiasis of vagina|Candidiasis of vagina
C0006852|T047|FN|72934000|SNOMEDCT_CORE|Candidiasis of vagina|Candidiasis of vagina
C0006852|T047|IS|72934000|SNOMEDCT_CORE|Monial infection of vagina|Candidiasis of vagina
C0006852|T047|SY|72934000|SNOMEDCT_CORE|Monilial infection of vagina|Candidiasis of vagina
C0006852|T047|SY|72934000|SNOMEDCT_CORE|Vaginal candida|Candidiasis of vagina
C0006852|T047|SY|72934000|SNOMEDCT_CORE|Vaginal candidiasis|Candidiasis of vagina
C0006852|T047|SY|72934000|SNOMEDCT_CORE|Vaginal candidosis|Candidiasis of vagina
C0006852|T047|SY|72934000|SNOMEDCT_CORE|Vaginal thrush|Candidiasis of vagina
C0006868|T048|PT|37344009|SNOMEDCT_CORE|Cannabis abuse|Cannabis abuse
C0006868|T048|FN|37344009|SNOMEDCT_CORE|Cannabis abuse|Cannabis abuse
C0006870|T048|PT|85005007|SNOMEDCT_CORE|Cannabis dependence|Cannabis dependence
C0006870|T048|FN|85005007|SNOMEDCT_CORE|Cannabis dependence|Cannabis dependence
C0007020|T037|SY|17383000|SNOMEDCT_CORE|Carbon monoxide poisoning|Carbon monoxide poisoning
C0007078|T047|PT|416893007|SNOMEDCT_CORE|Carbuncle|Carbuncle
C0007078|T047|FN|416893007|SNOMEDCT_CORE|Carbuncle|Carbuncle
C0007093|T047|PT|36222008|SNOMEDCT_CORE|Carcinoid heart disease|Carcinoid heart disease
C0007093|T047|FN|36222008|SNOMEDCT_CORE|Carcinoid heart disease|Carcinoid heart disease
C0007095|T191|SY|189607006|SNOMEDCT_CORE|Carcinoid|Carcinoid tumor - morphology
C0007095|T191|SY|189607006|SNOMEDCT_CORE|Carcinoid tumor|Carcinoid tumor - morphology
C0007095|T191|PT|443492008|SNOMEDCT_CORE|Carcinoid tumor|Carcinoid tumor - morphology
C0007095|T191|FN|443492008|SNOMEDCT_CORE|Carcinoid tumor|Carcinoid tumor - morphology
C0007095|T191|PT|189607006|SNOMEDCT_CORE|Carcinoid tumor - morphology|Carcinoid tumor - morphology
C0007095|T191|FN|189607006|SNOMEDCT_CORE|Carcinoid tumor - morphology|Carcinoid tumor - morphology
C0007095|T191|IS|189607006|SNOMEDCT_CORE|Carcinoid tumors|Carcinoid tumor - morphology
C0007095|T191|SYGB|189607006|SNOMEDCT_CORE|Carcinoid tumour|Carcinoid tumor - morphology
C0007095|T191|PTGB|443492008|SNOMEDCT_CORE|Carcinoid tumour|Carcinoid tumor - morphology
C0007095|T191|PTGB|189607006|SNOMEDCT_CORE|Carcinoid tumour - morphology|Carcinoid tumor - morphology
C0007095|T191|IS|189607006|SNOMEDCT_CORE|Carcinoid tumours|Carcinoid tumor - morphology
C0007102|T191|SY|363406005|SNOMEDCT_CORE|CA - Cancer of colon|Malignant tumor of colon
C0007102|T191|SY|363406005|SNOMEDCT_CORE|Cancer of colon|Malignant tumor of colon
C0007102|T191|SY|363406005|SNOMEDCT_CORE|Malignant neoplasm of colon|Malignant tumor of colon
C0007102|T191|FN|363406005|SNOMEDCT_CORE|Malignant neoplasm of colon|Malignant tumor of colon
C0007102|T191|PT|363406005|SNOMEDCT_CORE|Malignant tumor of colon|Malignant tumor of colon
C0007102|T191|OF|363406005|SNOMEDCT_CORE|Malignant tumor of colon|Malignant tumor of colon
C0007102|T191|PTGB|363406005|SNOMEDCT_CORE|Malignant tumour of colon|Malignant tumor of colon
C0007107|T191|SY|363429002|SNOMEDCT_CORE|CA - Cancer of larynx|Malignant tumor of larynx
C0007107|T191|SY|363429002|SNOMEDCT_CORE|Cancer of larynx|Malignant tumor of larynx
C0007107|T191|SY|363429002|SNOMEDCT_CORE|Laryngeal cancer|Malignant tumor of larynx
C0007107|T191|PT|363429002|SNOMEDCT_CORE|Malignant tumor of larynx|Malignant tumor of larynx
C0007107|T191|FN|363429002|SNOMEDCT_CORE|Malignant tumor of larynx|Malignant tumor of larynx
C0007107|T191|PTGB|363429002|SNOMEDCT_CORE|Malignant tumour of larynx|Malignant tumor of larynx
C0007112|T191|PT|399490008|SNOMEDCT_CORE|Adenocarcinoma of prostate|Adenocarcinoma of prostate
C0007112|T191|FN|399490008|SNOMEDCT_CORE|Adenocarcinoma of prostate|Adenocarcinoma of prostate
C0007113|T191|IS|254582000|SNOMEDCT_CORE|Carcinoma of rectum|Carcinoma of rectum
C0007113|T191|IS|254582000|SNOMEDCT_CORE|Rectal carcinoma|Carcinoma of rectum
C0007114|T191|SY|372130007|SNOMEDCT_CORE|Cancer of skin|Malignant neoplasm of skin
C0007114|T191|PT|372130007|SNOMEDCT_CORE|Malignant neoplasm of skin|Malignant neoplasm of skin
C0007114|T191|FN|372130007|SNOMEDCT_CORE|Malignant neoplasm of skin|Malignant neoplasm of skin
C0007114|T191|SY|372130007|SNOMEDCT_CORE|Skin cancer|Malignant neoplasm of skin
C0007115|T191|IS|94098005|SNOMEDCT_CORE|Malignant neoplasm of thyroid gland|Malignant tumor of thyroid gland
C0007115|T191|PT|363478007|SNOMEDCT_CORE|Malignant tumor of thyroid gland|Malignant tumor of thyroid gland
C0007115|T191|FN|363478007|SNOMEDCT_CORE|Malignant tumor of thyroid gland|Malignant tumor of thyroid gland
C0007115|T191|PTGB|363478007|SNOMEDCT_CORE|Malignant tumour of thyroid gland|Malignant tumor of thyroid gland
C0007115|T191|SY|363478007|SNOMEDCT_CORE|Thyroid Ca|Malignant tumor of thyroid gland
C0007115|T191|SY|363478007|SNOMEDCT_CORE|Thyroid cancer|Malignant tumor of thyroid gland
C0007121|T191|SY|254622008|SNOMEDCT_CORE|BC - Bronchogenic carcinoma|Bronchial carcinoma
C0007121|T191|SY|254622008|SNOMEDCT_CORE|Bronchial carcinoma|Bronchial carcinoma
C0007121|T191|SY|254622008|SNOMEDCT_CORE|Bronchogenic carcinoma|Bronchial carcinoma
C0007121|T191|SY|254622008|SNOMEDCT_CORE|CA - Carcinoma of bronchus|Bronchial carcinoma
C0007121|T191|SY|254622008|SNOMEDCT_CORE|Carcinoma of bronchus|Bronchial carcinoma
C0007124|T191|PT|109889007|SNOMEDCT_CORE|Intraductal carcinoma in situ of breast|Intraductal carcinoma in situ of breast
C0007124|T191|FN|109889007|SNOMEDCT_CORE|Intraductal carcinoma in situ of breast|Intraductal carcinoma in situ of breast
C0007129|T191|PT|253001006|SNOMEDCT_CORE|Merkel cell carcinoma|Merkel cell carcinoma
C0007129|T191|FN|253001006|SNOMEDCT_CORE|Merkel cell carcinoma|Merkel cell carcinoma
C0007129|T191|SY|253001006|SNOMEDCT_CORE|Merkel cell tumor|Merkel cell carcinoma
C0007129|T191|SYGB|253001006|SNOMEDCT_CORE|Merkel cell tumour|Merkel cell carcinoma
C0007129|T191|SY|253001006|SNOMEDCT_CORE|Trabecular cell carcinoma of skin|Merkel cell carcinoma
C0007131|T191|PT|254637007|SNOMEDCT_CORE|Non-small cell lung cancer|Non-small cell lung cancer
C0007131|T191|FN|254637007|SNOMEDCT_CORE|Non-small cell lung cancer|Non-small cell lung cancer
C0007131|T191|SY|254637007|SNOMEDCT_CORE|NSCLC - Non-small cell lung cancer|Non-small cell lung cancer
C0007134|T191|IS|254915003|SNOMEDCT_CORE|Adenocarcinoma of kidney|Renal cell adenocarcinoma
C0007134|T191|IS|254915003|SNOMEDCT_CORE|Renal cell adenocarcinoma|Renal cell adenocarcinoma
C0007134|T191|IS|254915003|SNOMEDCT_CORE|Renal cell carcinoma|Renal cell adenocarcinoma
C0007137|T191|PT|402815007|SNOMEDCT_CORE|Squamous cell carcinoma|Squamous cell carcinoma
C0007137|T191|FN|402815007|SNOMEDCT_CORE|Squamous cell carcinoma|Squamous cell carcinoma
C0007192|T047|SY|83521008|SNOMEDCT_CORE|Alcoholic cardiomyopathy|Dilated cardiomyopathy secondary to alcohol
C0007192|T047|FN|83521008|SNOMEDCT_CORE|Dilated cardiomyopathy caused by alcohol|Dilated cardiomyopathy secondary to alcohol
C0007192|T047|SY|83521008|SNOMEDCT_CORE|Dilated cardiomyopathy caused by alcohol|Dilated cardiomyopathy secondary to alcohol
C0007192|T047|PT|83521008|SNOMEDCT_CORE|Dilated cardiomyopathy secondary to alcohol|Dilated cardiomyopathy secondary to alcohol
C0007192|T047|OF|83521008|SNOMEDCT_CORE|Dilated cardiomyopathy secondary to alcohol|Dilated cardiomyopathy secondary to alcohol
C0007193|T047|SY|399020009|SNOMEDCT_CORE|CCM - Congestive cardiomyopathy|Dilated cardiomyopathy
C0007193|T047|SY|399020009|SNOMEDCT_CORE|COCM - Congestive cardiomyopathy|Dilated cardiomyopathy
C0007193|T047|SY|399020009|SNOMEDCT_CORE|Congestive cardiomyopathy|Dilated cardiomyopathy
C0007193|T047|FN|399020009|SNOMEDCT_CORE|Congestive cardiomyopathy|Dilated cardiomyopathy
C0007193|T047|SY|399020009|SNOMEDCT_CORE|Congestive dilated cardiomyopathy|Dilated cardiomyopathy
C0007193|T047|SY|399020009|SNOMEDCT_CORE|DCM - Dilated cardiomyopathy|Dilated cardiomyopathy
C0007193|T047|PT|399020009|SNOMEDCT_CORE|Dilated cardiomyopathy|Dilated cardiomyopathy
C0007194|T047|SY|233873004|SNOMEDCT_CORE|HCM - Hypertrophic cardiomyopathy|Hypertrophic cardiomyopathy
C0007194|T047|PT|233873004|SNOMEDCT_CORE|Hypertrophic cardiomyopathy|Hypertrophic cardiomyopathy
C0007194|T047|FN|233873004|SNOMEDCT_CORE|Hypertrophic cardiomyopathy|Hypertrophic cardiomyopathy
C0007196|T047|SY|415295002|SNOMEDCT_CORE|Constrictive cardiomyopathy|Restrictive cardiomyopathy
C0007196|T047|PT|415295002|SNOMEDCT_CORE|Restrictive cardiomyopathy|Restrictive cardiomyopathy
C0007196|T047|FN|415295002|SNOMEDCT_CORE|Restrictive cardiomyopathy|Restrictive cardiomyopathy
C0007222|T047|SY|49601007|SNOMEDCT_CORE|Cardiovascular disease|Disorder of cardiovascular system
C0007222|T047|IS|49601007|SNOMEDCT_CORE|Cardiovascular disease, NOS|Disorder of cardiovascular system
C0007222|T047|SY|49601007|SNOMEDCT_CORE|Cardiovascular disorder|Disorder of cardiovascular system
C0007222|T047|IS|49601007|SNOMEDCT_CORE|Cardiovascular disorder, NOS|Disorder of cardiovascular system
C0007222|T047|SY|49601007|SNOMEDCT_CORE|Cardiovascular system disease|Disorder of cardiovascular system
C0007222|T047|IS|49601007|SNOMEDCT_CORE|CVD|Disorder of cardiovascular system
C0007222|T047|SY|49601007|SNOMEDCT_CORE|CVD - cardiovascular disease|Disorder of cardiovascular system
C0007222|T047|IS|49601007|SNOMEDCT_CORE|CVD, NOS|Disorder of cardiovascular system
C0007222|T047|IS|49601007|SNOMEDCT_CORE|CVS disease|Disorder of cardiovascular system
C0007222|T047|SY|49601007|SNOMEDCT_CORE|CVS disease - cardiovascular system disease|Disorder of cardiovascular system
C0007222|T047|IS|49601007|SNOMEDCT_CORE|Disease of cardiovascular system|Disorder of cardiovascular system
C0007222|T047|OF|49601007|SNOMEDCT_CORE|Disease of cardiovascular system|Disorder of cardiovascular system
C0007222|T047|IS|49601007|SNOMEDCT_CORE|Disease of cardiovascular system, NOS|Disorder of cardiovascular system
C0007222|T047|FN|49601007|SNOMEDCT_CORE|Disorder of cardiovascular system|Disorder of cardiovascular system
C0007222|T047|PT|49601007|SNOMEDCT_CORE|Disorder of cardiovascular system|Disorder of cardiovascular system
C0007273|T047|SY|371160000|SNOMEDCT_CORE|Carotid artery disease|Disorder of carotid artery
C0007273|T047|SY|371160000|SNOMEDCT_CORE|Disease of carotid artery|Disorder of carotid artery
C0007273|T047|PT|371160000|SNOMEDCT_CORE|Disorder of carotid artery|Disorder of carotid artery
C0007273|T047|FN|371160000|SNOMEDCT_CORE|Disorder of carotid artery|Disorder of carotid artery
C0007280|T033|PT|419642000|SNOMEDCT_CORE|Carotid bruit|Carotid bruit
C0007280|T033|FN|419642000|SNOMEDCT_CORE|Carotid bruit|Carotid bruit
C0007282|T047|SY|64586002|SNOMEDCT_CORE|Carotid artery narrowing|Carotid artery stenosis
C0007282|T047|PT|64586002|SNOMEDCT_CORE|Carotid artery stenosis|Carotid artery stenosis
C0007282|T047|FN|64586002|SNOMEDCT_CORE|Carotid artery stenosis|Carotid artery stenosis
C0007286|T047|SY|57406009|SNOMEDCT_CORE|Carpal canal|Carpal tunnel syndrome
C0007286|T047|SY|57406009|SNOMEDCT_CORE|Carpal tunnel|Carpal tunnel syndrome
C0007286|T047|PT|57406009|SNOMEDCT_CORE|Carpal tunnel syndrome|Carpal tunnel syndrome
C0007286|T047|FN|57406009|SNOMEDCT_CORE|Carpal tunnel syndrome|Carpal tunnel syndrome
C0007286|T047|SY|57406009|SNOMEDCT_CORE|CTS - Carpal tunnel syndrome|Carpal tunnel syndrome
C0007286|T047|SY|57406009|SNOMEDCT_CORE|Distal median nerve compression|Carpal tunnel syndrome
C0007286|T047|SY|57406009|SNOMEDCT_CORE|Distal median nerve entrapment|Carpal tunnel syndrome
C0007286|T047|IS|57406009|SNOMEDCT_CORE|Median nerve compression|Carpal tunnel syndrome
C0007286|T047|IS|57406009|SNOMEDCT_CORE|Median nerve entrapment|Carpal tunnel syndrome
C0007459|T047|PT|12454008|SNOMEDCT_CORE|Cauda equina syndrome with neurogenic bladder|Cauda equina syndrome with neurogenic bladder
C0007459|T047|FN|12454008|SNOMEDCT_CORE|Cauda equina syndrome with neurogenic bladder|Cauda equina syndrome with neurogenic bladder
C0007570|T047|SY|396331005|SNOMEDCT_CORE|CD - Celiac disease|Celiac disease
C0007570|T047|SYGB|396331005|SNOMEDCT_CORE|CD - Coeliac disease|Celiac disease
C0007570|T047|PT|396331005|SNOMEDCT_CORE|Celiac disease|Celiac disease
C0007570|T047|FN|396331005|SNOMEDCT_CORE|Celiac disease|Celiac disease
C0007570|T047|SY|396331005|SNOMEDCT_CORE|Celiac sprue|Celiac disease
C0007570|T047|SY|396331005|SNOMEDCT_CORE|Celiac syndrome|Celiac disease
C0007570|T047|PTGB|396331005|SNOMEDCT_CORE|Coeliac disease|Celiac disease
C0007570|T047|SYGB|396331005|SNOMEDCT_CORE|Coeliac sprue|Celiac disease
C0007570|T047|SYGB|396331005|SNOMEDCT_CORE|Coeliac syndrome|Celiac disease
C0007570|T047|SY|396331005|SNOMEDCT_CORE|CS - Celiac sprue|Celiac disease
C0007570|T047|SYGB|396331005|SNOMEDCT_CORE|CS - Coeliac sprue|Celiac disease
C0007570|T047|SY|396331005|SNOMEDCT_CORE|Gluten enteropathy|Celiac disease
C0007570|T047|SY|396331005|SNOMEDCT_CORE|Gluten-induced enteropathy syndrome|Celiac disease
C0007570|T047|SY|396331005|SNOMEDCT_CORE|Gluten-responsive sprue|Celiac disease
C0007570|T047|SY|396331005|SNOMEDCT_CORE|Gluten-sensitive enteropathy|Celiac disease
C0007570|T047|SY|396331005|SNOMEDCT_CORE|GSE - Gluten-sensitive enteropathy|Celiac disease
C0007570|T047|SY|396331005|SNOMEDCT_CORE|Idiopathic steatorrhea|Celiac disease
C0007570|T047|SYGB|396331005|SNOMEDCT_CORE|Idiopathic steatorrhoea|Celiac disease
C0007570|T047|SY|396331005|SNOMEDCT_CORE|Non-tropical sprue|Celiac disease
C0007570|T047|SY|396331005|SNOMEDCT_CORE|Nontropical sprue|Celiac disease
C0007570|T047|IS|396331005|SNOMEDCT_CORE|Sprue|Celiac disease
C0007570|T047|SY|396331005|SNOMEDCT_CORE|Wheat-sensitive enteropathy|Celiac disease
C0007642|T046|PT|128045006|SNOMEDCT_CORE|Cellulitis|Cellulitis
C0007642|T046|FN|128045006|SNOMEDCT_CORE|Cellulitis|Cellulitis
C0007646|T047|PT|62837005|SNOMEDCT_CORE|Cellulitis of hand|Cellulitis of hand
C0007646|T047|FN|62837005|SNOMEDCT_CORE|Cellulitis of hand|Cellulitis of hand
C0007688|T047|PT|38742007|SNOMEDCT_CORE|Central retinal artery occlusion|Central retinal artery occlusion
C0007688|T047|FN|38742007|SNOMEDCT_CORE|Central retinal artery occlusion|Central retinal artery occlusion
C0007688|T047|SY|38742007|SNOMEDCT_CORE|CRA - Central retinal artery occlusion|Central retinal artery occlusion
C0007688|T047|SY|38742007|SNOMEDCT_CORE|CRAO - Central retinal artery occlusion|Central retinal artery occlusion
C0007722|T047|PTGB|206200000|SNOMEDCT_CORE|Cephalhaematoma due to birth trauma|Cephalhematoma due to birth trauma
C0007722|T047|PT|206200000|SNOMEDCT_CORE|Cephalhematoma due to birth trauma|Cephalhematoma due to birth trauma
C0007722|T047|FN|206200000|SNOMEDCT_CORE|Cephalhematoma due to birth trauma|Cephalhematoma due to birth trauma
C0007722|T047|SY|206200000|SNOMEDCT_CORE|Cephalohematoma due to birth trauma|Cephalhematoma due to birth trauma
C0007758|T047|PT|85102008|SNOMEDCT_CORE|Cerebellar ataxia|Cerebellar ataxia
C0007758|T047|FN|85102008|SNOMEDCT_CORE|Cerebellar ataxia|Cerebellar ataxia
C0007758|T047|IS|85102008|SNOMEDCT_CORE|Cerebellar ataxia, NOS|Cerebellar ataxia
C0007766|T047|PT|128609009|SNOMEDCT_CORE|Intracranial aneurysm|Intracranial aneurysm
C0007766|T047|FN|128609009|SNOMEDCT_CORE|Intracranial aneurysm|Intracranial aneurysm
C0007766|T047|IS|42994005|SNOMEDCT_CORE|Intracranial aneurysm, NOS|Intracranial aneurysm
C0007775|T047|SY|55382008|SNOMEDCT_CORE|Atherosclerosis of intracranial artery|Cerebral atherosclerosis
C0007775|T047|PT|55382008|SNOMEDCT_CORE|Cerebral atherosclerosis|Cerebral atherosclerosis
C0007775|T047|FN|55382008|SNOMEDCT_CORE|Cerebral atherosclerosis|Cerebral atherosclerosis
C0007775|T047|SY|55382008|SNOMEDCT_CORE|ICAD - intracranial atherosclerotic disease|Cerebral atherosclerosis
C0007775|T047|SY|55382008|SNOMEDCT_CORE|ICAS - intracranial atherosclerosis|Cerebral atherosclerosis
C0007780|T047|SY|75543006|SNOMEDCT_CORE|Cerebral arterial embolism|Cerebral embolism
C0007780|T047|PT|75543006|SNOMEDCT_CORE|Cerebral embolism|Cerebral embolism
C0007780|T047|FN|75543006|SNOMEDCT_CORE|Cerebral embolism|Cerebral embolism
C0007785|T047|PT|432504007|SNOMEDCT_CORE|Cerebral infarction|Cerebral infarction
C0007785|T047|FN|432504007|SNOMEDCT_CORE|Cerebral infarction|Cerebral infarction
C0007787|T047|SY|266257000|SNOMEDCT_CORE|Temporary cerebral vascular dysfunction|Transient cerebral ischemia
C0007787|T047|SY|266257000|SNOMEDCT_CORE|TIA|Transient cerebral ischemia
C0007787|T047|SYGB|266257000|SNOMEDCT_CORE|TIA - Transient ischaemic attack|Transient cerebral ischemia
C0007787|T047|PTGB|266257000|SNOMEDCT_CORE|Transient cerebral ischaemia|Transient cerebral ischemia
C0007787|T047|PT|266257000|SNOMEDCT_CORE|Transient cerebral ischemia|Transient cerebral ischemia
C0007787|T047|SYGB|266257000|SNOMEDCT_CORE|Transient ischaemic attack|Transient cerebral ischemia
C0007787|T047|SY|266257000|SNOMEDCT_CORE|Transient ischemic attack|Transient cerebral ischemia
C0007787|T047|FN|266257000|SNOMEDCT_CORE|Transient ischemic attack|Transient cerebral ischemia
C0007789|T047|PT|128188000|SNOMEDCT_CORE|Cerebral palsy|Cerebral palsy
C0007789|T047|SY|128188000|SNOMEDCT_CORE|Cerebral palsy|Cerebral palsy
C0007789|T047|FN|128188000|SNOMEDCT_CORE|Cerebral palsy|Cerebral palsy
C0007789|T047|IS|1178005|SNOMEDCT_CORE|Cerebral palsy, NOS|Cerebral palsy
C0007789|T047|SY|128188000|SNOMEDCT_CORE|Congenital cerebral palsy|Cerebral palsy
C0007789|T047|SY|128188000|SNOMEDCT_CORE|CP - Cerebral palsy|Cerebral palsy
C0007789|T047|SY|128188000|SNOMEDCT_CORE|Infantile cerebral palsy|Cerebral palsy
C0007820|T047|PT|62914000|SNOMEDCT_CORE|Cerebrovascular disease|Cerebrovascular disease
C0007820|T047|FN|62914000|SNOMEDCT_CORE|Cerebrovascular disease|Cerebrovascular disease
C0007820|T047|IS|62914000|SNOMEDCT_CORE|Cerebrovascular disease, NOS|Cerebrovascular disease
C0007820|T047|IS|62914000|SNOMEDCT_CORE|Cerebrovascular lesion|Cerebrovascular disease
C0007820|T047|IS|62914000|SNOMEDCT_CORE|Cerebrovascular lesion, NOS|Cerebrovascular disease
C0007820|T047|SY|62914000|SNOMEDCT_CORE|CVD - Cerebrovascular disease|Cerebrovascular disease
C0007847|T191|SY|363354003|SNOMEDCT_CORE|Cancer of the uterine cervix|Malignant tumor of cervix
C0007847|T191|SY|363354003|SNOMEDCT_CORE|Cervical cancer|Malignant tumor of cervix
C0007847|T191|SY|363354003|SNOMEDCT_CORE|Malignant neoplasm of cervix|Malignant tumor of cervix
C0007847|T191|SY|363354003|SNOMEDCT_CORE|Malignant neoplasm of cervix uteri|Malignant tumor of cervix
C0007847|T191|PT|363354003|SNOMEDCT_CORE|Malignant tumor of cervix|Malignant tumor of cervix
C0007847|T191|FN|363354003|SNOMEDCT_CORE|Malignant tumor of cervix|Malignant tumor of cervix
C0007847|T191|PTGB|363354003|SNOMEDCT_CORE|Malignant tumour of cervix|Malignant tumor of cervix
C0007855|T191|SY|65576009|SNOMEDCT_CORE|Cervical polyp|Polyp of cervix
C0007855|T191|PT|65576009|SNOMEDCT_CORE|Polyp of cervix|Polyp of cervix
C0007855|T191|FN|65576009|SNOMEDCT_CORE|Polyp of cervix|Polyp of cervix
C0007855|T191|IS|65576009|SNOMEDCT_CORE|Polyp of cervix, NOS|Polyp of cervix
C0007859|T184|SY|81680005|SNOMEDCT_CORE|Cervical pain|Neck pain
C0007859|T184|SY|81680005|SNOMEDCT_CORE|Cervicalgia|Neck pain
C0007859|T184|IS|81680005|SNOMEDCT_CORE|Cervicodynia|Neck pain
C0007859|T184|SY|81680005|SNOMEDCT_CORE|Neck ache|Neck pain
C0007859|T184|PT|81680005|SNOMEDCT_CORE|Neck pain|Neck pain
C0007859|T184|FN|81680005|SNOMEDCT_CORE|Neck pain|Neck pain
C0007859|T184|SY|81680005|SNOMEDCT_CORE|Nonspecific pain in the neck region|Neck pain
C0007859|T184|SY|81680005|SNOMEDCT_CORE|Painful neck|Neck pain
C0007860|T047|SY|37610005|SNOMEDCT_CORE|Cervicitis|Inflammation of cervix
C0007860|T047|PT|37610005|SNOMEDCT_CORE|Inflammation of cervix|Inflammation of cervix
C0007860|T047|FN|37610005|SNOMEDCT_CORE|Inflammation of cervix|Inflammation of cervix
C0007860|T047|SY|37610005|SNOMEDCT_CORE|Inflammatory disease of the cervix|Inflammation of cervix
C0007860|T047|IS|37610005|SNOMEDCT_CORE|Inflammatory disease of the uterine cervix|Inflammation of cervix
C0007860|T047|SY|37610005|SNOMEDCT_CORE|Trachelitis|Inflammation of cervix
C0007863|T047|PT|71760005|SNOMEDCT_CORE|Cervico-occipital neuralgia|Cervico-occipital neuralgia
C0007863|T047|FN|71760005|SNOMEDCT_CORE|Cervico-occipital neuralgia|Cervico-occipital neuralgia
C0007863|T047|SY|71760005|SNOMEDCT_CORE|Occipital neuralgia|Cervico-occipital neuralgia
C0007867|T047|SY|63339007|SNOMEDCT_CORE|Disease of cervix|Disorder of uterine cervix
C0007867|T047|IS|63339007|SNOMEDCT_CORE|Disease of cervix, NOS|Disorder of uterine cervix
C0007867|T047|IS|63339007|SNOMEDCT_CORE|Disease of uterine cervix|Disorder of uterine cervix
C0007867|T047|OF|63339007|SNOMEDCT_CORE|Disease of uterine cervix|Disorder of uterine cervix
C0007867|T047|IS|63339007|SNOMEDCT_CORE|Disease of uterine cervix, NOS|Disorder of uterine cervix
C0007867|T047|SY|63339007|SNOMEDCT_CORE|Disorder of cervix|Disorder of uterine cervix
C0007867|T047|IS|63339007|SNOMEDCT_CORE|Disorder of cervix, NOS|Disorder of uterine cervix
C0007867|T047|PT|63339007|SNOMEDCT_CORE|Disorder of uterine cervix|Disorder of uterine cervix
C0007867|T047|FN|63339007|SNOMEDCT_CORE|Disorder of uterine cervix|Disorder of uterine cervix
C0007867|T047|IS|63339007|SNOMEDCT_CORE|Disorder of uterine cervix, NOS|Disorder of uterine cervix
C0007868|T047|SY|73391008|SNOMEDCT_CORE|Cervical dysplasia|Dysplasia of cervix
C0007868|T047|PT|73391008|SNOMEDCT_CORE|Dysplasia of cervix|Dysplasia of cervix
C0007868|T047|FN|73391008|SNOMEDCT_CORE|Dysplasia of cervix|Dysplasia of cervix
C0007868|T047|SY|73391008|SNOMEDCT_CORE|Dysplasia of cervix uteri|Dysplasia of cervix
C0007871|T046|SY|17382005|SNOMEDCT_CORE|Abnormal dilatation of cervix before onset of labor|Cervical incompetence
C0007871|T046|SYGB|17382005|SNOMEDCT_CORE|Abnormal dilatation of cervix before onset of labour|Cervical incompetence
C0007871|T046|PT|17382005|SNOMEDCT_CORE|Cervical incompetence|Cervical incompetence
C0007871|T046|FN|17382005|SNOMEDCT_CORE|Cervical incompetence|Cervical incompetence
C0007871|T046|SY|17382005|SNOMEDCT_CORE|Cervical insufficiency|Cervical incompetence
C0007871|T046|SY|17382005|SNOMEDCT_CORE|CI - Cervical incompetence|Cervical incompetence
C0007871|T046|SY|17382005|SNOMEDCT_CORE|Incompetence of cervix|Cervical incompetence
C0007871|T046|SY|17382005|SNOMEDCT_CORE|Incompetent cervix|Cervical incompetence
C0007933|T047|PT|1482004|SNOMEDCT_CORE|Chalazion|Chalazion
C0007933|T047|OF|1482004|SNOMEDCT_CORE|Chalazion|Chalazion
C0007933|T047|SY|1482004|SNOMEDCT_CORE|Cyst of meibomian gland|Chalazion
C0007933|T047|FN|1482004|SNOMEDCT_CORE|Cyst of meibomian gland|Chalazion
C0007933|T047|SY|1482004|SNOMEDCT_CORE|Meibomian cyst|Chalazion
C0007933|T047|SY|1482004|SNOMEDCT_CORE|Meibomian gland cyst|Chalazion
C0007933|T047|SY|1482004|SNOMEDCT_CORE|Tarsal cyst|Chalazion
C0007959|T047|OAP|50548001|SNOMEDCT_CORE|Charcot-Marie-Tooth disease|Hereditary sensory-motor neuropathy, NOS
C0007959|T047|OAF|50548001|SNOMEDCT_CORE|Charcot-Marie-Tooth disease|Hereditary sensory-motor neuropathy, NOS
C0007959|T047|OAS|50548001|SNOMEDCT_CORE|CMT - Charcot-Marie-Tooth disease|Hereditary sensory-motor neuropathy, NOS
C0007959|T047|IS|50548001|SNOMEDCT_CORE|Hereditary sensory-motor neuropathy, NOS|Hereditary sensory-motor neuropathy, NOS
C0007959|T047|IS|50548001|SNOMEDCT_CORE|Neuropathic muscular atrophy|Hereditary sensory-motor neuropathy, NOS
C0007959|T047|OAS|50548001|SNOMEDCT_CORE|Peroneal muscular atrophy|Hereditary sensory-motor neuropathy, NOS
C0007971|T047|PT|7847004|SNOMEDCT_CORE|Cheilitis|Cheilitis
C0007971|T047|FN|7847004|SNOMEDCT_CORE|Cheilitis|Cheilitis
C0007971|T047|IS|7847004|SNOMEDCT_CORE|Cheilitis, NOS|Cheilitis
C0008031|T184|PT|29857009|SNOMEDCT_CORE|Chest pain|Chest pain
C0008031|T184|FN|29857009|SNOMEDCT_CORE|Chest pain|Chest pain
C0008031|T184|IS|29857009|SNOMEDCT_CORE|Chest pain, NOS|Chest pain
C0008033|T184|SY|2237002|SNOMEDCT_CORE|Pleural pain|Pleuritic pain
C0008033|T184|SY|2237002|SNOMEDCT_CORE|Pleuralgia|Pleuritic pain
C0008033|T184|IS|2237002|SNOMEDCT_CORE|Pleuritic chest pain|Pleuritic pain
C0008033|T184|PT|2237002|SNOMEDCT_CORE|Pleuritic pain|Pleuritic pain
C0008033|T184|FN|2237002|SNOMEDCT_CORE|Pleuritic pain|Pleuritic pain
C0008033|T184|SY|2237002|SNOMEDCT_CORE|Pleurodynia|Pleuritic pain
C0008035|T184|PT|102588006|SNOMEDCT_CORE|Chest wall pain|Chest wall pain
C0008035|T184|FN|102588006|SNOMEDCT_CORE|Chest wall pain|Chest wall pain
C0008049|T047|SY|38907003|SNOMEDCT_CORE|Chicken pox|Varicella
C0008049|T047|SY|38907003|SNOMEDCT_CORE|Chickenpox|Varicella
C0008049|T047|IS|38907003|SNOMEDCT_CORE|Chickenpox, NOS|Varicella
C0008049|T047|PT|38907003|SNOMEDCT_CORE|Varicella|Varicella
C0008049|T047|FN|38907003|SNOMEDCT_CORE|Varicella|Varicella
C0008049|T047|SY|38907003|SNOMEDCT_CORE|Varicella infection|Varicella
C0008049|T047|IS|38907003|SNOMEDCT_CORE|Varicella, NOS|Varicella
C0008060|T048|PT|418189009|SNOMEDCT_CORE|Child abuse|Child abuse
C0008060|T048|FN|418189009|SNOMEDCT_CORE|Child abuse|Child abuse
C0008062|T048|SY|95922009|SNOMEDCT_CORE|CSA - Child sexual abuse|CSA - Child sexual abuse
C0008073|T048|PT|5294002|SNOMEDCT_CORE|Developmental disorder|Developmental disorder
C0008073|T048|FN|5294002|SNOMEDCT_CORE|Developmental disorder|Developmental disorder
C0008073|T048|IS|5294002|SNOMEDCT_CORE|Developmental disorder, NOS|Developmental disorder
C0008149|T047|PT|105629000|SNOMEDCT_CORE|Chlamydial infection|Chlamydial infection
C0008149|T047|FN|105629000|SNOMEDCT_CORE|Chlamydial infection|Chlamydial infection
C0008272|T047|SYGB|87522002|SNOMEDCT_CORE|Asiderotic anaemia|Asiderotic anemia
C0008272|T047|SY|87522002|SNOMEDCT_CORE|Asiderotic anemia|Asiderotic anemia
C0008272|T047|SYGB|87522002|SNOMEDCT_CORE|Chlorotic anaemia|Asiderotic anemia
C0008272|T047|SY|87522002|SNOMEDCT_CORE|Chlorotic anemia|Asiderotic anemia
C0008298|T191|PT|373610002|SNOMEDCT_CORE|Polyp in nasopharynx|Polyp in nasopharynx
C0008298|T191|FN|373610002|SNOMEDCT_CORE|Polyp in nasopharynx|Polyp in nasopharynx
C0008301|T046|PT|249489001|SNOMEDCT_CORE|Choking|Choking
C0008301|T046|FN|249489001|SNOMEDCT_CORE|Choking|Choking
C0008311|T047|PT|82403002|SNOMEDCT_CORE|Cholangitis|Cholangitis
C0008311|T047|FN|82403002|SNOMEDCT_CORE|Cholangitis|Cholangitis
C0008311|T047|IS|82403002|SNOMEDCT_CORE|Cholangitis, NOS|Cholangitis
C0008312|T047|SY|1761006|SNOMEDCT_CORE|Chronic nonsuppurative destructive cholangitis|Primary biliary cholangitis
C0008312|T047|SY|31712002|SNOMEDCT_CORE|Hanot's cirrhosis|Primary biliary cholangitis
C0008312|T047|IS|31712002|SNOMEDCT_CORE|PBC- Primary biliary cirrhosis|Primary biliary cholangitis
C0008312|T047|PT|31712002|SNOMEDCT_CORE|Primary biliary cholangitis|Primary biliary cholangitis
C0008312|T047|FN|31712002|SNOMEDCT_CORE|Primary biliary cholangitis|Primary biliary cholangitis
C0008312|T047|SY|31712002|SNOMEDCT_CORE|Primary biliary cirrhosis|Primary biliary cholangitis
C0008312|T047|OF|31712002|SNOMEDCT_CORE|Primary biliary cirrhosis|Primary biliary cholangitis
C0008313|T047|PT|235917005|SNOMEDCT_CORE|Sclerosing cholangitis|Sclerosing cholangitis
C0008313|T047|FN|235917005|SNOMEDCT_CORE|Sclerosing cholangitis|Sclerosing cholangitis
C0008325|T047|PT|76581006|SNOMEDCT_CORE|Cholecystitis|Cholecystitis
C0008325|T047|FN|76581006|SNOMEDCT_CORE|Cholecystitis|Cholecystitis
C0008325|T047|IS|76581006|SNOMEDCT_CORE|Cholecystitis, NOS|Cholecystitis
C0008325|T047|SY|76581006|SNOMEDCT_CORE|Inflamed gallbladder|Cholecystitis
C0008350|T047|PT|266474003|SNOMEDCT_CORE|Biliary calculus|Biliary calculus
C0008350|T047|SY|266474003|SNOMEDCT_CORE|Calculus - biliary|Biliary calculus
C0008350|T047|SY|266474003|SNOMEDCT_CORE|Calculus in biliary tract|Biliary calculus
C0008350|T047|FN|266474003|SNOMEDCT_CORE|Calculus in biliary tract|Biliary calculus
C0008350|T047|SY|266474003|SNOMEDCT_CORE|Cholelithiasis|Biliary calculus
C0008350|T047|SY|266474003|SNOMEDCT_CORE|CL - Cholelithiasis|Biliary calculus
C0008350|T047|SY|266474003|SNOMEDCT_CORE|Stone - biliary|Biliary calculus
C0008370|T047|SY|33688009|SNOMEDCT_CORE|Bile stasis|Cholestasis
C0008370|T047|IS|33688009|SNOMEDCT_CORE|Bile stasis, NOS|Cholestasis
C0008370|T047|PT|33688009|SNOMEDCT_CORE|Cholestasis|Cholestasis
C0008370|T047|FN|33688009|SNOMEDCT_CORE|Cholestasis|Cholestasis
C0008370|T047|IS|33688009|SNOMEDCT_CORE|Cholestasis, NOS|Cholestasis
C0008373|T047|PT|363668000|SNOMEDCT_CORE|Cholesteatoma|Cholesteatoma
C0008373|T047|FN|363668000|SNOMEDCT_CORE|Cholesteatoma|Cholesteatoma
C0008475|T047|IS|36071006|SNOMEDCT_CORE|Buedinger-Ludloff-Laewen disease|Chondromalacia of patella
C0008475|T047|PT|36071006|SNOMEDCT_CORE|Chondromalacia of patella|Chondromalacia of patella
C0008475|T047|FN|36071006|SNOMEDCT_CORE|Chondromalacia of patella|Chondromalacia of patella
C0008475|T047|SY|36071006|SNOMEDCT_CORE|Chondromalacia patella|Chondromalacia of patella
C0008475|T047|SY|36071006|SNOMEDCT_CORE|Chondromalacia patellae|Chondromalacia of patella
C0008475|T047|SY|36071006|SNOMEDCT_CORE|Degeneration of articular cartilage of patella|Chondromalacia of patella
C0008479|T191|PT|443520009|SNOMEDCT_CORE|Chondrosarcoma|Chondrosarcoma
C0008479|T191|SY|14990007|SNOMEDCT_CORE|Chondrosarcoma|Chondrosarcoma
C0008479|T191|OF|14990007|SNOMEDCT_CORE|Chondrosarcoma|Chondrosarcoma
C0008479|T191|FN|443520009|SNOMEDCT_CORE|Chondrosarcoma|Chondrosarcoma
C0008479|T191|SY|14990007|SNOMEDCT_CORE|Chondrosarcoma morphology|Chondrosarcoma
C0008479|T191|PT|14990007|SNOMEDCT_CORE|Chondrosarcoma, no ICD-O subtype|Chondrosarcoma
C0008479|T191|OF|14990007|SNOMEDCT_CORE|Chondrosarcoma, no ICD-O subtype|Chondrosarcoma
C0008479|T191|FN|14990007|SNOMEDCT_CORE|Chondrosarcoma, no International Classification of Diseases for Oncology subtype|Chondrosarcoma
C0008479|T191|SY|14990007|SNOMEDCT_CORE|Chondrosarcoma, no International Classification of Diseases for Oncology subtype|Chondrosarcoma
C0008479|T191|IS|14990007|SNOMEDCT_CORE|Chondrosarcoma, NOS|Chondrosarcoma
C0008479|T191|SY|443520009|SNOMEDCT_CORE|Fibrochondrosarcoma|Chondrosarcoma
C0008489|T047|PT|271700006|SNOMEDCT_CORE|Chorea|Chorea
C0008489|T047|FN|271700006|SNOMEDCT_CORE|Chorea|Chorea
C0008489|T047|IS|271700006|SNOMEDCT_CORE|Choreaform movement|Chorea
C0008489|T047|SY|271700006|SNOMEDCT_CORE|Choreic movement|Chorea
C0008489|T047|SY|271700006|SNOMEDCT_CORE|Choreiform movement|Chorea
C0008495|T047|PT|11612004|SNOMEDCT_CORE|Chorioamnionitis|Chorioamnionitis
C0008495|T047|FN|11612004|SNOMEDCT_CORE|Chorioamnionitis|Chorioamnionitis
C0008495|T047|SY|11612004|SNOMEDCT_CORE|Membranitis|Chorioamnionitis
C0008512|T020|PT|53854005|SNOMEDCT_CORE|Chorioretinal scar|Chorioretinal scar
C0008512|T020|FN|53854005|SNOMEDCT_CORE|Chorioretinal scar|Chorioretinal scar
C0008512|T020|IS|53854005|SNOMEDCT_CORE|Chorioretinal scar, NOS|Chorioretinal scar
C0008533|T047|SY|41788008|SNOMEDCT_CORE|Christmas disease|Hereditary factor IX deficiency disease
C0008533|T047|SY|41788008|SNOMEDCT_CORE|Congenital factor IX deficiency|Hereditary factor IX deficiency disease
C0008533|T047|IS|41788008|SNOMEDCT_CORE|Factor IX deficiency|Hereditary factor IX deficiency disease
C0008533|T047|SYGB|41788008|SNOMEDCT_CORE|Haemophilia B|Hereditary factor IX deficiency disease
C0008533|T047|IS|41788008|SNOMEDCT_CORE|Haemophilia B, NOS|Hereditary factor IX deficiency disease
C0008533|T047|SY|41788008|SNOMEDCT_CORE|Hemophilia B|Hereditary factor IX deficiency disease
C0008533|T047|OF|41788008|SNOMEDCT_CORE|Hemophilia B|Hereditary factor IX deficiency disease
C0008533|T047|IS|41788008|SNOMEDCT_CORE|Hemophilia B, NOS|Hereditary factor IX deficiency disease
C0008533|T047|PT|41788008|SNOMEDCT_CORE|Hereditary factor IX deficiency disease|Hereditary factor IX deficiency disease
C0008533|T047|FN|41788008|SNOMEDCT_CORE|Hereditary factor IX deficiency disease|Hereditary factor IX deficiency disease
C0008533|T047|SY|41788008|SNOMEDCT_CORE|PTC deficiency disease|Hereditary factor IX deficiency disease
C0008533|T047|SY|41788008|SNOMEDCT_CORE|Sex-linked factor IX deficiency disease|Hereditary factor IX deficiency disease
C0008626|T019|SY|74345006|SNOMEDCT_CORE|Anomaly of chromosome|Congenital chromosomal disease
C0008626|T019|IS|74345006|SNOMEDCT_CORE|Anomaly of chromosome, NOS|Congenital chromosomal disease
C0008626|T019|SY|74345006|SNOMEDCT_CORE|Chromosomal abnormality syndrome|Congenital chromosomal disease
C0008626|T019|IS|74345006|SNOMEDCT_CORE|Chromosomal abnormality syndrome, NOS|Congenital chromosomal disease
C0008626|T019|IS|74345006|SNOMEDCT_CORE|Chromosomal disease, NOS|Congenital chromosomal disease
C0008626|T019|SY|74345006|SNOMEDCT_CORE|Chromosomal hereditary disorder|Congenital chromosomal disease
C0008626|T019|IS|74345006|SNOMEDCT_CORE|Chromosomal hereditary disorder, NOS|Congenital chromosomal disease
C0008626|T019|SY|74345006|SNOMEDCT_CORE|Chromosomal imbalance syndrome|Congenital chromosomal disease
C0008626|T019|IS|74345006|SNOMEDCT_CORE|Chromosomal imbalance syndrome, NOS|Congenital chromosomal disease
C0008626|T019|SY|74345006|SNOMEDCT_CORE|Chromosomopathy|Congenital chromosomal disease
C0008626|T019|IS|74345006|SNOMEDCT_CORE|Chromosomopathy, NOS|Congenital chromosomal disease
C0008626|T019|PT|74345006|SNOMEDCT_CORE|Congenital chromosomal disease|Congenital chromosomal disease
C0008626|T019|FN|74345006|SNOMEDCT_CORE|Congenital disorder due to abnormality of chromosome number OR structure|Congenital chromosomal disease
C0008626|T019|SY|74345006|SNOMEDCT_CORE|Congenital disorder due to abnormality of chromosome number OR structure|Congenital chromosomal disease
C0008677|T047|PT|63480004|SNOMEDCT_CORE|Chronic bronchitis|Chronic bronchitis
C0008677|T047|FN|63480004|SNOMEDCT_CORE|Chronic bronchitis|Chronic bronchitis
C0008677|T047|IS|63480004|SNOMEDCT_CORE|Chronic bronchitis, NOS|Chronic bronchitis
C0008681|T047|PT|73237007|SNOMEDCT_CORE|Chronic ethmoidal sinusitis|Chronic ethmoidal sinusitis
C0008681|T047|FN|73237007|SNOMEDCT_CORE|Chronic ethmoidal sinusitis|Chronic ethmoidal sinusitis
C0008681|T047|SY|73237007|SNOMEDCT_CORE|Chronic ethmoiditis|Chronic ethmoidal sinusitis
C0008684|T047|PT|72621003|SNOMEDCT_CORE|Chronic gingivitis|Chronic gingivitis
C0008684|T047|FN|72621003|SNOMEDCT_CORE|Chronic gingivitis|Chronic gingivitis
C0008690|T047|PT|398155003|SNOMEDCT_CORE|Chronic anterior uveitis|Chronic anterior uveitis
C0008690|T047|FN|398155003|SNOMEDCT_CORE|Chronic anterior uveitis|Chronic anterior uveitis
C0008690|T047|SY|398155003|SNOMEDCT_CORE|Chronic iritis|Chronic anterior uveitis
C0008698|T047|SY|35923002|SNOMEDCT_CORE|Chronic antritis|Chronic maxillary sinusitis
C0008698|T047|PT|35923002|SNOMEDCT_CORE|Chronic maxillary sinusitis|Chronic maxillary sinusitis
C0008698|T047|FN|35923002|SNOMEDCT_CORE|Chronic maxillary sinusitis|Chronic maxillary sinusitis
C0008707|T047|PT|40970001|SNOMEDCT_CORE|Chronic osteomyelitis|Chronic osteomyelitis
C0008707|T047|FN|40970001|SNOMEDCT_CORE|Chronic osteomyelitis|Chronic osteomyelitis
C0008707|T047|IS|40970001|SNOMEDCT_CORE|Chronic osteomyelitis with or without periostitis|Chronic osteomyelitis
C0008707|T047|IS|40970001|SNOMEDCT_CORE|Chronic osteomyelitis, NOS|Chronic osteomyelitis
C0008711|T047|PT|86094006|SNOMEDCT_CORE|Chronic rhinitis|Chronic rhinitis
C0008711|T047|FN|86094006|SNOMEDCT_CORE|Chronic rhinitis|Chronic rhinitis
C0008728|T047|SY|82275008|SNOMEDCT_CORE|Allergic granulomatosis angiitis|Eosinophilic granulomatosis with polyangiitis
C0008728|T047|FN|82275008|SNOMEDCT_CORE|Allergic granulomatosis angiitis|Eosinophilic granulomatosis with polyangiitis
C0008728|T047|SY|82275008|SNOMEDCT_CORE|Allergic granulomatous angiitis|Eosinophilic granulomatosis with polyangiitis
C0008728|T047|SY|82275008|SNOMEDCT_CORE|Churg Strauss syndrome|Eosinophilic granulomatosis with polyangiitis
C0008728|T047|SY|82275008|SNOMEDCT_CORE|Churg-Strauss syndrome|Eosinophilic granulomatosis with polyangiitis
C0008728|T047|SY|82275008|SNOMEDCT_CORE|CSS - Churg-Strauss syndrome|Eosinophilic granulomatosis with polyangiitis
C0008728|T047|SY|82275008|SNOMEDCT_CORE|EGPA - eosinophilic granulomatosis with polyangiitis|Eosinophilic granulomatosis with polyangiitis
C0008728|T047|PT|82275008|SNOMEDCT_CORE|Eosinophilic granulomatosis with polyangiitis|Eosinophilic granulomatosis with polyangiitis
C0008827|T047|IS|19943007|SNOMEDCT_CORE|Cirrhosis of liver without mention of alcohol|Cirrhosis of liver without mention of alcohol
C0008909|T048|PT|19887002|SNOMEDCT_CORE|Claustrophobia|Claustrophobia
C0008909|T048|FN|19887002|SNOMEDCT_CORE|Claustrophobia|Claustrophobia
C0008909|T048|SY|19887002|SNOMEDCT_CORE|Fear of confined spaces|Claustrophobia
C0008925|T019|PT|87979003|SNOMEDCT_CORE|Cleft palate|Cleft palate
C0008925|T019|FN|87979003|SNOMEDCT_CORE|Cleft palate|Cleft palate
C0008925|T019|IS|87979003|SNOMEDCT_CORE|Cleft palate, NOS|Cleft palate
C0008925|T019|SY|87979003|SNOMEDCT_CORE|CP - Cleft palate|Cleft palate
C0008925|T019|SY|87979003|SNOMEDCT_CORE|Palatoschisis|Cleft palate
C0008925|T019|SY|87979003|SNOMEDCT_CORE|Uranoschisis|Cleft palate
C0009041|T037|OAP|63079007|SNOMEDCT_CORE|Closed dislocation of hip|Closed dislocation of hip
C0009041|T037|IS|63079007|SNOMEDCT_CORE|Closed dislocation of hip, NOS|Closed dislocation of hip
C0009044|T037|OP|9468002|SNOMEDCT_CORE|Closed fracture carpal bone|Closed fracture of carpal bone
C0009044|T037|OF|9468002|SNOMEDCT_CORE|Closed fracture carpal bone|Closed fracture of carpal bone
C0009044|T037|IS|9468002|SNOMEDCT_CORE|Closed fracture carpal bone, NOS|Closed fracture of carpal bone
C0009044|T037|PT|9468002|SNOMEDCT_CORE|Closed fracture of carpal bone|Closed fracture of carpal bone
C0009044|T037|FN|9468002|SNOMEDCT_CORE|Closed fracture of carpal bone|Closed fracture of carpal bone
C0009044|T037|SY|9468002|SNOMEDCT_CORE|Closed fracture of carpal bone of wrist|Closed fracture of carpal bone
C0009044|T037|IS|9468002|SNOMEDCT_CORE|Closed fracture of wrist|Closed fracture of carpal bone
C0009044|T037|IS|9468002|SNOMEDCT_CORE|Closed fracture of wrist, NOS|Closed fracture of carpal bone
C0009045|T037|IS|34649000|SNOMEDCT_CORE|Closed fracture of malar and maxillary bones, NOS|Closed fracture of malar AND/OR maxillary bones
C0009045|T037|PT|34649000|SNOMEDCT_CORE|Closed fracture of malar AND/OR maxillary bones|Closed fracture of malar AND/OR maxillary bones
C0009045|T037|FN|34649000|SNOMEDCT_CORE|Closed fracture of malar AND/OR maxillary bones|Closed fracture of malar AND/OR maxillary bones
C0009081|T019|SY|397932003|SNOMEDCT_CORE|Clubfoot|Talipes equinovarus
C0009081|T019|IS|397932003|SNOMEDCT_CORE|Clubfoot - congenital|Talipes equinovarus
C0009081|T019|IS|397932003|SNOMEDCT_CORE|Congenital clubfoot|Talipes equinovarus
C0009081|T019|IS|397932003|SNOMEDCT_CORE|Congenital talipes equinovarus|Talipes equinovarus
C0009081|T019|SY|397932003|SNOMEDCT_CORE|Equinovarus deformity|Talipes equinovarus
C0009081|T019|PT|397932003|SNOMEDCT_CORE|Talipes equinovarus|Talipes equinovarus
C0009081|T019|FN|397932003|SNOMEDCT_CORE|Talipes equinovarus|Talipes equinovarus
C0009081|T019|SY|397932003|SNOMEDCT_CORE|TEV - Talipes equinovarus|Talipes equinovarus
C0009088|T047|PT|193031009|SNOMEDCT_CORE|Cluster headache|Cluster headache
C0009088|T047|SY|193031009|SNOMEDCT_CORE|Cluster headache syndrome|Cluster headache
C0009088|T047|FN|193031009|SNOMEDCT_CORE|Cluster headache syndrome|Cluster headache
C0009088|T047|SY|193031009|SNOMEDCT_CORE|Histamine cephalgia|Cluster headache
C0009088|T047|SY|193031009|SNOMEDCT_CORE|Histamine headache|Cluster headache
C0009088|T047|SY|193031009|SNOMEDCT_CORE|Horton's headache|Cluster headache
C0009088|T047|SY|193031009|SNOMEDCT_CORE|Horton's neuralgia|Cluster headache
C0009088|T047|SY|193031009|SNOMEDCT_CORE|Migrainous neuralgia|Cluster headache
C0009088|T047|SY|193031009|SNOMEDCT_CORE|Neuralgic migraine|Cluster headache
C0009088|T047|SY|193031009|SNOMEDCT_CORE|Vasomotor headache|Cluster headache
C0009171|T048|PT|78267003|SNOMEDCT_CORE|Cocaine abuse|Cocaine abuse
C0009171|T048|FN|78267003|SNOMEDCT_CORE|Cocaine abuse|Cocaine abuse
C0009186|T047|PT|60826002|SNOMEDCT_CORE|Coccidioidomycosis|Coccidioidomycosis
C0009186|T047|FN|60826002|SNOMEDCT_CORE|Coccidioidomycosis|Coccidioidomycosis
C0009186|T047|SY|60826002|SNOMEDCT_CORE|Coccidioidomycosis infection|Coccidioidomycosis
C0009186|T047|IS|60826002|SNOMEDCT_CORE|Coccidioidomycosis, NOS|Coccidioidomycosis
C0009186|T047|IS|60826002|SNOMEDCT_CORE|Infection by Coccidioides immitis|Coccidioidomycosis
C0009186|T047|SY|60826002|SNOMEDCT_CORE|Posadas-Wernicke disease|Coccidioidomycosis
C0009193|T184|SY|34789001|SNOMEDCT_CORE|Coccyalgia|Pain in the coccyx
C0009193|T184|SY|34789001|SNOMEDCT_CORE|Coccydynia|Pain in the coccyx
C0009193|T184|SY|34789001|SNOMEDCT_CORE|Coccygalgia|Pain in the coccyx
C0009193|T184|IS|34789001|SNOMEDCT_CORE|Coccygodynia|Pain in the coccyx
C0009193|T184|SY|34789001|SNOMEDCT_CORE|Coccyodynia|Pain in the coccyx
C0009193|T184|FN|34789001|SNOMEDCT_CORE|Pain in the coccyx|Pain in the coccyx
C0009193|T184|PT|34789001|SNOMEDCT_CORE|Pain in the coccyx|Pain in the coccyx
C0009241|T048|PT|443265004|SNOMEDCT_CORE|Cognitive disorder|Cognitive disorder
C0009241|T048|FN|443265004|SNOMEDCT_CORE|Cognitive disorder|Cognitive disorder
C0009250|T047|PT|308689002|SNOMEDCT_CORE|Coin lesion of lung|Coin lesion of lung
C0009250|T047|FN|308689002|SNOMEDCT_CORE|Coin lesion of lung|Coin lesion of lung
C0009269|T033|SY|80585000|SNOMEDCT_CORE|Chilly person|Intolerant of cold
C0009269|T033|IS|80585000|SNOMEDCT_CORE|Cold intolerance|Intolerant of cold
C0009269|T033|SY|80585000|SNOMEDCT_CORE|Cold sensitivity|Intolerant of cold
C0009269|T033|SY|80585000|SNOMEDCT_CORE|Feels the cold|Intolerant of cold
C0009269|T033|PT|80585000|SNOMEDCT_CORE|Intolerant of cold|Intolerant of cold
C0009269|T033|FN|80585000|SNOMEDCT_CORE|Intolerant of cold|Intolerant of cold
C0009269|T033|SY|80585000|SNOMEDCT_CORE|Sensitive to cold|Intolerant of cold
C0009319|T047|PT|64226004|SNOMEDCT_CORE|Colitis|Colitis
C0009319|T047|FN|64226004|SNOMEDCT_CORE|Colitis|Colitis
C0009319|T047|IS|64226004|SNOMEDCT_CORE|Colitis, NOS|Colitis
C0009319|T047|SY|64226004|SNOMEDCT_CORE|Colon inflammation|Colitis
C0009324|T047|SY|64766004|SNOMEDCT_CORE|Colitis gravis|Ulcerative colitis
C0009324|T047|IS|64766004|SNOMEDCT_CORE|Colitis gravis, NOS|Ulcerative colitis
C0009324|T047|SY|64766004|SNOMEDCT_CORE|Idiopathic proctocolitis|Ulcerative colitis
C0009324|T047|SY|64766004|SNOMEDCT_CORE|UC - Ulcerative colitis|Ulcerative colitis
C0009324|T047|PT|64766004|SNOMEDCT_CORE|Ulcerative colitis|Ulcerative colitis
C0009324|T047|FN|64766004|SNOMEDCT_CORE|Ulcerative colitis|Ulcerative colitis
C0009324|T047|IS|64766004|SNOMEDCT_CORE|Ulcerative colitis, NOS|Ulcerative colitis
C0009326|T047|PT|81573002|SNOMEDCT_CORE|Collagen disease|Collagen disease
C0009326|T047|FN|81573002|SNOMEDCT_CORE|Collagen disease|Collagen disease
C0009326|T047|IS|81573002|SNOMEDCT_CORE|Collagen disease, NOS|Collagen disease
C0009326|T047|SY|81573002|SNOMEDCT_CORE|Collagen disorder|Collagen disease
C0009326|T047|IS|81573002|SNOMEDCT_CORE|Collagen disorder, NOS|Collagen disease
C0009354|T037|PT|269083002|SNOMEDCT_CORE|Closed Colles' fracture|Closed Colles' fracture
C0009354|T037|FN|269083002|SNOMEDCT_CORE|Closed Colles' fracture|Closed Colles' fracture
C0009376|T190|SY|68496003|SNOMEDCT_CORE|Colonic polyp|Polyp of colon
C0009376|T190|IS|68496003|SNOMEDCT_CORE|Colonic polyp, NOS|Polyp of colon
C0009376|T190|SY|68496003|SNOMEDCT_CORE|Polyp colon|Polyp of colon
C0009376|T190|PT|68496003|SNOMEDCT_CORE|Polyp of colon|Polyp of colon
C0009376|T190|FN|68496003|SNOMEDCT_CORE|Polyp of colon|Polyp of colon
C0009376|T190|IS|68496003|SNOMEDCT_CORE|Polyp of colon, NOS|Polyp of colon
C0009377|T047|PT|35065006|SNOMEDCT_CORE|Primary chronic pseudo-obstruction of colon|Primary chronic pseudo-obstruction of colon
C0009377|T047|FN|35065006|SNOMEDCT_CORE|Primary chronic pseudo-obstruction of colon|Primary chronic pseudo-obstruction of colon
C0009443|T047|SY|82272006|SNOMEDCT_CORE|Acute coryza|Common cold
C0009443|T047|SY|82272006|SNOMEDCT_CORE|Acute infective rhinitis|Common cold
C0009443|T047|SY|82272006|SNOMEDCT_CORE|Acute nasal catarrh|Common cold
C0009443|T047|SY|82272006|SNOMEDCT_CORE|Acute nasopharyngitis|Common cold
C0009443|T047|IS|82272006|SNOMEDCT_CORE|Acute nasopharyngitis, NOS|Common cold
C0009443|T047|SY|82272006|SNOMEDCT_CORE|Acute rhinitis|Common cold
C0009443|T047|SY|82272006|SNOMEDCT_CORE|Cold|Common cold
C0009443|T047|PT|82272006|SNOMEDCT_CORE|Common cold|Common cold
C0009443|T047|FN|82272006|SNOMEDCT_CORE|Common cold|Common cold
C0009443|T047|SY|82272006|SNOMEDCT_CORE|Head cold|Common cold
C0009443|T047|IS|54150009|SNOMEDCT_CORE|Head cold, NOS|Common cold
C0009443|T047|SY|82272006|SNOMEDCT_CORE|Infective nasopharyngitis|Common cold
C0009443|T047|IS|82272006|SNOMEDCT_CORE|Infective nasopharyngitis, NOS|Common cold
C0009443|T047|SY|82272006|SNOMEDCT_CORE|Infective rhinitis|Common cold
C0009447|T047|PTGB|23238000|SNOMEDCT_CORE|Common variable agammaglobulinaemia|Common variable agammaglobulinemia
C0009447|T047|PT|23238000|SNOMEDCT_CORE|Common variable agammaglobulinemia|Common variable agammaglobulinemia
C0009447|T047|FN|23238000|SNOMEDCT_CORE|Common variable agammaglobulinemia|Common variable agammaglobulinemia
C0009447|T047|SYGB|23238000|SNOMEDCT_CORE|Common variable hypogammaglobulinaemia|Common variable agammaglobulinemia
C0009447|T047|SY|23238000|SNOMEDCT_CORE|Common variable hypogammaglobulinemia|Common variable agammaglobulinemia
C0009447|T047|SY|23238000|SNOMEDCT_CORE|Common variable immunodeficiency|Common variable agammaglobulinemia
C0009447|T047|SY|23238000|SNOMEDCT_CORE|CVAG|Common variable agammaglobulinemia
C0009447|T047|SY|23238000|SNOMEDCT_CORE|CVI - Common variable immunodeficiency|Common variable agammaglobulinemia
C0009447|T047|SY|23238000|SNOMEDCT_CORE|CVID - Common variable immunodeficiency|Common variable agammaglobulinemia
C0009447|T047|SY|23238000|SNOMEDCT_CORE|Late onset immunoglobulin deficiency|Common variable agammaglobulinemia
C0009450|T047|PT|191415002|SNOMEDCT_CORE|Communicable disease|Disorder due to infection
C0009450|T047|OF|191415002|SNOMEDCT_CORE|Communicable disease|Disorder due to infection
C0009450|T047|FN|191415002|SNOMEDCT_CORE|Communicable disease|Disorder due to infection
C0009450|T047|SY|40733004|SNOMEDCT_CORE|Disease due to infection|Disorder due to infection
C0009450|T047|PT|40733004|SNOMEDCT_CORE|Disorder due to infection|Disorder due to infection
C0009450|T047|SY|40733004|SNOMEDCT_CORE|Infection|Disorder due to infection
C0009450|T047|IS|40733004|SNOMEDCT_CORE|Infection, NOS|Disorder due to infection
C0009450|T047|SY|40733004|SNOMEDCT_CORE|Infectious disease|Disorder due to infection
C0009450|T047|FN|40733004|SNOMEDCT_CORE|Infectious disease|Disorder due to infection
C0009450|T047|IS|40733004|SNOMEDCT_CORE|Infectious disease, NOS|Disorder due to infection
C0009450|T047|SY|40733004|SNOMEDCT_CORE|Infective disorder|Disorder due to infection
C0009451|T047|PT|271569006|SNOMEDCT_CORE|Communicating hydrocephalus|Communicating hydrocephalus
C0009451|T047|FN|271569006|SNOMEDCT_CORE|Communicating hydrocephalus|Communicating hydrocephalus
C0009492|T047|PT|111245009|SNOMEDCT_CORE|Compartment syndrome|Compartment syndrome
C0009492|T047|FN|111245009|SNOMEDCT_CORE|Compartment syndrome|Compartment syndrome
C0009492|T047|IS|111245009|SNOMEDCT_CORE|Compartment syndrome, NOS|Compartment syndrome
C0009492|T047|IS|45781009|SNOMEDCT_CORE|Compartment syndrome, NOS|Compartment syndrome
C0009492|T047|IS|111245009|SNOMEDCT_CORE|Compartmental syndrome, NOS|Compartment syndrome
C0009492|T047|IS|45781009|SNOMEDCT_CORE|Compartmental syndrome, NOS|Compartment syndrome
C0009595|T048|SY|1376001|SNOMEDCT_CORE|Anancastic personality disorder|Obsessive compulsive personality disorder
C0009595|T048|SY|1376001|SNOMEDCT_CORE|Anankastic personality disorder|Obsessive compulsive personality disorder
C0009595|T048|IS|1376001|SNOMEDCT_CORE|Obsessional personality|Obsessive compulsive personality disorder
C0009595|T048|IS|1376001|SNOMEDCT_CORE|Obsessional personality disorder|Obsessive compulsive personality disorder
C0009595|T048|PT|1376001|SNOMEDCT_CORE|Obsessive compulsive personality disorder|Obsessive compulsive personality disorder
C0009595|T048|FN|1376001|SNOMEDCT_CORE|Obsessive compulsive personality disorder|Obsessive compulsive personality disorder
C0009663|T047|SY|240542006|SNOMEDCT_CORE|AGW - Anogenital warts|Genital warts
C0009663|T047|SY|240542006|SNOMEDCT_CORE|Anogenital wart|Genital warts
C0009663|T047|SY|240542006|SNOMEDCT_CORE|Anogenital warts|Genital warts
C0009663|T047|FN|240542006|SNOMEDCT_CORE|Anogenital warts|Genital warts
C0009663|T047|IS|240542006|SNOMEDCT_CORE|Condyloma acuminatum|Genital warts
C0009663|T047|PT|240542006|SNOMEDCT_CORE|Condyloma acuminatum of the anogenital region|Genital warts
C0009663|T047|IS|240542006|SNOMEDCT_CORE|Condylomata acuminata|Genital warts
C0009663|T047|IS|240542006|SNOMEDCT_CORE|Condylomata acuminatum|Genital warts
C0009663|T047|SY|240542006|SNOMEDCT_CORE|Condylomata acuminatum of the anogenital region|Genital warts
C0009663|T047|SY|266113007|SNOMEDCT_CORE|Genital wart|Genital warts
C0009663|T047|PT|266113007|SNOMEDCT_CORE|Genital warts|Genital warts
C0009663|T047|FN|266113007|SNOMEDCT_CORE|Genital warts|Genital warts
C0009663|T047|SY|240542006|SNOMEDCT_CORE|Venereal wart|Genital warts
C0009663|T047|SY|240542006|SNOMEDCT_CORE|Venereal warts|Genital warts
C0009663|T047|SY|240542006|SNOMEDCT_CORE|Verruca acuminata|Genital warts
C0009691|T019|PT|79410001|SNOMEDCT_CORE|Congenital cataract|Congenital cataract
C0009691|T019|FN|79410001|SNOMEDCT_CORE|Congenital cataract|Congenital cataract
C0009691|T019|IS|79410001|SNOMEDCT_CORE|Congenital cataract, NOS|Congenital cataract
C0009702|T019|OAP|33543001|SNOMEDCT_CORE|Unilateral congenital dislocation of hip|Unilateral congenital dislocation of hip
C0009702|T019|OF|33543001|SNOMEDCT_CORE|Unilateral congenital dislocation of hip|Unilateral congenital dislocation of hip
C0009702|T019|OAF|33543001|SNOMEDCT_CORE|Unilateral congenital dislocation of hip|Unilateral congenital dislocation of hip
C0009726|T019|SY|205564003|SNOMEDCT_CORE|Congenital pigmentary anomaly of skin|Congenital pigmentary skin anomalies
C0009726|T019|PT|205564003|SNOMEDCT_CORE|Congenital pigmentary skin anomalies|Congenital pigmentary skin anomalies
C0009726|T019|FN|205564003|SNOMEDCT_CORE|Congenital pigmentary skin anomalies|Congenital pigmentary skin anomalies
C0009759|T047|SY|59698003|SNOMEDCT_CORE|Disease of conjunctiva|Disorder of conjunctiva
C0009759|T047|PT|59698003|SNOMEDCT_CORE|Disorder of conjunctiva|Disorder of conjunctiva
C0009759|T047|FN|59698003|SNOMEDCT_CORE|Disorder of conjunctiva|Disorder of conjunctiva
C0009759|T047|IS|59698003|SNOMEDCT_CORE|Disorder of conjunctiva, NOS|Disorder of conjunctiva
C0009760|T046|PTGB|21117005|SNOMEDCT_CORE|Conjunctival haemorrhage|Conjunctival hemorrhage
C0009760|T046|PT|21117005|SNOMEDCT_CORE|Conjunctival hemorrhage|Conjunctival hemorrhage
C0009760|T046|FN|21117005|SNOMEDCT_CORE|Conjunctival hemorrhage|Conjunctival hemorrhage
C0009763|T047|PT|9826008|SNOMEDCT_CORE|Conjunctivitis|Conjunctivitis
C0009763|T047|FN|9826008|SNOMEDCT_CORE|Conjunctivitis|Conjunctivitis
C0009763|T047|IS|9826008|SNOMEDCT_CORE|Conjunctivitis, NOS|Conjunctivitis
C0009763|T047|SY|9826008|SNOMEDCT_CORE|Inflammation of conjunctiva|Conjunctivitis
C0009763|T047|SY|9826008|SNOMEDCT_CORE|Pink eye disease|Conjunctivitis
C0009766|T047|IS|231854006|SNOMEDCT_CORE|Allergic conjunctivitis|Atopic conjunctivitis
C0009766|T047|PT|231854006|SNOMEDCT_CORE|Atopic conjunctivitis|Atopic conjunctivitis
C0009766|T047|FN|231854006|SNOMEDCT_CORE|Atopic conjunctivitis|Atopic conjunctivitis
C0009768|T047|PT|128350005|SNOMEDCT_CORE|Bacterial conjunctivitis|Bacterial conjunctivitis
C0009768|T047|FN|128350005|SNOMEDCT_CORE|Bacterial conjunctivitis|Bacterial conjunctivitis
C0009769|T047|PT|231857004|SNOMEDCT_CORE|Giant papillary conjunctivitis|Giant papillary conjunctivitis
C0009769|T047|FN|231857004|SNOMEDCT_CORE|Giant papillary conjunctivitis|Giant papillary conjunctivitis
C0009769|T047|SY|231857004|SNOMEDCT_CORE|GPC - Giant papillary conjunctivitis|Giant papillary conjunctivitis
C0009773|T047|SY|318316003|SNOMEDCT_CORE|Spring conjunctivitis|Vernal conjunctivitis
C0009773|T047|SY|318316003|SNOMEDCT_CORE|Spring ophthalmia|Vernal conjunctivitis
C0009773|T047|PT|318316003|SNOMEDCT_CORE|Vernal conjunctivitis|Vernal conjunctivitis
C0009773|T047|FN|318316003|SNOMEDCT_CORE|Vernal conjunctivitis|Vernal conjunctivitis
C0009774|T047|PT|45261009|SNOMEDCT_CORE|Viral conjunctivitis|Viral conjunctivitis
C0009774|T047|FN|45261009|SNOMEDCT_CORE|Viral conjunctivitis|Viral conjunctivitis
C0009774|T047|IS|45261009|SNOMEDCT_CORE|Viral conjunctivitis, NOS|Viral conjunctivitis
C0009782|T047|SY|105969002|SNOMEDCT_CORE|Connective tissue disease|Disorder of connective tissue
C0009782|T047|IS|105969002|SNOMEDCT_CORE|Disease of connective tissues|Disorder of connective tissue
C0009782|T047|OF|105969002|SNOMEDCT_CORE|Disease of connective tissues|Disorder of connective tissue
C0009782|T047|PT|105969002|SNOMEDCT_CORE|Disorder of connective tissue|Disorder of connective tissue
C0009782|T047|FN|105969002|SNOMEDCT_CORE|Disorder of connective tissue|Disorder of connective tissue
C0009806|T184|SY|14760008|SNOMEDCT_CORE|CN - Constipation|Constipation
C0009806|T184|SY|14760008|SNOMEDCT_CORE|Constipated|Constipation
C0009806|T184|PT|14760008|SNOMEDCT_CORE|Constipation|Constipation
C0009806|T184|OF|14760008|SNOMEDCT_CORE|Constipation|Constipation
C0009806|T184|FN|14760008|SNOMEDCT_CORE|Constipation|Constipation
C0009806|T184|SY|14760008|SNOMEDCT_CORE|Costiveness|Constipation
C0009806|T184|SY|14760008|SNOMEDCT_CORE|Difficult passing motion|Constipation
C0009806|T184|SYGB|14760008|SNOMEDCT_CORE|Difficulty defaecating|Constipation
C0009806|T184|SY|14760008|SNOMEDCT_CORE|Difficulty defecating|Constipation
C0009806|T184|SY|14760008|SNOMEDCT_CORE|Difficulty opening bowels|Constipation
C0009806|T184|SY|14760008|SNOMEDCT_CORE|Difficulty passing stool|Constipation
C0009918|T190|PT|7890003|SNOMEDCT_CORE|Contracture of joint|Contracture of joint
C0009918|T190|FN|7890003|SNOMEDCT_CORE|Contracture of joint|Contracture of joint
C0009918|T190|IS|7890003|SNOMEDCT_CORE|Contracture of joint, NOS|Contracture of joint
C0009918|T190|SY|7890003|SNOMEDCT_CORE|Joint contraction|Contracture of joint
C0009938|T037|SY|125667009|SNOMEDCT_CORE|Bruise|Contusion
C0009938|T037|SY|125667009|SNOMEDCT_CORE|Bruising|Contusion
C0009938|T037|PT|125667009|SNOMEDCT_CORE|Contusion|Contusion
C0009938|T037|FN|125667009|SNOMEDCT_CORE|Contusion|Contusion
C0009946|T048|SY|20734000|SNOMEDCT_CORE|Conversion disorder|Psychologic conversion disorder
C0009946|T048|PT|20734000|SNOMEDCT_CORE|Psychologic conversion disorder|Psychologic conversion disorder
C0009946|T048|FN|20734000|SNOMEDCT_CORE|Psychologic conversion disorder|Psychologic conversion disorder
C0009946|T048|OF|20734000|SNOMEDCT_CORE|Psychologic conversion disorder|Psychologic conversion disorder
C0009946|T048|IS|20734000|SNOMEDCT_CORE|Psychologic conversion disorder, NOS|Psychologic conversion disorder
C0009952|T047|PT|41497008|SNOMEDCT_CORE|Febrile convulsion|Febrile convulsion
C0009952|T047|FN|41497008|SNOMEDCT_CORE|Febrile convulsion|Febrile convulsion
C0009952|T047|SY|41497008|SNOMEDCT_CORE|Febrile fit|Febrile convulsion
C0009952|T047|SY|41497008|SNOMEDCT_CORE|Febrile seizure|Febrile convulsion
C0009952|T047|SY|41497008|SNOMEDCT_CORE|Fever seizure|Febrile convulsion
C0009952|T047|SY|41497008|SNOMEDCT_CORE|Pyrexial convulsion|Febrile convulsion
C0010032|T037|SY|85848002|SNOMEDCT_CORE|CA - Corneal abrasion|Corneal abrasion
C0010032|T037|PT|85848002|SNOMEDCT_CORE|Corneal abrasion|Corneal abrasion
C0010032|T037|FN|85848002|SNOMEDCT_CORE|Corneal abrasion|Corneal abrasion
C0010032|T037|SY|85848002|SNOMEDCT_CORE|Scratch of cornea|Corneal abrasion
C0010032|T037|SY|85848002|SNOMEDCT_CORE|Scratch to cornea|Corneal abrasion
C0010034|T047|SY|15250008|SNOMEDCT_CORE|Corneal disorder|Disorder of cornea
C0010034|T047|IS|15250008|SNOMEDCT_CORE|Disease of cornea|Disorder of cornea
C0010034|T047|OF|15250008|SNOMEDCT_CORE|Disease of cornea|Disorder of cornea
C0010034|T047|IS|15250008|SNOMEDCT_CORE|Disease of cornea, NOS|Disorder of cornea
C0010034|T047|PT|15250008|SNOMEDCT_CORE|Disorder of cornea|Disorder of cornea
C0010034|T047|FN|15250008|SNOMEDCT_CORE|Disorder of cornea|Disorder of cornea
C0010034|T047|IS|15250008|SNOMEDCT_CORE|Disorder of cornea, NOS|Disorder of cornea
C0010035|T047|PT|77797009|SNOMEDCT_CORE|Hereditary corneal dystrophy|Hereditary corneal dystrophy
C0010035|T047|FN|77797009|SNOMEDCT_CORE|Hereditary corneal dystrophy|Hereditary corneal dystrophy
C0010035|T047|IS|77797009|SNOMEDCT_CORE|Hereditary corneal dystrophy, NOS|Hereditary corneal dystrophy
C0010037|T046|PT|27194006|SNOMEDCT_CORE|Corneal edema|Corneal edema
C0010037|T046|FN|27194006|SNOMEDCT_CORE|Corneal edema|Corneal edema
C0010037|T046|IS|27194006|SNOMEDCT_CORE|Corneal edema, NOS|Corneal edema
C0010037|T046|PTGB|27194006|SNOMEDCT_CORE|Corneal oedema|Corneal edema
C0010038|T033|PT|64634000|SNOMEDCT_CORE|Corneal opacity|Corneal opacity
C0010038|T033|FN|64634000|SNOMEDCT_CORE|Corneal opacity|Corneal opacity
C0010038|T033|IS|64634000|SNOMEDCT_CORE|Corneal opacity, NOS|Corneal opacity
C0010043|T047|PT|91514001|SNOMEDCT_CORE|Corneal ulcer|Corneal ulcer
C0010043|T047|FN|91514001|SNOMEDCT_CORE|Corneal ulcer|Corneal ulcer
C0010043|T047|IS|91514001|SNOMEDCT_CORE|Corneal ulcer, NOS|Corneal ulcer
C0010046|T020|IS|46014006|SNOMEDCT_CORE|Clavus|Corn of toe
C0010046|T020|SY|201038005|SNOMEDCT_CORE|Clavus|Corn of toe
C0010046|T020|SY|201038005|SNOMEDCT_CORE|Corn|Corn of toe
C0010046|T020|FN|201038005|SNOMEDCT_CORE|Corn - lesion|Corn of toe
C0010046|T020|PT|201038005|SNOMEDCT_CORE|Corn - lesion|Corn of toe
C0010046|T020|PT|46014006|SNOMEDCT_CORE|Corn of toe|Corn of toe
C0010046|T020|FN|46014006|SNOMEDCT_CORE|Corn of toe|Corn of toe
C0010054|T047|SY|53741008|SNOMEDCT_CORE|Arteriosclerotic heart disease|Coronary atherosclerosis
C0010054|T047|IS|53741008|SNOMEDCT_CORE|ASHD - Atherosclerotic heart disease|Coronary atherosclerosis
C0010054|T047|SY|443502000|SNOMEDCT_CORE|Atherosclerosis of coronary artery|Coronary atherosclerosis
C0010054|T047|FN|443502000|SNOMEDCT_CORE|Atherosclerosis of coronary artery|Coronary atherosclerosis
C0010054|T047|SY|443502000|SNOMEDCT_CORE|Atherosclerosis of native coronary artery|Coronary atherosclerosis
C0010054|T047|IS|53741008|SNOMEDCT_CORE|Atherosclerotic heart disease|Coronary atherosclerosis
C0010054|T047|PT|53741008|SNOMEDCT_CORE|Coronary arteriosclerosis|Coronary atherosclerosis
C0010054|T047|FN|53741008|SNOMEDCT_CORE|Coronary arteriosclerosis|Coronary atherosclerosis
C0010054|T047|PT|443502000|SNOMEDCT_CORE|Coronary atherosclerosis|Coronary atherosclerosis
C0010054|T047|SY|53741008|SNOMEDCT_CORE|Coronary sclerosis|Coronary atherosclerosis
C0010068|T047|SY|53741008|SNOMEDCT_CORE|CHD - Coronary heart disease|Coronary heart disease
C0010068|T047|SY|53741008|SNOMEDCT_CORE|Coronary heart disease|Coronary heart disease
C0010073|T047|PT|23687008|SNOMEDCT_CORE|Coronary artery spasm|Coronary artery spasm
C0010073|T047|FN|23687008|SNOMEDCT_CORE|Coronary artery spasm|Coronary artery spasm
C0010073|T047|SY|23687008|SNOMEDCT_CORE|Coronary spasm|Coronary artery spasm
C0010093|T047|PT|386762009|SNOMEDCT_CORE|Corpus luteum cyst|Corpus luteum cyst
C0010093|T047|FN|386762009|SNOMEDCT_CORE|Corpus luteum cyst|Corpus luteum cyst
C0010093|T047|SY|386762009|SNOMEDCT_CORE|Lutein cyst|Corpus luteum cyst
C0010200|T184|PT|49727002|SNOMEDCT_CORE|Cough|Cough
C0010200|T184|FN|49727002|SNOMEDCT_CORE|Cough|Cough
C0010200|T184|IS|49727002|SNOMEDCT_CORE|Cough, NOS|Cough
C0010200|T184|IS|49727002|SNOMEDCT_CORE|Finding of cough|Cough
C0010200|T184|SY|49727002|SNOMEDCT_CORE|Observation of cough|Cough
C0010201|T184|PT|68154008|SNOMEDCT_CORE|Chronic cough|Chronic cough
C0010201|T184|FN|68154008|SNOMEDCT_CORE|Chronic cough|Chronic cough
C0010246|T047|PT|186658007|SNOMEDCT_CORE|Coxsackie virus disease|Coxsackie virus disease
C0010246|T047|FN|186658007|SNOMEDCT_CORE|Coxsackie virus disease|Coxsackie virus disease
C0010263|T184|SY|424647005|SNOMEDCT_CORE|Cramp in extremity|Cramp in limb
C0010263|T184|PT|424647005|SNOMEDCT_CORE|Cramp in limb|Cramp in limb
C0010263|T184|FN|424647005|SNOMEDCT_CORE|Cramp in limb|Cramp in limb
C0010276|T191|PT|189179009|SNOMEDCT_CORE|Craniopharyngioma|Craniopharyngioma
C0010276|T191|FN|189179009|SNOMEDCT_CORE|Craniopharyngioma|Craniopharyngioma
C0010278|T047|SY|57219006|SNOMEDCT_CORE|Congenital ossification of cranial sutures|Craniosynostosis syndrome
C0010278|T047|SY|57219006|SNOMEDCT_CORE|Congenital ossification of sutures of skull|Craniosynostosis syndrome
C0010278|T047|SY|57219006|SNOMEDCT_CORE|Craniostenosis|Craniosynostosis syndrome
C0010278|T047|SY|57219006|SNOMEDCT_CORE|Craniostosis|Craniosynostosis syndrome
C0010278|T047|SY|57219006|SNOMEDCT_CORE|Craniosynostosis|Craniosynostosis syndrome
C0010278|T047|PT|57219006|SNOMEDCT_CORE|Craniosynostosis syndrome|Craniosynostosis syndrome
C0010278|T047|FN|57219006|SNOMEDCT_CORE|Craniosynostosis syndrome|Craniosynostosis syndrome
C0010278|T047|SY|57219006|SNOMEDCT_CORE|CSO - Craniosynostosis|Craniosynostosis syndrome
C0010278|T047|SY|57219006|SNOMEDCT_CORE|Premature closure of cranial sutures|Craniosynostosis syndrome
C0010278|T047|SY|57219006|SNOMEDCT_CORE|Premature cranial suture closure|Craniosynostosis syndrome
C0010308|T047|IS|217710005|SNOMEDCT_CORE|CHT - Congenital hypothyroidism|Cretinism
C0010308|T047|SY|217710005|SNOMEDCT_CORE|Congenital goiter|Cretinism
C0010308|T047|SYGB|217710005|SNOMEDCT_CORE|Congenital goitre|Cretinism
C0010308|T047|IS|217710005|SNOMEDCT_CORE|Congenital hypothyroidism|Cretinism
C0010308|T047|SY|217710005|SNOMEDCT_CORE|Congenital hypothyroidism not due to iodine deficiency|Cretinism
C0010308|T047|SY|217710005|SNOMEDCT_CORE|Cretinism|Cretinism
C0010308|T047|SY|217710005|SNOMEDCT_CORE|Infantile hypothyroidism|Cretinism
C0010346|T047|SY|34000006|SNOMEDCT_CORE|CD - Crohn's disease|Crohn's disease
C0010346|T047|SY|34000006|SNOMEDCT_CORE|Crohn disease|Crohn's disease
C0010346|T047|PT|34000006|SNOMEDCT_CORE|Crohn's disease|Crohn's disease
C0010346|T047|FN|34000006|SNOMEDCT_CORE|Crohn's disease|Crohn's disease
C0010346|T047|IS|34000006|SNOMEDCT_CORE|Crohn's disease, NOS|Crohn's disease
C0010346|T047|SY|34000006|SNOMEDCT_CORE|Crohn's regional enteritis|Crohn's disease
C0010346|T047|SY|34000006|SNOMEDCT_CORE|Crohns disease|Crohn's disease
C0010346|T047|SY|34000006|SNOMEDCT_CORE|Granulomatous enteritis|Crohn's disease
C0010346|T047|IS|34000006|SNOMEDCT_CORE|Granulomatous enteritis, NOS|Crohn's disease
C0010346|T047|SY|34000006|SNOMEDCT_CORE|RE - regional enteritis|Crohn's disease
C0010346|T047|IS|34000006|SNOMEDCT_CORE|RE - Regional enteritis|Crohn's disease
C0010346|T047|SY|34000006|SNOMEDCT_CORE|Regional enteritis|Crohn's disease
C0010346|T047|IS|34000006|SNOMEDCT_CORE|Regional enteritis, NOS|Crohn's disease
C0010380|T047|PT|71186008|SNOMEDCT_CORE|Croup|Croup
C0010380|T047|FN|71186008|SNOMEDCT_CORE|Croup|Croup
C0010380|T047|SY|71186008|SNOMEDCT_CORE|Croup syndrome|Croup
C0010403|T047|PTGB|30911005|SNOMEDCT_CORE|Cryoglobulinaemia|Cryoglobulinemia
C0010403|T047|IS|30911005|SNOMEDCT_CORE|Cryoglobulinaemia, NOS|Cryoglobulinemia
C0010403|T047|PT|30911005|SNOMEDCT_CORE|Cryoglobulinemia|Cryoglobulinemia
C0010403|T047|FN|30911005|SNOMEDCT_CORE|Cryoglobulinemia|Cryoglobulinemia
C0010403|T047|IS|30911005|SNOMEDCT_CORE|Cryoglobulinemia, NOS|Cryoglobulinemia
C0010403|T047|SYGB|30911005|SNOMEDCT_CORE|Cryoimmunoglobulinaemia|Cryoglobulinemia
C0010403|T047|SY|30911005|SNOMEDCT_CORE|Cryoimmunoglobulinemia|Cryoglobulinemia
C0010403|T047|IS|30911005|SNOMEDCT_CORE|Cryoimmunoglobulinemia, NOS|Cryoglobulinemia
C0010417|T019|SY|204878001|SNOMEDCT_CORE|Cryptorchidism|Undescended testicle
C0010417|T019|SY|204878001|SNOMEDCT_CORE|Cryptorchism|Undescended testicle
C0010417|T019|SY|204878001|SNOMEDCT_CORE|IDT - Imperfectly descended testis|Undescended testicle
C0010417|T019|SY|204878001|SNOMEDCT_CORE|Imperfectly descended testis|Undescended testicle
C0010417|T019|SY|204878001|SNOMEDCT_CORE|Maldescent of testis|Undescended testicle
C0010417|T019|SY|204878001|SNOMEDCT_CORE|UDT - Undescended testes|Undescended testicle
C0010417|T019|PT|204878001|SNOMEDCT_CORE|Undescended testicle|Undescended testicle
C0010417|T019|FN|204878001|SNOMEDCT_CORE|Undescended testicle|Undescended testicle
C0010417|T019|SY|204878001|SNOMEDCT_CORE|Undescended testis|Undescended testicle
C0010481|T047|SY|47270006|SNOMEDCT_CORE|Cushing's syndrome|Cushing's syndrome III
C0010481|T047|SY|47270006|SNOMEDCT_CORE|Cushing's syndrome III|Cushing's syndrome III
C0010481|T047|SY|47270006|SNOMEDCT_CORE|Itsenko disease|Cushing's syndrome III
C0010481|T047|SY|47270006|SNOMEDCT_CORE|Itsenko-Cushing syndrome|Cushing's syndrome III
C0010481|T047|SY|47270006|SNOMEDCT_CORE|Suprarenogenic syndrome|Cushing's syndrome III
C0010495|T047|SY|58588007|SNOMEDCT_CORE|Chalazodermia|Cutis laxa
C0010495|T047|PT|58588007|SNOMEDCT_CORE|Cutis laxa|Cutis laxa
C0010495|T047|FN|58588007|SNOMEDCT_CORE|Cutis laxa|Cutis laxa
C0010495|T047|IS|58588007|SNOMEDCT_CORE|Cutis laxa, NOS|Cutis laxa
C0010495|T047|IS|58588007|SNOMEDCT_CORE|Dermatochalasia|Cutis laxa
C0010495|T047|IS|58588007|SNOMEDCT_CORE|Dermatochalasis|Cutis laxa
C0010495|T047|SY|58588007|SNOMEDCT_CORE|Dermatolysis|Cutis laxa
C0010495|T047|IS|58588007|SNOMEDCT_CORE|Dermatolysis, NOS|Cutis laxa
C0010495|T047|SY|58588007|SNOMEDCT_CORE|Dermatomegaly|Cutis laxa
C0010495|T047|IS|58588007|SNOMEDCT_CORE|Generalised dermatochalasis|Cutis laxa
C0010495|T047|IS|58588007|SNOMEDCT_CORE|Generalized dermatochalasis|Cutis laxa
C0010495|T047|SY|58588007|SNOMEDCT_CORE|Primary elastolysis|Cutis laxa
C0010520|T184|PT|3415004|SNOMEDCT_CORE|Cyanosis|Cyanosis
C0010520|T184|FN|3415004|SNOMEDCT_CORE|Cyanosis|Cyanosis
C0010598|T048|SY|76105009|SNOMEDCT_CORE|Affective personality disorder|Cyclothymia
C0010598|T048|PT|76105009|SNOMEDCT_CORE|Cyclothymia|Cyclothymia
C0010598|T048|FN|76105009|SNOMEDCT_CORE|Cyclothymia|Cyclothymia
C0010598|T048|SY|76105009|SNOMEDCT_CORE|Cyclothymic disorder|Cyclothymia
C0010623|T190|PT|197464001|SNOMEDCT_CORE|Cyst and pseudocyst of pancreas|Cyst and pseudocyst of pancreas
C0010623|T190|FN|197464001|SNOMEDCT_CORE|Cyst and pseudocyst of pancreas|Cyst and pseudocyst of pancreas
C0010666|T047|SY|13277001|SNOMEDCT_CORE|Acne cystica|Cystic acne
C0010666|T047|PT|13277001|SNOMEDCT_CORE|Cystic acne|Cystic acne
C0010666|T047|FN|13277001|SNOMEDCT_CORE|Cystic acne|Cystic acne
C0010666|T047|SY|13277001|SNOMEDCT_CORE|Cystic acne vulgaris|Cystic acne
C0010673|T191|PT|198321009|SNOMEDCT_CORE|Endometrial cystic hyperplasia|Endometrial cystic hyperplasia
C0010673|T191|FN|198321009|SNOMEDCT_CORE|Endometrial cystic hyperplasia|Endometrial cystic hyperplasia
C0010673|T191|SY|198321009|SNOMEDCT_CORE|Swiss cheese hyperplasia of the endometrium|Endometrial cystic hyperplasia
C0010674|T047|SY|190905008|SNOMEDCT_CORE|CF - Cystic fibrosis|Cystic fibrosis
C0010674|T047|PT|190905008|SNOMEDCT_CORE|Cystic fibrosis|Cystic fibrosis
C0010674|T047|FN|190905008|SNOMEDCT_CORE|Cystic fibrosis|Cystic fibrosis
C0010674|T047|SY|190905008|SNOMEDCT_CORE|Fibrocystic disease|Cystic fibrosis
C0010674|T047|SY|190905008|SNOMEDCT_CORE|Mucoviscidosis|Cystic fibrosis
C0010692|T047|SY|38822007|SNOMEDCT_CORE|Bladder infection|Cystitis
C0010692|T047|PT|38822007|SNOMEDCT_CORE|Cystitis|Cystitis
C0010692|T047|FN|38822007|SNOMEDCT_CORE|Cystitis|Cystitis
C0010692|T047|IS|38822007|SNOMEDCT_CORE|Cystitis, NOS|Cystitis
C0010709|T047|PT|441457006|SNOMEDCT_CORE|Cyst|Cyst
C0010709|T047|FN|441457006|SNOMEDCT_CORE|Cyst|Cyst
C0010823|T047|SY|28944009|SNOMEDCT_CORE|CMV - Cytomegalovirus infection|Cytomegalovirus infection
C0010823|T047|SY|28944009|SNOMEDCT_CORE|Cytomegalic inclusion disease|Cytomegalovirus infection
C0010823|T047|SY|28944009|SNOMEDCT_CORE|Cytomegalovirus disease|Cytomegalovirus infection
C0010823|T047|PT|28944009|SNOMEDCT_CORE|Cytomegalovirus infection|Cytomegalovirus infection
C0010823|T047|FN|28944009|SNOMEDCT_CORE|Cytomegalovirus infection|Cytomegalovirus infection
C0010823|T047|IS|28944009|SNOMEDCT_CORE|Cytomegalovirus infection, NOS|Cytomegalovirus infection
C0010823|T047|SY|28944009|SNOMEDCT_CORE|Disease due to Cytomegalovirus|Cytomegalovirus infection
C0010823|T047|IS|28944009|SNOMEDCT_CORE|Salivary gland virus disease|Cytomegalovirus infection
C0010930|T047|PT|85777005|SNOMEDCT_CORE|Dacryocystitis|Dacryocystitis
C0010930|T047|FN|85777005|SNOMEDCT_CORE|Dacryocystitis|Dacryocystitis
C0010930|T047|IS|85777005|SNOMEDCT_CORE|Dacryocystitis, NOS|Dacryocystitis
C0011053|T033|IS|15188001|SNOMEDCT_CORE|Deafness|Deafness
C0011053|T033|IS|15188001|SNOMEDCT_CORE|Deafness, NOS|Deafness
C0011057|T033|PT|79471008|SNOMEDCT_CORE|Sudden hearing loss|Sudden hearing loss
C0011057|T033|OF|79471008|SNOMEDCT_CORE|Sudden hearing loss|Sudden hearing loss
C0011057|T033|FN|79471008|SNOMEDCT_CORE|Sudden hearing loss|Sudden hearing loss
C0011057|T033|IS|79471008|SNOMEDCT_CORE|Sudden hearing loss, NOS|Sudden hearing loss
C0011071|T046|PT|26636000|SNOMEDCT_CORE|Sudden death|Sudden death
C0011071|T046|OF|26636000|SNOMEDCT_CORE|Sudden death|Sudden death
C0011071|T046|FN|26636000|SNOMEDCT_CORE|Sudden death|Sudden death
C0011071|T046|IS|26636000|SNOMEDCT_CORE|Sudden death, NOS|Sudden death
C0011124|T033|IS|8357008|SNOMEDCT_CORE|Decreased libido|Reduced libido
C0011124|T033|SY|8357008|SNOMEDCT_CORE|Low libido|Reduced libido
C0011124|T033|PT|8357008|SNOMEDCT_CORE|Reduced libido|Reduced libido
C0011124|T033|FN|8357008|SNOMEDCT_CORE|Reduced libido|Reduced libido
C0011127|T047|OAS|400192002|SNOMEDCT_CORE|Bed sore|Pressure ulcer
C0011127|T047|SY|399912005|SNOMEDCT_CORE|Contact ulcer|Pressure ulcer
C0011127|T047|OAS|400192002|SNOMEDCT_CORE|Decubitus pressure sore|Pressure ulcer
C0011127|T047|OAP|400192002|SNOMEDCT_CORE|Decubitus ulcer|Pressure ulcer
C0011127|T047|OAF|400192002|SNOMEDCT_CORE|Decubitus ulcer|Pressure ulcer
C0011127|T047|SY|399912005|SNOMEDCT_CORE|Pressure sore|Pressure ulcer
C0011127|T047|OF|399912005|SNOMEDCT_CORE|Pressure sore|Pressure ulcer
C0011127|T047|PT|399912005|SNOMEDCT_CORE|Pressure ulcer|Pressure ulcer
C0011127|T047|FN|399912005|SNOMEDCT_CORE|Pressure ulcer|Pressure ulcer
C0011168|T047|SY|40739000|SNOMEDCT_CORE|Can't get food down|Dysphagia
C0011168|T047|SY|40739000|SNOMEDCT_CORE|Cannot get food down|Dysphagia
C0011168|T047|SY|40739000|SNOMEDCT_CORE|Difficulty in swallowing|Dysphagia
C0011168|T047|PT|40739000|SNOMEDCT_CORE|Dysphagia|Dysphagia
C0011168|T047|FN|40739000|SNOMEDCT_CORE|Dysphagia|Dysphagia
C0011168|T047|IS|40739000|SNOMEDCT_CORE|Dysphagia, NOS|Dysphagia
C0011168|T047|SY|40739000|SNOMEDCT_CORE|Swallowing difficult|Dysphagia
C0011175|T047|OAS|37472003|SNOMEDCT_CORE|Deficient fluid volume|Dehydration
C0011175|T047|PT|34095006|SNOMEDCT_CORE|Dehydration|Dehydration
C0011175|T047|FN|34095006|SNOMEDCT_CORE|Dehydration|Dehydration
C0011175|T047|SY|34095006|SNOMEDCT_CORE|Pure water depletion syndrome|Dehydration
C0011206|T048|SY|2776000|SNOMEDCT_CORE|ABS - Acute brain syndrome|Delirium
C0011206|T048|SY|2776000|SNOMEDCT_CORE|Acute brain syndrome|Delirium
C0011206|T048|IS|2776000|SNOMEDCT_CORE|Acute brain syndrome, NOS|Delirium
C0011206|T048|PT|419567006|SNOMEDCT_CORE|Delirious|Delirium
C0011206|T048|FN|419567006|SNOMEDCT_CORE|Delirious|Delirium
C0011206|T048|PT|2776000|SNOMEDCT_CORE|Delirium|Delirium
C0011206|T048|FN|2776000|SNOMEDCT_CORE|Delirium|Delirium
C0011206|T048|IS|2776000|SNOMEDCT_CORE|Delirium, NOS|Delirium
C0011251|T048|PT|48500005|SNOMEDCT_CORE|Delusional disorder|Delusional disorder
C0011251|T048|FN|48500005|SNOMEDCT_CORE|Delusional disorder|Delusional disorder
C0011251|T048|IS|48500005|SNOMEDCT_CORE|Delusional disorder, NOS|Delusional disorder
C0011253|T048|IS|2073000|SNOMEDCT_CORE|Delusion|Delusions
C0011253|T048|IS|2073000|SNOMEDCT_CORE|Delusion, NOS|Delusions
C0011253|T048|SY|2073000|SNOMEDCT_CORE|Delusional ideas|Delusions
C0011253|T048|SY|2073000|SNOMEDCT_CORE|Delusional thoughts|Delusions
C0011253|T048|PT|2073000|SNOMEDCT_CORE|Delusions|Delusions
C0011253|T048|FN|2073000|SNOMEDCT_CORE|Delusions|Delusions
C0011263|T047|SY|56267009|SNOMEDCT_CORE|MID - Multi-infarct dementia|Multi-infarct dementia
C0011263|T047|SY|56267009|SNOMEDCT_CORE|Multi infarct dementia|Multi-infarct dementia
C0011263|T047|PT|56267009|SNOMEDCT_CORE|Multi-infarct dementia|Multi-infarct dementia
C0011263|T047|FN|56267009|SNOMEDCT_CORE|Multi-infarct dementia|Multi-infarct dementia
C0011263|T047|IS|56267009|SNOMEDCT_CORE|Multi-infarct dementia, NOS|Multi-infarct dementia
C0011268|T048|SY|15662003|SNOMEDCT_CORE|SD - Senile dementia|Senile dementia
C0011268|T048|PT|15662003|SNOMEDCT_CORE|Senile dementia|Senile dementia
C0011268|T048|FN|15662003|SNOMEDCT_CORE|Senile dementia|Senile dementia
C0011268|T048|IS|15662003|SNOMEDCT_CORE|Senile dementia, NOS|Senile dementia
C0011269|T047|SY|56267009|SNOMEDCT_CORE|VAD - Vascular dementia|Vascular dementia
C0011269|T047|IS|56267009|SNOMEDCT_CORE|Vascular dementia|Vascular dementia
C0011269|T047|PT|429998004|SNOMEDCT_CORE|Vascular dementia|Vascular dementia
C0011269|T047|FN|429998004|SNOMEDCT_CORE|Vascular dementia|Vascular dementia
C0011269|T047|IS|56267009|SNOMEDCT_CORE|Vascular dementia, NOS|Vascular dementia
C0011302|T047|SY|6118003|SNOMEDCT_CORE|Demyelinating CNS disease|Demyelinating disease of central nervous system
C0011302|T047|SY|6118003|SNOMEDCT_CORE|Demyelinating disease central nervous system|Demyelinating disease of central nervous system
C0011302|T047|PT|6118003|SNOMEDCT_CORE|Demyelinating disease of central nervous system|Demyelinating disease of central nervous system
C0011302|T047|FN|6118003|SNOMEDCT_CORE|Demyelinating disease of central nervous system|Demyelinating disease of central nervous system
C0011302|T047|IS|6118003|SNOMEDCT_CORE|Demyelinating disease of central nervous system, NOS|Demyelinating disease of central nervous system
C0011302|T047|SY|6118003|SNOMEDCT_CORE|Demyelinating disorders of the central nervous system|Demyelinating disease of central nervous system
C0011330|T033|PT|17552000|SNOMEDCT_CORE|Dental calculus|Dental calculus
C0011330|T033|FN|17552000|SNOMEDCT_CORE|Dental calculus|Dental calculus
C0011330|T033|IS|17552000|SNOMEDCT_CORE|Dental calculus, NOS|Dental calculus
C0011330|T033|SY|17552000|SNOMEDCT_CORE|Odontolith|Dental calculus
C0011330|T033|SY|17552000|SNOMEDCT_CORE|Tartar|Dental calculus
C0011334|T047|SY|80967001|SNOMEDCT_CORE|Carious lesion|Dental caries
C0011334|T047|PT|80967001|SNOMEDCT_CORE|Dental caries|Dental caries
C0011334|T047|FN|80967001|SNOMEDCT_CORE|Dental caries|Dental caries
C0011334|T047|IS|80967001|SNOMEDCT_CORE|Dental caries, NOS|Dental caries
C0011334|T047|SY|80967001|SNOMEDCT_CORE|Dental cavity|Dental caries
C0011334|T047|IS|80967001|SNOMEDCT_CORE|Dental cavity, NOS|Dental caries
C0011334|T047|SY|80967001|SNOMEDCT_CORE|Dental decay|Dental caries
C0011334|T047|IS|80967001|SNOMEDCT_CORE|Saprodontia|Dental caries
C0011334|T047|SY|80967001|SNOMEDCT_CORE|Teeth decayed|Dental caries
C0011334|T047|SY|80967001|SNOMEDCT_CORE|Tooth caries|Dental caries
C0011334|T047|SY|80967001|SNOMEDCT_CORE|Tooth decay|Dental caries
C0011334|T047|SY|80967001|SNOMEDCT_CORE|Tooth decayed|Dental caries
C0011548|T048|PT|84466009|SNOMEDCT_CORE|Dependent personality disorder|Dependent personality disorder
C0011548|T048|FN|84466009|SNOMEDCT_CORE|Dependent personality disorder|Dependent personality disorder
C0011570|T048|OAP|41006004|SNOMEDCT_CORE|Depression|Depression
C0011570|T048|OAF|41006004|SNOMEDCT_CORE|Depression|Depression
C0011570|T048|IS|41006004|SNOMEDCT_CORE|Depression, NOS|Depression
C0011573|T048|PT|300706003|SNOMEDCT_CORE|Endogenous depression|Endogenous depression
C0011573|T048|FN|300706003|SNOMEDCT_CORE|Endogenous depression|Endogenous depression
C0011579|T048|SY|87414006|SNOMEDCT_CORE|Reactive depression|Reactive depression
C0011579|T048|PT|87414006|SNOMEDCT_CORE|Reactive depression|Reactive depression
C0011579|T048|OF|87414006|SNOMEDCT_CORE|Reactive depression|Reactive depression
C0011579|T048|FN|87414006|SNOMEDCT_CORE|Reactive depression|Reactive depression
C0011581|T048|SY|35489007|SNOMEDCT_CORE|Depression|Depressive disorder
C0011581|T048|PT|35489007|SNOMEDCT_CORE|Depressive disorder|Depressive disorder
C0011581|T048|FN|35489007|SNOMEDCT_CORE|Depressive disorder|Depressive disorder
C0011581|T048|IS|35489007|SNOMEDCT_CORE|Depressive disorder, NOS|Depressive disorder
C0011581|T048|SY|35489007|SNOMEDCT_CORE|Depressive illness|Depressive disorder
C0011581|T048|SY|78667006|SNOMEDCT_CORE|Depressive neurosis|Depressive disorder
C0011581|T048|SY|35489007|SNOMEDCT_CORE|Mood disorder of depressed type|Depressive disorder
C0011603|T047|OAP|182782007|SNOMEDCT_CORE|Dermatitis|Dermatitis
C0011603|T047|IS|43116000|SNOMEDCT_CORE|Dermatitis|Dermatitis
C0011603|T047|SY|703938007|SNOMEDCT_CORE|Dermatitis|Dermatitis
C0011603|T047|OAF|182782007|SNOMEDCT_CORE|Dermatitis|Dermatitis
C0011603|T047|OAS|182782007|SNOMEDCT_CORE|Inflammation of skin|Dermatitis
C0011606|T047|PT|399992009|SNOMEDCT_CORE|Erythroderma|Erythroderma
C0011606|T047|FN|399992009|SNOMEDCT_CORE|Erythroderma|Erythroderma
C0011606|T047|SY|399992009|SNOMEDCT_CORE|Erythrodermatitis|Erythroderma
C0011606|T047|SY|399992009|SNOMEDCT_CORE|Exfoliative dermatitis|Erythroderma
C0011606|T047|OAP|396350005|SNOMEDCT_CORE|Generalised exfoliative dermatitis|Erythroderma
C0011606|T047|SYGB|399992009|SNOMEDCT_CORE|Generalised exfoliative dermatitis|Erythroderma
C0011606|T047|OAP|396350005|SNOMEDCT_CORE|Generalized exfoliative dermatitis|Erythroderma
C0011606|T047|SY|399992009|SNOMEDCT_CORE|Generalized exfoliative dermatitis|Erythroderma
C0011606|T047|OAF|396350005|SNOMEDCT_CORE|Generalized exfoliative dermatitis|Erythroderma
C0011606|T047|OAS|396350005|SNOMEDCT_CORE|Pityriasis rubra of Hebra|Erythroderma
C0011608|T047|PT|111196000|SNOMEDCT_CORE|Dermatitis herpetiformis|Dermatitis herpetiformis
C0011608|T047|FN|111196000|SNOMEDCT_CORE|Dermatitis herpetiformis|Dermatitis herpetiformis
C0011608|T047|SY|111196000|SNOMEDCT_CORE|Dermatosis herpetiformis|Dermatitis herpetiformis
C0011608|T047|SY|111196000|SNOMEDCT_CORE|DH - Dermatitis herpetiformis|Dermatitis herpetiformis
C0011608|T047|SY|111196000|SNOMEDCT_CORE|Duhring-Brocq disease|Dermatitis herpetiformis
C0011608|T047|SY|111196000|SNOMEDCT_CORE|Duhring's disease|Dermatitis herpetiformis
C0011609|T047|SY|28926001|SNOMEDCT_CORE|Dermatitis medicamentosa|Eruption due to drug
C0011609|T047|SY|28926001|SNOMEDCT_CORE|Drug eruption|Eruption due to drug
C0011609|T047|IS|28926001|SNOMEDCT_CORE|Drug eruption, NOS|Eruption due to drug
C0011609|T047|SY|28926001|SNOMEDCT_CORE|Drug rash|Eruption due to drug
C0011609|T047|IS|28926001|SNOMEDCT_CORE|Drug rash, NOS|Eruption due to drug
C0011609|T047|SY|28926001|SNOMEDCT_CORE|Drug-induced rash|Eruption due to drug
C0011609|T047|FN|28926001|SNOMEDCT_CORE|Eruption caused by drug|Eruption due to drug
C0011609|T047|SY|28926001|SNOMEDCT_CORE|Eruption caused by drug|Eruption due to drug
C0011609|T047|PT|28926001|SNOMEDCT_CORE|Eruption due to drug|Eruption due to drug
C0011609|T047|OF|28926001|SNOMEDCT_CORE|Eruption due to drug|Eruption due to drug
C0011609|T047|IS|28926001|SNOMEDCT_CORE|Eruption due to drug, NOS|Eruption due to drug
C0011615|T047|SY|24079001|SNOMEDCT_CORE|AD - Atopic dermatitis|Atopic dermatitis
C0011615|T047|SY|24079001|SNOMEDCT_CORE|Allergic dermatitis|Atopic dermatitis
C0011615|T047|SY|24079001|SNOMEDCT_CORE|Allergic eczema|Atopic dermatitis
C0011615|T047|PT|24079001|SNOMEDCT_CORE|Atopic dermatitis|Atopic dermatitis
C0011615|T047|FN|24079001|SNOMEDCT_CORE|Atopic dermatitis|Atopic dermatitis
C0011615|T047|IS|24079001|SNOMEDCT_CORE|Atopic dermatitis, NOS|Atopic dermatitis
C0011615|T047|SY|24079001|SNOMEDCT_CORE|Atopic eczema|Atopic dermatitis
C0011615|T047|IS|24079001|SNOMEDCT_CORE|Atopic neurodermatitis|Atopic dermatitis
C0011615|T047|IS|24079001|SNOMEDCT_CORE|Canine atopy|Atopic dermatitis
C0011615|T047|SY|24079001|SNOMEDCT_CORE|Constitutional eczema|Atopic dermatitis
C0011615|T047|SY|24079001|SNOMEDCT_CORE|Disseminated neurodermatitis|Atopic dermatitis
C0011616|T047|SY|40275004|SNOMEDCT_CORE|CD - Contact dermatitis|Contact dermatitis
C0011616|T047|PT|40275004|SNOMEDCT_CORE|Contact dermatitis|Contact dermatitis
C0011616|T047|FN|40275004|SNOMEDCT_CORE|Contact dermatitis|Contact dermatitis
C0011616|T047|IS|40275004|SNOMEDCT_CORE|Contact dermatitis, NOS|Contact dermatitis
C0011616|T047|SY|40275004|SNOMEDCT_CORE|Contact eczema|Contact dermatitis
C0011616|T047|SY|40275004|SNOMEDCT_CORE|Dermatitis venenata|Contact dermatitis
C0011620|T047|SY|35498005|SNOMEDCT_CORE|Gravitational eczema|Stasis dermatitis
C0011620|T047|PT|35498005|SNOMEDCT_CORE|Stasis dermatitis|Stasis dermatitis
C0011620|T047|FN|35498005|SNOMEDCT_CORE|Stasis dermatitis|Stasis dermatitis
C0011620|T047|IS|35498005|SNOMEDCT_CORE|Stasis dermatitis, NOS|Stasis dermatitis
C0011620|T047|SY|35498005|SNOMEDCT_CORE|Stasis eczema|Stasis dermatitis
C0011620|T047|IS|35498005|SNOMEDCT_CORE|Varicose eczema|Stasis dermatitis
C0011620|T047|IS|35498005|SNOMEDCT_CORE|Venous eczema|Stasis dermatitis
C0011630|T047|SY|14560005|SNOMEDCT_CORE|Cutaneous mycosis|Dermal mycosis
C0011630|T047|IS|14560005|SNOMEDCT_CORE|Cutaneous mycosis, NOS|Dermal mycosis
C0011630|T047|PT|14560005|SNOMEDCT_CORE|Dermal mycosis|Dermal mycosis
C0011630|T047|FN|14560005|SNOMEDCT_CORE|Dermal mycosis|Dermal mycosis
C0011630|T047|IS|14560005|SNOMEDCT_CORE|Dermal mycosis, NOS|Dermal mycosis
C0011630|T047|IS|47382004|SNOMEDCT_CORE|Dermatomycosis|Dermal mycosis
C0011630|T047|SY|14560005|SNOMEDCT_CORE|Dermatomycosis|Dermal mycosis
C0011630|T047|SY|14560005|SNOMEDCT_CORE|Fungal dermatitis|Dermal mycosis
C0011630|T047|IS|14560005|SNOMEDCT_CORE|Fungal dermatitis, NOS|Dermal mycosis
C0011630|T047|SY|14560005|SNOMEDCT_CORE|Fungal dermatosis|Dermal mycosis
C0011633|T047|PT|396230008|SNOMEDCT_CORE|Dermatomyositis|Dermatomyositis
C0011633|T047|FN|396230008|SNOMEDCT_CORE|Dermatomyositis|Dermatomyositis
C0011633|T047|SY|396230008|SNOMEDCT_CORE|DM - Dermatomyositis|Dermatomyositis
C0011633|T047|SY|396230008|SNOMEDCT_CORE|Polymyositis with skin involvement|Dermatomyositis
C0011633|T047|SY|396230008|SNOMEDCT_CORE|Wagner-Unverricht syndrome|Dermatomyositis
C0011636|T047|PT|47382004|SNOMEDCT_CORE|Dermatophytosis|Dermatophytosis
C0011636|T047|FN|47382004|SNOMEDCT_CORE|Dermatophytosis|Dermatophytosis
C0011644|T047|OAP|201441006|SNOMEDCT_CORE|Scleroderma|Scleroderma
C0011644|T047|IS|89155008|SNOMEDCT_CORE|Scleroderma|Scleroderma
C0011644|T047|OF|201441006|SNOMEDCT_CORE|Scleroderma|Scleroderma
C0011644|T047|OAF|201441006|SNOMEDCT_CORE|Scleroderma|Scleroderma
C0011649|T191|OAP|439575008|SNOMEDCT_CORE|Mature cystic teratoma|Mature cystic teratoma
C0011649|T191|OAF|439575008|SNOMEDCT_CORE|Mature cystic teratoma|Mature cystic teratoma
C0011848|T047|SY|15771004|SNOMEDCT_CORE|DI - Diabetes insipidus|Diabetes insipidus
C0011848|T047|PT|15771004|SNOMEDCT_CORE|Diabetes insipidus|Diabetes insipidus
C0011848|T047|FN|15771004|SNOMEDCT_CORE|Diabetes insipidus|Diabetes insipidus
C0011848|T047|IS|15771004|SNOMEDCT_CORE|Diabetes insipidus, NOS|Diabetes insipidus
C0011849|T047|PT|73211009|SNOMEDCT_CORE|Diabetes mellitus|Diabetes mellitus
C0011849|T047|FN|73211009|SNOMEDCT_CORE|Diabetes mellitus|Diabetes mellitus
C0011849|T047|IS|73211009|SNOMEDCT_CORE|Diabetes mellitus, NOS|Diabetes mellitus
C0011849|T047|SY|73211009|SNOMEDCT_CORE|DM - Diabetes mellitus|Diabetes mellitus
C0011854|T047|SY|46635009|SNOMEDCT_CORE|Diabetes mellitus type 1|Type 1 diabetes mellitus
C0011854|T047|FN|46635009|SNOMEDCT_CORE|Diabetes mellitus type 1|Type 1 diabetes mellitus
C0011854|T047|SY|46635009|SNOMEDCT_CORE|Diabetes mellitus type I|Type 1 diabetes mellitus
C0011854|T047|IS|46635009|SNOMEDCT_CORE|IDDM|Type 1 diabetes mellitus
C0011854|T047|IS|46635009|SNOMEDCT_CORE|IDDM - Insulin-dependent diabetes mellitus|Type 1 diabetes mellitus
C0011854|T047|IS|46635009|SNOMEDCT_CORE|Insulin dependent diabetes mellitus|Type 1 diabetes mellitus
C0011854|T047|IS|46635009|SNOMEDCT_CORE|Insulin-dependent diabetes mellitus|Type 1 diabetes mellitus
C0011854|T047|IS|46635009|SNOMEDCT_CORE|Juvenile onset diabetes mellitus|Type 1 diabetes mellitus
C0011854|T047|PT|46635009|SNOMEDCT_CORE|Type 1 diabetes mellitus|Type 1 diabetes mellitus
C0011854|T047|SY|46635009|SNOMEDCT_CORE|Type I diabetes mellitus|Type 1 diabetes mellitus
C0011859|T047|IS|71325002|SNOMEDCT_CORE|Lipoatrophic diabetes, NOS|Lipoatrophic diabetes, NOS
C0011859|T047|IS|71325002|SNOMEDCT_CORE|Lipodystrophic diabetes, NOS|Lipodystrophic diabetes, NOS
C0011860|T047|IS|44054006|SNOMEDCT_CORE|Diabetes mellitus - adult onset|Type 2 diabetes mellitus
C0011860|T047|SY|44054006|SNOMEDCT_CORE|Diabetes mellitus type 2|Type 2 diabetes mellitus
C0011860|T047|FN|44054006|SNOMEDCT_CORE|Diabetes mellitus type 2|Type 2 diabetes mellitus
C0011860|T047|SY|44054006|SNOMEDCT_CORE|Diabetes mellitus type II|Type 2 diabetes mellitus
C0011860|T047|IS|44054006|SNOMEDCT_CORE|Maturity onset diabetes mellitus|Type 2 diabetes mellitus
C0011860|T047|IS|44054006|SNOMEDCT_CORE|NCDMM|Type 2 diabetes mellitus
C0011860|T047|IS|44054006|SNOMEDCT_CORE|NIDDM|Type 2 diabetes mellitus
C0011860|T047|IS|44054006|SNOMEDCT_CORE|NIDDM - Non-insulin dependent diabetes mellitus|Type 2 diabetes mellitus
C0011860|T047|IS|44054006|SNOMEDCT_CORE|Non-insulin dependent diabetes mellitus|Type 2 diabetes mellitus
C0011860|T047|IS|44054006|SNOMEDCT_CORE|Non-insulin-dependent diabetes mellitus|Type 2 diabetes mellitus
C0011860|T047|PT|44054006|SNOMEDCT_CORE|Type 2 diabetes mellitus|Type 2 diabetes mellitus
C0011860|T047|SY|44054006|SNOMEDCT_CORE|Type II diabetes mellitus|Type 2 diabetes mellitus
C0011871|T047|SY|127014009|SNOMEDCT_CORE|Diabetes with peripheral circulatory disorder|Peripheral angiopathy due to diabetes mellitus
C0011871|T047|IS|127014009|SNOMEDCT_CORE|Diabetes with peripheral circulatory disorders|Peripheral angiopathy due to diabetes mellitus
C0011871|T047|SY|127014009|SNOMEDCT_CORE|Diabetic peripheral angiopathy|Peripheral angiopathy due to diabetes mellitus
C0011871|T047|OF|127014009|SNOMEDCT_CORE|Diabetic peripheral angiopathy|Peripheral angiopathy due to diabetes mellitus
C0011871|T047|SY|127014009|SNOMEDCT_CORE|Diabetic peripheral vascular disease|Peripheral angiopathy due to diabetes mellitus
C0011871|T047|PT|127014009|SNOMEDCT_CORE|Peripheral angiopathy due to diabetes mellitus|Peripheral angiopathy due to diabetes mellitus
C0011871|T047|FN|127014009|SNOMEDCT_CORE|Peripheral angiopathy due to diabetes mellitus|Peripheral angiopathy due to diabetes mellitus
C0011876|T047|OF|43959009|SNOMEDCT_CORE|Cataract co-occurrent and due to diabetes mellitus|Cataract due to diabetes mellitus
C0011876|T047|OP|43959009|SNOMEDCT_CORE|Cataract co-occurrent and due to diabetes mellitus|Cataract due to diabetes mellitus
C0011876|T047|PT|43959009|SNOMEDCT_CORE|Cataract due to diabetes mellitus|Cataract due to diabetes mellitus
C0011876|T047|SY|43959009|SNOMEDCT_CORE|Cataract of eye due to diabetes mellitus|Cataract due to diabetes mellitus
C0011876|T047|FN|43959009|SNOMEDCT_CORE|Cataract of eye due to diabetes mellitus|Cataract due to diabetes mellitus
C0011876|T047|SY|43959009|SNOMEDCT_CORE|Diabetic cataract|Cataract due to diabetes mellitus
C0011876|T047|OF|43959009|SNOMEDCT_CORE|Diabetic cataract|Cataract due to diabetes mellitus
C0011880|T047|SY|420422005|SNOMEDCT_CORE|Diabetes mellitus with ketoacidosis|Diabetic ketoacidosis
C0011880|T047|SY|420422005|SNOMEDCT_CORE|Diabetic acidosis|Diabetic ketoacidosis
C0011880|T047|PT|420422005|SNOMEDCT_CORE|Diabetic ketoacidosis|Diabetic ketoacidosis
C0011880|T047|SY|420422005|SNOMEDCT_CORE|DKA - diabetic ketoacidosis|Diabetic ketoacidosis
C0011880|T047|FN|420422005|SNOMEDCT_CORE|Ketoacidosis due to diabetes mellitus|Diabetic ketoacidosis
C0011880|T047|SY|420422005|SNOMEDCT_CORE|Ketoacidosis due to diabetes mellitus|Diabetic ketoacidosis
C0011880|T047|SY|420422005|SNOMEDCT_CORE|Ketoacidosis in diabetes mellitus|Diabetic ketoacidosis
C0011880|T047|OF|420422005|SNOMEDCT_CORE|Ketoacidosis in diabetes mellitus|Diabetic ketoacidosis
C0011881|T047|SY|127013003|SNOMEDCT_CORE|Diabetic nephropathy|Disorder of kidney due to diabetes mellitus
C0011881|T047|SY|127013003|SNOMEDCT_CORE|Diabetic renal disease|Disorder of kidney due to diabetes mellitus
C0011881|T047|OF|127013003|SNOMEDCT_CORE|Diabetic renal disease|Disorder of kidney due to diabetes mellitus
C0011881|T047|OF|127013003|SNOMEDCT_CORE|Disorder of kidney co-occurrent and due to diabetes mellitus|Disorder of kidney due to diabetes mellitus
C0011881|T047|IS|127013003|SNOMEDCT_CORE|Disorder of kidney co-occurrent and due to diabetes mellitus|Disorder of kidney due to diabetes mellitus
C0011881|T047|PT|127013003|SNOMEDCT_CORE|Disorder of kidney due to diabetes mellitus|Disorder of kidney due to diabetes mellitus
C0011881|T047|FN|127013003|SNOMEDCT_CORE|Disorder of kidney due to diabetes mellitus|Disorder of kidney due to diabetes mellitus
C0011881|T047|SY|127013003|SNOMEDCT_CORE|Kidney disorder due to diabetes mellitus|Disorder of kidney due to diabetes mellitus
C0011881|T047|SY|127013003|SNOMEDCT_CORE|Renal disorder associated with diabetes mellitus|Disorder of kidney due to diabetes mellitus
C0011882|T047|SY|230572002|SNOMEDCT_CORE|Diabetes mellitus with neuropathy|Neuropathy due to diabetes mellitus
C0011882|T047|SY|230572002|SNOMEDCT_CORE|Diabetic neuropathy|Neuropathy due to diabetes mellitus
C0011882|T047|OF|230572002|SNOMEDCT_CORE|Diabetic neuropathy|Neuropathy due to diabetes mellitus
C0011882|T047|OF|230572002|SNOMEDCT_CORE|Neuropathy co-occurrent and due to diabetes mellitus|Neuropathy due to diabetes mellitus
C0011882|T047|IS|230572002|SNOMEDCT_CORE|Neuropathy co-occurrent and due to diabetes mellitus|Neuropathy due to diabetes mellitus
C0011882|T047|FN|230572002|SNOMEDCT_CORE|Neuropathy due to diabetes mellitus|Neuropathy due to diabetes mellitus
C0011882|T047|PT|230572002|SNOMEDCT_CORE|Neuropathy due to diabetes mellitus|Neuropathy due to diabetes mellitus
C0011884|T047|SY|4855003|SNOMEDCT_CORE|Diabetic retinopathy|Retinopathy due to diabetes mellitus
C0011884|T047|OF|4855003|SNOMEDCT_CORE|Diabetic retinopathy|Retinopathy due to diabetes mellitus
C0011884|T047|IS|4855003|SNOMEDCT_CORE|Diabetic retinopathy, NOS|Retinopathy due to diabetes mellitus
C0011884|T047|SY|4855003|SNOMEDCT_CORE|DR - Diabetic retinopathy|Retinopathy due to diabetes mellitus
C0011884|T047|SY|4855003|SNOMEDCT_CORE|Retinal abnormality - diabetes-related|Retinopathy due to diabetes mellitus
C0011884|T047|OF|4855003|SNOMEDCT_CORE|Retinopathy co-occurrent and due to diabetes mellitus|Retinopathy due to diabetes mellitus
C0011884|T047|IS|4855003|SNOMEDCT_CORE|Retinopathy co-occurrent and due to diabetes mellitus|Retinopathy due to diabetes mellitus
C0011884|T047|PT|4855003|SNOMEDCT_CORE|Retinopathy due to diabetes mellitus|Retinopathy due to diabetes mellitus
C0011884|T047|FN|4855003|SNOMEDCT_CORE|Retinopathy due to diabetes mellitus|Retinopathy due to diabetes mellitus
C0011974|T047|SY|91487003|SNOMEDCT_CORE|Ammonia dermatitis|Diaper rash
C0011974|T047|SYGB|91487003|SNOMEDCT_CORE|Ammoniacal napkin dermatitis|Diaper rash
C0011974|T047|SY|91487003|SNOMEDCT_CORE|Diaper dermatitis|Diaper rash
C0011974|T047|SY|91487003|SNOMEDCT_CORE|Diaper erythema|Diaper rash
C0011974|T047|PT|91487003|SNOMEDCT_CORE|Diaper rash|Diaper rash
C0011974|T047|FN|91487003|SNOMEDCT_CORE|Diaper rash|Diaper rash
C0011974|T047|SYGB|91487003|SNOMEDCT_CORE|Irritant napkin dermatitis|Diaper rash
C0011974|T047|SY|91487003|SNOMEDCT_CORE|Jacquet's dermatitis|Diaper rash
C0011974|T047|SY|91487003|SNOMEDCT_CORE|Jacquet's erythema|Diaper rash
C0011974|T047|IS|91487003|SNOMEDCT_CORE|Napkin rash|Diaper rash
C0011974|T047|PTGB|91487003|SNOMEDCT_CORE|Nappy rash|Diaper rash
C0011974|T047|SYGB|91487003|SNOMEDCT_CORE|Nappy rash - irritant|Diaper rash
C0011991|T184|SY|62315008|SNOMEDCT_CORE|D - Diarrhea|Diarrhea
C0011991|T184|SYGB|62315008|SNOMEDCT_CORE|D - Diarrhoea|Diarrhea
C0011991|T184|PT|62315008|SNOMEDCT_CORE|Diarrhea|Diarrhea
C0011991|T184|FN|62315008|SNOMEDCT_CORE|Diarrhea|Diarrhea
C0011991|T184|IS|62315008|SNOMEDCT_CORE|Diarrhea, NOS|Diarrhea
C0011991|T184|PTGB|62315008|SNOMEDCT_CORE|Diarrhoea|Diarrhea
C0011991|T184|IS|62315008|SNOMEDCT_CORE|Loose bowel motions|Diarrhea
C0011991|T184|IS|62315008|SNOMEDCT_CORE|Loose bowel movement|Diarrhea
C0011991|T184|SY|62315008|SNOMEDCT_CORE|Observation of diarrhea|Diarrhea
C0011991|T184|SYGB|62315008|SNOMEDCT_CORE|Observation of diarrhoea|Diarrhea
C0012569|T033|PT|24982008|SNOMEDCT_CORE|Diplopia|Diplopia
C0012569|T033|FN|24982008|SNOMEDCT_CORE|Diplopia|Diplopia
C0012569|T033|SY|24982008|SNOMEDCT_CORE|Double vision|Diplopia
C0012569|T033|SY|24982008|SNOMEDCT_CORE|Seeing double|Diplopia
C0012624|T047|PT|2304001|SNOMEDCT_CORE|Discitis|Discitis
C0012624|T047|FN|2304001|SNOMEDCT_CORE|Discitis|Discitis
C0012624|T047|IS|2304001|SNOMEDCT_CORE|Discitis, NOS|Discitis
C0012624|T047|SY|2304001|SNOMEDCT_CORE|Intervertebral discitis|Discitis
C0012715|T047|PT|30913008|SNOMEDCT_CORE|Disorder of iron metabolism|Disorder of iron metabolism
C0012715|T047|FN|30913008|SNOMEDCT_CORE|Disorder of iron metabolism|Disorder of iron metabolism
C0012715|T047|IS|30913008|SNOMEDCT_CORE|Disorder of iron metabolism, NOS|Disorder of iron metabolism
C0012716|T047|PT|60853003|SNOMEDCT_CORE|Disorder of magnesium metabolism|Disorder of magnesium metabolism
C0012716|T047|FN|60853003|SNOMEDCT_CORE|Disorder of magnesium metabolism|Disorder of magnesium metabolism
C0012716|T047|IS|60853003|SNOMEDCT_CORE|Disorder of magnesium metabolism, NOS|Disorder of magnesium metabolism
C0012734|T048|PT|54319003|SNOMEDCT_CORE|Disruptive behavior disorder|Disruptive behavior disorder
C0012734|T048|FN|54319003|SNOMEDCT_CORE|Disruptive behavior disorder|Disruptive behavior disorder
C0012734|T048|IS|54319003|SNOMEDCT_CORE|Disruptive behavior disorder, NOS|Disruptive behavior disorder
C0012734|T048|PTGB|54319003|SNOMEDCT_CORE|Disruptive behaviour disorder|Disruptive behavior disorder
C0012736|T047|IS|308546005|SNOMEDCT_CORE|Dissecting aortic aneurysm|Dissecting aortic aneurysm
C0012739|T047|SY|67406007|SNOMEDCT_CORE|Consumptive coagulopathy|Disseminated intravascular coagulation
C0012739|T047|SYGB|67406007|SNOMEDCT_CORE|Consumptive thrombohaemorrhagic disorder|Disseminated intravascular coagulation
C0012739|T047|SY|67406007|SNOMEDCT_CORE|Consumptive thrombohemorrhagic disorder|Disseminated intravascular coagulation
C0012739|T047|IS|67406007|SNOMEDCT_CORE|Consumptive thrombohemorrhagic disorder, NOS|Disseminated intravascular coagulation
C0012739|T047|SY|67406007|SNOMEDCT_CORE|Defibrination syndrome|Disseminated intravascular coagulation
C0012739|T047|SY|67406007|SNOMEDCT_CORE|DIC - Disseminated intravascular coagulation|Disseminated intravascular coagulation
C0012739|T047|SY|67406007|SNOMEDCT_CORE|DIC syndrome|Disseminated intravascular coagulation
C0012739|T047|PT|67406007|SNOMEDCT_CORE|Disseminated intravascular coagulation|Disseminated intravascular coagulation
C0012739|T047|FN|67406007|SNOMEDCT_CORE|Disseminated intravascular coagulation|Disseminated intravascular coagulation
C0012739|T047|SYGB|67406007|SNOMEDCT_CORE|Haemorrhagic fibrinogenolysis|Disseminated intravascular coagulation
C0012739|T047|SY|67406007|SNOMEDCT_CORE|Hemorrhagic fibrinogenolysis|Disseminated intravascular coagulation
C0012766|T184|IS|80910005|SNOMEDCT_CORE|Abnormal skin sensitivity|Skin sensation disturbance
C0012766|T184|PT|80910005|SNOMEDCT_CORE|Skin sensation disturbance|Skin sensation disturbance
C0012766|T184|FN|80910005|SNOMEDCT_CORE|Skin sensation disturbance|Skin sensation disturbance
C0012767|T047|SY|234949000|SNOMEDCT_CORE|Abnormal tooth eruption|Tooth eruption disorder
C0012767|T047|SY|234949000|SNOMEDCT_CORE|Anomaly of tooth eruption|Tooth eruption disorder
C0012767|T047|PT|234949000|SNOMEDCT_CORE|Tooth eruption disorder|Tooth eruption disorder
C0012767|T047|FN|234949000|SNOMEDCT_CORE|Tooth eruption disorder|Tooth eruption disorder
C0012767|T047|IS|234949000|SNOMEDCT_CORE|Tooth eruption disorders|Tooth eruption disorder
C0012767|T047|OF|234949000|SNOMEDCT_CORE|Tooth eruption disorders|Tooth eruption disorder
C0012767|T047|SY|234949000|SNOMEDCT_CORE|Tooth eruption disturbance|Tooth eruption disorder
C0012767|T047|IS|234949000|SNOMEDCT_CORE|Tooth eruption disturbances|Tooth eruption disorder
C0012813|T047|PT|307496006|SNOMEDCT_CORE|Diverticulitis|Diverticulitis
C0012813|T047|FN|307496006|SNOMEDCT_CORE|Diverticulitis|Diverticulitis
C0012814|T047|PT|111359004|SNOMEDCT_CORE|Diverticulitis of colon|Diverticulitis of colon
C0012814|T047|FN|111359004|SNOMEDCT_CORE|Diverticulitis of colon|Diverticulitis of colon
C0012818|T047|SY|429430001|SNOMEDCT_CORE|Asymptomatic diverticulosis of sigmoid colon|Diverticulosis of sigmoid colon
C0012818|T047|SY|429430001|SNOMEDCT_CORE|Diverticulosis of sigmoid|Diverticulosis of sigmoid colon
C0012818|T047|PT|429430001|SNOMEDCT_CORE|Diverticulosis of sigmoid colon|Diverticulosis of sigmoid colon
C0012818|T047|FN|429430001|SNOMEDCT_CORE|Diverticulosis of sigmoid colon|Diverticulosis of sigmoid colon
C0012818|T047|OF|429430001|SNOMEDCT_CORE|Diverticulosis of sigmoid colon|Diverticulosis of sigmoid colon
C0012819|T047|PT|398050005|SNOMEDCT_CORE|Diverticular disease of colon|Diverticular disease of colon
C0012819|T047|FN|398050005|SNOMEDCT_CORE|Diverticular disease of colon|Diverticular disease of colon
C0012819|T047|IS|398050005|SNOMEDCT_CORE|Diverticulosis of colon|Diverticular disease of colon
C0012819|T047|IS|398050005|SNOMEDCT_CORE|Diverticulosis of the colon|Diverticular disease of colon
C0012819|T047|SY|398050005|SNOMEDCT_CORE|Symptomatic diverticulosis of colon|Diverticular disease of colon
C0012833|T184|PT|404640003|SNOMEDCT_CORE|Dizziness|Dizziness
C0012833|T184|FN|404640003|SNOMEDCT_CORE|Dizziness|Dizziness
C0012833|T184|SY|271789005|SNOMEDCT_CORE|Dizzy|Dizziness
C0013069|T019|IS|7484005|SNOMEDCT_CORE|Dextratransposition of aorta|Double outlet right ventricle
C0013069|T019|SY|7484005|SNOMEDCT_CORE|DORV - Double outlet right ventricle|Double outlet right ventricle
C0013069|T019|PT|7484005|SNOMEDCT_CORE|Double outlet right ventricle|Double outlet right ventricle
C0013069|T019|FN|7484005|SNOMEDCT_CORE|Double outlet right ventricle|Double outlet right ventricle
C0013069|T019|SY|7484005|SNOMEDCT_CORE|Origin of both great vessels from right ventricle|Double outlet right ventricle
C0013069|T019|SY|7484005|SNOMEDCT_CORE|Transposition of great vessels, interventricular septal defect AND overriding aorta|Double outlet right ventricle
C0013069|T019|IS|7484005|SNOMEDCT_CORE|Transposition of great vessels, interventricular septal defect and overriding aorta|Double outlet right ventricle
C0013080|T047|PT|41040004|SNOMEDCT_CORE|Complete trisomy 21 syndrome|Complete trisomy 21 syndrome
C0013080|T047|FN|41040004|SNOMEDCT_CORE|Complete trisomy 21 syndrome|Complete trisomy 21 syndrome
C0013080|T047|SY|41040004|SNOMEDCT_CORE|Down syndrome|Complete trisomy 21 syndrome
C0013080|T047|SY|41040004|SNOMEDCT_CORE|Downs syndrome|Complete trisomy 21 syndrome
C0013080|T047|IS|41040004|SNOMEDCT_CORE|Mongolism|Complete trisomy 21 syndrome
C0013080|T047|SY|41040004|SNOMEDCT_CORE|T21 - Trisomy 21|Complete trisomy 21 syndrome
C0013143|T037|PT|212962007|SNOMEDCT_CORE|Drowning and non-fatal immersion|Drowning and non-fatal immersion
C0013143|T037|FN|212962007|SNOMEDCT_CORE|Drowning and non-fatal immersion|Drowning and non-fatal immersion
C0013143|T037|SY|212962007|SNOMEDCT_CORE|Drowning and non-fatal submersion|Drowning and non-fatal immersion
C0013144|T033|SY|271782001|SNOMEDCT_CORE|Drowsiness|Drowsy
C0013144|T033|PT|271782001|SNOMEDCT_CORE|Drowsy|Drowsy
C0013144|T033|FN|271782001|SNOMEDCT_CORE|Drowsy|Drowsy
C0013144|T033|SY|271782001|SNOMEDCT_CORE|Mental status, drowsy|Drowsy
C0013144|T033|SY|271782001|SNOMEDCT_CORE|Sleepiness|Drowsy
C0013144|T033|SY|271782001|SNOMEDCT_CORE|Sleepy|Drowsy
C0013144|T033|SY|271782001|SNOMEDCT_CORE|Somnolence|Drowsy
C0013146|T048|PT|26416006|SNOMEDCT_CORE|Drug abuse|Drug abuse
C0013146|T048|FN|26416006|SNOMEDCT_CORE|Drug abuse|Drug abuse
C0013146|T048|IS|26416006|SNOMEDCT_CORE|Drug abuse, NOS|Drug abuse
C0013146|T048|SY|26416006|SNOMEDCT_CORE|Medication abuse|Drug abuse
C0013182|T046|PT|416098002|SNOMEDCT_CORE|Allergy to drug|Allergy to drug
C0013182|T046|FN|416098002|SNOMEDCT_CORE|Allergy to drug|Allergy to drug
C0013182|T046|SY|416098002|SNOMEDCT_CORE|Drug allergy|Allergy to drug
C0013182|T046|OF|416098002|SNOMEDCT_CORE|Drug allergy|Allergy to drug
C0013182|T046|SY|416098002|SNOMEDCT_CORE|Medication allergy|Allergy to drug
C0013182|T046|SY|416098002|SNOMEDCT_CORE|Medicine allergy|Allergy to drug
C0013221|T037|SY|7895008|SNOMEDCT_CORE|Drug poisoning|Poisoning by drug AND/OR medicinal substance
C0013221|T037|IS|7895008|SNOMEDCT_CORE|Drug poisoning, NOS|Poisoning by drug AND/OR medicinal substance
C0013221|T037|SY|7895008|SNOMEDCT_CORE|Drug toxicity|Poisoning by drug AND/OR medicinal substance
C0013221|T037|SY|7895008|SNOMEDCT_CORE|Intoxication by drug|Poisoning by drug AND/OR medicinal substance
C0013221|T037|SY|7895008|SNOMEDCT_CORE|Intoxication caused by drug|Poisoning by drug AND/OR medicinal substance
C0013221|T037|SY|7895008|SNOMEDCT_CORE|Medicament poisoning|Poisoning by drug AND/OR medicinal substance
C0013221|T037|SY|7895008|SNOMEDCT_CORE|Medicinal poisoning|Poisoning by drug AND/OR medicinal substance
C0013221|T037|IS|7895008|SNOMEDCT_CORE|Overdose of drug with toxic effect|Poisoning by drug AND/OR medicinal substance
C0013221|T037|OF|7895008|SNOMEDCT_CORE|Poisoning by drug AND/OR medicinal substance|Poisoning by drug AND/OR medicinal substance
C0013221|T037|PT|7895008|SNOMEDCT_CORE|Poisoning by drug AND/OR medicinal substance|Poisoning by drug AND/OR medicinal substance
C0013221|T037|SY|7895008|SNOMEDCT_CORE|Poisoning by drug or medicinal substance|Poisoning by drug AND/OR medicinal substance
C0013221|T037|FN|7895008|SNOMEDCT_CORE|Poisoning caused by drug AND/OR medicinal substance|Poisoning by drug AND/OR medicinal substance
C0013221|T037|SY|7895008|SNOMEDCT_CORE|Poisoning caused by drug AND/OR medicinal substance|Poisoning by drug AND/OR medicinal substance
C0013221|T037|SY|7895008|SNOMEDCT_CORE|Poisoning caused by drug or medicinal substance|Poisoning by drug AND/OR medicinal substance
C0013221|T037|SY|7895008|SNOMEDCT_CORE|Therapeutic agent toxicity|Poisoning by drug AND/OR medicinal substance
C0013238|T047|SY|46152009|SNOMEDCT_CORE|Dry eye syndrome|Dry eye syndrome
C0013240|T047|PT|251331003|SNOMEDCT_CORE|Alveolar periostitis|Alveolar periostitis
C0013240|T047|FN|251331003|SNOMEDCT_CORE|Alveolar periostitis|Alveolar periostitis
C0013274|T019|SY|83330001|SNOMEDCT_CORE|Patent arterial duct|Patent ductus arteriosus
C0013274|T019|PT|83330001|SNOMEDCT_CORE|Patent ductus arteriosus|Patent ductus arteriosus
C0013274|T019|FN|83330001|SNOMEDCT_CORE|Patent ductus arteriosus|Patent ductus arteriosus
C0013274|T019|IS|83330001|SNOMEDCT_CORE|Patent ductus arteriosus - persisting type|Patent ductus arteriosus
C0013274|T019|SY|83330001|SNOMEDCT_CORE|Patent ductus Botalli|Patent ductus arteriosus
C0013274|T019|SY|83330001|SNOMEDCT_CORE|PDA - Patent ductus arteriosus|Patent ductus arteriosus
C0013274|T019|IS|83330001|SNOMEDCT_CORE|Persistent ductus arteriosus|Patent ductus arteriosus
C0013288|T047|SY|80193009|SNOMEDCT_CORE|Dumping syndrome|Dumping syndrome
C0013292|T047|PT|95532008|SNOMEDCT_CORE|Obstruction of duodenum|Obstruction of duodenum
C0013292|T047|FN|95532008|SNOMEDCT_CORE|Obstruction of duodenum|Obstruction of duodenum
C0013295|T047|SY|51868009|SNOMEDCT_CORE|DU - Duodenal ulcer|Ulcer of duodenum
C0013295|T047|SY|51868009|SNOMEDCT_CORE|DUD - Duodenal ulcer disease|Ulcer of duodenum
C0013295|T047|SY|51868009|SNOMEDCT_CORE|Duodenal ulcer|Ulcer of duodenum
C0013295|T047|SY|51868009|SNOMEDCT_CORE|Duodenal ulcer disease|Ulcer of duodenum
C0013295|T047|OF|51868009|SNOMEDCT_CORE|Duodenal ulcer disease|Ulcer of duodenum
C0013295|T047|IS|51868009|SNOMEDCT_CORE|Duodenal ulcer disease, NOS|Ulcer of duodenum
C0013295|T047|PT|51868009|SNOMEDCT_CORE|Ulcer of duodenum|Ulcer of duodenum
C0013295|T047|FN|51868009|SNOMEDCT_CORE|Ulcer of duodenum|Ulcer of duodenum
C0013298|T047|PT|72007001|SNOMEDCT_CORE|Duodenitis|Duodenitis
C0013298|T047|FN|72007001|SNOMEDCT_CORE|Duodenitis|Duodenitis
C0013298|T047|IS|72007001|SNOMEDCT_CORE|Duodenitis, NOS|Duodenitis
C0013312|T047|SY|274142002|SNOMEDCT_CORE|Dupuytren contracture|Dupuytren's contracture
C0013312|T047|PT|274142002|SNOMEDCT_CORE|Dupuytren's contracture|Dupuytren's contracture
C0013312|T047|FN|274142002|SNOMEDCT_CORE|Dupuytren's contracture|Dupuytren's contracture
C0013312|T047|SY|274142002|SNOMEDCT_CORE|Dupuytrens contracture|Dupuytren's contracture
C0013336|T019|SY|422065006|SNOMEDCT_CORE|Constitutional dwarfism|Constitutional short stature
C0013336|T019|PT|422065006|SNOMEDCT_CORE|Constitutional short stature|Constitutional short stature
C0013336|T019|FN|422065006|SNOMEDCT_CORE|Constitutional short stature|Constitutional short stature
C0013336|T019|IS|237836003|SNOMEDCT_CORE|Dwarf|Constitutional short stature
C0013336|T019|IS|237836003|SNOMEDCT_CORE|Dwarfism|Constitutional short stature
C0013336|T019|SY|422065006|SNOMEDCT_CORE|Physiologic dwarfism|Constitutional short stature
C0013336|T019|SY|237836003|SNOMEDCT_CORE|Short stature|Constitutional short stature
C0013336|T019|PT|237836003|SNOMEDCT_CORE|Short stature disorder|Constitutional short stature
C0013336|T019|FN|237836003|SNOMEDCT_CORE|Short stature disorder|Constitutional short stature
C0013338|T047|SY|367460001|SNOMEDCT_CORE|Hypopituitary dwarfism|Pituitary dwarfism
C0013338|T047|SY|367460001|SNOMEDCT_CORE|Hyposomatotropic dwarfism|Pituitary dwarfism
C0013338|T047|SY|367460001|SNOMEDCT_CORE|Isolated deficiency of growth hormone in children|Pituitary dwarfism
C0013338|T047|SY|367460001|SNOMEDCT_CORE|Lorain - Levi dwarfism|Pituitary dwarfism
C0013338|T047|PT|367460001|SNOMEDCT_CORE|Pituitary dwarfism|Pituitary dwarfism
C0013338|T047|FN|367460001|SNOMEDCT_CORE|Pituitary dwarfism|Pituitary dwarfism
C0013338|T047|SY|367460001|SNOMEDCT_CORE|Pituitary nanism|Pituitary dwarfism
C0013338|T047|SY|367460001|SNOMEDCT_CORE|Prepuberal dwarfism|Pituitary dwarfism
C0013338|T047|SY|367460001|SNOMEDCT_CORE|Prepubertal dwarfism|Pituitary dwarfism
C0013362|T048|PT|8011004|SNOMEDCT_CORE|Dysarthria|Dysarthria
C0013362|T048|FN|8011004|SNOMEDCT_CORE|Dysarthria|Dysarthria
C0013363|T047|SY|15241006|SNOMEDCT_CORE|Dysautonomia|Dysautonomia
C0013363|T047|IS|15241006|SNOMEDCT_CORE|Dysautonomia, NOS|Dysautonomia
C0013369|T047|OAP|111939009|SNOMEDCT_CORE|Dysentery|Dysentery
C0013369|T047|OAF|111939009|SNOMEDCT_CORE|Dysentery|Dysentery
C0013369|T047|IS|111939009|SNOMEDCT_CORE|Dysentery, NOS|Dysentery
C0013384|T047|PT|9748009|SNOMEDCT_CORE|Dyskinesia|Dyskinesia
C0013384|T047|FN|9748009|SNOMEDCT_CORE|Dyskinesia|Dyskinesia
C0013386|T047|IS|38941006|SNOMEDCT_CORE|Drug-induced dyskinesia|Drug-induced dyskinesia
C0013390|T047|PT|266599000|SNOMEDCT_CORE|Dysmenorrhea|Dysmenorrhea
C0013390|T047|FN|266599000|SNOMEDCT_CORE|Dysmenorrhea|Dysmenorrhea
C0013390|T047|PTGB|266599000|SNOMEDCT_CORE|Dysmenorrhoea|Dysmenorrhea
C0013390|T047|SY|266599000|SNOMEDCT_CORE|Menorrhalgia|Dysmenorrhea
C0013390|T047|SY|266599000|SNOMEDCT_CORE|Menstrual cramps|Dysmenorrhea
C0013390|T047|IS|266599000|SNOMEDCT_CORE|Painful menstruation|Dysmenorrhea
C0013390|T047|SY|266599000|SNOMEDCT_CORE|Period pain|Dysmenorrhea
C0013394|T047|IS|81712001|SNOMEDCT_CORE|Dyspareunia|Pain in female genitalia on intercourse
C0013394|T047|SY|81712001|SNOMEDCT_CORE|Female coitalgia|Pain in female genitalia on intercourse
C0013394|T047|PT|81712001|SNOMEDCT_CORE|Pain in female genitalia on intercourse|Pain in female genitalia on intercourse
C0013394|T047|FN|81712001|SNOMEDCT_CORE|Pain in female genitalia on intercourse|Pain in female genitalia on intercourse
C0013394|T047|IS|81712001|SNOMEDCT_CORE|Painful sexual act of female|Pain in female genitalia on intercourse
C0013395|T184|SY|162031009|SNOMEDCT_CORE|Dyspepsia|Indigestion
C0013395|T184|PT|162031009|SNOMEDCT_CORE|Indigestion|Indigestion
C0013395|T184|FN|162031009|SNOMEDCT_CORE|Indigestion|Indigestion
C0013403|T191|SY|254819008|SNOMEDCT_CORE|Atypical mole syndrome|B-K mole syndrome
C0013403|T191|FN|254819008|SNOMEDCT_CORE|Atypical mole syndrome|B-K mole syndrome
C0013403|T191|PT|254819008|SNOMEDCT_CORE|B-K mole syndrome|B-K mole syndrome
C0013403|T191|SY|254819008|SNOMEDCT_CORE|Familial atypical mole malignant melanoma syndrome|B-K mole syndrome
C0013403|T191|SY|254819008|SNOMEDCT_CORE|FAMMM - Familial atypical mole malignant melanoma syndrome|B-K mole syndrome
C0013404|T184|SY|267036007|SNOMEDCT_CORE|Breathless|Dyspnea
C0013404|T184|SY|267036007|SNOMEDCT_CORE|Breathlessness|Dyspnea
C0013404|T184|PT|267036007|SNOMEDCT_CORE|Dyspnea|Dyspnea
C0013404|T184|FN|267036007|SNOMEDCT_CORE|Dyspnea|Dyspnea
C0013404|T184|PTGB|267036007|SNOMEDCT_CORE|Dyspnoea|Dyspnea
C0013404|T184|SY|267036007|SNOMEDCT_CORE|Shortness of breath|Dyspnea
C0013404|T184|SY|267036007|SNOMEDCT_CORE|SOB - Shortness of breath|Dyspnea
C0013415|T048|PT|78667006|SNOMEDCT_CORE|Dysthymia|Dysthymia
C0013415|T048|FN|78667006|SNOMEDCT_CORE|Dysthymia|Dysthymia
C0013415|T048|IS|78667006|SNOMEDCT_CORE|Dysthymia, NOS|Dysthymia
C0013426|T047|PT|51689003|SNOMEDCT_CORE|Dystrophy of vulva|Dystrophy of vulva
C0013426|T047|FN|51689003|SNOMEDCT_CORE|Dystrophy of vulva|Dystrophy of vulva
C0013428|T184|PT|49650001|SNOMEDCT_CORE|Dysuria|Dysuria
C0013428|T184|FN|49650001|SNOMEDCT_CORE|Dysuria|Dysuria
C0013428|T184|IS|49650001|SNOMEDCT_CORE|Dysuria, NOS|Dysuria
C0013428|T184|SY|49650001|SNOMEDCT_CORE|Pain emptying bladder|Dysuria
C0013428|T184|SY|49650001|SNOMEDCT_CORE|Pain on micturition|Dysuria
C0013428|T184|SY|49650001|SNOMEDCT_CORE|Pain on voiding|Dysuria
C0013428|T184|SY|49650001|SNOMEDCT_CORE|Pain passing urine|Dysuria
C0013428|T184|SY|49650001|SNOMEDCT_CORE|Pain passing water|Dysuria
C0013428|T184|SY|49650001|SNOMEDCT_CORE|Painful micturition|Dysuria
C0013428|T184|SY|49650001|SNOMEDCT_CORE|Passing water hurts|Dysuria
C0013428|T184|SY|49650001|SNOMEDCT_CORE|Urination painful|Dysuria
C0013456|T184|SY|16001004|SNOMEDCT_CORE|Ear ache|Otalgia
C0013456|T184|SY|16001004|SNOMEDCT_CORE|Ear pain|Otalgia
C0013456|T184|SY|16001004|SNOMEDCT_CORE|Earache|Otalgia
C0013456|T184|IS|16001004|SNOMEDCT_CORE|Earache, NOS|Otalgia
C0013456|T184|PT|16001004|SNOMEDCT_CORE|Otalgia|Otalgia
C0013456|T184|OF|16001004|SNOMEDCT_CORE|Otalgia|Otalgia
C0013456|T184|FN|16001004|SNOMEDCT_CORE|Otalgia|Otalgia
C0013456|T184|IS|16001004|SNOMEDCT_CORE|Otalgia, NOS|Otalgia
C0013456|T184|SY|16001004|SNOMEDCT_CORE|Pain in ear|Otalgia
C0013456|T184|IS|16001004|SNOMEDCT_CORE|Pain in ear, NOS|Otalgia
C0013473|T048|PT|72366004|SNOMEDCT_CORE|Eating disorder|Eating disorder
C0013473|T048|FN|72366004|SNOMEDCT_CORE|Eating disorder|Eating disorder
C0013473|T048|IS|72366004|SNOMEDCT_CORE|Eating disorder, NOS|Eating disorder
C0013481|T019|SY|204357006|SNOMEDCT_CORE|Ebstein anomaly of tricuspid valve|Ebstein's anomaly
C0013481|T019|PT|204357006|SNOMEDCT_CORE|Ebstein's anomaly|Ebstein's anomaly
C0013481|T019|SY|204357006|SNOMEDCT_CORE|Ebstein's anomaly of tricuspid valve|Ebstein's anomaly
C0013481|T019|FN|204357006|SNOMEDCT_CORE|Ebstein's anomaly of tricuspid valve|Ebstein's anomaly
C0013481|T019|SY|204357006|SNOMEDCT_CORE|Ebstein's malformation of tricuspid valve|Ebstein's anomaly
C0013481|T019|SY|204357006|SNOMEDCT_CORE|Ebsteins anomaly|Ebstein's anomaly
C0013491|T046|PT|302227002|SNOMEDCT_CORE|Ecchymosis|Ecchymosis
C0013491|T046|FN|302227002|SNOMEDCT_CORE|Ecchymosis|Ecchymosis
C0013592|T047|PT|62909004|SNOMEDCT_CORE|Ectropion|Ectropion
C0013592|T047|SY|62909004|SNOMEDCT_CORE|Ectropion of eyelid|Ectropion
C0013592|T047|FN|62909004|SNOMEDCT_CORE|Ectropion of eyelid|Ectropion
C0013592|T047|IS|62909004|SNOMEDCT_CORE|Ectropion, NOS|Ectropion
C0013592|T047|SY|62909004|SNOMEDCT_CORE|Eversion of the eyelid|Ectropion
C0013592|T047|SY|62909004|SNOMEDCT_CORE|Eyelashes turned out|Ectropion
C0013592|T047|SY|62909004|SNOMEDCT_CORE|Eyelid everted|Ectropion
C0013592|T047|SY|62909004|SNOMEDCT_CORE|Eyelid turned out|Ectropion
C0013595|T047|PT|43116000|SNOMEDCT_CORE|Eczema|Eczema
C0013595|T047|OF|43116000|SNOMEDCT_CORE|Eczema|Eczema
C0013595|T047|FN|43116000|SNOMEDCT_CORE|Eczema|Eczema
C0013595|T047|IS|43116000|SNOMEDCT_CORE|Eczema, NOS|Eczema
C0013595|T047|IS|43116000|SNOMEDCT_CORE|Eczematous dermatitis|Eczema
C0013595|T047|IS|43116000|SNOMEDCT_CORE|Eczematous dermatitis, NOS|Eczema
C0013604|T046|PT|267038008|SNOMEDCT_CORE|Edema|Edema
C0013604|T046|FN|267038008|SNOMEDCT_CORE|Edema|Edema
C0013604|T046|SY|267038008|SNOMEDCT_CORE|Interstitial edema|Edema
C0013604|T046|SYGB|267038008|SNOMEDCT_CORE|Interstitial oedema|Edema
C0013604|T046|PTGB|267038008|SNOMEDCT_CORE|Oedema|Edema
C0013609|T046|PTGB|274724004|SNOMEDCT_CORE|Localised oedema|Localized edema
C0013609|T046|PT|274724004|SNOMEDCT_CORE|Localized edema|Localized edema
C0013609|T046|FN|274724004|SNOMEDCT_CORE|Localized edema|Localized edema
C0013720|T047|SY|398114001|SNOMEDCT_CORE|Cutis elastica|Ehlers-Danlos syndrome
C0013720|T047|SY|398114001|SNOMEDCT_CORE|Cutis hyperelastica|Ehlers-Danlos syndrome
C0013720|T047|SY|398114001|SNOMEDCT_CORE|Cutis hyperelastica dermatorrhexis|Ehlers-Danlos syndrome
C0013720|T047|SY|398114001|SNOMEDCT_CORE|Danlos disease|Ehlers-Danlos syndrome
C0013720|T047|SY|398114001|SNOMEDCT_CORE|Dystrophia mesodermalis congenita|Ehlers-Danlos syndrome
C0013720|T047|PT|398114001|SNOMEDCT_CORE|Ehlers-Danlos syndrome|Ehlers-Danlos syndrome
C0013720|T047|FN|398114001|SNOMEDCT_CORE|Ehlers-Danlos syndrome|Ehlers-Danlos syndrome
C0013720|T047|SY|398114001|SNOMEDCT_CORE|Fibrodysplasia elastica generalisata|Ehlers-Danlos syndrome
C0013720|T047|SY|398114001|SNOMEDCT_CORE|Hereditary collagen dysplasia|Ehlers-Danlos syndrome
C0013720|T047|SY|398114001|SNOMEDCT_CORE|India rubber skin|Ehlers-Danlos syndrome
C0013720|T047|SY|398114001|SNOMEDCT_CORE|Meekeren-Ehlers-Danlos syndrome|Ehlers-Danlos syndrome
C0014009|T047|PT|312682007|SNOMEDCT_CORE|Empyema|Empyema
C0014009|T047|FN|312682007|SNOMEDCT_CORE|Empyema|Empyema
C0014012|T047|PT|73125001|SNOMEDCT_CORE|Empyema of gallbladder|Empyema of gallbladder
C0014012|T047|FN|73125001|SNOMEDCT_CORE|Empyema of gallbladder|Empyema of gallbladder
C0014013|T047|PT|58554001|SNOMEDCT_CORE|Empyema of pleura|Empyema of pleura
C0014013|T047|FN|58554001|SNOMEDCT_CORE|Empyema of pleura|Empyema of pleura
C0014013|T047|IS|58554001|SNOMEDCT_CORE|Empyema of pleura, NOS|Empyema of pleura
C0014013|T047|SY|58554001|SNOMEDCT_CORE|Empyema thoracis|Empyema of pleura
C0014013|T047|SY|58554001|SNOMEDCT_CORE|Purulent pleurisy|Empyema of pleura
C0014013|T047|SY|58554001|SNOMEDCT_CORE|Pyothorax|Empyema of pleura
C0014013|T047|SY|58554001|SNOMEDCT_CORE|Suppurative pleurisy|Empyema of pleura
C0014038|T047|PT|45170000|SNOMEDCT_CORE|Encephalitis|Encephalitis
C0014038|T047|FN|45170000|SNOMEDCT_CORE|Encephalitis|Encephalitis
C0014038|T047|IS|45170000|SNOMEDCT_CORE|Encephalitis, NOS|Encephalitis
C0014060|T047|FN|417192005|SNOMEDCT_CORE|Saint Louis encephalitis virus infection|St. Louis encephalitis virus infection
C0014060|T047|SY|417192005|SNOMEDCT_CORE|Saint Louis encephalitis virus infection|St. Louis encephalitis virus infection
C0014060|T047|PT|417192005|SNOMEDCT_CORE|St. Louis encephalitis virus infection|St. Louis encephalitis virus infection
C0014060|T047|OF|417192005|SNOMEDCT_CORE|St. Louis encephalitis virus infection|St. Louis encephalitis virus infection
C0014060|T047|SY|417192005|SNOMEDCT_CORE|St. Louis viral disease|St. Louis encephalitis virus infection
C0014118|T047|PT|56819008|SNOMEDCT_CORE|Endocarditis|Endocarditis
C0014118|T047|FN|56819008|SNOMEDCT_CORE|Endocarditis|Endocarditis
C0014118|T047|IS|56819008|SNOMEDCT_CORE|Endocarditis, NOS|Endocarditis
C0014121|T047|PT|301183007|SNOMEDCT_CORE|Bacterial endocarditis|Bacterial endocarditis
C0014121|T047|FN|301183007|SNOMEDCT_CORE|Bacterial endocarditis|Bacterial endocarditis
C0014121|T047|SY|301183007|SNOMEDCT_CORE|BE - Bacterial endocarditis|Bacterial endocarditis
C0014122|T047|SY|73774007|SNOMEDCT_CORE|Endocarditis lenta|Subacute bacterial endocarditis
C0014122|T047|SY|73774007|SNOMEDCT_CORE|SBE|Subacute bacterial endocarditis
C0014122|T047|SY|73774007|SNOMEDCT_CORE|SBE - Subacute bacterial endocarditis|Subacute bacterial endocarditis
C0014122|T047|PT|73774007|SNOMEDCT_CORE|Subacute bacterial endocarditis|Subacute bacterial endocarditis
C0014122|T047|FN|73774007|SNOMEDCT_CORE|Subacute bacterial endocarditis|Subacute bacterial endocarditis
C0014126|T191|PT|8220004|SNOMEDCT_CORE|Endocervical polyp|Endocervical polyp
C0014126|T191|FN|8220004|SNOMEDCT_CORE|Endocervical polyp|Endocervical polyp
C0014130|T047|SY|362969004|SNOMEDCT_CORE|Disease of endocrine gland|Disorder of endocrine system
C0014130|T047|SY|362969004|SNOMEDCT_CORE|Disorder of endocrine gland|Disorder of endocrine system
C0014130|T047|FN|362969004|SNOMEDCT_CORE|Disorder of endocrine system|Disorder of endocrine system
C0014130|T047|PT|362969004|SNOMEDCT_CORE|Disorder of endocrine system|Disorder of endocrine system
C0014130|T047|SY|362969004|SNOMEDCT_CORE|Endocrine disease|Disorder of endocrine system
C0014130|T047|SY|362969004|SNOMEDCT_CORE|Endocrine disorder|Disorder of endocrine system
C0014130|T047|SY|362969004|SNOMEDCT_CORE|Endocrine disturbance|Disorder of endocrine system
C0014130|T047|SY|362969004|SNOMEDCT_CORE|Endocrine system disease|Disorder of endocrine system
C0014130|T047|SY|362969004|SNOMEDCT_CORE|Endocrinopathy|Disorder of endocrine system
C0014130|T047|SY|362969004|SNOMEDCT_CORE|Hormone disturbance|Disorder of endocrine system
C0014173|T047|PT|237072009|SNOMEDCT_CORE|Endometrial hyperplasia|Endometrial hyperplasia
C0014173|T047|FN|237072009|SNOMEDCT_CORE|Endometrial hyperplasia|Endometrial hyperplasia
C0014175|T047|SY|129103003|SNOMEDCT_CORE|Endometriosis|Endometriosis
C0014175|T047|PT|129103003|SNOMEDCT_CORE|Endometriosis|Endometriosis
C0014175|T047|FN|129103003|SNOMEDCT_CORE|Endometriosis|Endometriosis
C0014179|T047|PT|78623009|SNOMEDCT_CORE|Endometritis|Endometritis
C0014179|T047|FN|78623009|SNOMEDCT_CORE|Endometritis|Endometritis
C0014179|T047|IS|78623009|SNOMEDCT_CORE|Endometritis, NOS|Endometritis
C0014236|T047|PT|1847009|SNOMEDCT_CORE|Endophthalmitis|Endophthalmitis
C0014236|T047|FN|1847009|SNOMEDCT_CORE|Endophthalmitis|Endophthalmitis
C0014236|T047|IS|1847009|SNOMEDCT_CORE|Endophthalmitis, NOS|Endophthalmitis
C0014306|T047|SY|80093006|SNOMEDCT_CORE|Enophthalmia|Enophthalmos
C0014306|T047|PT|80093006|SNOMEDCT_CORE|Enophthalmos|Enophthalmos
C0014306|T047|FN|80093006|SNOMEDCT_CORE|Enophthalmos|Enophthalmos
C0014306|T047|IS|80093006|SNOMEDCT_CORE|Enophthalmos, NOS|Enophthalmos
C0014335|T047|SY|64613007|SNOMEDCT_CORE|Enteritis|Enteritis of small intestine
C0014335|T047|PT|64613007|SNOMEDCT_CORE|Enteritis of small intestine|Enteritis of small intestine
C0014335|T047|OF|64613007|SNOMEDCT_CORE|Enteritis, inflammatory disorder of small intestine|Enteritis of small intestine
C0014335|T047|SY|64613007|SNOMEDCT_CORE|Enteritis, inflammatory disorder of small intestine|Enteritis of small intestine
C0014335|T047|IS|64613007|SNOMEDCT_CORE|Enteritis, NOS|Enteritis of small intestine
C0014335|T047|SY|64613007|SNOMEDCT_CORE|Inflammation of small intestine|Enteritis of small intestine
C0014335|T047|FN|64613007|SNOMEDCT_CORE|Inflammation of small intestine|Enteritis of small intestine
C0014358|T047|OAP|397683000|SNOMEDCT_CORE|Pseudomembranous enterocolitis|Pseudomembranous enterocolitis
C0014358|T047|OAF|397683000|SNOMEDCT_CORE|Pseudomembranous enterocolitis|Pseudomembranous enterocolitis
C0014390|T047|PT|33168009|SNOMEDCT_CORE|Entropion|Entropion
C0014390|T047|OF|33168009|SNOMEDCT_CORE|Entropion|Entropion
C0014390|T047|SY|33168009|SNOMEDCT_CORE|Entropion of eyelid|Entropion
C0014390|T047|FN|33168009|SNOMEDCT_CORE|Entropion of eyelid|Entropion
C0014390|T047|IS|33168009|SNOMEDCT_CORE|Entropion, NOS|Entropion
C0014390|T047|SY|33168009|SNOMEDCT_CORE|Eyelashes turned in|Entropion
C0014390|T047|SY|33168009|SNOMEDCT_CORE|Eyelid inverted|Entropion
C0014390|T047|SY|33168009|SNOMEDCT_CORE|Eyelid turned in|Entropion
C0014390|T047|SY|33168009|SNOMEDCT_CORE|Folded in eyelid|Entropion
C0014394|T047|IS|8009008|SNOMEDCT_CORE|Enuresis|Enuresis
C0014474|T191|PT|443643007|SNOMEDCT_CORE|Ependymoma|Ependymoma
C0014474|T191|PT|57706008|SNOMEDCT_CORE|Ependymoma|Ependymoma
C0014474|T191|FN|443643007|SNOMEDCT_CORE|Ependymoma|Ependymoma
C0014474|T191|OF|57706008|SNOMEDCT_CORE|Ependymoma, no ICD-O subtype|Ependymoma
C0014474|T191|SY|57706008|SNOMEDCT_CORE|Ependymoma, no ICD-O subtype|Ependymoma
C0014474|T191|FN|57706008|SNOMEDCT_CORE|Ependymoma, no International Classification of Diseases for Oncology subtype|Ependymoma
C0014474|T191|SY|57706008|SNOMEDCT_CORE|Ependymoma, no International Classification of Diseases for Oncology subtype|Ependymoma
C0014474|T191|IS|57706008|SNOMEDCT_CORE|Ependymoma, NOS|Ependymoma
C0014474|T191|SY|57706008|SNOMEDCT_CORE|Epithelial ependymoma|Ependymoma
C0014488|T047|PT|73583000|SNOMEDCT_CORE|Epicondylitis|Epicondylitis
C0014488|T047|FN|73583000|SNOMEDCT_CORE|Epicondylitis|Epicondylitis
C0014488|T047|IS|73583000|SNOMEDCT_CORE|Epicondylitis, NOS|Epicondylitis
C0014511|T190|SY|419893006|SNOMEDCT_CORE|Epidermal cyst|Epidermoid cyst
C0014511|T190|IS|419603000|SNOMEDCT_CORE|Epidermal cyst|Epidermoid cyst
C0014511|T190|PT|419893006|SNOMEDCT_CORE|Epidermoid cyst|Epidermoid cyst
C0014511|T190|FN|419893006|SNOMEDCT_CORE|Epidermoid cyst|Epidermoid cyst
C0014511|T190|FN|419603000|SNOMEDCT_CORE|Epidermoid cyst of skin|Epidermoid cyst
C0014511|T190|PT|419603000|SNOMEDCT_CORE|Epidermoid cyst of skin|Epidermoid cyst
C0014511|T190|IS|419603000|SNOMEDCT_CORE|Epithelial cyst|Epidermoid cyst
C0014511|T190|IS|419603000|SNOMEDCT_CORE|Keratinous cyst|Epidermoid cyst
C0014511|T190|IS|419603000|SNOMEDCT_CORE|Sebaceous cyst|Epidermoid cyst
C0014534|T047|PT|31070006|SNOMEDCT_CORE|Epididymitis|Epididymitis
C0014534|T047|FN|31070006|SNOMEDCT_CORE|Epididymitis|Epididymitis
C0014534|T047|IS|31070006|SNOMEDCT_CORE|Epididymitis, NOS|Epididymitis
C0014544|T047|SY|84757009|SNOMEDCT_CORE|EP - Epilepsy|Epilepsy
C0014544|T047|IS|84757009|SNOMEDCT_CORE|Epilectic attack, NOS|Epilepsy
C0014544|T047|FN|84757009|SNOMEDCT_CORE|Epilepsy|Epilepsy
C0014544|T047|PT|84757009|SNOMEDCT_CORE|Epilepsy|Epilepsy
C0014544|T047|IS|84757009|SNOMEDCT_CORE|Epilepsy, NOS|Epilepsy
C0014544|T047|SY|84757009|SNOMEDCT_CORE|Epileptic|Epilepsy
C0014544|T047|IS|84757009|SNOMEDCT_CORE|Epileptic attack|Epilepsy
C0014544|T047|IS|84757009|SNOMEDCT_CORE|Epileptic attack, NOS|Epilepsy
C0014544|T047|IS|84757009|SNOMEDCT_CORE|Epileptic convulsions|Epilepsy
C0014544|T047|IS|84757009|SNOMEDCT_CORE|Epileptic convulsions, NOS|Epilepsy
C0014544|T047|SY|84757009|SNOMEDCT_CORE|Epileptic disorder|Epilepsy
C0014544|T047|IS|84757009|SNOMEDCT_CORE|Epileptic disorder, NOS|Epilepsy
C0014544|T047|IS|84757009|SNOMEDCT_CORE|Epileptic fits|Epilepsy
C0014544|T047|IS|84757009|SNOMEDCT_CORE|Epileptic fits, NOS|Epilepsy
C0014544|T047|IS|84757009|SNOMEDCT_CORE|Epileptic seizures|Epilepsy
C0014544|T047|IS|84757009|SNOMEDCT_CORE|Epileptic seizures, NOS|Epilepsy
C0014544|T047|FN|128613002|SNOMEDCT_CORE|Seizure disorder|Epilepsy
C0014544|T047|PT|128613002|SNOMEDCT_CORE|Seizure disorder|Epilepsy
C0014547|T047|IS|29753000|SNOMEDCT_CORE|Focal epilepsy|Localization-related epilepsy
C0014547|T047|SY|230381009|SNOMEDCT_CORE|Focal epilepsy|Localization-related epilepsy
C0014547|T047|SY|230381009|SNOMEDCT_CORE|Local epilepsy|Localization-related epilepsy
C0014547|T047|PTGB|230381009|SNOMEDCT_CORE|Localisation-related epilepsy|Localization-related epilepsy
C0014547|T047|PT|230381009|SNOMEDCT_CORE|Localization-related epilepsy|Localization-related epilepsy
C0014547|T047|FN|230381009|SNOMEDCT_CORE|Localization-related epilepsy|Localization-related epilepsy
C0014547|T047|SY|230381009|SNOMEDCT_CORE|Partial epilepsy|Localization-related epilepsy
C0014548|T047|PTGB|19598007|SNOMEDCT_CORE|Generalised epilepsy|Generalized epilepsy
C0014548|T047|PT|19598007|SNOMEDCT_CORE|Generalized epilepsy|Generalized epilepsy
C0014548|T047|FN|19598007|SNOMEDCT_CORE|Generalized epilepsy|Generalized epilepsy
C0014548|T047|IS|19598007|SNOMEDCT_CORE|Generalized epilepsy, NOS|Generalized epilepsy
C0014549|T047|SY|352818000|SNOMEDCT_CORE|Grand mal epilepsy|Tonic-clonic epilepsy
C0014549|T047|PT|352818000|SNOMEDCT_CORE|Tonic-clonic epilepsy|Tonic-clonic epilepsy
C0014549|T047|FN|352818000|SNOMEDCT_CORE|Tonic-clonic epilepsy|Tonic-clonic epilepsy
C0014553|T047|PT|79631006|SNOMEDCT_CORE|Absence seizure|Absence seizure
C0014553|T047|FN|79631006|SNOMEDCT_CORE|Absence seizure|Absence seizure
C0014553|T047|IS|79631006|SNOMEDCT_CORE|Absence seizures|Absence seizure
C0014553|T047|SY|79631006|SNOMEDCT_CORE|Petit mal|Absence seizure
C0014553|T047|SY|79631006|SNOMEDCT_CORE|Petit-mal seizure|Absence seizure
C0014583|T047|PT|815008|SNOMEDCT_CORE|Episcleritis|Episcleritis
C0014583|T047|FN|815008|SNOMEDCT_CORE|Episcleritis|Episcleritis
C0014583|T047|IS|815008|SNOMEDCT_CORE|Episcleritis, NOS|Episcleritis
C0014591|T046|PT|249366005|SNOMEDCT_CORE|Bleeding from nose|Bleeding from nose
C0014591|T046|FN|249366005|SNOMEDCT_CORE|Bleeding from nose|Bleeding from nose
C0014591|T046|SY|249366005|SNOMEDCT_CORE|Epistaxis|Bleeding from nose
C0014591|T046|OAP|12441001|SNOMEDCT_CORE|Epistaxis|Bleeding from nose
C0014591|T046|OAF|12441001|SNOMEDCT_CORE|Epistaxis|Bleeding from nose
C0014591|T046|SY|249366005|SNOMEDCT_CORE|Finding of bleeding of nose|Bleeding from nose
C0014591|T046|OAS|12441001|SNOMEDCT_CORE|Nasal haemorrhage|Bleeding from nose
C0014591|T046|SYGB|249366005|SNOMEDCT_CORE|Nasal haemorrhage|Bleeding from nose
C0014591|T046|OAS|12441001|SNOMEDCT_CORE|Nasal hemorrhage|Bleeding from nose
C0014591|T046|SY|249366005|SNOMEDCT_CORE|Nasal hemorrhage|Bleeding from nose
C0014591|T046|OAS|12441001|SNOMEDCT_CORE|Nose bleed|Bleeding from nose
C0014591|T046|OAS|12441001|SNOMEDCT_CORE|Nosebleed|Bleeding from nose
C0014591|T046|SY|249366005|SNOMEDCT_CORE|Nosebleed|Bleeding from nose
C0014591|T046|SY|249366005|SNOMEDCT_CORE|Observation of bleeding of nose|Bleeding from nose
C0014718|T047|SY|266158001|SNOMEDCT_CORE|Candida infection of flexural skin|Candidal intertrigo
C0014718|T047|SY|266158001|SNOMEDCT_CORE|Candida intertrigo|Candidal intertrigo
C0014718|T047|FN|266158001|SNOMEDCT_CORE|Candida intertrigo|Candidal intertrigo
C0014718|T047|PT|266158001|SNOMEDCT_CORE|Candidal intertrigo|Candidal intertrigo
C0014718|T047|SY|266158001|SNOMEDCT_CORE|Flexural candidosis|Candidal intertrigo
C0014724|T184|SY|271834000|SNOMEDCT_CORE|Belching|Burping
C0014724|T184|PT|271834000|SNOMEDCT_CORE|Burping|Burping
C0014724|T184|FN|271834000|SNOMEDCT_CORE|Burping|Burping
C0014724|T184|SY|271834000|SNOMEDCT_CORE|Eructation|Burping
C0014733|T047|PT|44653001|SNOMEDCT_CORE|Erysipelas|Erysipelas
C0014733|T047|FN|44653001|SNOMEDCT_CORE|Erysipelas|Erysipelas
C0014733|T047|SY|44653001|SNOMEDCT_CORE|Patch of erysipelas|Erysipelas
C0014742|T047|SY|36715001|SNOMEDCT_CORE|EM - Erythema multiforme|Erythema multiforme
C0014742|T047|PT|36715001|SNOMEDCT_CORE|Erythema multiforme|Erythema multiforme
C0014742|T047|FN|36715001|SNOMEDCT_CORE|Erythema multiforme|Erythema multiforme
C0014742|T047|IS|36715001|SNOMEDCT_CORE|Erythema multiforme, NOS|Erythema multiforme
C0014742|T047|SY|36715001|SNOMEDCT_CORE|Target lesion|Erythema multiforme
C0014743|T047|SY|32861005|SNOMEDCT_CORE|EN - Erythema nodosum|Erythema nodosum
C0014743|T047|PT|32861005|SNOMEDCT_CORE|Erythema nodosum|Erythema nodosum
C0014743|T047|FN|32861005|SNOMEDCT_CORE|Erythema nodosum|Erythema nodosum
C0014743|T047|IS|32861005|SNOMEDCT_CORE|Erythema nodosum, NOS|Erythema nodosum
C0014804|T047|SY|37151006|SNOMEDCT_CORE|Erythermalgia|Erythromelalgia
C0014804|T047|SY|37151006|SNOMEDCT_CORE|Erythralgia|Erythromelalgia
C0014804|T047|PT|37151006|SNOMEDCT_CORE|Erythromelalgia|Erythromelalgia
C0014804|T047|FN|37151006|SNOMEDCT_CORE|Erythromelalgia|Erythromelalgia
C0014804|T047|SY|37151006|SNOMEDCT_CORE|Weir Mitchell's disease|Erythromelalgia
C0014836|T047|SY|71057007|SNOMEDCT_CORE|Bacterial infection caused by E. coli|Infection due to Escherichia coli
C0014836|T047|SY|71057007|SNOMEDCT_CORE|Bacterial infection due to E. coli|Infection due to Escherichia coli
C0014836|T047|IS|71057007|SNOMEDCT_CORE|Bacterial infection due to E. coli, NOS|Infection due to Escherichia coli
C0014836|T047|SY|71057007|SNOMEDCT_CORE|Colibacillosis|Infection due to Escherichia coli
C0014836|T047|SY|71057007|SNOMEDCT_CORE|E. coli infection|Infection due to Escherichia coli
C0014836|T047|SY|71057007|SNOMEDCT_CORE|Escherichia coli infection|Infection due to Escherichia coli
C0014836|T047|SY|71057007|SNOMEDCT_CORE|Infection caused by Escherichia coli|Infection due to Escherichia coli
C0014836|T047|FN|71057007|SNOMEDCT_CORE|Infection caused by Escherichia coli|Infection due to Escherichia coli
C0014836|T047|PT|71057007|SNOMEDCT_CORE|Infection due to Escherichia coli|Infection due to Escherichia coli
C0014836|T047|OF|71057007|SNOMEDCT_CORE|Infection due to Escherichia coli|Infection due to Escherichia coli
C0014836|T047|IS|71057007|SNOMEDCT_CORE|Infection due to Escherichia coli, NOS|Infection due to Escherichia coli
C0014848|T047|SY|45564002|SNOMEDCT_CORE|Achalasia of cardia|Achalasia of esophagus
C0014848|T047|PT|45564002|SNOMEDCT_CORE|Achalasia of esophagus|Achalasia of esophagus
C0014848|T047|FN|45564002|SNOMEDCT_CORE|Achalasia of esophagus|Achalasia of esophagus
C0014848|T047|PTGB|45564002|SNOMEDCT_CORE|Achalasia of oesophagus|Achalasia of esophagus
C0014848|T047|SY|45564002|SNOMEDCT_CORE|Cardiospasm|Achalasia of esophagus
C0014848|T047|IS|45564002|SNOMEDCT_CORE|Cardiospasm, NOS|Achalasia of esophagus
C0014848|T047|IS|45564002|SNOMEDCT_CORE|Hypertensive lower esophageal sphincter|Achalasia of esophagus
C0014848|T047|IS|45564002|SNOMEDCT_CORE|Hypertensive lower oesophageal sphincter|Achalasia of esophagus
C0014848|T047|SY|45564002|SNOMEDCT_CORE|Lack of reflex relaxation of lower esophageal sphincter|Achalasia of esophagus
C0014848|T047|SYGB|45564002|SNOMEDCT_CORE|Lack of reflex relaxation of lower oesophageal sphincter|Achalasia of esophagus
C0014848|T047|IS|45564002|SNOMEDCT_CORE|Megaoesophagus|Achalasia of esophagus
C0014852|T047|IS|37657006|SNOMEDCT_CORE|Disease of esophagus|Disorder of esophagus
C0014852|T047|OF|37657006|SNOMEDCT_CORE|Disease of esophagus|Disorder of esophagus
C0014852|T047|IS|37657006|SNOMEDCT_CORE|Disease of esophagus, NOS|Disorder of esophagus
C0014852|T047|IS|37657006|SNOMEDCT_CORE|Disease of oesophagus|Disorder of esophagus
C0014852|T047|PT|37657006|SNOMEDCT_CORE|Disorder of esophagus|Disorder of esophagus
C0014852|T047|FN|37657006|SNOMEDCT_CORE|Disorder of esophagus|Disorder of esophagus
C0014852|T047|IS|37657006|SNOMEDCT_CORE|Disorder of esophagus, NOS|Disorder of esophagus
C0014852|T047|PTGB|37657006|SNOMEDCT_CORE|Disorder of oesophagus|Disorder of esophagus
C0014858|T047|SY|79962008|SNOMEDCT_CORE|Dyskinesia of esophagus|Esophageal dysmotility
C0014858|T047|SYGB|79962008|SNOMEDCT_CORE|Dyskinesia of oesophagus|Esophageal dysmotility
C0014858|T047|IS|79962008|SNOMEDCT_CORE|Esophageal dysmotility|Esophageal dysmotility
C0014858|T047|PT|266434009|SNOMEDCT_CORE|Esophageal dysmotility|Esophageal dysmotility
C0014858|T047|FN|266434009|SNOMEDCT_CORE|Esophageal dysmotility|Esophageal dysmotility
C0014858|T047|SY|79962008|SNOMEDCT_CORE|Esophageal motility disorder|Esophageal dysmotility
C0014858|T047|SY|79962008|SNOMEDCT_CORE|Esophageal motor disorder|Esophageal dysmotility
C0014858|T047|IS|79962008|SNOMEDCT_CORE|Oesophageal dysmotility|Esophageal dysmotility
C0014858|T047|PTGB|266434009|SNOMEDCT_CORE|Oesophageal dysmotility|Esophageal dysmotility
C0014858|T047|SYGB|79962008|SNOMEDCT_CORE|Oesophageal motility disorder|Esophageal dysmotility
C0014858|T047|SYGB|79962008|SNOMEDCT_CORE|Oesophageal motor disorder|Esophageal dysmotility
C0014863|T047|SY|79962008|SNOMEDCT_CORE|Diffuse esophageal spasm|Diffuse spasm of esophagus
C0014863|T047|SYGB|79962008|SNOMEDCT_CORE|Diffuse oesophageal spasm|Diffuse spasm of esophagus
C0014863|T047|PT|79962008|SNOMEDCT_CORE|Diffuse spasm of esophagus|Diffuse spasm of esophagus
C0014863|T047|FN|79962008|SNOMEDCT_CORE|Diffuse spasm of esophagus|Diffuse spasm of esophagus
C0014863|T047|PTGB|79962008|SNOMEDCT_CORE|Diffuse spasm of oesophagus|Diffuse spasm of esophagus
C0014863|T047|SY|79962008|SNOMEDCT_CORE|DOS - Diffuse esophageal spasm|Diffuse spasm of esophagus
C0014863|T047|SYGB|79962008|SNOMEDCT_CORE|DOS - Diffuse oesophageal spasm|Diffuse spasm of esophagus
C0014863|T047|SY|79962008|SNOMEDCT_CORE|ES - Esophageal spasm|Diffuse spasm of esophagus
C0014863|T047|SYGB|79962008|SNOMEDCT_CORE|ES - Oesophageal spasm|Diffuse spasm of esophagus
C0014863|T047|SY|79962008|SNOMEDCT_CORE|Esophageal spasm|Diffuse spasm of esophagus
C0014863|T047|SY|79962008|SNOMEDCT_CORE|Esophagism|Diffuse spasm of esophagus
C0014863|T047|SY|79962008|SNOMEDCT_CORE|Esophagospasm|Diffuse spasm of esophagus
C0014863|T047|SYGB|79962008|SNOMEDCT_CORE|Oesophageal spasm|Diffuse spasm of esophagus
C0014863|T047|SYGB|79962008|SNOMEDCT_CORE|Oesophagism|Diffuse spasm of esophagus
C0014863|T047|SYGB|79962008|SNOMEDCT_CORE|Oesophagospasm|Diffuse spasm of esophagus
C0014863|T047|IS|79962008|SNOMEDCT_CORE|OS - Esophageal spasm|Diffuse spasm of esophagus
C0014863|T047|SYGB|79962008|SNOMEDCT_CORE|OS - Oesophageal spasm|Diffuse spasm of esophagus
C0014863|T047|SY|79962008|SNOMEDCT_CORE|Spasm of esophagus|Diffuse spasm of esophagus
C0014863|T047|SYGB|79962008|SNOMEDCT_CORE|Spasm of oesophagus|Diffuse spasm of esophagus
C0014866|T047|OAS|33282003|SNOMEDCT_CORE|Esophageal stenosis|Esophagostenosis
C0014866|T047|IS|63305008|SNOMEDCT_CORE|Esophagostenosis|Esophagostenosis
C0014866|T047|OAS|33282003|SNOMEDCT_CORE|Oesophageal stenosis|Esophagostenosis
C0014866|T047|IS|63305008|SNOMEDCT_CORE|Oesophagostenosis|Esophagostenosis
C0014866|T047|OAP|33282003|SNOMEDCT_CORE|Stenosis of esophagus|Esophagostenosis
C0014866|T047|IS|63305008|SNOMEDCT_CORE|Stenosis of esophagus|Esophagostenosis
C0014866|T047|OAF|33282003|SNOMEDCT_CORE|Stenosis of esophagus|Esophagostenosis
C0014866|T047|OAP|33282003|SNOMEDCT_CORE|Stenosis of oesophagus|Esophagostenosis
C0014866|T047|IS|63305008|SNOMEDCT_CORE|Stenosis of oesophagus|Esophagostenosis
C0014867|T047|PT|28670008|SNOMEDCT_CORE|Esophageal varices|Esophageal varices
C0014867|T047|FN|28670008|SNOMEDCT_CORE|Esophageal varices|Esophageal varices
C0014867|T047|IS|28670008|SNOMEDCT_CORE|Esophageal varices, NOS|Esophageal varices
C0014867|T047|SY|28670008|SNOMEDCT_CORE|Esophageal varix|Esophageal varices
C0014867|T047|PTGB|28670008|SNOMEDCT_CORE|Oesophageal varices|Esophageal varices
C0014867|T047|IS|28670008|SNOMEDCT_CORE|Oesophageal varices, NOS|Esophageal varices
C0014867|T047|SYGB|28670008|SNOMEDCT_CORE|Oesophageal varix|Esophageal varices
C0014867|T047|SY|28670008|SNOMEDCT_CORE|OV - Esophageal varices|Esophageal varices
C0014867|T047|SYGB|28670008|SNOMEDCT_CORE|OV - Oesophageal varices|Esophageal varices
C0014868|T047|PT|16761005|SNOMEDCT_CORE|Esophagitis|Esophagitis
C0014868|T047|FN|16761005|SNOMEDCT_CORE|Esophagitis|Esophagitis
C0014868|T047|IS|16761005|SNOMEDCT_CORE|Esophagitis, NOS|Esophagitis
C0014868|T047|PTGB|16761005|SNOMEDCT_CORE|Oesophagitis|Esophagitis
C0014868|T047|IS|16761005|SNOMEDCT_CORE|Oesophagitis, NOS|Esophagitis
C0014869|T047|IS|57643001|SNOMEDCT_CORE|Peptic esophagitis|Peptic reflux disease
C0014869|T047|IS|57643001|SNOMEDCT_CORE|Peptic oesophagitis|Peptic reflux disease
C0014869|T047|OAP|57643001|SNOMEDCT_CORE|Peptic reflux disease|Peptic reflux disease
C0014869|T047|OAF|57643001|SNOMEDCT_CORE|Peptic reflux disease|Peptic reflux disease
C0014869|T047|OAS|57643001|SNOMEDCT_CORE|Peptic reflux esophagitis|Peptic reflux disease
C0014869|T047|OAS|57643001|SNOMEDCT_CORE|Peptic reflux oesophagitis|Peptic reflux disease
C0014877|T047|SY|16596007|SNOMEDCT_CORE|Convergent squint|Esotropia
C0014877|T047|SY|16596007|SNOMEDCT_CORE|Convergent strabismus|Esotropia
C0014877|T047|SY|16596007|SNOMEDCT_CORE|Cross-eye|Esotropia
C0014877|T047|PT|16596007|SNOMEDCT_CORE|Esotropia|Esotropia
C0014877|T047|FN|16596007|SNOMEDCT_CORE|Esotropia|Esotropia
C0014877|T047|IS|16596007|SNOMEDCT_CORE|Esotropia, NOS|Esotropia
C0015029|T047|PT|18643000|SNOMEDCT_CORE|Ethmoidal sinusitis|Ethmoidal sinusitis
C0015029|T047|FN|18643000|SNOMEDCT_CORE|Ethmoidal sinusitis|Ethmoidal sinusitis
C0015029|T047|IS|18643000|SNOMEDCT_CORE|Ethmoidal sinusitis, NOS|Ethmoidal sinusitis
C0015230|T184|SY|271807003|SNOMEDCT_CORE|Breaking out - eruption|Eruption
C0015230|T184|PT|271807003|SNOMEDCT_CORE|Eruption|Eruption
C0015230|T184|OF|271807003|SNOMEDCT_CORE|Eruption|Eruption
C0015230|T184|SY|271807003|SNOMEDCT_CORE|Eruption of skin|Eruption
C0015230|T184|FN|271807003|SNOMEDCT_CORE|Eruption of skin|Eruption
C0015230|T184|SY|271807003|SNOMEDCT_CORE|Exanthem|Eruption
C0015230|T184|SY|271807003|SNOMEDCT_CORE|Rash|Eruption
C0015230|T184|SY|271807003|SNOMEDCT_CORE|Skin eruption|Eruption
C0015230|T184|SY|271807003|SNOMEDCT_CORE|Skin rash|Eruption
C0015231|T047|SY|54385001|SNOMEDCT_CORE|Exanthem subitum|Exanthema subitum
C0015231|T047|PT|54385001|SNOMEDCT_CORE|Exanthema subitum|Exanthema subitum
C0015231|T047|FN|54385001|SNOMEDCT_CORE|Exanthema subitum|Exanthema subitum
C0015231|T047|SY|54385001|SNOMEDCT_CORE|Pseudorubella|Exanthema subitum
C0015231|T047|SY|54385001|SNOMEDCT_CORE|Roseola infantum|Exanthema subitum
C0015231|T047|SY|54385001|SNOMEDCT_CORE|Sixth disease|Exanthema subitum
C0015231|T047|SY|54385001|SNOMEDCT_CORE|Three day fever|Exanthema subitum
C0015256|T037|PT|247444006|SNOMEDCT_CORE|Excoriation of skin|Excoriation of skin
C0015256|T037|FN|247444006|SNOMEDCT_CORE|Excoriation of skin|Excoriation of skin
C0015300|T047|SY|18265008|SNOMEDCT_CORE|Exophthalmia|Exophthalmos
C0015300|T047|PT|18265008|SNOMEDCT_CORE|Exophthalmos|Exophthalmos
C0015300|T047|FN|18265008|SNOMEDCT_CORE|Exophthalmos|Exophthalmos
C0015300|T047|IS|18265008|SNOMEDCT_CORE|Exophthalmos, NOS|Exophthalmos
C0015300|T047|SY|18265008|SNOMEDCT_CORE|Eye displaced forwards|Exophthalmos
C0015300|T047|SY|18265008|SNOMEDCT_CORE|Proptosis|Exophthalmos
C0015300|T047|IS|18265008|SNOMEDCT_CORE|Proptosis, NOS|Exophthalmos
C0015310|T047|SY|399054005|SNOMEDCT_CORE|Divergent squint|Exotropia
C0015310|T047|SY|399054005|SNOMEDCT_CORE|Divergent strabismus|Exotropia
C0015310|T047|PT|399054005|SNOMEDCT_CORE|Exotropia|Exotropia
C0015310|T047|FN|399054005|SNOMEDCT_CORE|Exotropia|Exotropia
C0015310|T047|SY|399054005|SNOMEDCT_CORE|External strabismus|Exotropia
C0015310|T047|SY|399054005|SNOMEDCT_CORE|XT - Exotropia|Exotropia
C0015371|T047|PT|76349003|SNOMEDCT_CORE|Extrapyramidal disease|Extrapyramidal disease
C0015371|T047|FN|76349003|SNOMEDCT_CORE|Extrapyramidal disease|Extrapyramidal disease
C0015371|T047|IS|76349003|SNOMEDCT_CORE|Extrapyramidal disease, NOS|Extrapyramidal disease
C0015371|T047|SY|76349003|SNOMEDCT_CORE|Extrapyramidal disorder|Extrapyramidal disease
C0015371|T047|IS|76349003|SNOMEDCT_CORE|Extrapyramidal disorder, NOS|Extrapyramidal disease
C0015393|T019|SY|19416009|SNOMEDCT_CORE|Congenital abnormality of eye|Congenital anomaly of eye
C0015393|T019|IS|19416009|SNOMEDCT_CORE|Congenital anolmaly of eye|Congenital anomaly of eye
C0015393|T019|IS|19416009|SNOMEDCT_CORE|Congenital anolmaly of the globe|Congenital anomaly of eye
C0015393|T019|PT|19416009|SNOMEDCT_CORE|Congenital anomaly of eye|Congenital anomaly of eye
C0015393|T019|FN|19416009|SNOMEDCT_CORE|Congenital anomaly of eye|Congenital anomaly of eye
C0015393|T019|IS|19416009|SNOMEDCT_CORE|Congenital anomaly of eye, NOS|Congenital anomaly of eye
C0015393|T019|SY|19416009|SNOMEDCT_CORE|Congenital anomaly of the globe|Congenital anomaly of eye
C0015393|T019|SY|19416009|SNOMEDCT_CORE|Congenital deformity of eye|Congenital anomaly of eye
C0015393|T019|IS|19416009|SNOMEDCT_CORE|Congenital deformity of eye, NOS|Congenital anomaly of eye
C0015393|T019|SY|19416009|SNOMEDCT_CORE|Congenital eye anomalies|Congenital anomaly of eye
C0015393|T019|SY|19416009|SNOMEDCT_CORE|Congenital malformation of eye|Congenital anomaly of eye
C0015397|T047|SY|371405004|SNOMEDCT_CORE|Disease of eyeball|Disorder of eye
C0015397|T047|IS|371409005|SNOMEDCT_CORE|Disorder of eye|Disorder of eye
C0015397|T047|PT|371405004|SNOMEDCT_CORE|Disorder of eye|Disorder of eye
C0015397|T047|FN|371405004|SNOMEDCT_CORE|Disorder of eye proper|Disorder of eye
C0015397|T047|SY|371405004|SNOMEDCT_CORE|Disorder of eye proper|Disorder of eye
C0015397|T047|FN|371409005|SNOMEDCT_CORE|Disorder of eye region|Disorder of eye
C0015397|T047|PT|371409005|SNOMEDCT_CORE|Disorder of eye region|Disorder of eye
C0015397|T047|SY|371405004|SNOMEDCT_CORE|Disorder of eyeball|Disorder of eye
C0015397|T047|SY|371405004|SNOMEDCT_CORE|Disorder of globe|Disorder of eye
C0015397|T047|SY|371409005|SNOMEDCT_CORE|Disorder of orbital region|Disorder of eye
C0015397|T047|IS|371409005|SNOMEDCT_CORE|Eye disorder|Disorder of eye
C0015397|T047|SY|371405004|SNOMEDCT_CORE|Eye disorder|Disorder of eye
C0015397|T047|SY|371409005|SNOMEDCT_CORE|Ophthalmological disorder|Disorder of eye
C0015401|T037|SY|82576008|SNOMEDCT_CORE|Foreign body in eye|Retained foreign body in eye
C0015401|T037|SY|82576008|SNOMEDCT_CORE|Foreign body in eyeball|Retained foreign body in eye
C0015401|T037|SY|82576008|SNOMEDCT_CORE|Intraocular foreign body|Retained foreign body in eye
C0015401|T037|SY|82576008|SNOMEDCT_CORE|IOFB - Intraocular foreign body|Retained foreign body in eye
C0015401|T037|PT|82576008|SNOMEDCT_CORE|Retained foreign body in eye|Retained foreign body in eye
C0015401|T037|FN|82576008|SNOMEDCT_CORE|Retained foreign body in eye|Retained foreign body in eye
C0015401|T037|IS|82576008|SNOMEDCT_CORE|Retained foreign body in eye, NOS|Retained foreign body in eye
C0015401|T037|SY|82576008|SNOMEDCT_CORE|Retained intraocular foreign body|Retained foreign body in eye
C0015401|T037|IS|82576008|SNOMEDCT_CORE|Retained intraocular foreign body, NOS|Retained foreign body in eye
C0015403|T047|PT|128351009|SNOMEDCT_CORE|Eye infection|Eye infection
C0015403|T047|FN|128351009|SNOMEDCT_CORE|Eye infection|Eye infection
C0015403|T047|IS|128351009|SNOMEDCT_CORE|Periocular infection|Eye infection
C0015408|T037|IS|367423000|SNOMEDCT_CORE|Injury of eye, NOS|Injury of eye, NOS
C0015423|T047|PT|60113004|SNOMEDCT_CORE|Disorder of eyelid|Disorder of eyelid
C0015423|T047|FN|60113004|SNOMEDCT_CORE|Disorder of eyelid|Disorder of eyelid
C0015423|T047|IS|60113004|SNOMEDCT_CORE|Disorder of eyelid, NOS|Disorder of eyelid
C0015459|T037|SY|125593007|SNOMEDCT_CORE|Face injury|Injury of face
C0015459|T037|SY|125593007|SNOMEDCT_CORE|Facial injury|Injury of face
C0015459|T037|PT|125593007|SNOMEDCT_CORE|Injury of face|Injury of face
C0015459|T037|FN|125593007|SNOMEDCT_CORE|Injury of face|Injury of face
C0015464|T047|SY|422426003|SNOMEDCT_CORE|Disorder of facial nerve|Facial nerve disorder
C0015464|T047|SY|422426003|SNOMEDCT_CORE|Disorder of seventh cranial nerve|Facial nerve disorder
C0015464|T047|SY|422426003|SNOMEDCT_CORE|Disorders of the seventh nerve|Facial nerve disorder
C0015464|T047|SY|422426003|SNOMEDCT_CORE|Disorders of the VIIth cranial nerve|Facial nerve disorder
C0015464|T047|PT|422426003|SNOMEDCT_CORE|Facial nerve disorder|Facial nerve disorder
C0015464|T047|FN|422426003|SNOMEDCT_CORE|Facial nerve disorder|Facial nerve disorder
C0015464|T047|SY|422426003|SNOMEDCT_CORE|Facial neuropathy|Facial nerve disorder
C0015468|T184|SY|95668009|SNOMEDCT_CORE|Facial pain|Pain in face
C0015468|T184|IS|95668009|SNOMEDCT_CORE|Facial pain, NOS|Pain in face
C0015468|T184|PT|95668009|SNOMEDCT_CORE|Pain in face|Pain in face
C0015468|T184|FN|95668009|SNOMEDCT_CORE|Pain in face|Pain in face
C0015468|T184|SY|95668009|SNOMEDCT_CORE|Pain of face|Pain in face
C0015468|T184|IS|95668009|SNOMEDCT_CORE|Pain of face, NOS|Pain in face
C0015469|T047|SY|280816001|SNOMEDCT_CORE|Facial nerve paralysis|Facial palsy
C0015469|T047|PT|280816001|SNOMEDCT_CORE|Facial palsy|Facial palsy
C0015469|T047|FN|280816001|SNOMEDCT_CORE|Facial palsy|Facial palsy
C0015544|T047|PT|54840006|SNOMEDCT_CORE|Failure to thrive|Failure to thrive
C0015544|T047|FN|54840006|SNOMEDCT_CORE|Failure to thrive|Failure to thrive
C0015544|T047|IS|54840006|SNOMEDCT_CORE|Failure to thrive syndrome|Failure to thrive
C0015544|T047|SY|54840006|SNOMEDCT_CORE|Faltering growth|Failure to thrive
C0015544|T047|SY|54840006|SNOMEDCT_CORE|FTT - failure to thrive|Failure to thrive
C0015544|T047|IS|54840006|SNOMEDCT_CORE|FTT - Failure to thrive|Failure to thrive
C0015582|T033|PT|28332004|SNOMEDCT_CORE|Family disruption|Family disruption
C0015582|T033|FN|28332004|SNOMEDCT_CORE|Family disruption|Family disruption
C0015643|T047|SY|6374002|SNOMEDCT_CORE|Fascicular block|Fascicular block
C0015644|T184|IS|82470000|SNOMEDCT_CORE|Fasciculation|Muscle fasciculation
C0015644|T184|SY|82470000|SNOMEDCT_CORE|Flickering muscles|Muscle fasciculation
C0015644|T184|SY|82470000|SNOMEDCT_CORE|Fluttering muscles|Muscle fasciculation
C0015644|T184|PT|82470000|SNOMEDCT_CORE|Muscle fasciculation|Muscle fasciculation
C0015644|T184|FN|82470000|SNOMEDCT_CORE|Muscle fasciculation|Muscle fasciculation
C0015644|T184|SY|82470000|SNOMEDCT_CORE|Muscular fasciculation|Muscle fasciculation
C0015644|T184|SY|82470000|SNOMEDCT_CORE|Spontaneous contraction of muscle|Muscle fasciculation
C0015644|T184|SY|82470000|SNOMEDCT_CORE|Writhing muscles|Muscle fasciculation
C0015645|T047|PT|36948007|SNOMEDCT_CORE|Fasciitis|Fasciitis
C0015645|T047|FN|36948007|SNOMEDCT_CORE|Fasciitis|Fasciitis
C0015645|T047|IS|36948007|SNOMEDCT_CORE|Fasciitis, NOS|Fasciitis
C0015672|T184|PT|84229001|SNOMEDCT_CORE|Fatigue|Fatigue
C0015672|T184|FN|84229001|SNOMEDCT_CORE|Fatigue|Fatigue
C0015672|T184|IS|84229001|SNOMEDCT_CORE|Tiredness|Fatigue
C0015672|T184|SY|84229001|SNOMEDCT_CORE|Weariness|Fatigue
C0015674|T047|IS|52702003|SNOMEDCT_CORE|Akureyri disease|Chronic fatigue syndrome
C0015674|T047|SY|52702003|SNOMEDCT_CORE|Benign myalgic encephalomyelitis|Chronic fatigue syndrome
C0015674|T047|SY|52702003|SNOMEDCT_CORE|CFS - Chronic fatigue syndrome|Chronic fatigue syndrome
C0015674|T047|PT|52702003|SNOMEDCT_CORE|Chronic fatigue syndrome|Chronic fatigue syndrome
C0015674|T047|FN|52702003|SNOMEDCT_CORE|Chronic fatigue syndrome|Chronic fatigue syndrome
C0015674|T047|IS|52702003|SNOMEDCT_CORE|Epidemic neuromyasthenia|Chronic fatigue syndrome
C0015674|T047|SY|52702003|SNOMEDCT_CORE|Iceland disease|Chronic fatigue syndrome
C0015674|T047|SY|52702003|SNOMEDCT_CORE|ME - Myalgic encephalomyelitis|Chronic fatigue syndrome
C0015674|T047|SY|52702003|SNOMEDCT_CORE|Myalgic encephalomyelitis|Chronic fatigue syndrome
C0015674|T047|SY|52702003|SNOMEDCT_CORE|Myalgic encephalomyelitis syndrome|Chronic fatigue syndrome
C0015674|T047|IS|52702003|SNOMEDCT_CORE|Postviral fatigue syndrome|Chronic fatigue syndrome
C0015674|T047|IS|52702003|SNOMEDCT_CORE|PVFS - Postviral fatigue syndrome|Chronic fatigue syndrome
C0015695|T047|OAP|371330000|SNOMEDCT_CORE|Fatty liver|Hepatic lipidosis
C0015695|T047|SY|197321007|SNOMEDCT_CORE|Fatty liver|Hepatic lipidosis
C0015695|T047|OAF|371330000|SNOMEDCT_CORE|Fatty liver|Hepatic lipidosis
C0015695|T047|OAS|371330000|SNOMEDCT_CORE|Hepatic lipidosis|Hepatic lipidosis
C0015695|T047|SY|197321007|SNOMEDCT_CORE|Hepatic lipidosis|Hepatic lipidosis
C0015696|T047|PT|50325005|SNOMEDCT_CORE|Alcoholic fatty liver|Alcoholic fatty liver
C0015696|T047|FN|50325005|SNOMEDCT_CORE|Alcoholic fatty liver|Alcoholic fatty liver
C0015696|T047|SY|50325005|SNOMEDCT_CORE|Alcoholic fatty liver disease|Alcoholic fatty liver
C0015732|T047|IS|72042002|SNOMEDCT_CORE|Alteration in bowel elimination: incontinence|Incontinence of feces
C0015732|T047|SY|72042002|SNOMEDCT_CORE|Bowel incontinence|Incontinence of feces
C0015732|T047|SY|72042002|SNOMEDCT_CORE|Bowels: incontinent|Incontinence of feces
C0015732|T047|PTGB|72042002|SNOMEDCT_CORE|Incontinence of faeces|Incontinence of feces
C0015732|T047|PT|72042002|SNOMEDCT_CORE|Incontinence of feces|Incontinence of feces
C0015732|T047|FN|72042002|SNOMEDCT_CORE|Incontinence of feces|Incontinence of feces
C0015732|T047|SYGB|72042002|SNOMEDCT_CORE|Incontinent of faeces|Incontinence of feces
C0015732|T047|SY|72042002|SNOMEDCT_CORE|Incontinent of feces|Incontinence of feces
C0015732|T047|SY|72042002|SNOMEDCT_CORE|Involuntary stool|Incontinence of feces
C0015734|T033|PTGB|44635007|SNOMEDCT_CORE|Faecal impaction|Fecal impaction
C0015734|T033|SYGB|44635007|SNOMEDCT_CORE|Faecal impaction of rectum|Fecal impaction
C0015734|T033|SYGB|44635007|SNOMEDCT_CORE|Faeces - impacted|Fecal impaction
C0015734|T033|PT|44635007|SNOMEDCT_CORE|Fecal impaction|Fecal impaction
C0015734|T033|FN|44635007|SNOMEDCT_CORE|Fecal impaction|Fecal impaction
C0015734|T033|SY|44635007|SNOMEDCT_CORE|Fecal impaction in rectum|Fecal impaction
C0015734|T033|SY|44635007|SNOMEDCT_CORE|Fecal impaction of rectum|Fecal impaction
C0015734|T033|SY|44635007|SNOMEDCT_CORE|Feces - impacted|Fecal impaction
C0015734|T033|SYGB|44635007|SNOMEDCT_CORE|Impacted faeces|Fecal impaction
C0015734|T033|SY|44635007|SNOMEDCT_CORE|Impacted feces|Fecal impaction
C0015734|T033|SY|44635007|SNOMEDCT_CORE|Impacted stool in rectum|Fecal impaction
C0015802|T037|PT|71620000|SNOMEDCT_CORE|Fracture of femur|Fracture of femur
C0015802|T037|FN|71620000|SNOMEDCT_CORE|Fracture of femur|Fracture of femur
C0015802|T037|IS|71620000|SNOMEDCT_CORE|Fracture of femur, NOS|Fracture of femur
C0015802|T037|SY|71620000|SNOMEDCT_CORE|Fracture of thigh|Fracture of femur
C0015802|T037|IS|71620000|SNOMEDCT_CORE|Fracture of thigh, NOS|Fracture of femur
C0015802|T037|SY|71620000|SNOMEDCT_CORE|Fracture of upper leg|Fracture of femur
C0015802|T037|IS|71620000|SNOMEDCT_CORE|Fracture of upper leg, NOS|Fracture of femur
C0015806|T037|SY|5913000|SNOMEDCT_CORE|Femoral neck fracture|Fracture of neck of femur
C0015806|T037|PT|5913000|SNOMEDCT_CORE|Fracture of neck of femur|Fracture of neck of femur
C0015806|T037|FN|5913000|SNOMEDCT_CORE|Fracture of neck of femur|Fracture of neck of femur
C0015806|T037|SY|5913000|SNOMEDCT_CORE|NOF - Fracture of neck of femur|Fracture of neck of femur
C0015927|T046|PT|276507005|SNOMEDCT_CORE|Fetal death|Fetal death
C0015927|T046|OF|276507005|SNOMEDCT_CORE|Fetal death|Fetal death
C0015927|T046|FN|276507005|SNOMEDCT_CORE|Fetal death|Fetal death
C0015927|T046|SYGB|276507005|SNOMEDCT_CORE|Foetal death|Fetal death
C0015931|T047|SY|12867002|SNOMEDCT_CORE|Abnormal foetal heart rate AND/OR rhythm affecting management of mother|Fetal distress affecting management of mother
C0015931|T047|PT|12867002|SNOMEDCT_CORE|Fetal distress affecting management of mother|Fetal distress affecting management of mother
C0015931|T047|FN|12867002|SNOMEDCT_CORE|Fetal distress affecting management of mother|Fetal distress affecting management of mother
C0015931|T047|SY|12867002|SNOMEDCT_CORE|Foetal distress affecting management of mother|Fetal distress affecting management of mother
C0015934|T047|PT|22033007|SNOMEDCT_CORE|Fetal growth restriction|Fetal growth restriction
C0015934|T047|SY|22033007|SNOMEDCT_CORE|Fetal growth retardation|Fetal growth restriction
C0015934|T047|FN|22033007|SNOMEDCT_CORE|Fetal growth retardation|Fetal growth restriction
C0015934|T047|IS|22033007|SNOMEDCT_CORE|Fetal growth retardation, NOS|Fetal growth restriction
C0015934|T047|SY|22033007|SNOMEDCT_CORE|FGR - Fetal growth retardation|Fetal growth restriction
C0015934|T047|SY|22033007|SNOMEDCT_CORE|FGR - Foetal growth retardation|Fetal growth restriction
C0015934|T047|SY|22033007|SNOMEDCT_CORE|Foetal growth retardation|Fetal growth restriction
C0015934|T047|IS|22033007|SNOMEDCT_CORE|Foetal growth retardation, NOS|Fetal growth restriction
C0015934|T047|SY|22033007|SNOMEDCT_CORE|Intrauterine growth retardation|Fetal growth restriction
C0015934|T047|IS|22033007|SNOMEDCT_CORE|Intrauterine growth retardation, NOS|Fetal growth restriction
C0015934|T047|SY|22033007|SNOMEDCT_CORE|IUGR - Intrauterine growth retardation|Fetal growth restriction
C0015934|T047|SY|22033007|SNOMEDCT_CORE|Microsomia|Fetal growth restriction
C0015934|T047|SY|22033007|SNOMEDCT_CORE|Microsomic baby|Fetal growth restriction
C0015934|T047|SY|22033007|SNOMEDCT_CORE|Poor fetal growth|Fetal growth restriction
C0015934|T047|SY|22033007|SNOMEDCT_CORE|Poor fetal growth state|Fetal growth restriction
C0015934|T047|SY|22033007|SNOMEDCT_CORE|Poor foetal growth|Fetal growth restriction
C0015934|T047|SY|22033007|SNOMEDCT_CORE|Poor foetal growth state|Fetal growth restriction
C0015944|T046|PT|44223004|SNOMEDCT_CORE|Premature rupture of membranes|Premature rupture of membranes
C0015944|T046|FN|44223004|SNOMEDCT_CORE|Premature rupture of membranes|Premature rupture of membranes
C0015944|T046|OAP|237266003|SNOMEDCT_CORE|Preterm rupture of membranes|Premature rupture of membranes
C0015944|T046|OAF|237266003|SNOMEDCT_CORE|Preterm rupture of membranes|Premature rupture of membranes
C0015944|T046|SY|44223004|SNOMEDCT_CORE|PROM - Premature rupture of membranes|Premature rupture of membranes
C0015944|T046|SY|44223004|SNOMEDCT_CORE|Rupture of amniotic sac under 24 hours before onset of labor|Premature rupture of membranes
C0015944|T046|SYGB|44223004|SNOMEDCT_CORE|Rupture of amniotic sac under 24 hours before onset of labour|Premature rupture of membranes
C0015944|T046|SY|44223004|SNOMEDCT_CORE|Rupture of membranes prior to onset of labor|Premature rupture of membranes
C0015967|T184|SY|386661006|SNOMEDCT_CORE|Febrile|Fever
C0015967|T184|PT|386661006|SNOMEDCT_CORE|Fever|Fever
C0015967|T184|FN|386661006|SNOMEDCT_CORE|Fever|Fever
C0015967|T184|SY|386661006|SNOMEDCT_CORE|Pyrexia|Fever
C0015967|T184|SY|386661006|SNOMEDCT_CORE|Pyrexial|Fever
C0015970|T184|SY|7520000|SNOMEDCT_CORE|F.U.O.|Pyrexia of unknown origin
C0015970|T184|SY|7520000|SNOMEDCT_CORE|Fever of unknown origin|Pyrexia of unknown origin
C0015970|T184|SY|7520000|SNOMEDCT_CORE|PUO - Pyrexia of unknown origin|Pyrexia of unknown origin
C0015970|T184|PT|7520000|SNOMEDCT_CORE|Pyrexia of unknown origin|Pyrexia of unknown origin
C0015970|T184|FN|7520000|SNOMEDCT_CORE|Pyrexia of unknown origin|Pyrexia of unknown origin
C0016034|T047|SY|27431007|SNOMEDCT_CORE|Diffuse cystic mastopathy|Fibrocystic disease of breast
C0016034|T047|SY|27431007|SNOMEDCT_CORE|Fibrocystic breast changes|Fibrocystic disease of breast
C0016034|T047|FN|27431007|SNOMEDCT_CORE|Fibrocystic breast changes|Fibrocystic disease of breast
C0016034|T047|SY|27431007|SNOMEDCT_CORE|Fibrocystic change of breast|Fibrocystic disease of breast
C0016034|T047|PT|27431007|SNOMEDCT_CORE|Fibrocystic disease of breast|Fibrocystic disease of breast
C0016034|T047|OF|27431007|SNOMEDCT_CORE|Fibrocystic disease of breast|Fibrocystic disease of breast
C0016034|T047|SY|27431007|SNOMEDCT_CORE|Fibrocystic mastopathy|Fibrocystic disease of breast
C0016034|T047|SY|27431007|SNOMEDCT_CORE|Gross cystic disease of breast|Fibrocystic disease of breast
C0016034|T047|SY|27431007|SNOMEDCT_CORE|Schimmelbusch's disease|Fibrocystic disease of breast
C0016045|T191|PT|424568000|SNOMEDCT_CORE|Fibroma|Fibroma
C0016045|T191|FN|424568000|SNOMEDCT_CORE|Fibroma|Fibroma
C0016052|T047|OAS|359553002|SNOMEDCT_CORE|Arterial fibromuscular dysplasia|Fibromuscular dysplasia of wall of artery
C0016052|T047|FN|783729004|SNOMEDCT_CORE|Fibromuscular dysplasia of wall of artery|Fibromuscular dysplasia of wall of artery
C0016052|T047|PT|783729004|SNOMEDCT_CORE|Fibromuscular dysplasia of wall of artery|Fibromuscular dysplasia of wall of artery
C0016052|T047|OAP|359553002|SNOMEDCT_CORE|Fibromuscular hyperplasia of artery|Fibromuscular dysplasia of wall of artery
C0016052|T047|SY|783729004|SNOMEDCT_CORE|Fibromuscular hyperplasia of artery|Fibromuscular dysplasia of wall of artery
C0016052|T047|OAF|359553002|SNOMEDCT_CORE|Fibromuscular hyperplasia of artery|Fibromuscular dysplasia of wall of artery
C0016052|T047|OAS|359553002|SNOMEDCT_CORE|FMD - Fibromuscular dysplasia|Fibromuscular dysplasia of wall of artery
C0016053|T047|IS|24693007|SNOMEDCT_CORE|Diffuse myofascial pain syndrome|Fibrositis
C0016053|T047|IS|24693007|SNOMEDCT_CORE|Fibromyalgia|Fibrositis
C0016053|T047|IS|24693007|SNOMEDCT_CORE|Fibromyalgia, NOS|Fibrositis
C0016053|T047|PT|24693007|SNOMEDCT_CORE|Fibromyositis|Fibrositis
C0016053|T047|FN|24693007|SNOMEDCT_CORE|Fibromyositis|Fibrositis
C0016053|T047|IS|24693007|SNOMEDCT_CORE|Fibromyositis, NOS|Fibrositis
C0016053|T047|IS|24693007|SNOMEDCT_CORE|Fibrositis|Fibrositis
C0016053|T047|PT|56557000|SNOMEDCT_CORE|Fibrositis|Fibrositis
C0016053|T047|FN|56557000|SNOMEDCT_CORE|Fibrositis|Fibrositis
C0016053|T047|IS|56557000|SNOMEDCT_CORE|Fibrositis, NOS|Fibrositis
C0016053|T047|IS|24693007|SNOMEDCT_CORE|MPDS - Myofacial pain dysfunction syndrome|Fibrositis
C0016053|T047|IS|24693007|SNOMEDCT_CORE|Myofacial pain dysfunction syndrome|Fibrositis
C0016053|T047|IS|24693007|SNOMEDCT_CORE|Myofascial pain dysfunction syndrome|Fibrositis
C0016053|T047|IS|24693007|SNOMEDCT_CORE|Myofascial pain syndrome|Fibrositis
C0016057|T191|SY|443250000|SNOMEDCT_CORE|Fibrosarcoma|Fibrosarcoma
C0016057|T191|PT|53654007|SNOMEDCT_CORE|Fibrosarcoma|Fibrosarcoma
C0016057|T191|FN|53654007|SNOMEDCT_CORE|Fibrosarcoma|Fibrosarcoma
C0016057|T191|IS|53654007|SNOMEDCT_CORE|Fibrosarcoma NOS|Fibrosarcoma
C0016057|T191|IS|53654007|SNOMEDCT_CORE|Fibrosarcoma, NOS|Fibrosarcoma
C0016124|T037|SY|52011008|SNOMEDCT_CORE|Finger injury|Injury of finger
C0016124|T037|PT|52011008|SNOMEDCT_CORE|Injury of finger|Injury of finger
C0016124|T037|FN|52011008|SNOMEDCT_CORE|Injury of finger|Injury of finger
C0016167|T047|PT|30037006|SNOMEDCT_CORE|Anal fissure|Anal fissure
C0016167|T047|FN|30037006|SNOMEDCT_CORE|Anal fissure|Anal fissure
C0016167|T047|SY|30037006|SNOMEDCT_CORE|Fissure in ano|Anal fissure
C0016167|T047|SY|30037006|SNOMEDCT_CORE|Nontraumatic tear of anus|Anal fissure
C0016169|T190|PT|428794004|SNOMEDCT_CORE|Fistula|Fistula
C0016169|T190|FN|428794004|SNOMEDCT_CORE|Fistula|Fistula
C0016199|T184|PT|247355005|SNOMEDCT_CORE|Flank pain|Flank pain
C0016199|T184|FN|247355005|SNOMEDCT_CORE|Flank pain|Flank pain
C0016204|T184|IS|162076009|SNOMEDCT_CORE|Flatulence|Flatulence symptom
C0016204|T184|PT|308698004|SNOMEDCT_CORE|Flatulence symptom|Flatulence symptom
C0016204|T184|OF|308698004|SNOMEDCT_CORE|Flatulence symptom|Flatulence symptom
C0016204|T184|FN|308698004|SNOMEDCT_CORE|Flatulence symptom|Flatulence symptom
C0016204|T184|SY|162076009|SNOMEDCT_CORE|Full of wind|Flatulence symptom
C0016204|T184|SY|308698004|SNOMEDCT_CORE|Wind symptom|Flatulence symptom
C0016205|T184|PT|271832001|SNOMEDCT_CORE|Flatulence, eructation and gas pain|Flatulence, eructation and gas pain
C0016205|T184|FN|271832001|SNOMEDCT_CORE|Flatulence, eructation and gas pain|Flatulence, eructation and gas pain
C0016242|T033|SY|15013002|SNOMEDCT_CORE|Musca volitans|Vitreous floaters
C0016242|T033|SY|15013002|SNOMEDCT_CORE|Muscae volitantes|Vitreous floaters
C0016242|T033|PT|15013002|SNOMEDCT_CORE|Vitreous floaters|Vitreous floaters
C0016242|T033|FN|15013002|SNOMEDCT_CORE|Vitreous floaters|Vitreous floaters
C0016382|T184|PT|238810007|SNOMEDCT_CORE|Flushing|Flushing
C0016382|T184|FN|238810007|SNOMEDCT_CORE|Flushing|Flushing
C0016429|T047|SY|2615004|SNOMEDCT_CORE|Cyst of graafian follicle|Follicular cyst of ovary
C0016429|T047|PT|2615004|SNOMEDCT_CORE|Follicular cyst of ovary|Follicular cyst of ovary
C0016429|T047|FN|2615004|SNOMEDCT_CORE|Follicular cyst of ovary|Follicular cyst of ovary
C0016429|T047|SY|2615004|SNOMEDCT_CORE|Follicular cystic ovary disease|Follicular cyst of ovary
C0016429|T047|SY|2615004|SNOMEDCT_CORE|Graafian follicle cyst|Follicular cyst of ovary
C0016436|T047|PT|13600006|SNOMEDCT_CORE|Folliculitis|Folliculitis
C0016436|T047|FN|13600006|SNOMEDCT_CORE|Folliculitis|Folliculitis
C0016470|T046|PT|414285001|SNOMEDCT_CORE|Allergy to food|Allergy to food
C0016470|T046|FN|414285001|SNOMEDCT_CORE|Allergy to food|Allergy to food
C0016470|T046|SY|414285001|SNOMEDCT_CORE|Food allergy|Allergy to food
C0016470|T046|OF|414285001|SNOMEDCT_CORE|Food allergy|Allergy to food
C0016479|T037|PT|75258004|SNOMEDCT_CORE|Food poisoning|Food poisoning
C0016479|T037|FN|75258004|SNOMEDCT_CORE|Food poisoning|Food poisoning
C0016479|T037|IS|75258004|SNOMEDCT_CORE|Food poisoning, NOS|Food poisoning
C0016479|T037|SY|75258004|SNOMEDCT_CORE|FP - Food poisoning|Food poisoning
C0016506|T190|PT|229844004|SNOMEDCT_CORE|Deformity of foot|Deformity of foot
C0016506|T190|FN|229844004|SNOMEDCT_CORE|Deformity of foot|Deformity of foot
C0016507|T020|SY|240244006|SNOMEDCT_CORE|Acquired deformity of the foot|Acquired deformity of the foot
C0016508|T019|PT|302297009|SNOMEDCT_CORE|Congenital deformity of foot|Congenital deformity of foot
C0016508|T019|FN|302297009|SNOMEDCT_CORE|Congenital deformity of foot|Congenital deformity of foot
C0016512|T184|PT|47933007|SNOMEDCT_CORE|Foot pain|Foot pain
C0016512|T184|FN|47933007|SNOMEDCT_CORE|Foot pain|Foot pain
C0016512|T184|IS|47933007|SNOMEDCT_CORE|Podalgia|Foot pain
C0016522|T019|PT|204317008|SNOMEDCT_CORE|Patent foramen ovale|Patent foramen ovale
C0016522|T019|FN|204317008|SNOMEDCT_CORE|Patent foramen ovale|Patent foramen ovale
C0016522|T019|SY|204317008|SNOMEDCT_CORE|PFO - Patent foramen ovale|Patent foramen ovale
C0016537|T037|SY|125597008|SNOMEDCT_CORE|Forearm injury|Injury of forearm
C0016537|T037|PT|125597008|SNOMEDCT_CORE|Injury of forearm|Injury of forearm
C0016537|T037|FN|125597008|SNOMEDCT_CORE|Injury of forearm|Injury of forearm
C0016542|T037|SY|125670008|SNOMEDCT_CORE|Disorder due to presence of foreign body|Foreign body
C0016542|T037|SY|125670008|SNOMEDCT_CORE|FB - Foreign body of body structure|Foreign body
C0016542|T037|PT|125670008|SNOMEDCT_CORE|Foreign body|Foreign body
C0016542|T037|FN|125670008|SNOMEDCT_CORE|Foreign body|Foreign body
C0016542|T037|SY|125670008|SNOMEDCT_CORE|Foreign body of body structure|Foreign body
C0016546|T037|SY|33334006|SNOMEDCT_CORE|Foreign body in alimentary tract|Foreign body in digestive tract
C0016546|T037|IS|33334006|SNOMEDCT_CORE|Foreign body in alimentary tract, NOS|Foreign body in digestive tract
C0016546|T037|IS|33334006|SNOMEDCT_CORE|Foreign body in digestive system, NOS|Foreign body in digestive tract
C0016546|T037|PT|33334006|SNOMEDCT_CORE|Foreign body in digestive tract|Foreign body in digestive tract
C0016546|T037|FN|33334006|SNOMEDCT_CORE|Foreign body in digestive tract|Foreign body in digestive tract
C0016546|T037|SY|33334006|SNOMEDCT_CORE|Foreign body of digestive structure|Foreign body in digestive tract
C0016547|T037|SY|93458008|SNOMEDCT_CORE|FB - Foreign body in skin|Foreign body in skin
C0016547|T037|PT|93458008|SNOMEDCT_CORE|Foreign body in skin|Foreign body in skin
C0016547|T037|FN|93458008|SNOMEDCT_CORE|Foreign body in skin|Foreign body in skin
C0016547|T037|IS|93458008|SNOMEDCT_CORE|Foreign body in skin, NOS|Foreign body in skin
C0016658|T037|SY|125605004|SNOMEDCT_CORE|Broken bone|Fracture of bone
C0016658|T037|SY|125605004|SNOMEDCT_CORE|Fracture|Fracture of bone
C0016658|T037|PT|125605004|SNOMEDCT_CORE|Fracture of bone|Fracture of bone
C0016658|T037|FN|125605004|SNOMEDCT_CORE|Fracture of bone|Fracture of bone
C0016659|T037|PT|423125000|SNOMEDCT_CORE|Closed fracture|Closed fracture
C0016659|T037|SY|423125000|SNOMEDCT_CORE|Closed fracture of bone|Closed fracture
C0016659|T037|FN|423125000|SNOMEDCT_CORE|Closed fracture of bone|Closed fracture
C0016664|T037|SY|23382007|SNOMEDCT_CORE|Fatigue fracture|Stress fracture
C0016664|T037|PT|240197007|SNOMEDCT_CORE|Stress fracture|Stress fracture
C0016664|T037|OF|240197007|SNOMEDCT_CORE|Stress fracture|Stress fracture
C0016664|T037|PT|23382007|SNOMEDCT_CORE|Stress fracture|Stress fracture
C0016664|T037|IS|23382007|SNOMEDCT_CORE|Stress fracture|Stress fracture
C0016664|T037|FN|23382007|SNOMEDCT_CORE|Stress fracture|Stress fracture
C0016664|T037|FN|240197007|SNOMEDCT_CORE|Stress fracture|Stress fracture
C0016665|T046|PT|302941001|SNOMEDCT_CORE|Nonunion of fracture|Nonunion of fracture
C0016665|T046|FN|302941001|SNOMEDCT_CORE|Nonunion of fracture|Nonunion of fracture
C0016735|T047|PT|78737005|SNOMEDCT_CORE|Frontal sinusitis|Frontal sinusitis
C0016735|T047|FN|78737005|SNOMEDCT_CORE|Frontal sinusitis|Frontal sinusitis
C0016735|T047|IS|78737005|SNOMEDCT_CORE|Frontal sinusitis, NOS|Frontal sinusitis
C0016781|T047|SY|193839007|SNOMEDCT_CORE|Fuch's endothelial corneal dystrophy|Fuchs' corneal dystrophy
C0016781|T047|SY|193839007|SNOMEDCT_CORE|Fuchs corneal dystrophy|Fuchs' corneal dystrophy
C0016781|T047|PT|193839007|SNOMEDCT_CORE|Fuchs' corneal dystrophy|Fuchs' corneal dystrophy
C0016781|T047|FN|193839007|SNOMEDCT_CORE|Fuchs' corneal dystrophy|Fuchs' corneal dystrophy
C0016781|T047|SY|193839007|SNOMEDCT_CORE|Fuchs' endothelial dystrophy|Fuchs' corneal dystrophy
C0016782|T047|SY|11226001|SNOMEDCT_CORE|Fuchs uveitis syndrome|Fuchs' heterochromic cyclitis
C0016782|T047|PT|11226001|SNOMEDCT_CORE|Fuchs' heterochromic cyclitis|Fuchs' heterochromic cyclitis
C0016782|T047|FN|11226001|SNOMEDCT_CORE|Fuchs' heterochromic cyclitis|Fuchs' heterochromic cyclitis
C0016782|T047|SY|11226001|SNOMEDCT_CORE|Fuchs' heterochromic iridocyclitis|Fuchs' heterochromic cyclitis
C0016782|T047|SY|11226001|SNOMEDCT_CORE|Fuchs' heterochromic uveitis|Fuchs' heterochromic cyclitis
C0016807|T047|PT|81120009|SNOMEDCT_CORE|Functional disorder of intestine|Functional disorder of intestine
C0016807|T047|FN|81120009|SNOMEDCT_CORE|Functional disorder of intestine|Functional disorder of intestine
C0016807|T047|IS|81120009|SNOMEDCT_CORE|Functional disorder of intestine, NOS|Functional disorder of intestine
C0016842|T019|SY|391982004|SNOMEDCT_CORE|Congenital funnel chest|Congenital pectus excavatum
C0016842|T019|PT|391982004|SNOMEDCT_CORE|Congenital pectus excavatum|Congenital pectus excavatum
C0016842|T019|FN|391982004|SNOMEDCT_CORE|Congenital pectus excavatum|Congenital pectus excavatum
C0016842|T019|IS|391982004|SNOMEDCT_CORE|Funnel chest|Congenital pectus excavatum
C0016842|T019|IS|391982004|SNOMEDCT_CORE|Pectus recurvatum|Congenital pectus excavatum
C0016842|T019|IS|391982004|SNOMEDCT_CORE|Trichterbrust|Congenital pectus excavatum
C0016977|T047|OF|39621005|SNOMEDCT_CORE|Disease of gallbladder|Disorder of gallbladder
C0016977|T047|IS|39621005|SNOMEDCT_CORE|Disease of gallbladder|Disorder of gallbladder
C0016977|T047|IS|39621005|SNOMEDCT_CORE|Disease of gallbladder, NOS|Disorder of gallbladder
C0016977|T047|PT|39621005|SNOMEDCT_CORE|Disorder of gallbladder|Disorder of gallbladder
C0016977|T047|FN|39621005|SNOMEDCT_CORE|Disorder of gallbladder|Disorder of gallbladder
C0016977|T047|SY|39621005|SNOMEDCT_CORE|Gallbladder disease|Disorder of gallbladder
C0016977|T047|SY|39621005|SNOMEDCT_CORE|Gallbladder disorder|Disorder of gallbladder
C0016977|T047|IS|39621005|SNOMEDCT_CORE|Gallbladder disorder, NOS|Disorder of gallbladder
C0017086|T047|SY|372070002|SNOMEDCT_CORE|Gangrene|Gangrenous disorder
C0017086|T047|FN|372070002|SNOMEDCT_CORE|Gangrenous disorder|Gangrenous disorder
C0017086|T047|PT|372070002|SNOMEDCT_CORE|Gangrenous disorder|Gangrenous disorder
C0017145|T047|PT|91109007|SNOMEDCT_CORE|Gastric varices|Gastric varices
C0017145|T047|FN|91109007|SNOMEDCT_CORE|Gastric varices|Gastric varices
C0017145|T047|SY|91109007|SNOMEDCT_CORE|Gastric varix|Gastric varices
C0017152|T047|SY|4556007|SNOMEDCT_CORE|Gastric catarrh|Gastritis
C0017152|T047|PT|4556007|SNOMEDCT_CORE|Gastritis|Gastritis
C0017152|T047|FN|4556007|SNOMEDCT_CORE|Gastritis|Gastritis
C0017152|T047|IS|4556007|SNOMEDCT_CORE|Gastritis, NOS|Gastritis
C0017154|T047|SY|84568007|SNOMEDCT_CORE|AG - Atrophic gastritis|Atrophic gastritis
C0017154|T047|PT|84568007|SNOMEDCT_CORE|Atrophic gastritis|Atrophic gastritis
C0017154|T047|FN|84568007|SNOMEDCT_CORE|Atrophic gastritis|Atrophic gastritis
C0017154|T047|SY|84568007|SNOMEDCT_CORE|CAG - Chronic atrophic gastritis|Atrophic gastritis
C0017154|T047|SY|84568007|SNOMEDCT_CORE|Chronic atrophic gastritis|Atrophic gastritis
C0017154|T047|SY|84568007|SNOMEDCT_CORE|Gastric atrophy|Atrophic gastritis
C0017160|T047|PT|25374005|SNOMEDCT_CORE|Gastroenteritis|Gastroenteritis
C0017160|T047|FN|25374005|SNOMEDCT_CORE|Gastroenteritis|Gastroenteritis
C0017160|T047|IS|25374005|SNOMEDCT_CORE|Gastroenteritis, NOS|Gastroenteritis
C0017160|T047|SY|25374005|SNOMEDCT_CORE|GE - Gastroenteritis|Gastroenteritis
C0017168|T047|IS|235595009|SNOMEDCT_CORE|Acid reflux|Gastroesophageal reflux disease
C0017168|T047|IS|235595009|SNOMEDCT_CORE|Esophageal reflux|Gastroesophageal reflux disease
C0017168|T047|IS|235595009|SNOMEDCT_CORE|Gastresophageal reflux disease|Gastroesophageal reflux disease
C0017168|T047|SY|235595009|SNOMEDCT_CORE|Gastro-esophageal reflux|Gastroesophageal reflux disease
C0017168|T047|SY|235595009|SNOMEDCT_CORE|Gastro-esophageal reflux disease|Gastroesophageal reflux disease
C0017168|T047|SYGB|235595009|SNOMEDCT_CORE|Gastro-oesophageal reflux|Gastroesophageal reflux disease
C0017168|T047|SYGB|235595009|SNOMEDCT_CORE|Gastro-oesophageal reflux disease|Gastroesophageal reflux disease
C0017168|T047|PT|235595009|SNOMEDCT_CORE|Gastroesophageal reflux disease|Gastroesophageal reflux disease
C0017168|T047|FN|235595009|SNOMEDCT_CORE|Gastroesophageal reflux disease|Gastroesophageal reflux disease
C0017168|T047|PTGB|235595009|SNOMEDCT_CORE|Gastrooesophageal reflux disease|Gastroesophageal reflux disease
C0017168|T047|SY|235595009|SNOMEDCT_CORE|GERD - Gastro-esophageal reflux disease|Gastroesophageal reflux disease
C0017168|T047|SY|235595009|SNOMEDCT_CORE|GOR - Gastro-esophageal reflux|Gastroesophageal reflux disease
C0017168|T047|SYGB|235595009|SNOMEDCT_CORE|GOR - Gastro-oesophageal reflux|Gastroesophageal reflux disease
C0017168|T047|SY|235595009|SNOMEDCT_CORE|GORD - Gastro-esophageal reflux disease|Gastroesophageal reflux disease
C0017168|T047|SYGB|235595009|SNOMEDCT_CORE|GORD - Gastro-oesophageal reflux disease|Gastroesophageal reflux disease
C0017168|T047|IS|235595009|SNOMEDCT_CORE|Oesophageal reflux|Gastroesophageal reflux disease
C0017178|T047|SY|25374005|SNOMEDCT_CORE|Gastroenteropathy|Gastroenteropathy
C0017181|T046|SY|74474003|SNOMEDCT_CORE|Gastrointestinal bleed|Gastrointestinal hemorrhage
C0017181|T046|SY|74474003|SNOMEDCT_CORE|Gastrointestinal bleeding|Gastrointestinal hemorrhage
C0017181|T046|IS|74474003|SNOMEDCT_CORE|Gastrointestinal bleeding, NOS|Gastrointestinal hemorrhage
C0017181|T046|PTGB|74474003|SNOMEDCT_CORE|Gastrointestinal haemorrhage|Gastrointestinal hemorrhage
C0017181|T046|PT|74474003|SNOMEDCT_CORE|Gastrointestinal hemorrhage|Gastrointestinal hemorrhage
C0017181|T046|FN|74474003|SNOMEDCT_CORE|Gastrointestinal hemorrhage|Gastrointestinal hemorrhage
C0017181|T046|IS|74474003|SNOMEDCT_CORE|Gastrointestinal hemorrhage, NOS|Gastrointestinal hemorrhage
C0017181|T046|SY|74474003|SNOMEDCT_CORE|GI - Gastrointestinal bleed|Gastrointestinal hemorrhage
C0017181|T046|SYGB|74474003|SNOMEDCT_CORE|GI - Gastrointestinal haemorrhage|Gastrointestinal hemorrhage
C0017181|T046|SY|74474003|SNOMEDCT_CORE|GI - Gastrointestinal hemorrhage|Gastrointestinal hemorrhage
C0017181|T046|SY|74474003|SNOMEDCT_CORE|GI bleeding|Gastrointestinal hemorrhage
C0017181|T046|IS|74474003|SNOMEDCT_CORE|GI bleeding, NOS|Gastrointestinal hemorrhage
C0017181|T046|SYGB|74474003|SNOMEDCT_CORE|GI haemorrhage|Gastrointestinal hemorrhage
C0017181|T046|SY|74474003|SNOMEDCT_CORE|GI hemorrhage|Gastrointestinal hemorrhage
C0017181|T046|IS|74474003|SNOMEDCT_CORE|GI hemorrhage, NOS|Gastrointestinal hemorrhage
C0017181|T046|SYGB|74474003|SNOMEDCT_CORE|GIH - Gastrointestinal haemorrhage|Gastrointestinal hemorrhage
C0017181|T046|SY|74474003|SNOMEDCT_CORE|GIH - Gastrointestinal hemorrhage|Gastrointestinal hemorrhage
C0017181|T046|SYGB|74474003|SNOMEDCT_CORE|GIT - Gastrointestinal tract haemorrhage|Gastrointestinal hemorrhage
C0017181|T046|SY|74474003|SNOMEDCT_CORE|GIT - Gastrointestinal tract hemorrhage|Gastrointestinal hemorrhage
C0017327|T047|PTGB|39823006|SNOMEDCT_CORE|Generalised atherosclerosis|Generalized atherosclerosis
C0017327|T047|IS|39823006|SNOMEDCT_CORE|Generalized and unspecified atherosclerosis|Generalized atherosclerosis
C0017327|T047|PT|39823006|SNOMEDCT_CORE|Generalized atherosclerosis|Generalized atherosclerosis
C0017327|T047|FN|39823006|SNOMEDCT_CORE|Generalized atherosclerosis|Generalized atherosclerosis
C0017332|T047|PTGB|192979009|SNOMEDCT_CORE|Generalised non-convulsive epilepsy|Generalized non-convulsive epilepsy
C0017332|T047|SYGB|192979009|SNOMEDCT_CORE|Generalised nonconvulsive epilepsy|Generalized non-convulsive epilepsy
C0017332|T047|PT|192979009|SNOMEDCT_CORE|Generalized non-convulsive epilepsy|Generalized non-convulsive epilepsy
C0017332|T047|FN|192979009|SNOMEDCT_CORE|Generalized non-convulsive epilepsy|Generalized non-convulsive epilepsy
C0017332|T047|SY|192979009|SNOMEDCT_CORE|Generalized nonconvulsive epilepsy|Generalized non-convulsive epilepsy
C0017525|T191|PT|443790001|SNOMEDCT_CORE|Giant cell tumor|Giant cell tumor
C0017525|T191|PT|115238001|SNOMEDCT_CORE|Giant cell tumor|Giant cell tumor
C0017525|T191|FN|115238001|SNOMEDCT_CORE|Giant cell tumor|Giant cell tumor
C0017525|T191|FN|443790001|SNOMEDCT_CORE|Giant cell tumor|Giant cell tumor
C0017525|T191|PTGB|443790001|SNOMEDCT_CORE|Giant cell tumour|Giant cell tumor
C0017525|T191|PTGB|115238001|SNOMEDCT_CORE|Giant cell tumour|Giant cell tumor
C0017551|T047|SYGB|27503000|SNOMEDCT_CORE|Benign unconjugated bilirubinaemia syndrome|Gilbert's syndrome
C0017551|T047|SY|27503000|SNOMEDCT_CORE|Benign unconjugated bilirubinemia syndrome|Gilbert's syndrome
C0017551|T047|SYGB|27503000|SNOMEDCT_CORE|Cholaemia familiaris simplex|Gilbert's syndrome
C0017551|T047|SY|27503000|SNOMEDCT_CORE|Cholemia familiaris simplex|Gilbert's syndrome
C0017551|T047|SY|27503000|SNOMEDCT_CORE|Chronic intermittent juvenile jaundice|Gilbert's syndrome
C0017551|T047|SYGB|27503000|SNOMEDCT_CORE|Congenital familial cholaemia|Gilbert's syndrome
C0017551|T047|SY|27503000|SNOMEDCT_CORE|Congenital familial cholemia|Gilbert's syndrome
C0017551|T047|SY|27503000|SNOMEDCT_CORE|Constitutional hepatic dysfunction|Gilbert's syndrome
C0017551|T047|SYGB|27503000|SNOMEDCT_CORE|Familial nonhaemolytic bilirubinaemia|Gilbert's syndrome
C0017551|T047|SYGB|27503000|SNOMEDCT_CORE|Familial nonhaemolytic jaundice|Gilbert's syndrome
C0017551|T047|SY|27503000|SNOMEDCT_CORE|Familial nonhemolytic bilirubinemia|Gilbert's syndrome
C0017551|T047|SY|27503000|SNOMEDCT_CORE|Familial nonhemolytic jaundice|Gilbert's syndrome
C0017551|T047|SY|27503000|SNOMEDCT_CORE|Gilbert syndrome|Gilbert's syndrome
C0017551|T047|SY|27503000|SNOMEDCT_CORE|Gilbert-Lereboullet syndrome|Gilbert's syndrome
C0017551|T047|SY|27503000|SNOMEDCT_CORE|Gilbert's disease|Gilbert's syndrome
C0017551|T047|PT|27503000|SNOMEDCT_CORE|Gilbert's syndrome|Gilbert's syndrome
C0017551|T047|FN|27503000|SNOMEDCT_CORE|Gilbert's syndrome|Gilbert's syndrome
C0017551|T047|SY|27503000|SNOMEDCT_CORE|Gilberts syndrome|Gilbert's syndrome
C0017551|T047|SYGB|27503000|SNOMEDCT_CORE|Hereditary nonhaemolytic jaundice|Gilbert's syndrome
C0017551|T047|SY|27503000|SNOMEDCT_CORE|Hereditary nonhemolytic jaundice|Gilbert's syndrome
C0017551|T047|SYGB|27503000|SNOMEDCT_CORE|Low-grade chronic hyperbilirubinaemia syndrome|Gilbert's syndrome
C0017551|T047|SY|27503000|SNOMEDCT_CORE|Low-grade chronic hyperbilirubinemia syndrome|Gilbert's syndrome
C0017551|T047|SY|27503000|SNOMEDCT_CORE|Meulengracht syndrome|Gilbert's syndrome
C0017565|T046|PT|86276007|SNOMEDCT_CORE|Bleeding gums|Bleeding gums
C0017565|T046|FN|86276007|SNOMEDCT_CORE|Bleeding gums|Bleeding gums
C0017565|T046|SY|86276007|SNOMEDCT_CORE|Gingival bleeding|Bleeding gums
C0017565|T046|SYGB|86276007|SNOMEDCT_CORE|Gingival haemorrhage|Bleeding gums
C0017565|T046|SY|86276007|SNOMEDCT_CORE|Gingival hemorrhage|Bleeding gums
C0017574|T047|PT|66383009|SNOMEDCT_CORE|Gingivitis|Gingivitis
C0017574|T047|FN|66383009|SNOMEDCT_CORE|Gingivitis|Gingivitis
C0017574|T047|IS|66383009|SNOMEDCT_CORE|Gingivitis, NOS|Gingivitis
C0017601|T047|PT|23986001|SNOMEDCT_CORE|Glaucoma|Glaucoma
C0017601|T047|FN|23986001|SNOMEDCT_CORE|Glaucoma|Glaucoma
C0017601|T047|IS|23986001|SNOMEDCT_CORE|Glaucoma, NOS|Glaucoma
C0017605|T047|SY|392291006|SNOMEDCT_CORE|ACG - Angle closure glaucoma|Angle-closure glaucoma
C0017605|T047|IS|33647009|SNOMEDCT_CORE|Angle-closure glaucoma|Angle-closure glaucoma
C0017605|T047|PT|392291006|SNOMEDCT_CORE|Angle-closure glaucoma|Angle-closure glaucoma
C0017605|T047|FN|392291006|SNOMEDCT_CORE|Angle-closure glaucoma|Angle-closure glaucoma
C0017605|T047|SY|392291006|SNOMEDCT_CORE|Narrow angle glaucoma|Angle-closure glaucoma
C0017605|T047|SY|33647009|SNOMEDCT_CORE|Narrow cleft glaucoma|Angle-closure glaucoma
C0017605|T047|SY|392291006|SNOMEDCT_CORE|Narrow-angle glaucoma|Angle-closure glaucoma
C0017606|T047|PT|392288006|SNOMEDCT_CORE|Primary angle-closure glaucoma|Primary angle-closure glaucoma
C0017606|T047|FN|392288006|SNOMEDCT_CORE|Primary angle-closure glaucoma|Primary angle-closure glaucoma
C0017609|T047|PT|232086000|SNOMEDCT_CORE|Neovascular glaucoma|Neovascular glaucoma
C0017609|T047|FN|232086000|SNOMEDCT_CORE|Neovascular glaucoma|Neovascular glaucoma
C0017609|T047|SY|232086000|SNOMEDCT_CORE|Rubeotic glaucoma|Neovascular glaucoma
C0017609|T047|SY|232086000|SNOMEDCT_CORE|Secondary angle closure glaucoma with rubeosis|Neovascular glaucoma
C0017612|T047|SY|84494001|SNOMEDCT_CORE|OAG - Open-angle glaucoma|Open-angle glaucoma
C0017612|T047|SY|84494001|SNOMEDCT_CORE|Open angle glaucoma|Open-angle glaucoma
C0017612|T047|SY|84494001|SNOMEDCT_CORE|Open cleft glaucoma|Open-angle glaucoma
C0017612|T047|PT|84494001|SNOMEDCT_CORE|Open-angle glaucoma|Open-angle glaucoma
C0017612|T047|FN|84494001|SNOMEDCT_CORE|Open-angle glaucoma|Open-angle glaucoma
C0017612|T047|IS|84494001|SNOMEDCT_CORE|Open-angle glaucoma, NOS|Open-angle glaucoma
C0017612|T047|SY|84494001|SNOMEDCT_CORE|Wide-angle glaucoma|Open-angle glaucoma
C0017612|T047|IS|84494001|SNOMEDCT_CORE|Wide-angle glaucoma, NOS|Open-angle glaucoma
C0017614|T047|PT|232079008|SNOMEDCT_CORE|Glaucoma suspect|Glaucoma suspect
C0017614|T047|OF|232079008|SNOMEDCT_CORE|Glaucoma suspect|Glaucoma suspect
C0017614|T047|FN|232079008|SNOMEDCT_CORE|Glaucoma suspect|Glaucoma suspect
C0017636|T191|PT|63634009|SNOMEDCT_CORE|Glioblastoma|Glioblastoma
C0017636|T191|OF|63634009|SNOMEDCT_CORE|Glioblastoma|Glioblastoma
C0017636|T191|SY|63634009|SNOMEDCT_CORE|Glioblastoma, no ICD-O subtype|Glioblastoma
C0017636|T191|OF|63634009|SNOMEDCT_CORE|Glioblastoma, no ICD-O subtype|Glioblastoma
C0017636|T191|SY|63634009|SNOMEDCT_CORE|Glioblastoma, no International Classification of Diseases for Oncology subtype|Glioblastoma
C0017636|T191|FN|63634009|SNOMEDCT_CORE|Glioblastoma, no International Classification of Diseases for Oncology subtype|Glioblastoma
C0017636|T191|IS|63634009|SNOMEDCT_CORE|Glioblastoma, NOS|Glioblastoma
C0017650|T184|PT|267103008|SNOMEDCT_CORE|Feeling of lump in throat|Feeling of lump in throat
C0017650|T184|FN|267103008|SNOMEDCT_CORE|Feeling of lump in throat|Feeling of lump in throat
C0017650|T184|OAP|44037003|SNOMEDCT_CORE|Globus hystericus|Feeling of lump in throat
C0017650|T184|SY|267103008|SNOMEDCT_CORE|Globus hystericus|Feeling of lump in throat
C0017650|T184|OAF|44037003|SNOMEDCT_CORE|Globus hystericus|Feeling of lump in throat
C0017650|T184|OAS|44037003|SNOMEDCT_CORE|Globus pharyngeus|Feeling of lump in throat
C0017650|T184|SY|267103008|SNOMEDCT_CORE|Globus pharyngeus|Feeling of lump in throat
C0017650|T184|OAP|88889000|SNOMEDCT_CORE|Globus sensation|Feeling of lump in throat
C0017650|T184|SY|267103008|SNOMEDCT_CORE|Globus sensation|Feeling of lump in throat
C0017650|T184|OAF|88889000|SNOMEDCT_CORE|Globus sensation|Feeling of lump in throat
C0017650|T184|OAS|44037003|SNOMEDCT_CORE|Globus syndrome|Feeling of lump in throat
C0017650|T184|OAS|44037003|SNOMEDCT_CORE|Idiopathic globus|Feeling of lump in throat
C0017658|T047|PT|36171008|SNOMEDCT_CORE|Glomerulonephritis|Glomerulonephritis
C0017658|T047|FN|36171008|SNOMEDCT_CORE|Glomerulonephritis|Glomerulonephritis
C0017658|T047|IS|36171008|SNOMEDCT_CORE|Glomerulonephritis, NOS|Glomerulonephritis
C0017658|T047|SY|36171008|SNOMEDCT_CORE|GN - Glomerulonephritis|Glomerulonephritis
C0017661|T047|SY|236407003|SNOMEDCT_CORE|IgA glomerulonephritis|IgA nephropathy
C0017661|T047|PT|236407003|SNOMEDCT_CORE|IgA nephropathy|IgA nephropathy
C0017661|T047|OF|236407003|SNOMEDCT_CORE|IgA nephropathy|IgA nephropathy
C0017661|T047|SY|236407003|SNOMEDCT_CORE|IgAN - IgA nephropathy|IgA nephropathy
C0017661|T047|FN|236407003|SNOMEDCT_CORE|Immunoglobulin A nephropathy|IgA nephropathy
C0017661|T047|SY|236407003|SNOMEDCT_CORE|Immunoglobulin A nephropathy|IgA nephropathy
C0017662|T047|SY|80321008|SNOMEDCT_CORE|Lobular glomerulonephritis|Mesangiocapillary glomerulonephritis
C0017662|T047|SY|80321008|SNOMEDCT_CORE|MCGN - Mesangiocapillary glomerulonephritis|Mesangiocapillary glomerulonephritis
C0017662|T047|SY|80321008|SNOMEDCT_CORE|Membranoproliferative glomerulonephritis|Mesangiocapillary glomerulonephritis
C0017662|T047|PT|80321008|SNOMEDCT_CORE|Mesangiocapillary glomerulonephritis|Mesangiocapillary glomerulonephritis
C0017662|T047|FN|80321008|SNOMEDCT_CORE|Mesangiocapillary glomerulonephritis|Mesangiocapillary glomerulonephritis
C0017662|T047|IS|80321008|SNOMEDCT_CORE|Mesangiocapillary glomerulonephritis, NOS|Mesangiocapillary glomerulonephritis
C0017662|T047|SY|80321008|SNOMEDCT_CORE|MPGN - Membranoproliferative glomerulonephritis|Mesangiocapillary glomerulonephritis
C0017665|T047|SY|77182004|SNOMEDCT_CORE|Chronic nephritic syndrome, diffuse membranous glomerulonephritis|Membranous glomerulonephritis
C0017665|T047|IS|77182004|SNOMEDCT_CORE|Chronic nephritic syndrome, diffuse membranous glomerulonephritis|Membranous glomerulonephritis
C0017665|T047|PT|77182004|SNOMEDCT_CORE|Membranous glomerulonephritis|Membranous glomerulonephritis
C0017665|T047|FN|77182004|SNOMEDCT_CORE|Membranous glomerulonephritis|Membranous glomerulonephritis
C0017665|T047|SY|77182004|SNOMEDCT_CORE|MGN - Membranous glomerulonephritis|Membranous glomerulonephritis
C0017668|T047|SY|25821008|SNOMEDCT_CORE|FGS - Focal glomerulosclerosis|Focal glomerular sclerosis
C0017668|T047|PT|25821008|SNOMEDCT_CORE|Focal glomerular sclerosis|Focal glomerular sclerosis
C0017668|T047|FN|25821008|SNOMEDCT_CORE|Focal glomerular sclerosis|Focal glomerular sclerosis
C0017668|T047|SY|25821008|SNOMEDCT_CORE|Focal glomerulosclerosis|Focal glomerular sclerosis
C0017672|T184|SY|30731004|SNOMEDCT_CORE|Glossalgia|Glossodynia
C0017672|T184|IS|399044006|SNOMEDCT_CORE|Glossodynia|Glossodynia
C0017672|T184|PT|30731004|SNOMEDCT_CORE|Glossodynia|Glossodynia
C0017672|T184|FN|30731004|SNOMEDCT_CORE|Glossodynia|Glossodynia
C0017672|T184|IS|399044006|SNOMEDCT_CORE|Painful tongue|Glossodynia
C0017672|T184|SY|30731004|SNOMEDCT_CORE|Painful tongue|Glossodynia
C0017672|T184|SY|30731004|SNOMEDCT_CORE|Soreness of tongue|Glossodynia
C0017675|T047|PT|45534005|SNOMEDCT_CORE|Glossitis|Glossitis
C0017675|T047|FN|45534005|SNOMEDCT_CORE|Glossitis|Glossitis
C0017675|T047|IS|45534005|SNOMEDCT_CORE|Glossitis, NOS|Glossitis
C0017675|T047|SY|45534005|SNOMEDCT_CORE|Inflammation of tongue|Glossitis
C0017979|T033|SY|45154002|SNOMEDCT_CORE|Glucosuria|Glycosuria
C0017979|T033|PT|45154002|SNOMEDCT_CORE|Glycosuria|Glycosuria
C0017979|T033|FN|45154002|SNOMEDCT_CORE|Glycosuria|Glycosuria
C0018021|T047|SY|3716002|SNOMEDCT_CORE|Enlargement of thyroid|Goiter
C0018021|T047|PT|3716002|SNOMEDCT_CORE|Goiter|Goiter
C0018021|T047|FN|3716002|SNOMEDCT_CORE|Goiter|Goiter
C0018021|T047|IS|3716002|SNOMEDCT_CORE|Goiter, NOS|Goiter
C0018021|T047|PTGB|3716002|SNOMEDCT_CORE|Goitre|Goiter
C0018021|T047|IS|3716002|SNOMEDCT_CORE|Goitre, NOS|Goiter
C0018021|T047|SY|3716002|SNOMEDCT_CORE|Struma - goiter|Goiter
C0018021|T047|SYGB|3716002|SNOMEDCT_CORE|Struma - goitre|Goiter
C0018021|T047|SY|3716002|SNOMEDCT_CORE|Struma of thyroid|Goiter
C0018021|T047|SY|3716002|SNOMEDCT_CORE|Swelling of thyroid gland|Goiter
C0018021|T047|SY|3716002|SNOMEDCT_CORE|Thyroid enlargement|Goiter
C0018021|T047|SY|3716002|SNOMEDCT_CORE|Thyroid goiter|Goiter
C0018021|T047|SYGB|3716002|SNOMEDCT_CORE|Thyroid goitre|Goiter
C0018022|T047|PT|56805008|SNOMEDCT_CORE|Endemic goiter|Endemic goiter
C0018022|T047|FN|56805008|SNOMEDCT_CORE|Endemic goiter|Endemic goiter
C0018022|T047|PTGB|56805008|SNOMEDCT_CORE|Endemic goitre|Endemic goiter
C0018022|T047|IS|56805008|SNOMEDCT_CORE|Simple goiter|Endemic goiter
C0018022|T047|PT|267369002|SNOMEDCT_CORE|Simple goiter|Endemic goiter
C0018022|T047|FN|267369002|SNOMEDCT_CORE|Simple goiter|Endemic goiter
C0018022|T047|IS|56805008|SNOMEDCT_CORE|Simple goitre|Endemic goiter
C0018022|T047|PTGB|267369002|SNOMEDCT_CORE|Simple goitre|Endemic goiter
C0018022|T047|SY|56805008|SNOMEDCT_CORE|Simple iodine deficiency goiter|Endemic goiter
C0018022|T047|SYGB|56805008|SNOMEDCT_CORE|Simple iodine deficiency goitre|Endemic goiter
C0018023|T047|IS|237570007|SNOMEDCT_CORE|Nodular goiter|Nodular goiter
C0018023|T047|IS|190236006|SNOMEDCT_CORE|Nodular goiter|Nodular goiter
C0018023|T047|PT|419153005|SNOMEDCT_CORE|Nodular goiter|Nodular goiter
C0018023|T047|FN|419153005|SNOMEDCT_CORE|Nodular goiter|Nodular goiter
C0018023|T047|IS|237570007|SNOMEDCT_CORE|Nodular goitre|Nodular goiter
C0018023|T047|IS|190236006|SNOMEDCT_CORE|Nodular goitre|Nodular goiter
C0018023|T047|PTGB|419153005|SNOMEDCT_CORE|Nodular goitre|Nodular goiter
C0018023|T047|SY|419153005|SNOMEDCT_CORE|Nodular hyperplasia of thyroid|Nodular goiter
C0018051|T019|SY|38804009|SNOMEDCT_CORE|Gonadal dysgenesis syndrome|Gonadal dysgenesis syndrome
C0018081|T047|SY|15628003|SNOMEDCT_CORE|Clap|Gonorrhea
C0018081|T047|SY|15628003|SNOMEDCT_CORE|GC - Gonococcus infection|Gonorrhea
C0018081|T047|SY|15628003|SNOMEDCT_CORE|GCI - Gonococcal infection|Gonorrhea
C0018081|T047|SY|15628003|SNOMEDCT_CORE|Gonococcal infection|Gonorrhea
C0018081|T047|IS|15628003|SNOMEDCT_CORE|Gonococcal infection, NOS|Gonorrhea
C0018081|T047|PT|15628003|SNOMEDCT_CORE|Gonorrhea|Gonorrhea
C0018081|T047|FN|15628003|SNOMEDCT_CORE|Gonorrhea|Gonorrhea
C0018081|T047|IS|15628003|SNOMEDCT_CORE|Gonorrhea, NOS|Gonorrhea
C0018081|T047|PTGB|15628003|SNOMEDCT_CORE|Gonorrhoea|Gonorrhea
C0018081|T047|IS|15628003|SNOMEDCT_CORE|Infection due to Neisseria gonorrheae|Gonorrhea
C0018081|T047|SYGB|15628003|SNOMEDCT_CORE|Infection due to Neisseria gonorrhoeae|Gonorrhea
C0018099|T047|PT|90560007|SNOMEDCT_CORE|Gout|Gout
C0018099|T047|OF|90560007|SNOMEDCT_CORE|Gout|Gout
C0018099|T047|IS|90560007|SNOMEDCT_CORE|Gout, NOS|Gout
C0018099|T047|SY|90560007|SNOMEDCT_CORE|Inflammatory disorder due to increased blood urate level|Gout
C0018099|T047|FN|90560007|SNOMEDCT_CORE|Inflammatory disorder due to increased blood urate level|Gout
C0018133|T047|PT|234646005|SNOMEDCT_CORE|Graft versus host disease|Graft versus host disease
C0018133|T047|SY|234646005|SNOMEDCT_CORE|Graft-versus-host disease|Graft versus host disease
C0018133|T047|FN|234646005|SNOMEDCT_CORE|Graft-versus-host disease|Graft versus host disease
C0018133|T047|SY|234646005|SNOMEDCT_CORE|GVHD - Graft-versus-host disease|Graft versus host disease
C0018213|T047|SY|353295004|SNOMEDCT_CORE|Basedow disease|Graves' disease
C0018213|T047|SY|353295004|SNOMEDCT_CORE|Basedow's disease|Graves' disease
C0018213|T047|SY|353295004|SNOMEDCT_CORE|Exophthalmic goiter|Graves' disease
C0018213|T047|SYGB|353295004|SNOMEDCT_CORE|Exophthalmic goitre|Graves' disease
C0018213|T047|SY|353295004|SNOMEDCT_CORE|Graves disease|Graves' disease
C0018213|T047|PT|353295004|SNOMEDCT_CORE|Graves' disease|Graves' disease
C0018213|T047|FN|353295004|SNOMEDCT_CORE|Graves' disease|Graves' disease
C0018378|T047|IS|40956001|SNOMEDCT_CORE|GBS - Guillain-Barre syndrome|Guillain-Barré syndrome
C0018378|T047|SY|40956001|SNOMEDCT_CORE|Guillain Barre syndrome|Guillain-Barré syndrome
C0018378|T047|SY|40956001|SNOMEDCT_CORE|Guillain-Barre syndrome|Guillain-Barré syndrome
C0018378|T047|PT|40956001|SNOMEDCT_CORE|Guillain-Barré syndrome|Guillain-Barré syndrome
C0018378|T047|FN|40956001|SNOMEDCT_CORE|Guillain-Barré syndrome|Guillain-Barré syndrome
C0018378|T047|OF|40956001|SNOMEDCT_CORE|Guillain-Barre syndrome|Guillain-Barré syndrome
C0018378|T047|SY|40956001|SNOMEDCT_CORE|Landry-Guillain-Barre syndrome|Guillain-Barré syndrome
C0018418|T047|PTGB|4754008|SNOMEDCT_CORE|Gynaecomastia|Gynecomastia
C0018418|T047|SYGB|4754008|SNOMEDCT_CORE|Gynaecomazia|Gynecomastia
C0018418|T047|PT|4754008|SNOMEDCT_CORE|Gynecomastia|Gynecomastia
C0018418|T047|FN|4754008|SNOMEDCT_CORE|Gynecomastia|Gynecomastia
C0018418|T047|SY|4754008|SNOMEDCT_CORE|Gynecomazia|Gynecomastia
C0018418|T047|SY|4754008|SNOMEDCT_CORE|Hypertrophy of male breast|Gynecomastia
C0018520|T184|SY|79879001|SNOMEDCT_CORE|Bad breath|Breath smells unpleasant
C0018520|T184|SY|79879001|SNOMEDCT_CORE|Bad breath - halitosis|Breath smells unpleasant
C0018520|T184|SY|79879001|SNOMEDCT_CORE|Breath smells offensive|Breath smells unpleasant
C0018520|T184|PT|79879001|SNOMEDCT_CORE|Breath smells unpleasant|Breath smells unpleasant
C0018520|T184|FN|79879001|SNOMEDCT_CORE|Breath smells unpleasant|Breath smells unpleasant
C0018520|T184|SY|79879001|SNOMEDCT_CORE|Fetor ex ore|Breath smells unpleasant
C0018520|T184|SY|79879001|SNOMEDCT_CORE|Fetor oris|Breath smells unpleasant
C0018520|T184|SY|79879001|SNOMEDCT_CORE|Foul breath|Breath smells unpleasant
C0018520|T184|IS|79879001|SNOMEDCT_CORE|Halitosis|Breath smells unpleasant
C0018520|T184|SY|79879001|SNOMEDCT_CORE|Smelly breath|Breath smells unpleasant
C0018520|T184|SY|79879001|SNOMEDCT_CORE|Stomatodysodia|Breath smells unpleasant
C0018524|T048|IS|7011001|SNOMEDCT_CORE|Hallucination|Hallucinations
C0018524|T048|IS|7011001|SNOMEDCT_CORE|Hallucination, NOS|Hallucinations
C0018524|T048|PT|7011001|SNOMEDCT_CORE|Hallucinations|Hallucinations
C0018524|T048|FN|7011001|SNOMEDCT_CORE|Hallucinations|Hallucinations
C0018536|T190|SY|122480009|SNOMEDCT_CORE|Hallux abductovalgus|Hallux valgus
C0018536|T190|PT|122480009|SNOMEDCT_CORE|Hallux valgus|Hallux valgus
C0018536|T190|FN|122480009|SNOMEDCT_CORE|Hallux valgus|Hallux valgus
C0018536|T190|SY|122480009|SNOMEDCT_CORE|HAV - Hallux abductovalgus|Hallux valgus
C0018536|T190|SY|122480009|SNOMEDCT_CORE|HV - Hallux valgus|Hallux valgus
C0018564|T190|PT|299033004|SNOMEDCT_CORE|Deformity of hand|Deformity of hand
C0018564|T190|FN|299033004|SNOMEDCT_CORE|Deformity of hand|Deformity of hand
C0018571|T037|SY|125599006|SNOMEDCT_CORE|Hand injury|Injury of hand
C0018571|T037|PT|125599006|SNOMEDCT_CORE|Injury of hand|Injury of hand
C0018571|T037|FN|125599006|SNOMEDCT_CORE|Injury of hand|Injury of hand
C0018572|T047|PT|266108008|SNOMEDCT_CORE|Enteroviral vesicular stomatitis with exanthem|Enteroviral vesicular stomatitis with exanthem
C0018572|T047|SY|266108008|SNOMEDCT_CORE|Hand foot and mouth disease|Enteroviral vesicular stomatitis with exanthem
C0018572|T047|FN|266108008|SNOMEDCT_CORE|Hand foot and mouth disease|Enteroviral vesicular stomatitis with exanthem
C0018572|T047|SY|266108008|SNOMEDCT_CORE|Hand, foot and mouth disease|Enteroviral vesicular stomatitis with exanthem
C0018572|T047|SY|266108008|SNOMEDCT_CORE|Vesicular stomatitis with xanthem|Enteroviral vesicular stomatitis with exanthem
C0018621|T047|FN|21719001|SNOMEDCT_CORE|Allergic rhinitis caused by pollen|Seasonal allergic rhinitis
C0018621|T047|SY|21719001|SNOMEDCT_CORE|Allergic rhinitis caused by pollen|Seasonal allergic rhinitis
C0018621|T047|SY|21719001|SNOMEDCT_CORE|Allergic rhinitis caused by pollens|Seasonal allergic rhinitis
C0018621|T047|PT|21719001|SNOMEDCT_CORE|Allergic rhinitis due to pollen|Seasonal allergic rhinitis
C0018621|T047|OF|21719001|SNOMEDCT_CORE|Allergic rhinitis due to pollen|Seasonal allergic rhinitis
C0018621|T047|SY|21719001|SNOMEDCT_CORE|Allergic rhinitis due to pollens|Seasonal allergic rhinitis
C0018621|T047|SY|21719001|SNOMEDCT_CORE|Hay fever|Seasonal allergic rhinitis
C0018621|T047|SY|21719001|SNOMEDCT_CORE|Hayfever|Seasonal allergic rhinitis
C0018621|T047|SY|21719001|SNOMEDCT_CORE|Pollinosis|Seasonal allergic rhinitis
C0018621|T047|PT|367498001|SNOMEDCT_CORE|Seasonal allergic rhinitis|Seasonal allergic rhinitis
C0018621|T047|FN|367498001|SNOMEDCT_CORE|Seasonal allergic rhinitis|Seasonal allergic rhinitis
C0018621|T047|SY|367498001|SNOMEDCT_CORE|Spasmodic rhinorrhea|Seasonal allergic rhinitis
C0018621|T047|SYGB|367498001|SNOMEDCT_CORE|Spasmodic rhinorrhoea|Seasonal allergic rhinitis
C0018674|T037|SY|82271004|SNOMEDCT_CORE|Head injury|Injury of head
C0018674|T037|IS|82271004|SNOMEDCT_CORE|Head injury, NOS|Injury of head
C0018674|T037|SY|82271004|SNOMEDCT_CORE|HI - Head injury|Injury of head
C0018674|T037|PT|82271004|SNOMEDCT_CORE|Injury of head|Injury of head
C0018674|T037|FN|82271004|SNOMEDCT_CORE|Injury of head|Injury of head
C0018674|T037|SY|82271004|SNOMEDCT_CORE|Injury of head region|Injury of head
C0018674|T037|IS|82271004|SNOMEDCT_CORE|Injury of head, NOS|Injury of head
C0018681|T184|SY|25064002|SNOMEDCT_CORE|Cephalalgia|Headache
C0018681|T184|SY|25064002|SNOMEDCT_CORE|Cephalgia|Headache
C0018681|T184|SY|25064002|SNOMEDCT_CORE|Cephalodynia|Headache
C0018681|T184|SY|25064002|SNOMEDCT_CORE|HA - Headache|Headache
C0018681|T184|SY|25064002|SNOMEDCT_CORE|Head pain|Headache
C0018681|T184|PT|25064002|SNOMEDCT_CORE|Headache|Headache
C0018681|T184|FN|25064002|SNOMEDCT_CORE|Headache|Headache
C0018681|T184|IS|25064002|SNOMEDCT_CORE|Headache, NOS|Headache
C0018681|T184|SY|25064002|SNOMEDCT_CORE|Pain in head|Headache
C0018772|T033|PT|343087000|SNOMEDCT_CORE|Partial deafness|Partial deafness
C0018772|T033|OF|343087000|SNOMEDCT_CORE|Partial deafness|Partial deafness
C0018772|T033|FN|343087000|SNOMEDCT_CORE|Partial deafness|Partial deafness
C0018775|T047|PT|95820000|SNOMEDCT_CORE|Bilateral hearing loss|Bilateral hearing loss
C0018775|T047|OF|95820000|SNOMEDCT_CORE|Bilateral hearing loss|Bilateral hearing loss
C0018775|T047|FN|95820000|SNOMEDCT_CORE|Bilateral hearing loss|Bilateral hearing loss
C0018777|T047|SY|44057004|SNOMEDCT_CORE|CD - Conductive deafness|Conductive hearing loss
C0018777|T047|SY|44057004|SNOMEDCT_CORE|CHL - Conductive hearing loss|Conductive hearing loss
C0018777|T047|SY|44057004|SNOMEDCT_CORE|Conductive deafness|Conductive hearing loss
C0018777|T047|IS|44057004|SNOMEDCT_CORE|Conductive deafness, NOS|Conductive hearing loss
C0018777|T047|PT|44057004|SNOMEDCT_CORE|Conductive hearing loss|Conductive hearing loss
C0018777|T047|OF|44057004|SNOMEDCT_CORE|Conductive hearing loss|Conductive hearing loss
C0018777|T047|FN|44057004|SNOMEDCT_CORE|Conductive hearing loss|Conductive hearing loss
C0018777|T047|IS|44057004|SNOMEDCT_CORE|Conductive hearing loss, NOS|Conductive hearing loss
C0018780|T047|PT|232326009|SNOMEDCT_CORE|High frequency deafness|High frequency deafness
C0018780|T047|OF|232326009|SNOMEDCT_CORE|High frequency deafness|High frequency deafness
C0018780|T047|FN|232326009|SNOMEDCT_CORE|High frequency deafness|High frequency deafness
C0018784|T047|SY|60700002|SNOMEDCT_CORE|Neurosensory deafness|Sensorineural hearing loss
C0018784|T047|SY|60700002|SNOMEDCT_CORE|PD - Perceptive deafness|Sensorineural hearing loss
C0018784|T047|SY|60700002|SNOMEDCT_CORE|Perceptive deafness|Sensorineural hearing loss
C0018784|T047|IS|60700002|SNOMEDCT_CORE|Perceptive deafness, NOS|Sensorineural hearing loss
C0018784|T047|SY|60700002|SNOMEDCT_CORE|Perceptive hearing loss|Sensorineural hearing loss
C0018784|T047|IS|60700002|SNOMEDCT_CORE|Perceptive hearing loss, NOS|Sensorineural hearing loss
C0018784|T047|SY|60700002|SNOMEDCT_CORE|Sensorineural deafness|Sensorineural hearing loss
C0018784|T047|FN|60700002|SNOMEDCT_CORE|Sensorineural hearing loss|Sensorineural hearing loss
C0018784|T047|PT|60700002|SNOMEDCT_CORE|Sensorineural hearing loss|Sensorineural hearing loss
C0018784|T047|OF|60700002|SNOMEDCT_CORE|Sensorineural hearing loss|Sensorineural hearing loss
C0018784|T047|IS|60700002|SNOMEDCT_CORE|Sensorineural hearing loss, NOS|Sensorineural hearing loss
C0018784|T047|SY|60700002|SNOMEDCT_CORE|Sensory-neural deafness|Sensorineural hearing loss
C0018784|T047|SY|60700002|SNOMEDCT_CORE|Sensory-neural hearing loss|Sensorineural hearing loss
C0018784|T047|SY|60700002|SNOMEDCT_CORE|SND - Sensorineural deafness|Sensorineural hearing loss
C0018784|T047|SY|60700002|SNOMEDCT_CORE|SNHL - Sensorineural hearing loss|Sensorineural hearing loss
C0018790|T047|PT|410429000|SNOMEDCT_CORE|Cardiac arrest|Cardiac arrest
C0018790|T047|FN|410429000|SNOMEDCT_CORE|Cardiac arrest|Cardiac arrest
C0018794|T047|SY|233916004|SNOMEDCT_CORE|HB - Heart block|Heart block
C0018794|T047|PT|233916004|SNOMEDCT_CORE|Heart block|Heart block
C0018794|T047|FN|233916004|SNOMEDCT_CORE|Heart block|Heart block
C0018798|T019|SY|13213009|SNOMEDCT_CORE|Congenital anomaly of heart|Congenital anomaly of heart
C0018798|T019|IS|13213009|SNOMEDCT_CORE|Congenital anomaly of heart, NOS|Congenital anomaly of heart
C0018799|T047|SY|56265001|SNOMEDCT_CORE|Cardiac disorder|Heart disease
C0018799|T047|SY|56265001|SNOMEDCT_CORE|Cardiopathy|Heart disease
C0018799|T047|IS|56265001|SNOMEDCT_CORE|Cardiopathy, NOS|Heart disease
C0018799|T047|SY|56265001|SNOMEDCT_CORE|Disorder of heart|Heart disease
C0018799|T047|PT|56265001|SNOMEDCT_CORE|Heart disease|Heart disease
C0018799|T047|FN|56265001|SNOMEDCT_CORE|Heart disease|Heart disease
C0018799|T047|IS|56265001|SNOMEDCT_CORE|Heart disease, NOS|Heart disease
C0018799|T047|SY|56265001|SNOMEDCT_CORE|Morbus cordis|Heart disease
C0018799|T047|IS|56265001|SNOMEDCT_CORE|Morbus cordis, NOS|Heart disease
C0018800|T033|PT|8186001|SNOMEDCT_CORE|Cardiomegaly|Cardiomegaly
C0018800|T033|FN|8186001|SNOMEDCT_CORE|Cardiomegaly|Cardiomegaly
C0018800|T033|SY|8186001|SNOMEDCT_CORE|Enlarged heart|Cardiomegaly
C0018801|T047|SY|84114007|SNOMEDCT_CORE|Cardiac failure|Heart failure
C0018801|T047|IS|84114007|SNOMEDCT_CORE|Cardiac failure, NOS|Heart failure
C0018801|T047|SY|84114007|SNOMEDCT_CORE|Cardiac insufficiency|Heart failure
C0018801|T047|PT|84114007|SNOMEDCT_CORE|Heart failure|Heart failure
C0018801|T047|FN|84114007|SNOMEDCT_CORE|Heart failure|Heart failure
C0018801|T047|IS|84114007|SNOMEDCT_CORE|Heart failure, NOS|Heart failure
C0018801|T047|SY|84114007|SNOMEDCT_CORE|HF - Heart failure|Heart failure
C0018801|T047|SY|84114007|SNOMEDCT_CORE|Weak heart|Heart failure
C0018801|T047|IS|84114007|SNOMEDCT_CORE|Weak heart, NOS|Heart failure
C0018802|T047|SY|42343007|SNOMEDCT_CORE|CCF - Congestive cardiac failure|Congestive heart failure
C0018802|T047|SY|42343007|SNOMEDCT_CORE|CHF - Congestive heart failure|Congestive heart failure
C0018802|T047|SY|42343007|SNOMEDCT_CORE|Congestive cardiac failure|Congestive heart failure
C0018802|T047|SY|42343007|SNOMEDCT_CORE|Congestive heart disease|Congestive heart failure
C0018802|T047|PT|42343007|SNOMEDCT_CORE|Congestive heart failure|Congestive heart failure
C0018802|T047|FN|42343007|SNOMEDCT_CORE|Congestive heart failure|Congestive heart failure
C0018808|T033|IS|88610006|SNOMEDCT_CORE|Cardiac murmur|Heart murmur
C0018808|T033|IS|88610006|SNOMEDCT_CORE|Cardiac murmur, NOS|Heart murmur
C0018808|T033|SY|88610006|SNOMEDCT_CORE|Finding of heart murmur|Heart murmur
C0018808|T033|PT|88610006|SNOMEDCT_CORE|Heart murmur|Heart murmur
C0018808|T033|FN|88610006|SNOMEDCT_CORE|Heart murmur|Heart murmur
C0018808|T033|IS|88610006|SNOMEDCT_CORE|Heart murmur, NOS|Heart murmur
C0018808|T033|IS|88610006|SNOMEDCT_CORE|Murmur|Heart murmur
C0018808|T033|IS|88610006|SNOMEDCT_CORE|Murmur, NOS|Heart murmur
C0018808|T033|SY|88610006|SNOMEDCT_CORE|Observation of heart murmur|Heart murmur
C0018817|T019|SY|70142008|SNOMEDCT_CORE|ASD - Atrial septal defect|Atrial septal defect
C0018817|T019|PT|70142008|SNOMEDCT_CORE|Atrial septal defect|Atrial septal defect
C0018817|T019|FN|70142008|SNOMEDCT_CORE|Atrial septal defect|Atrial septal defect
C0018817|T019|SY|70142008|SNOMEDCT_CORE|Interatrial septal defect|Atrial septal defect
C0018818|T019|SY|30288003|SNOMEDCT_CORE|Interventricular septal defect|Ventricular septal defect
C0018818|T019|IS|30288003|SNOMEDCT_CORE|Ventricular septal abnormality|Ventricular septal defect
C0018818|T019|PT|30288003|SNOMEDCT_CORE|Ventricular septal defect|Ventricular septal defect
C0018818|T019|FN|30288003|SNOMEDCT_CORE|Ventricular septal defect|Ventricular septal defect
C0018818|T019|SY|30288003|SNOMEDCT_CORE|VSD - Ventricular septal defect|Ventricular septal defect
C0018824|T047|SY|368009|SNOMEDCT_CORE|Disorder of heart valve|Heart valve disorder
C0018824|T047|SY|368009|SNOMEDCT_CORE|Heart valve disease|Heart valve disorder
C0018824|T047|PT|368009|SNOMEDCT_CORE|Heart valve disorder|Heart valve disorder
C0018824|T047|FN|368009|SNOMEDCT_CORE|Heart valve disorder|Heart valve disorder
C0018824|T047|IS|368009|SNOMEDCT_CORE|Heart valve disorder, NOS|Heart valve disorder
C0018824|T047|SY|368009|SNOMEDCT_CORE|Valvular heart disease|Heart valve disorder
C0018824|T047|IS|368009|SNOMEDCT_CORE|Valvular heart disease, NOS|Heart valve disorder
C0018834|T184|SY|16331000|SNOMEDCT_CORE|Burning reflux|Heartburn
C0018834|T184|PT|16331000|SNOMEDCT_CORE|Heartburn|Heartburn
C0018834|T184|FN|16331000|SNOMEDCT_CORE|Heartburn|Heartburn
C0018834|T184|SY|16331000|SNOMEDCT_CORE|Heartburn symptom|Heartburn
C0018834|T184|SY|16331000|SNOMEDCT_CORE|Pyrosis|Heartburn
C0018916|T191|PTGB|400210000|SNOMEDCT_CORE|Haemangioma|Hemangioma
C0018916|T191|PT|400210000|SNOMEDCT_CORE|Hemangioma|Hemangioma
C0018916|T191|FN|400210000|SNOMEDCT_CORE|Hemangioma|Hemangioma
C0018924|T046|SY|81808003|SNOMEDCT_CORE|Bleeding into joint|Hemarthrosis
C0018924|T046|PTGB|81808003|SNOMEDCT_CORE|Haemarthrosis|Hemarthrosis
C0018924|T046|IS|81808003|SNOMEDCT_CORE|Haemarthrosis, NOS|Hemarthrosis
C0018924|T046|PT|81808003|SNOMEDCT_CORE|Hemarthrosis|Hemarthrosis
C0018924|T046|FN|81808003|SNOMEDCT_CORE|Hemarthrosis|Hemarthrosis
C0018924|T046|IS|81808003|SNOMEDCT_CORE|Hemarthrosis, NOS|Hemarthrosis
C0018926|T184|PTGB|8765009|SNOMEDCT_CORE|Haematemesis|Hematemesis
C0018926|T184|PT|8765009|SNOMEDCT_CORE|Hematemesis|Hematemesis
C0018926|T184|FN|8765009|SNOMEDCT_CORE|Hematemesis|Hematemesis
C0018926|T184|SY|8765009|SNOMEDCT_CORE|Vomiting blood|Hematemesis
C0018926|T184|SY|8765009|SNOMEDCT_CORE|Vomiting of blood|Hematemesis
C0018932|T047|SYGB|405729008|SNOMEDCT_CORE|Blood in faeces|Hematochezia
C0018932|T047|SY|405729008|SNOMEDCT_CORE|Blood in feces|Hematochezia
C0018932|T047|SY|405729008|SNOMEDCT_CORE|Blood in stool|Hematochezia
C0018932|T047|SY|405729008|SNOMEDCT_CORE|Bloody stool|Hematochezia
C0018932|T047|IS|405729008|SNOMEDCT_CORE|BRBPR|Hematochezia
C0018932|T047|SY|405729008|SNOMEDCT_CORE|BRBPR - Bright red blood per rectum|Hematochezia
C0018932|T047|SY|405729008|SNOMEDCT_CORE|Bright red blood in stool|Hematochezia
C0018932|T047|SY|405729008|SNOMEDCT_CORE|Bright red blood per rectum|Hematochezia
C0018932|T047|SYGB|405729008|SNOMEDCT_CORE|Faeces: blood|Hematochezia
C0018932|T047|SY|405729008|SNOMEDCT_CORE|Feces: blood|Hematochezia
C0018932|T047|SY|405729008|SNOMEDCT_CORE|Fresh blood passed per rectum|Hematochezia
C0018932|T047|PTGB|405729008|SNOMEDCT_CORE|Haematochezia|Hematochezia
C0018932|T047|PT|405729008|SNOMEDCT_CORE|Hematochezia|Hematochezia
C0018932|T047|FN|405729008|SNOMEDCT_CORE|Hematochezia|Hematochezia
C0018932|T047|SY|405729008|SNOMEDCT_CORE|Passage of bloody stools|Hematochezia
C0018944|T046|PTGB|385494008|SNOMEDCT_CORE|Haematoma|Hematoma
C0018944|T046|PT|385494008|SNOMEDCT_CORE|Hematoma|Hematoma
C0018944|T046|FN|385494008|SNOMEDCT_CORE|Hematoma|Hematoma
C0018946|T046|PTGB|35486000|SNOMEDCT_CORE|Subdural haemorrhage|Subdural hemorrhage
C0018946|T046|PT|35486000|SNOMEDCT_CORE|Subdural hemorrhage|Subdural hemorrhage
C0018946|T046|OF|35486000|SNOMEDCT_CORE|Subdural hemorrhage|Subdural hemorrhage
C0018946|T046|IS|35486000|SNOMEDCT_CORE|Subdural hemorrhage, NOS|Subdural hemorrhage
C0018946|T046|SYGB|35486000|SNOMEDCT_CORE|Subdural intracranial haemorrhage|Subdural hemorrhage
C0018946|T046|SY|35486000|SNOMEDCT_CORE|Subdural intracranial hemorrhage|Subdural hemorrhage
C0018946|T046|FN|35486000|SNOMEDCT_CORE|Subdural intracranial hemorrhage|Subdural hemorrhage
C0018948|T046|PTGB|38280009|SNOMEDCT_CORE|Haematometra|Hematometra
C0018948|T046|SYGB|38280009|SNOMEDCT_CORE|Haemometra|Hematometra
C0018948|T046|PT|38280009|SNOMEDCT_CORE|Hematometra|Hematometra
C0018948|T046|FN|38280009|SNOMEDCT_CORE|Hematometra|Hematometra
C0018948|T046|SY|38280009|SNOMEDCT_CORE|Hemometra|Hematometra
C0018965|T047|PT|34436003|SNOMEDCT_CORE|Blood in urine|Blood in urine
C0018965|T047|FN|34436003|SNOMEDCT_CORE|Blood in urine|Blood in urine
C0018965|T047|SYGB|53298000|SNOMEDCT_CORE|Blood in urine - haematuria|Blood in urine
C0018965|T047|SY|53298000|SNOMEDCT_CORE|Blood in urine - hematuria|Blood in urine
C0018965|T047|SYGB|34436003|SNOMEDCT_CORE|Haematuria|Blood in urine
C0018965|T047|PTGB|53298000|SNOMEDCT_CORE|Haematuria syndrome|Blood in urine
C0018965|T047|SY|34436003|SNOMEDCT_CORE|Hematuria|Blood in urine
C0018965|T047|PT|53298000|SNOMEDCT_CORE|Hematuria syndrome|Blood in urine
C0018965|T047|FN|53298000|SNOMEDCT_CORE|Hematuria syndrome|Blood in urine
C0018965|T047|IS|53298000|SNOMEDCT_CORE|Hematuria syndrome, NOS|Blood in urine
C0018979|T047|PT|77674003|SNOMEDCT_CORE|Hemianopia|Hemianopia
C0018979|T047|FN|77674003|SNOMEDCT_CORE|Hemianopia|Hemianopia
C0018979|T047|IS|77674003|SNOMEDCT_CORE|Hemianopia, NOS|Hemianopia
C0018979|T047|IS|77674003|SNOMEDCT_CORE|Hemianopsia|Hemianopia
C0018979|T047|IS|77674003|SNOMEDCT_CORE|Hemianopsia, NOS|Hemianopia
C0018989|T184|PT|20022000|SNOMEDCT_CORE|Hemiparesis|Hemiparesis
C0018989|T184|FN|20022000|SNOMEDCT_CORE|Hemiparesis|Hemiparesis
C0018989|T184|SY|20022000|SNOMEDCT_CORE|Weakness of one side of body|Hemiparesis
C0018991|T184|PT|50582007|SNOMEDCT_CORE|Hemiplegia|Hemiplegia
C0018991|T184|FN|50582007|SNOMEDCT_CORE|Hemiplegia|Hemiplegia
C0018991|T184|IS|50582007|SNOMEDCT_CORE|Hemiplegia, NOS|Hemiplegia
C0018995|T047|PTGB|399187006|SNOMEDCT_CORE|Haemochromatosis|Hemochromatosis
C0018995|T047|PT|399187006|SNOMEDCT_CORE|Hemochromatosis|Hemochromatosis
C0018995|T047|FN|399187006|SNOMEDCT_CORE|Hemochromatosis|Hemochromatosis
C0018995|T047|SY|399187006|SNOMEDCT_CORE|Iron storage disease|Hemochromatosis
C0019045|T047|SY|80141007|SNOMEDCT_CORE|Globin abnormality|Hemoglobinopathy
C0019045|T047|IS|80141007|SNOMEDCT_CORE|Globin abnormality, NOS|Hemoglobinopathy
C0019045|T047|SYGB|80141007|SNOMEDCT_CORE|Haemoglobin disease|Hemoglobinopathy
C0019045|T047|IS|80141007|SNOMEDCT_CORE|Haemoglobin disease, NOS|Hemoglobinopathy
C0019045|T047|SYGB|80141007|SNOMEDCT_CORE|Haemoglobin disorder|Hemoglobinopathy
C0019045|T047|IS|80141007|SNOMEDCT_CORE|Haemoglobin disorder, NOS|Hemoglobinopathy
C0019045|T047|PTGB|80141007|SNOMEDCT_CORE|Haemoglobinopathy|Hemoglobinopathy
C0019045|T047|IS|80141007|SNOMEDCT_CORE|Haemoglobinopathy, NOS|Hemoglobinopathy
C0019045|T047|SY|80141007|SNOMEDCT_CORE|Hemoglobin disease|Hemoglobinopathy
C0019045|T047|IS|80141007|SNOMEDCT_CORE|Hemoglobin disease, NOS|Hemoglobinopathy
C0019045|T047|SY|80141007|SNOMEDCT_CORE|Hemoglobin disorder|Hemoglobinopathy
C0019045|T047|IS|80141007|SNOMEDCT_CORE|Hemoglobin disorder, NOS|Hemoglobinopathy
C0019045|T047|PT|80141007|SNOMEDCT_CORE|Hemoglobinopathy|Hemoglobinopathy
C0019045|T047|FN|80141007|SNOMEDCT_CORE|Hemoglobinopathy|Hemoglobinopathy
C0019045|T047|IS|80141007|SNOMEDCT_CORE|Hemoglobinopathy, NOS|Hemoglobinopathy
C0019061|T047|SY|111407006|SNOMEDCT_CORE|Gasser's syndrome|Hemolytic uremic syndrome
C0019061|T047|PTGB|111407006|SNOMEDCT_CORE|Haemolytic uraemic syndrome|Hemolytic uremic syndrome
C0019061|T047|IS|111407006|SNOMEDCT_CORE|Haemolytic uraemic syndrome, NOS|Hemolytic uremic syndrome
C0019061|T047|PT|111407006|SNOMEDCT_CORE|Hemolytic uremic syndrome|Hemolytic uremic syndrome
C0019061|T047|FN|111407006|SNOMEDCT_CORE|Hemolytic uremic syndrome|Hemolytic uremic syndrome
C0019061|T047|IS|111407006|SNOMEDCT_CORE|Hemolytic uremic syndrome, NOS|Hemolytic uremic syndrome
C0019061|T047|SYGB|111407006|SNOMEDCT_CORE|HUS - Haemolytic uraemic syndrome|Hemolytic uremic syndrome
C0019061|T047|SY|111407006|SNOMEDCT_CORE|HUS - Hemolytic uremic syndrome|Hemolytic uremic syndrome
C0019065|T046|SY|45626005|SNOMEDCT_CORE|Abdominal apoplexy|Hemoperitoneum
C0019065|T046|SYGB|45626005|SNOMEDCT_CORE|Haemoperitoneum|Hemoperitoneum
C0019065|T046|SY|45626005|SNOMEDCT_CORE|Hemoperitoneum|Hemoperitoneum
C0019065|T046|IS|45626005|SNOMEDCT_CORE|Hemoperitoneum, NOS|Hemoperitoneum
C0019065|T046|SYGB|45626005|SNOMEDCT_CORE|Peritoneal haemorrhage|Hemoperitoneum
C0019065|T046|SY|45626005|SNOMEDCT_CORE|Peritoneal hemorrhage|Hemoperitoneum
C0019065|T046|IS|45626005|SNOMEDCT_CORE|Peritoneal hemorrhage, NOS|Hemoperitoneum
C0019066|T046|SYGB|45626005|SNOMEDCT_CORE|Haemoperitoneum - non-traumatic|Nontraumatic hemoperitoneum
C0019066|T046|SY|45626005|SNOMEDCT_CORE|Hemoperitoneum - non-traumatic|Nontraumatic hemoperitoneum
C0019066|T046|PTGB|45626005|SNOMEDCT_CORE|Nontraumatic haemoperitoneum|Nontraumatic hemoperitoneum
C0019066|T046|PT|45626005|SNOMEDCT_CORE|Nontraumatic hemoperitoneum|Nontraumatic hemoperitoneum
C0019066|T046|FN|45626005|SNOMEDCT_CORE|Nontraumatic hemoperitoneum|Nontraumatic hemoperitoneum
C0019066|T046|SYGB|45626005|SNOMEDCT_CORE|Spontaneous intraperitoneal haemorrhage|Nontraumatic hemoperitoneum
C0019066|T046|SY|45626005|SNOMEDCT_CORE|Spontaneous intraperitoneal hemorrhage|Nontraumatic hemoperitoneum
C0019069|T047|SY|28293008|SNOMEDCT_CORE|AHG deficiency disease|Hereditary factor VIII deficiency disease
C0019069|T047|SYGB|28293008|SNOMEDCT_CORE|Classical haemophilia|Hereditary factor VIII deficiency disease
C0019069|T047|SY|28293008|SNOMEDCT_CORE|Classical hemophilia|Hereditary factor VIII deficiency disease
C0019069|T047|SY|28293008|SNOMEDCT_CORE|Congenital factor VIII deficiency|Hereditary factor VIII deficiency disease
C0019069|T047|SY|28293008|SNOMEDCT_CORE|Congenital factor VIII deficiency disease|Hereditary factor VIII deficiency disease
C0019069|T047|SYGB|28293008|SNOMEDCT_CORE|Haemophilia A|Hereditary factor VIII deficiency disease
C0019069|T047|IS|28293008|SNOMEDCT_CORE|Haemophilia A, NOS|Hereditary factor VIII deficiency disease
C0019069|T047|SY|28293008|SNOMEDCT_CORE|Hemophilia A|Hereditary factor VIII deficiency disease
C0019069|T047|OF|28293008|SNOMEDCT_CORE|Hemophilia A|Hereditary factor VIII deficiency disease
C0019069|T047|IS|28293008|SNOMEDCT_CORE|Hemophilia A, NOS|Hereditary factor VIII deficiency disease
C0019069|T047|PT|28293008|SNOMEDCT_CORE|Hereditary factor VIII deficiency disease|Hereditary factor VIII deficiency disease
C0019069|T047|FN|28293008|SNOMEDCT_CORE|Hereditary factor VIII deficiency disease|Hereditary factor VIII deficiency disease
C0019069|T047|SY|28293008|SNOMEDCT_CORE|Sex-linked factor VIII deficiency|Hereditary factor VIII deficiency disease
C0019079|T184|SY|66857006|SNOMEDCT_CORE|Coughing up blood|Hemoptysis
C0019079|T184|PTGB|66857006|SNOMEDCT_CORE|Haemoptysis|Hemoptysis
C0019079|T184|PT|66857006|SNOMEDCT_CORE|Hemoptysis|Hemoptysis
C0019079|T184|FN|66857006|SNOMEDCT_CORE|Hemoptysis|Hemoptysis
C0019079|T184|OF|66857006|SNOMEDCT_CORE|Hemoptysis|Hemoptysis
C0019080|T046|PT|131148009|SNOMEDCT_CORE|Bleeding|Bleeding
C0019080|T046|FN|131148009|SNOMEDCT_CORE|Bleeding|Bleeding
C0019080|T046|SYGB|131148009|SNOMEDCT_CORE|Haemorrhage|Bleeding
C0019080|T046|SY|131148009|SNOMEDCT_CORE|Hemorrhage|Bleeding
C0019081|T046|PTGB|266464001|SNOMEDCT_CORE|Haemorrhage of rectum and anus|Hemorrhage of rectum and anus
C0019081|T046|PT|266464001|SNOMEDCT_CORE|Hemorrhage of rectum and anus|Hemorrhage of rectum and anus
C0019081|T046|FN|266464001|SNOMEDCT_CORE|Hemorrhage of rectum and anus|Hemorrhage of rectum and anus
C0019112|T047|SYGB|70153002|SNOMEDCT_CORE|Haemorrhoid|Hemorrhoids
C0019112|T047|PTGB|70153002|SNOMEDCT_CORE|Haemorrhoids|Hemorrhoids
C0019112|T047|IS|70153002|SNOMEDCT_CORE|Haemorrhoids, NOS|Hemorrhoids
C0019112|T047|SY|70153002|SNOMEDCT_CORE|Hemorrhoid|Hemorrhoids
C0019112|T047|PT|70153002|SNOMEDCT_CORE|Hemorrhoids|Hemorrhoids
C0019112|T047|FN|70153002|SNOMEDCT_CORE|Hemorrhoids|Hemorrhoids
C0019112|T047|IS|70153002|SNOMEDCT_CORE|Hemorrhoids, NOS|Hemorrhoids
C0019112|T047|SY|70153002|SNOMEDCT_CORE|Piles|Hemorrhoids
C0019112|T047|SYGB|70153002|SNOMEDCT_CORE|Piles - haemorrhoids|Hemorrhoids
C0019112|T047|SY|70153002|SNOMEDCT_CORE|Piles - hemorrhoids|Hemorrhoids
C0019112|T047|IS|70153002|SNOMEDCT_CORE|Piles, NOS|Hemorrhoids
C0019123|T046|PTGB|31892009|SNOMEDCT_CORE|Haemothorax|Hemothorax
C0019123|T046|PT|31892009|SNOMEDCT_CORE|Hemothorax|Hemothorax
C0019123|T046|FN|31892009|SNOMEDCT_CORE|Hemothorax|Hemothorax
C0019123|T046|SYGB|31892009|SNOMEDCT_CORE|Pleural haemorrhage|Hemothorax
C0019123|T046|SY|31892009|SNOMEDCT_CORE|Pleural hemorrhage|Hemothorax
C0019151|T047|IS|13920009|SNOMEDCT_CORE|Gaustad's syndrome|Hepatic encephalopathy
C0019151|T047|SY|13920009|SNOMEDCT_CORE|HE - Hepatic encephalopathy|Hepatic encephalopathy
C0019151|T047|PT|13920009|SNOMEDCT_CORE|Hepatic encephalopathy|Hepatic encephalopathy
C0019151|T047|FN|13920009|SNOMEDCT_CORE|Hepatic encephalopathy|Hepatic encephalopathy
C0019151|T047|SY|13920009|SNOMEDCT_CORE|Hepatocerebral encephalopathy|Hepatic encephalopathy
C0019151|T047|IS|13920009|SNOMEDCT_CORE|Portal-systemic encephalopathy|Hepatic encephalopathy
C0019151|T047|IS|13920009|SNOMEDCT_CORE|Transient hepatargy syndrome|Hepatic encephalopathy
C0019154|T047|PT|38739001|SNOMEDCT_CORE|Hepatic vein thrombosis|Hepatic vein thrombosis
C0019154|T047|FN|38739001|SNOMEDCT_CORE|Hepatic vein thrombosis|Hepatic vein thrombosis
C0019158|T047|SY|128241005|SNOMEDCT_CORE|Hepatitis|Inflammatory disease of liver
C0019158|T047|PT|128241005|SNOMEDCT_CORE|Inflammatory disease of liver|Inflammatory disease of liver
C0019158|T047|FN|128241005|SNOMEDCT_CORE|Inflammatory disease of liver|Inflammatory disease of liver
C0019158|T047|SY|128241005|SNOMEDCT_CORE|Inflammatory disorder of liver|Inflammatory disease of liver
C0019158|T047|SY|128241005|SNOMEDCT_CORE|Inflammatory liver disease|Inflammatory disease of liver
C0019159|T047|SY|40468003|SNOMEDCT_CORE|Hepatitis A|Viral hepatitis, type A
C0019159|T047|SY|40468003|SNOMEDCT_CORE|IH - Infectious hepatitis|Viral hepatitis, type A
C0019159|T047|SY|40468003|SNOMEDCT_CORE|Infectious hepatitis|Viral hepatitis, type A
C0019159|T047|PT|40468003|SNOMEDCT_CORE|Viral hepatitis, type A|Viral hepatitis, type A
C0019159|T047|FN|40468003|SNOMEDCT_CORE|Viral hepatitis, type A|Viral hepatitis, type A
C0019163|T047|SY|66071002|SNOMEDCT_CORE|Hepatitis B|Type B viral hepatitis
C0019163|T047|SY|66071002|SNOMEDCT_CORE|Hepatitis B infection|Type B viral hepatitis
C0019163|T047|SY|66071002|SNOMEDCT_CORE|Serum hepatitis|Type B viral hepatitis
C0019163|T047|SY|66071002|SNOMEDCT_CORE|SH - Serum hepatitis|Type B viral hepatitis
C0019163|T047|PT|66071002|SNOMEDCT_CORE|Type B viral hepatitis|Type B viral hepatitis
C0019163|T047|OF|66071002|SNOMEDCT_CORE|Type B viral hepatitis|Type B viral hepatitis
C0019163|T047|SY|66071002|SNOMEDCT_CORE|Viral hepatitis type B|Type B viral hepatitis
C0019163|T047|FN|66071002|SNOMEDCT_CORE|Viral hepatitis type B|Type B viral hepatitis
C0019187|T047|SY|235875008|SNOMEDCT_CORE|AH - Alcoholic hepatitis|Alcoholic hepatitis
C0019187|T047|PT|235875008|SNOMEDCT_CORE|Alcoholic hepatitis|Alcoholic hepatitis
C0019187|T047|FN|235875008|SNOMEDCT_CORE|Alcoholic hepatitis|Alcoholic hepatitis
C0019189|T047|SY|76783007|SNOMEDCT_CORE|CH - Chronic hepatitis|Chronic hepatitis
C0019189|T047|PT|76783007|SNOMEDCT_CORE|Chronic hepatitis|Chronic hepatitis
C0019189|T047|FN|76783007|SNOMEDCT_CORE|Chronic hepatitis|Chronic hepatitis
C0019189|T047|IS|76783007|SNOMEDCT_CORE|Chronic hepatitis, NOS|Chronic hepatitis
C0019196|T047|SY|50711007|SNOMEDCT_CORE|Hepatitis C|Viral hepatitis C
C0019196|T047|IS|50711007|SNOMEDCT_CORE|Non-A, non-B hepatitis|Viral hepatitis C
C0019196|T047|SY|50711007|SNOMEDCT_CORE|Type C viral hepatitis|Viral hepatitis C
C0019196|T047|PT|50711007|SNOMEDCT_CORE|Viral hepatitis C|Viral hepatitis C
C0019196|T047|OF|50711007|SNOMEDCT_CORE|Viral hepatitis C|Viral hepatitis C
C0019196|T047|SY|50711007|SNOMEDCT_CORE|Viral hepatitis type C|Viral hepatitis C
C0019196|T047|FN|50711007|SNOMEDCT_CORE|Viral hepatitis type C|Viral hepatitis C
C0019196|T047|IS|50711007|SNOMEDCT_CORE|Viral hepatitis, non-A, non-B|Viral hepatitis C
C0019209|T033|SY|80515008|SNOMEDCT_CORE|Hepatomegaly|Large liver
C0019209|T033|PT|80515008|SNOMEDCT_CORE|Large liver|Large liver
C0019209|T033|FN|80515008|SNOMEDCT_CORE|Large liver|Large liver
C0019212|T047|SY|51292008|SNOMEDCT_CORE|Hepatorenal failure|Hepatorenal syndrome
C0019212|T047|PT|51292008|SNOMEDCT_CORE|Hepatorenal syndrome|Hepatorenal syndrome
C0019212|T047|FN|51292008|SNOMEDCT_CORE|Hepatorenal syndrome|Hepatorenal syndrome
C0019212|T047|SY|51292008|SNOMEDCT_CORE|HRF - Hepatorenal failure|Hepatorenal syndrome
C0019214|T184|PT|36760000|SNOMEDCT_CORE|Hepatosplenomegaly|Hepatosplenomegaly
C0019214|T184|FN|36760000|SNOMEDCT_CORE|Hepatosplenomegaly|Hepatosplenomegaly
C0019270|T190|SY|52515009|SNOMEDCT_CORE|Hernia|Hernia
C0019284|T047|PT|39839004|SNOMEDCT_CORE|Diaphragmatic hernia|Diaphragmatic hernia
C0019284|T047|FN|39839004|SNOMEDCT_CORE|Diaphragmatic hernia|Diaphragmatic hernia
C0019284|T047|IS|39839004|SNOMEDCT_CORE|Diaphragmatic hernia, NOS|Diaphragmatic hernia
C0019294|T190|SY|396232000|SNOMEDCT_CORE|IH - Inguinal hernia|Inguinal hernia
C0019294|T190|PT|396232000|SNOMEDCT_CORE|Inguinal hernia|Inguinal hernia
C0019294|T190|FN|396232000|SNOMEDCT_CORE|Inguinal hernia|Inguinal hernia
C0019311|T047|PT|29862005|SNOMEDCT_CORE|Paraumbilical hernia|Paraumbilical hernia
C0019311|T047|FN|29862005|SNOMEDCT_CORE|Paraumbilical hernia|Paraumbilical hernia
C0019311|T047|IS|29862005|SNOMEDCT_CORE|Paraumbilical hernia, NOS|Paraumbilical hernia
C0019322|T047|PT|396347007|SNOMEDCT_CORE|Umbilical hernia|Umbilical hernia
C0019322|T047|FN|396347007|SNOMEDCT_CORE|Umbilical hernia|Umbilical hernia
C0019326|T190|FN|414396006|SNOMEDCT_CORE|Hernia of anterior abdominal wall|Hernia of anterior abdominal wall
C0019326|T190|PT|414396006|SNOMEDCT_CORE|Hernia of anterior abdominal wall|Hernia of anterior abdominal wall
C0019326|T190|IS|414474001|SNOMEDCT_CORE|Ventral hernia|Hernia of anterior abdominal wall
C0019326|T190|SY|414396006|SNOMEDCT_CORE|Ventral hernia|Hernia of anterior abdominal wall
C0019337|T048|SY|231477003|SNOMEDCT_CORE|Heroin addiction|Heroin dependence
C0019337|T048|PT|231477003|SNOMEDCT_CORE|Heroin dependence|Heroin dependence
C0019337|T048|FN|231477003|SNOMEDCT_CORE|Heroin dependence|Heroin dependence
C0019338|T047|SY|186659004|SNOMEDCT_CORE|Enteroviral vesicular pharyngitis|Herpangina
C0019338|T047|PT|186659004|SNOMEDCT_CORE|Herpangina|Herpangina
C0019338|T047|FN|186659004|SNOMEDCT_CORE|Herpangina|Herpangina
C0019342|T047|PT|33839006|SNOMEDCT_CORE|Genital herpes simplex|Genital herpes simplex
C0019342|T047|FN|33839006|SNOMEDCT_CORE|Genital herpes simplex|Genital herpes simplex
C0019342|T047|IS|33839006|SNOMEDCT_CORE|Genital herpes simplex, NOS|Genital herpes simplex
C0019342|T047|SY|33839006|SNOMEDCT_CORE|Herpes genitalis|Genital herpes simplex
C0019345|T047|SY|1475003|SNOMEDCT_CORE|Cold sore|Herpes labialis
C0019345|T047|SY|1475003|SNOMEDCT_CORE|Cold sores|Herpes labialis
C0019345|T047|SY|1475003|SNOMEDCT_CORE|Fever blister|Herpes labialis
C0019345|T047|PT|1475003|SNOMEDCT_CORE|Herpes labialis|Herpes labialis
C0019345|T047|FN|1475003|SNOMEDCT_CORE|Herpes labialis|Herpes labialis
C0019345|T047|SY|1475003|SNOMEDCT_CORE|Herpes simplex labialis|Herpes labialis
C0019348|T047|PT|88594005|SNOMEDCT_CORE|Herpes simplex|Herpes simplex
C0019348|T047|FN|88594005|SNOMEDCT_CORE|Herpes simplex|Herpes simplex
C0019348|T047|SY|88594005|SNOMEDCT_CORE|Herpes simplex complex|Herpes simplex
C0019348|T047|SY|88594005|SNOMEDCT_CORE|Herpes simplex infection|Herpes simplex
C0019348|T047|SY|88594005|SNOMEDCT_CORE|Herpes simplex viral infection|Herpes simplex
C0019348|T047|IS|88594005|SNOMEDCT_CORE|Herpes simplex, NOS|Herpes simplex
C0019357|T047|PT|9389005|SNOMEDCT_CORE|Herpes simplex keratitis|Herpes simplex keratitis
C0019357|T047|FN|9389005|SNOMEDCT_CORE|Herpes simplex keratitis|Herpes simplex keratitis
C0019357|T047|SY|9389005|SNOMEDCT_CORE|Herpetic keratitis|Herpes simplex keratitis
C0019357|T047|SY|9389005|SNOMEDCT_CORE|HSV keratitis|Herpes simplex keratitis
C0019360|T047|PT|4740000|SNOMEDCT_CORE|Herpes zoster|Herpes zoster
C0019360|T047|FN|4740000|SNOMEDCT_CORE|Herpes zoster|Herpes zoster
C0019360|T047|SY|4740000|SNOMEDCT_CORE|Herpes zoster infection|Herpes zoster
C0019360|T047|IS|4740000|SNOMEDCT_CORE|Herpes zoster, NOS|Herpes zoster
C0019360|T047|SY|4740000|SNOMEDCT_CORE|Shingles|Herpes zoster
C0019360|T047|SY|4740000|SNOMEDCT_CORE|Zona|Herpes zoster
C0019360|T047|SY|4740000|SNOMEDCT_CORE|Zoster|Herpes zoster
C0019364|T047|PT|87513003|SNOMEDCT_CORE|Herpes zoster ophthalmicus|Herpes zoster ophthalmicus
C0019364|T047|FN|87513003|SNOMEDCT_CORE|Herpes zoster ophthalmicus|Herpes zoster ophthalmicus
C0019364|T047|SY|87513003|SNOMEDCT_CORE|Herpes zoster with ophthalmic complications|Herpes zoster ophthalmicus
C0019364|T047|SY|87513003|SNOMEDCT_CORE|Zoster ocular disease|Herpes zoster ophthalmicus
C0019364|T047|SY|87513003|SNOMEDCT_CORE|Zoster ophthalmicus|Herpes zoster ophthalmicus
C0019366|T047|IS|4740000|SNOMEDCT_CORE|Herpes zoster without mention of complication|Herpes zoster without mention of complication
C0019372|T047|SY|23513009|SNOMEDCT_CORE|Herpes infection|Herpesvirus infection
C0019372|T047|IS|23513009|SNOMEDCT_CORE|Herpes infection, NOS|Herpesvirus infection
C0019372|T047|PT|23513009|SNOMEDCT_CORE|Herpesvirus infection|Herpesvirus infection
C0019372|T047|FN|23513009|SNOMEDCT_CORE|Herpesvirus infection|Herpesvirus infection
C0019372|T047|IS|23513009|SNOMEDCT_CORE|Herpesvirus infection, NOS|Herpesvirus infection
C0019521|T033|SY|65958008|SNOMEDCT_CORE|Finding of hiccoughs|Hiccoughs
C0019521|T033|SY|65958008|SNOMEDCT_CORE|Hiccough|Hiccoughs
C0019521|T033|PT|65958008|SNOMEDCT_CORE|Hiccoughs|Hiccoughs
C0019521|T033|FN|65958008|SNOMEDCT_CORE|Hiccoughs|Hiccoughs
C0019521|T033|IS|65958008|SNOMEDCT_CORE|Hiccup|Hiccoughs
C0019521|T033|SY|65958008|SNOMEDCT_CORE|Hiccups|Hiccoughs
C0019521|T033|SY|65958008|SNOMEDCT_CORE|Observation of hiccoughs|Hiccoughs
C0019521|T033|SY|65958008|SNOMEDCT_CORE|Singultus|Hiccoughs
C0019555|T019|SY|48334007|SNOMEDCT_CORE|CDH - Congenital dislocation of the hip|Congenital dislocation of hip
C0019555|T019|PT|48334007|SNOMEDCT_CORE|Congenital dislocation of hip|Congenital dislocation of hip
C0019555|T019|FN|48334007|SNOMEDCT_CORE|Congenital dislocation of hip|Congenital dislocation of hip
C0019555|T019|IS|48334007|SNOMEDCT_CORE|Congenital dislocation of hip, NOS|Congenital dislocation of hip
C0019555|T019|SY|48334007|SNOMEDCT_CORE|Developmental dislocation of hip|Congenital dislocation of hip
C0019555|T019|SY|48334007|SNOMEDCT_CORE|Developmental displacement of the hip|Congenital dislocation of hip
C0019557|T037|SY|5913000|SNOMEDCT_CORE|Fracture of hip|Fracture of hip
C0019557|T037|IS|5913000|SNOMEDCT_CORE|Fracture of hip, NOS|Fracture of hip, NOS
C0019557|T037|SY|263225007|SNOMEDCT_CORE|Hip fracture|Hip fracture
C0019559|T184|SY|49218002|SNOMEDCT_CORE|Arthralgia of hip|Hip pain
C0019559|T184|IS|49218002|SNOMEDCT_CORE|Coxalgia|Hip pain
C0019559|T184|SY|49218002|SNOMEDCT_CORE|Hip joint pain|Hip pain
C0019559|T184|PT|49218002|SNOMEDCT_CORE|Hip pain|Hip pain
C0019559|T184|FN|49218002|SNOMEDCT_CORE|Hip pain|Hip pain
C0019562|T047|SY|46659004|SNOMEDCT_CORE|Cerebroretinal angiomatosis|Von Hippel-Lindau syndrome
C0019562|T047|SY|46659004|SNOMEDCT_CORE|Familial cerebello-retinal angiomatosis|Von Hippel-Lindau syndrome
C0019562|T047|SY|46659004|SNOMEDCT_CORE|Lindau' disease|Von Hippel-Lindau syndrome
C0019562|T047|SY|46659004|SNOMEDCT_CORE|Lindau's disease|Von Hippel-Lindau syndrome
C0019562|T047|SY|46659004|SNOMEDCT_CORE|VHL - von Hippel-Lindau syndrome|Von Hippel-Lindau syndrome
C0019562|T047|PT|46659004|SNOMEDCT_CORE|Von Hippel-Lindau syndrome|Von Hippel-Lindau syndrome
C0019562|T047|SY|46659004|SNOMEDCT_CORE|von Hippel-Lindau syndrome|Von Hippel-Lindau syndrome
C0019562|T047|FN|46659004|SNOMEDCT_CORE|Von Hippel-Lindau syndrome|Von Hippel-Lindau syndrome
C0019572|T033|SY|399939002|SNOMEDCT_CORE|Hirsutes|Hirsutism
C0019572|T033|SY|399939002|SNOMEDCT_CORE|Hirsuties|Hirsutism
C0019572|T033|PT|399939002|SNOMEDCT_CORE|Hirsutism|Hirsutism
C0019572|T033|FN|399939002|SNOMEDCT_CORE|Hirsutism|Hirsutism
C0019572|T033|SY|399939002|SNOMEDCT_CORE|Pilosis|Hirsutism
C0019621|T191|SY|65399007|SNOMEDCT_CORE|Differentiated progressive histiocytosis|Langerhans cell histiocytosis
C0019621|T191|SY|65399007|SNOMEDCT_CORE|Histiocytosis X|Langerhans cell histiocytosis
C0019621|T191|IS|65399007|SNOMEDCT_CORE|Histiocytosis X, NOS|Langerhans cell histiocytosis
C0019621|T191|SY|65399007|SNOMEDCT_CORE|Langerhan's cell histiocytosis|Langerhans cell histiocytosis
C0019621|T191|SY|65399007|SNOMEDCT_CORE|Langerhans cell disease|Langerhans cell histiocytosis
C0019621|T191|PT|65399007|SNOMEDCT_CORE|Langerhans cell histiocytosis|Langerhans cell histiocytosis
C0019621|T191|FN|65399007|SNOMEDCT_CORE|Langerhans cell histiocytosis|Langerhans cell histiocytosis
C0019621|T191|SY|65399007|SNOMEDCT_CORE|LCH - Langerhan's cell histiocytosis|Langerhans cell histiocytosis
C0019655|T047|PT|12962009|SNOMEDCT_CORE|Histoplasmosis|Histoplasmosis
C0019655|T047|FN|12962009|SNOMEDCT_CORE|Histoplasmosis|Histoplasmosis
C0019655|T047|IS|12962009|SNOMEDCT_CORE|Histoplasmosis, NOS|Histoplasmosis
C0019693|T047|SY|86406008|SNOMEDCT_CORE|HIV - Human immunodeficiency virus infection|Human immunodeficiency virus infection
C0019693|T047|SY|86406008|SNOMEDCT_CORE|HIV infection|Human immunodeficiency virus infection
C0019693|T047|PT|86406008|SNOMEDCT_CORE|Human immunodeficiency virus infection|Human immunodeficiency virus infection
C0019693|T047|FN|86406008|SNOMEDCT_CORE|Human immunodeficiency virus infection|Human immunodeficiency virus infection
C0019693|T047|IS|86406008|SNOMEDCT_CORE|Human immunodeficiency virus infection, NOS|Human immunodeficiency virus infection
C0019825|T184|SY|50219008|SNOMEDCT_CORE|Croaky voice|Hoarse
C0019825|T184|PT|50219008|SNOMEDCT_CORE|Hoarse|Hoarse
C0019825|T184|FN|50219008|SNOMEDCT_CORE|Hoarse|Hoarse
C0019825|T184|IS|50219008|SNOMEDCT_CORE|Hoarse voice quality|Hoarse
C0019825|T184|SY|50219008|SNOMEDCT_CORE|Hoarseness|Hoarse
C0019825|T184|SY|50219008|SNOMEDCT_CORE|Hoarseness - throat symptom|Hoarse
C0019825|T184|SY|50219008|SNOMEDCT_CORE|Hoarseness symptom|Hoarse
C0019825|T184|SY|50219008|SNOMEDCT_CORE|Husky voice|Hoarse
C0019825|T184|SY|50219008|SNOMEDCT_CORE|Voice hoarseness|Hoarse
C0019829|T191|SY|118599009|SNOMEDCT_CORE|HD - Hodgkin's disease|Hodgkin's disease
C0019829|T191|SY|118599009|SNOMEDCT_CORE|Hodgkin disease|Hodgkin's disease
C0019829|T191|SY|118599009|SNOMEDCT_CORE|Hodgkin's disease|Hodgkin's disease
C0019829|T191|PT|118599009|SNOMEDCT_CORE|Hodgkin's disease|Hodgkin's disease
C0019829|T191|FN|118599009|SNOMEDCT_CORE|Hodgkin's disease|Hodgkin's disease
C0019829|T191|SY|118599009|SNOMEDCT_CORE|Lymphoma, Hodgkins|Hodgkin's disease
C0019829|T191|SY|118599009|SNOMEDCT_CORE|Malignant Hodgkin's lymphoma|Hodgkin's disease
C0019917|T047|PT|397513003|SNOMEDCT_CORE|Hordeolum|Hordeolum
C0019917|T047|FN|397513003|SNOMEDCT_CORE|Hordeolum|Hordeolum
C0019937|T047|OAS|12731000|SNOMEDCT_CORE|Horner's syndrome|Horner's syndrome
C0020162|T037|PT|66308002|SNOMEDCT_CORE|Fracture of humerus|Fracture of humerus
C0020162|T037|FN|66308002|SNOMEDCT_CORE|Fracture of humerus|Fracture of humerus
C0020162|T037|IS|66308002|SNOMEDCT_CORE|Fracture of humerus, NOS|Fracture of humerus
C0020162|T037|SY|66308002|SNOMEDCT_CORE|Fracture of upper arm|Fracture of humerus
C0020162|T037|IS|66308002|SNOMEDCT_CORE|Fracture of upper arm, NOS|Fracture of humerus
C0020179|T047|SY|58756001|SNOMEDCT_CORE|Chronic progressive chorea|Huntington's chorea
C0020179|T047|SY|58756001|SNOMEDCT_CORE|Chronic progressive hereditary chorea|Huntington's chorea
C0020179|T047|SY|58756001|SNOMEDCT_CORE|HC - Huntington chorea|Huntington's chorea
C0020179|T047|SY|58756001|SNOMEDCT_CORE|HD - Huntington chorea|Huntington's chorea
C0020179|T047|SY|58756001|SNOMEDCT_CORE|Huntington chorea|Huntington's chorea
C0020179|T047|PT|58756001|SNOMEDCT_CORE|Huntington's chorea|Huntington's chorea
C0020179|T047|FN|58756001|SNOMEDCT_CORE|Huntington's chorea|Huntington's chorea
C0020192|T047|SY|46775006|SNOMEDCT_CORE|HMD - Hyaline membrane disease|HMD - Hyaline membrane disease
C0020192|T047|SY|46775006|SNOMEDCT_CORE|Hyaline membrane disease|HMD - Hyaline membrane disease
C0020217|T191|SY|417044008|SNOMEDCT_CORE|Hydatid mole|Hydatid mole
C0020217|T191|SY|417044008|SNOMEDCT_CORE|Hydatidiform mole|Hydatid mole
C0020217|T191|SY|417044008|SNOMEDCT_CORE|Molar pregnancy with hydatid mole|Hydatid mole
C0020217|T191|SY|417044008|SNOMEDCT_CORE|Molar pregnancy with vesicular mole|Hydatid mole
C0020224|T046|SY|86203003|SNOMEDCT_CORE|Excessive liquor|Polyhydramnios
C0020224|T046|SY|86203003|SNOMEDCT_CORE|Hydramnios|Polyhydramnios
C0020224|T046|PT|86203003|SNOMEDCT_CORE|Polyhydramnios|Polyhydramnios
C0020224|T046|FN|86203003|SNOMEDCT_CORE|Polyhydramnios|Polyhydramnios
C0020255|T047|PT|230745008|SNOMEDCT_CORE|Hydrocephalus|Hydrocephalus
C0020255|T047|FN|230745008|SNOMEDCT_CORE|Hydrocephalus|Hydrocephalus
C0020255|T047|SY|230745008|SNOMEDCT_CORE|Hydrocephaly|Hydrocephalus
C0020256|T019|SY|47032000|SNOMEDCT_CORE|Congenital dilatation of cerebral ventricles|Congenital hydrocephalus
C0020256|T019|SY|47032000|SNOMEDCT_CORE|Congenital hydrencephalus|Congenital hydrocephalus
C0020256|T019|SY|47032000|SNOMEDCT_CORE|Congenital hydrencephaly|Congenital hydrocephalus
C0020256|T019|PT|47032000|SNOMEDCT_CORE|Congenital hydrocephalus|Congenital hydrocephalus
C0020256|T019|FN|47032000|SNOMEDCT_CORE|Congenital hydrocephalus|Congenital hydrocephalus
C0020256|T019|SY|47032000|SNOMEDCT_CORE|Congenital hydrocephaly|Congenital hydrocephalus
C0020256|T019|SY|47032000|SNOMEDCT_CORE|Hydrocephalus in newborn|Congenital hydrocephalus
C0020256|T019|SY|47032000|SNOMEDCT_CORE|Primary hydrocephalus|Congenital hydrocephalus
C0020256|T019|SY|47032000|SNOMEDCT_CORE|Primary hydrocephaly|Congenital hydrocephalus
C0020258|T047|SY|30753002|SNOMEDCT_CORE|Low pressure hydrocephalus|Normal pressure hydrocephalus
C0020258|T047|PT|30753002|SNOMEDCT_CORE|Normal pressure hydrocephalus|Normal pressure hydrocephalus
C0020258|T047|FN|30753002|SNOMEDCT_CORE|Normal pressure hydrocephalus|Normal pressure hydrocephalus
C0020258|T047|SY|30753002|SNOMEDCT_CORE|NPH - Normal pressure hydrocephalus|Normal pressure hydrocephalus
C0020295|T047|PT|43064006|SNOMEDCT_CORE|Hydronephrosis|Hydronephrosis
C0020295|T047|FN|43064006|SNOMEDCT_CORE|Hydronephrosis|Hydronephrosis
C0020433|T047|SYGB|14783006|SNOMEDCT_CORE|Bilirubinaemia|Hyperbilirubinemia
C0020433|T047|SY|14783006|SNOMEDCT_CORE|Bilirubinemia|Hyperbilirubinemia
C0020433|T047|PTGB|14783006|SNOMEDCT_CORE|Hyperbilirubinaemia|Hyperbilirubinemia
C0020433|T047|PT|14783006|SNOMEDCT_CORE|Hyperbilirubinemia|Hyperbilirubinemia
C0020433|T047|FN|14783006|SNOMEDCT_CORE|Hyperbilirubinemia|Hyperbilirubinemia
C0020433|T047|IS|14783006|SNOMEDCT_CORE|Hyperbilirubinemia, NOS|Hyperbilirubinemia
C0020437|T047|PTGB|66931009|SNOMEDCT_CORE|Hypercalcaemia|Hypercalcemia
C0020437|T047|SYGB|66931009|SNOMEDCT_CORE|Hypercalcaemia syndrome|Hypercalcemia
C0020437|T047|PT|66931009|SNOMEDCT_CORE|Hypercalcemia|Hypercalcemia
C0020437|T047|FN|66931009|SNOMEDCT_CORE|Hypercalcemia|Hypercalcemia
C0020437|T047|SY|66931009|SNOMEDCT_CORE|Hypercalcemia syndrome|Hypercalcemia
C0020437|T047|PT|166702002|SNOMEDCT_CORE|Raised serum calcium level|Hypercalcemia
C0020437|T047|FN|166702002|SNOMEDCT_CORE|Raised serum calcium level|Hypercalcemia
C0020438|T033|PT|71938000|SNOMEDCT_CORE|Hypercalciuria|Hypercalciuria
C0020438|T033|FN|71938000|SNOMEDCT_CORE|Hypercalciuria|Hypercalciuria
C0020438|T033|SY|71938000|SNOMEDCT_CORE|Hypercalcuria|Hypercalciuria
C0020443|T047|SY|13644009|SNOMEDCT_CORE|High cholesterol|Hypercholesterolemia
C0020443|T047|PTGB|13644009|SNOMEDCT_CORE|Hypercholesterolaemia|Hypercholesterolemia
C0020443|T047|IS|13644009|SNOMEDCT_CORE|Hypercholesterolaemia, NOS|Hypercholesterolemia
C0020443|T047|PT|13644009|SNOMEDCT_CORE|Hypercholesterolemia|Hypercholesterolemia
C0020443|T047|FN|13644009|SNOMEDCT_CORE|Hypercholesterolemia|Hypercholesterolemia
C0020443|T047|IS|13644009|SNOMEDCT_CORE|Hypercholesterolemia, NOS|Hypercholesterolemia
C0020445|T047|SYGB|398036000|SNOMEDCT_CORE|Essential familial hypercholesterolaemia|Familial hypercholesterolemia
C0020445|T047|SY|398036000|SNOMEDCT_CORE|Essential familial hypercholesterolemia|Familial hypercholesterolemia
C0020445|T047|SYGB|398036000|SNOMEDCT_CORE|Familial hyperbetalipoproteinaemia|Familial hypercholesterolemia
C0020445|T047|SY|398036000|SNOMEDCT_CORE|Familial hyperbetalipoproteinemia|Familial hypercholesterolemia
C0020445|T047|PTGB|398036000|SNOMEDCT_CORE|Familial hypercholesterolaemia|Familial hypercholesterolemia
C0020445|T047|PT|398036000|SNOMEDCT_CORE|Familial hypercholesterolemia|Familial hypercholesterolemia
C0020445|T047|FN|398036000|SNOMEDCT_CORE|Familial hypercholesterolemia|Familial hypercholesterolemia
C0020445|T047|SY|398036000|SNOMEDCT_CORE|LDL - Low density lipoprotein receptor disorder|Familial hypercholesterolemia
C0020445|T047|SY|398036000|SNOMEDCT_CORE|LDL receptor disorder|Familial hypercholesterolemia
C0020445|T047|SY|398036000|SNOMEDCT_CORE|Low density lipoprotein catabolic defect|Familial hypercholesterolemia
C0020450|T184|SY|14094001|SNOMEDCT_CORE|Excessive pregnancy vomiting|Hyperemesis gravidarum
C0020450|T184|SY|14094001|SNOMEDCT_CORE|Excessive vomiting in pregnancy|Hyperemesis gravidarum
C0020450|T184|FN|14094001|SNOMEDCT_CORE|Excessive vomiting in pregnancy|Hyperemesis gravidarum
C0020450|T184|SY|14094001|SNOMEDCT_CORE|Hyperemesis arising during pregnancy|Hyperemesis gravidarum
C0020450|T184|PT|14094001|SNOMEDCT_CORE|Hyperemesis gravidarum|Hyperemesis gravidarum
C0020450|T184|SY|14094001|SNOMEDCT_CORE|Hyperemesis in pregnancy|Hyperemesis gravidarum
C0020450|T184|SY|14094001|SNOMEDCT_CORE|Hyperemesis of pregnancy|Hyperemesis gravidarum
C0020450|T184|SY|14094001|SNOMEDCT_CORE|Persistent AND/OR vicious vomiting arising during pregnancy|Hyperemesis gravidarum
C0020450|T184|IS|14094001|SNOMEDCT_CORE|Persistent or vicious vomiting arising during pregnancy|Hyperemesis gravidarum
C0020452|T047|IS|247441003|SNOMEDCT_CORE|Hyperaemia|Hyperemia
C0020452|T047|IS|247441003|SNOMEDCT_CORE|Hyperemia|Hyperemia
C0020456|T047|PTGB|80394007|SNOMEDCT_CORE|Hyperglycaemia|Hyperglycemia
C0020456|T047|IS|80394007|SNOMEDCT_CORE|Hyperglycaemia, NOS|Hyperglycemia
C0020456|T047|PT|80394007|SNOMEDCT_CORE|Hyperglycemia|Hyperglycemia
C0020456|T047|FN|80394007|SNOMEDCT_CORE|Hyperglycemia|Hyperglycemia
C0020456|T047|IS|80394007|SNOMEDCT_CORE|Hyperglycemia, NOS|Hyperglycemia
C0020458|T033|FN|312230002|SNOMEDCT_CORE|Hyperhidrosis|Hyperhidrosis
C0020458|T033|IS|52613005|SNOMEDCT_CORE|Hyperhidrosis|Hyperhidrosis
C0020458|T033|PT|312230002|SNOMEDCT_CORE|Hyperhidrosis|Hyperhidrosis
C0020458|T033|IS|312230002|SNOMEDCT_CORE|Hyperhydrosis disorder|Hyperhidrosis
C0020458|T033|OF|312230002|SNOMEDCT_CORE|Hyperhydrosis disorder|Hyperhidrosis
C0020459|T047|SYGB|83469008|SNOMEDCT_CORE|Hyperinsulinaemia|Hyperinsulinism
C0020459|T047|SY|83469008|SNOMEDCT_CORE|Hyperinsulinemia|Hyperinsulinism
C0020459|T047|PT|83469008|SNOMEDCT_CORE|Hyperinsulinism|Hyperinsulinism
C0020459|T047|FN|83469008|SNOMEDCT_CORE|Hyperinsulinism|Hyperinsulinism
C0020459|T047|IS|83469008|SNOMEDCT_CORE|Hyperinsulinism, NOS|Hyperinsulinism
C0020461|T033|PTGB|14140009|SNOMEDCT_CORE|Hyperkalaemia|Hyperkalemia
C0020461|T033|SYGB|14140009|SNOMEDCT_CORE|Hyperkalaemic syndrome|Hyperkalemia
C0020461|T033|PT|14140009|SNOMEDCT_CORE|Hyperkalemia|Hyperkalemia
C0020461|T033|FN|14140009|SNOMEDCT_CORE|Hyperkalemia|Hyperkalemia
C0020461|T033|SY|14140009|SNOMEDCT_CORE|Hyperkalemic syndrome|Hyperkalemia
C0020461|T033|SYGB|14140009|SNOMEDCT_CORE|Hyperpotassaemia|Hyperkalemia
C0020461|T033|SY|14140009|SNOMEDCT_CORE|Hyperpotassemia|Hyperkalemia
C0020461|T033|SY|14140009|SNOMEDCT_CORE|K excess|Hyperkalemia
C0020461|T033|SY|14140009|SNOMEDCT_CORE|K overload|Hyperkalemia
C0020461|T033|SY|14140009|SNOMEDCT_CORE|Potassium excess|Hyperkalemia
C0020473|T047|SYGB|55822004|SNOMEDCT_CORE|HLD - Hyperlipidaemia|Hyperlipidemia
C0020473|T047|SY|55822004|SNOMEDCT_CORE|HLD - Hyperlipidemia|Hyperlipidemia
C0020473|T047|PTGB|55822004|SNOMEDCT_CORE|Hyperlipidaemia|Hyperlipidemia
C0020473|T047|IS|55822004|SNOMEDCT_CORE|Hyperlipidaemia, NOS|Hyperlipidemia
C0020473|T047|PT|55822004|SNOMEDCT_CORE|Hyperlipidemia|Hyperlipidemia
C0020473|T047|FN|55822004|SNOMEDCT_CORE|Hyperlipidemia|Hyperlipidemia
C0020473|T047|IS|55822004|SNOMEDCT_CORE|Hyperlipidemia, NOS|Hyperlipidemia
C0020473|T047|SYGB|55822004|SNOMEDCT_CORE|Lipidaemia|Hyperlipidemia
C0020473|T047|SY|55822004|SNOMEDCT_CORE|Lipidemia|Hyperlipidemia
C0020474|T047|PTGB|238040008|SNOMEDCT_CORE|Familial combined hyperlipidaemia|Familial combined hyperlipidemia
C0020474|T047|PT|238040008|SNOMEDCT_CORE|Familial combined hyperlipidemia|Familial combined hyperlipidemia
C0020474|T047|FN|238040008|SNOMEDCT_CORE|Familial combined hyperlipidemia|Familial combined hyperlipidemia
C0020476|T047|PTGB|3744001|SNOMEDCT_CORE|Hyperlipoproteinaemia|Hyperlipoproteinemia
C0020476|T047|IS|3744001|SNOMEDCT_CORE|Hyperlipoproteinaemia, NOS|Hyperlipoproteinemia
C0020476|T047|PT|3744001|SNOMEDCT_CORE|Hyperlipoproteinemia|Hyperlipoproteinemia
C0020476|T047|FN|3744001|SNOMEDCT_CORE|Hyperlipoproteinemia|Hyperlipoproteinemia
C0020476|T047|IS|3744001|SNOMEDCT_CORE|Hyperlipoproteinemia, NOS|Hyperlipoproteinemia
C0020480|T047|PTGB|238085009|SNOMEDCT_CORE|Fredrickson type IV hyperlipoproteinaemia|Pure hyperglyceridemia
C0020480|T047|PT|238085009|SNOMEDCT_CORE|Fredrickson type IV hyperlipoproteinemia|Pure hyperglyceridemia
C0020480|T047|FN|238085009|SNOMEDCT_CORE|Fredrickson type IV hyperlipoproteinemia|Pure hyperglyceridemia
C0020480|T047|SYGB|238085009|SNOMEDCT_CORE|Fredrickson type IV lipidaemia|Pure hyperglyceridemia
C0020480|T047|SY|238085009|SNOMEDCT_CORE|Fredrickson type IV lipidemia|Pure hyperglyceridemia
C0020480|T047|PTGB|267433009|SNOMEDCT_CORE|Pure hyperglyceridaemia|Pure hyperglyceridemia
C0020480|T047|PT|267433009|SNOMEDCT_CORE|Pure hyperglyceridemia|Pure hyperglyceridemia
C0020480|T047|FN|267433009|SNOMEDCT_CORE|Pure hyperglyceridemia|Pure hyperglyceridemia
C0020488|T047|OAP|39355002|SNOMEDCT_CORE|Hypernatraemia|Hypernatremia
C0020488|T047|PTGB|771115008|SNOMEDCT_CORE|Hypernatraemia|Hypernatremia
C0020488|T047|IS|39355002|SNOMEDCT_CORE|Hypernatraemia, NOS|Hypernatremia
C0020488|T047|PT|771115008|SNOMEDCT_CORE|Hypernatremia|Hypernatremia
C0020488|T047|OAP|39355002|SNOMEDCT_CORE|Hypernatremia|Hypernatremia
C0020488|T047|OAF|39355002|SNOMEDCT_CORE|Hypernatremia|Hypernatremia
C0020488|T047|FN|771115008|SNOMEDCT_CORE|Hypernatremia|Hypernatremia
C0020488|T047|IS|39355002|SNOMEDCT_CORE|Hypernatremia, NOS|Hypernatremia
C0020488|T047|OAS|39355002|SNOMEDCT_CORE|Na excess|Hypernatremia
C0020488|T047|SY|771115008|SNOMEDCT_CORE|Na excess|Hypernatremia
C0020488|T047|OAS|39355002|SNOMEDCT_CORE|Na overload|Hypernatremia
C0020488|T047|SY|771115008|SNOMEDCT_CORE|Na overload|Hypernatremia
C0020488|T047|OAS|39355002|SNOMEDCT_CORE|Sodium overload|Hypernatremia
C0020488|T047|SY|771115008|SNOMEDCT_CORE|Sodium overload|Hypernatremia
C0020488|T047|OAS|39355002|SNOMEDCT_CORE|Sodium retention|Hypernatremia
C0020490|T047|SY|38101003|SNOMEDCT_CORE|Farsightedness|Hypermetropia
C0020490|T047|PT|38101003|SNOMEDCT_CORE|Hypermetropia|Hypermetropia
C0020490|T047|FN|38101003|SNOMEDCT_CORE|Hypermetropia|Hypermetropia
C0020490|T047|SY|38101003|SNOMEDCT_CORE|Hyperopia|Hypermetropia
C0020490|T047|SY|38101003|SNOMEDCT_CORE|Longsighted|Hypermetropia
C0020490|T047|SY|38101003|SNOMEDCT_CORE|Longsightedness|Hypermetropia
C0020498|T047|SY|31487001|SNOMEDCT_CORE|Ankylosing hyperostosis|Disseminated idiopathic skeletal hyperostosis
C0020498|T047|IS|31487001|SNOMEDCT_CORE|Ankylosing vertebral hyperostosis|Disseminated idiopathic skeletal hyperostosis
C0020498|T047|SY|31487001|SNOMEDCT_CORE|Diffuse idiopathic skeletal hyperostosis|Disseminated idiopathic skeletal hyperostosis
C0020498|T047|IS|31487001|SNOMEDCT_CORE|DISH|Disseminated idiopathic skeletal hyperostosis
C0020498|T047|SY|31487001|SNOMEDCT_CORE|DISH - Diffuse idiopathic skeletal hyperostosis|Disseminated idiopathic skeletal hyperostosis
C0020498|T047|PT|31487001|SNOMEDCT_CORE|Disseminated idiopathic skeletal hyperostosis|Disseminated idiopathic skeletal hyperostosis
C0020498|T047|FN|31487001|SNOMEDCT_CORE|Disseminated idiopathic skeletal hyperostosis|Disseminated idiopathic skeletal hyperostosis
C0020498|T047|SY|31487001|SNOMEDCT_CORE|Forestier's disease|Disseminated idiopathic skeletal hyperostosis
C0020501|T047|PT|17901006|SNOMEDCT_CORE|Primary hyperoxaluria|Primary hyperoxaluria
C0020501|T047|FN|17901006|SNOMEDCT_CORE|Primary hyperoxaluria|Primary hyperoxaluria
C0020501|T047|IS|17901006|SNOMEDCT_CORE|Primary hyperoxaluria, NOS|Primary hyperoxaluria
C0020501|T047|SY|17901006|SNOMEDCT_CORE|Primary oxalosis|Primary hyperoxaluria
C0020501|T047|IS|17901006|SNOMEDCT_CORE|Primary oxalosis, NOS|Primary hyperoxaluria
C0020502|T047|SY|66999008|SNOMEDCT_CORE|HPTH - Hyperparathyroidism|Hyperparathyroidism
C0020502|T047|PT|66999008|SNOMEDCT_CORE|Hyperparathyroidism|Hyperparathyroidism
C0020502|T047|FN|66999008|SNOMEDCT_CORE|Hyperparathyroidism|Hyperparathyroidism
C0020502|T047|IS|66999008|SNOMEDCT_CORE|Hyperparathyroidism, NOS|Hyperparathyroidism
C0020503|T047|PT|91478007|SNOMEDCT_CORE|Secondary hyperparathyroidism|Secondary hyperparathyroidism
C0020503|T047|FN|91478007|SNOMEDCT_CORE|Secondary hyperparathyroidism|Secondary hyperparathyroidism
C0020503|T047|IS|91478007|SNOMEDCT_CORE|Secondary hyperparathyroidism, NOS|Secondary hyperparathyroidism
C0020505|T033|IS|267023007|SNOMEDCT_CORE|:: Polyphagia|Excessive eating - polyphagia
C0020505|T033|SY|267023007|SNOMEDCT_CORE|Excessive eating|Excessive eating - polyphagia
C0020505|T033|PT|267023007|SNOMEDCT_CORE|Excessive eating - polyphagia|Excessive eating - polyphagia
C0020505|T033|FN|267023007|SNOMEDCT_CORE|Excessive eating - polyphagia|Excessive eating - polyphagia
C0020505|T033|SY|267023007|SNOMEDCT_CORE|Gluttony|Excessive eating - polyphagia
C0020505|T033|SY|267023007|SNOMEDCT_CORE|Hyperphagia|Excessive eating - polyphagia
C0020505|T033|SY|267023007|SNOMEDCT_CORE|Polyphagia|Excessive eating - polyphagia
C0020514|T047|PTGB|237662005|SNOMEDCT_CORE|Hyperprolactinaemia|Hyperprolactinemia
C0020514|T047|PT|237662005|SNOMEDCT_CORE|Hyperprolactinemia|Hyperprolactinemia
C0020514|T047|FN|237662005|SNOMEDCT_CORE|Hyperprolactinemia|Hyperprolactinemia
C0020517|T046|OAS|106190000|SNOMEDCT_CORE|Allergic state|Hypersensitivity reaction
C0020517|T046|OAF|106190000|SNOMEDCT_CORE|Allergic state|Hypersensitivity reaction
C0020517|T046|OAP|106190000|SNOMEDCT_CORE|Allergy|Hypersensitivity reaction
C0020517|T046|OF|106190000|SNOMEDCT_CORE|Allergy|Hypersensitivity reaction
C0020517|T046|OAS|106190000|SNOMEDCT_CORE|Atopic AND/OR hypersensitivity state|Hypersensitivity reaction
C0020517|T046|PT|421961002|SNOMEDCT_CORE|Hypersensitivity reaction|Hypersensitivity reaction
C0020517|T046|FN|421961002|SNOMEDCT_CORE|Hypersensitivity reaction|Hypersensitivity reaction
C0020530|T184|PT|79280005|SNOMEDCT_CORE|Hypersomnia with sleep apnea|Hypersomnia with sleep apnea
C0020530|T184|FN|79280005|SNOMEDCT_CORE|Hypersomnia with sleep apnea|Hypersomnia with sleep apnea
C0020530|T184|PTGB|79280005|SNOMEDCT_CORE|Hypersomnia with sleep apnoea|Hypersomnia with sleep apnea
C0020532|T047|SY|58381000|SNOMEDCT_CORE|Big spleen syndrome|Hypersplenism
C0020532|T047|SY|58381000|SNOMEDCT_CORE|Hypersplenia|Hypersplenism
C0020532|T047|PT|58381000|SNOMEDCT_CORE|Hypersplenism|Hypersplenism
C0020532|T047|FN|58381000|SNOMEDCT_CORE|Hypersplenism|Hypersplenism
C0020532|T047|IS|58381000|SNOMEDCT_CORE|Hypersplenism, NOS|Hypersplenism
C0020538|T047|SY|38341003|SNOMEDCT_CORE|BP - High blood pressure|Hypertensive disorder
C0020538|T047|SY|38341003|SNOMEDCT_CORE|BP+ - Hypertension|Hypertensive disorder
C0020538|T047|SY|38341003|SNOMEDCT_CORE|HBP - High blood pressure|Hypertensive disorder
C0020538|T047|SY|38341003|SNOMEDCT_CORE|High blood pressure|Hypertensive disorder
C0020538|T047|SY|38341003|SNOMEDCT_CORE|High blood pressure disorder|Hypertensive disorder
C0020538|T047|SY|38341003|SNOMEDCT_CORE|HT - Hypertension|Hypertensive disorder
C0020538|T047|SY|38341003|SNOMEDCT_CORE|HTN - Hypertension|Hypertensive disorder
C0020538|T047|IS|38341003|SNOMEDCT_CORE|Hyperpiesia|Hypertensive disorder
C0020538|T047|IS|38341003|SNOMEDCT_CORE|Hyperpiesis|Hypertensive disorder
C0020538|T047|SY|38341003|SNOMEDCT_CORE|Hypertension|Hypertensive disorder
C0020538|T047|IS|38341003|SNOMEDCT_CORE|Hypertension, NOS|Hypertensive disorder
C0020538|T047|IS|38341003|SNOMEDCT_CORE|Hypertensive disease|Hypertensive disorder
C0020538|T047|IS|38341003|SNOMEDCT_CORE|Hypertensive disease, NOS|Hypertensive disorder
C0020538|T047|PT|38341003|SNOMEDCT_CORE|Hypertensive disorder|Hypertensive disorder
C0020538|T047|FN|38341003|SNOMEDCT_CORE|Hypertensive disorder, systemic arterial|Hypertensive disorder
C0020538|T047|SY|38341003|SNOMEDCT_CORE|Hypertensive disorder, systemic arterial|Hypertensive disorder
C0020538|T047|SY|38341003|SNOMEDCT_CORE|Hypertensive vascular degeneration|Hypertensive disorder
C0020538|T047|SY|38341003|SNOMEDCT_CORE|Hypertensive vascular disease|Hypertensive disorder
C0020538|T047|OF|38341003|SNOMEDCT_CORE|Raised blood pressure|Hypertensive disorder
C0020538|T047|SY|38341003|SNOMEDCT_CORE|Systemic arterial hypertension|Hypertensive disorder
C0020540|T047|PT|70272006|SNOMEDCT_CORE|Malignant hypertension|Malignant hypertension
C0020540|T047|FN|70272006|SNOMEDCT_CORE|Malignant hypertension|Malignant hypertension
C0020541|T047|SY|34742003|SNOMEDCT_CORE|PHT - Portal hypertension|Portal hypertension
C0020541|T047|PT|34742003|SNOMEDCT_CORE|Portal hypertension|Portal hypertension
C0020541|T047|FN|34742003|SNOMEDCT_CORE|Portal hypertension|Portal hypertension
C0020542|T046|SY|70995007|SNOMEDCT_CORE|PHT - Pulmonary hypertension|Pulmonary hypertension
C0020542|T046|PT|70995007|SNOMEDCT_CORE|Pulmonary hypertension|Pulmonary hypertension
C0020542|T046|FN|70995007|SNOMEDCT_CORE|Pulmonary hypertension|Pulmonary hypertension
C0020542|T046|IS|70995007|SNOMEDCT_CORE|Pulmonary hypertension, NOS|Pulmonary hypertension
C0020544|T047|PT|28119000|SNOMEDCT_CORE|Renal hypertension|Renal hypertension
C0020544|T047|FN|28119000|SNOMEDCT_CORE|Renal hypertension|Renal hypertension
C0020545|T047|SY|123799005|SNOMEDCT_CORE|Hypertension due to renovascular disease|Renovascular hypertension
C0020545|T047|PT|123799005|SNOMEDCT_CORE|Renovascular hypertension|Renovascular hypertension
C0020545|T047|FN|123799005|SNOMEDCT_CORE|Renovascular hypertension|Renovascular hypertension
C0020550|T047|PT|34486009|SNOMEDCT_CORE|Hyperthyroidism|Hyperthyroidism
C0020550|T047|FN|34486009|SNOMEDCT_CORE|Hyperthyroidism|Hyperthyroidism
C0020550|T047|IS|34486009|SNOMEDCT_CORE|Hyperthyroidism, NOS|Hyperthyroidism
C0020557|T047|PTGB|302870006|SNOMEDCT_CORE|Hypertriglyceridaemia|Hypertriglyceridemia
C0020557|T047|PT|302870006|SNOMEDCT_CORE|Hypertriglyceridemia|Hypertriglyceridemia
C0020557|T047|FN|302870006|SNOMEDCT_CORE|Hypertriglyceridemia|Hypertriglyceridemia
C0020565|T046|PT|372281005|SNOMEDCT_CORE|Hypertrophy of breast|Hypertrophy of breast
C0020565|T046|FN|372281005|SNOMEDCT_CORE|Hypertrophy of breast|Hypertrophy of breast
C0020575|T047|PT|40608009|SNOMEDCT_CORE|Hypertropia|Hypertropia
C0020575|T047|FN|40608009|SNOMEDCT_CORE|Hypertropia|Hypertropia
C0020578|T033|SY|68978004|SNOMEDCT_CORE|HV - Hyperventilation|Hyperventilation
C0020578|T033|SY|68978004|SNOMEDCT_CORE|Hyperventilating|Hyperventilation
C0020578|T033|PT|68978004|SNOMEDCT_CORE|Hyperventilation|Hyperventilation
C0020578|T033|FN|68978004|SNOMEDCT_CORE|Hyperventilation|Hyperventilation
C0020578|T033|IS|68978004|SNOMEDCT_CORE|Hyperventilation, NOS|Hyperventilation
C0020578|T033|SY|68978004|SNOMEDCT_CORE|Overbreathing|Hyperventilation
C0020580|T033|PT|397974008|SNOMEDCT_CORE|Hypesthesia|Hypesthesia
C0020580|T033|FN|397974008|SNOMEDCT_CORE|Hypesthesia|Hypesthesia
C0020580|T033|SYGB|397974008|SNOMEDCT_CORE|Hypoaesthesia|Hypesthesia
C0020580|T033|PTGB|397974008|SNOMEDCT_CORE|Hypoesthesia|Hypesthesia
C0020580|T033|SY|397974008|SNOMEDCT_CORE|Hypoesthesia|Hypesthesia
C0020580|T033|SY|397974008|SNOMEDCT_CORE|Impaired sensation|Hypesthesia
C0020580|T033|SY|397974008|SNOMEDCT_CORE|Limited sensation|Hypesthesia
C0020580|T033|SY|397974008|SNOMEDCT_CORE|Reduced sensation|Hypesthesia
C0020581|T046|SY|75229002|SNOMEDCT_CORE|Blood in anterior chamber|Hyphema
C0020581|T046|PTGB|75229002|SNOMEDCT_CORE|Hyphaema|Hyphema
C0020581|T046|SYGB|75229002|SNOMEDCT_CORE|Hyphaemia|Hyphema
C0020581|T046|PT|75229002|SNOMEDCT_CORE|Hyphema|Hyphema
C0020581|T046|FN|75229002|SNOMEDCT_CORE|Hyphema|Hyphema
C0020581|T046|SY|75229002|SNOMEDCT_CORE|Hyphemia|Hyphema
C0020598|T047|SY|5291005|SNOMEDCT_CORE|Calcium deficiency disease|Hypocalcemia
C0020598|T047|PTGB|5291005|SNOMEDCT_CORE|Hypocalcaemia|Hypocalcemia
C0020598|T047|SYGB|5291005|SNOMEDCT_CORE|Hypocalcaemia syndrome|Hypocalcemia
C0020598|T047|PT|5291005|SNOMEDCT_CORE|Hypocalcemia|Hypocalcemia
C0020598|T047|FN|5291005|SNOMEDCT_CORE|Hypocalcemia|Hypocalcemia
C0020598|T047|SY|5291005|SNOMEDCT_CORE|Hypocalcemia syndrome|Hypocalcemia
C0020604|T048|SY|18193002|SNOMEDCT_CORE|Hypochondria|Hypochondriasis
C0020604|T048|SY|18193002|SNOMEDCT_CORE|Hypochondriacal neurosis|Hypochondriasis
C0020604|T048|PT|18193002|SNOMEDCT_CORE|Hypochondriasis|Hypochondriasis
C0020604|T048|FN|18193002|SNOMEDCT_CORE|Hypochondriasis|Hypochondriasis
C0020615|T047|PTGB|302866003|SNOMEDCT_CORE|Hypoglycaemia|Hypoglycemia
C0020615|T047|PT|302866003|SNOMEDCT_CORE|Hypoglycemia|Hypoglycemia
C0020615|T047|FN|302866003|SNOMEDCT_CORE|Hypoglycemia|Hypoglycemia
C0020619|T047|PT|48130008|SNOMEDCT_CORE|Hypogonadism|Hypogonadism
C0020619|T047|FN|48130008|SNOMEDCT_CORE|Hypogonadism|Hypogonadism
C0020619|T047|IS|48130008|SNOMEDCT_CORE|Hypogonadism, NOS|Hypogonadism
C0020621|T033|PTGB|43339004|SNOMEDCT_CORE|Hypokalaemia|Hypokalemia
C0020621|T033|SYGB|43339004|SNOMEDCT_CORE|Hypokalaemic syndrome|Hypokalemia
C0020621|T033|PT|43339004|SNOMEDCT_CORE|Hypokalemia|Hypokalemia
C0020621|T033|FN|43339004|SNOMEDCT_CORE|Hypokalemia|Hypokalemia
C0020621|T033|SY|43339004|SNOMEDCT_CORE|Hypokalemic syndrome|Hypokalemia
C0020621|T033|SYGB|43339004|SNOMEDCT_CORE|Hypopotassaemia|Hypokalemia
C0020621|T033|SYGB|43339004|SNOMEDCT_CORE|Hypopotassaemia syndrome|Hypokalemia
C0020621|T033|SY|43339004|SNOMEDCT_CORE|Hypopotassemia|Hypokalemia
C0020621|T033|SY|43339004|SNOMEDCT_CORE|Hypopotassemia syndrome|Hypokalemia
C0020625|T047|PTGB|89627008|SNOMEDCT_CORE|Hyponatraemia|Hyponatremia
C0020625|T047|IS|89627008|SNOMEDCT_CORE|Hyponatraemia, NOS|Hyponatremia
C0020625|T047|PT|89627008|SNOMEDCT_CORE|Hyponatremia|Hyponatremia
C0020625|T047|FN|89627008|SNOMEDCT_CORE|Hyponatremia|Hyponatremia
C0020625|T047|IS|89627008|SNOMEDCT_CORE|Hyponatremia, NOS|Hyponatremia
C0020626|T047|SY|36976004|SNOMEDCT_CORE|Deficiency of parathyrin|Hypoparathyroidism
C0020626|T047|SY|36976004|SNOMEDCT_CORE|Deficiency of parathyroid hormone|Hypoparathyroidism
C0020626|T047|SY|36976004|SNOMEDCT_CORE|Deficiency of PTH|Hypoparathyroidism
C0020626|T047|PT|36976004|SNOMEDCT_CORE|Hypoparathyroidism|Hypoparathyroidism
C0020626|T047|FN|36976004|SNOMEDCT_CORE|Hypoparathyroidism|Hypoparathyroidism
C0020626|T047|IS|36976004|SNOMEDCT_CORE|Hypoparathyroidism, NOS|Hypoparathyroidism
C0020635|T047|SY|74728003|SNOMEDCT_CORE|Deficient secretion of one OR more pituitary hormones|Hypopituitarism
C0020635|T047|IS|74728003|SNOMEDCT_CORE|Deficient secretion of one or more pituitary hormones|Hypopituitarism
C0020635|T047|PT|74728003|SNOMEDCT_CORE|Hypopituitarism|Hypopituitarism
C0020635|T047|FN|74728003|SNOMEDCT_CORE|Hypopituitarism|Hypopituitarism
C0020635|T047|IS|74728003|SNOMEDCT_CORE|Hypopituitarism, NOS|Hypopituitarism
C0020635|T047|SY|74728003|SNOMEDCT_CORE|Pituitary deficiency|Hypopituitarism
C0020635|T047|SY|74728003|SNOMEDCT_CORE|Pituitary failure|Hypopituitarism
C0020635|T047|SY|74728003|SNOMEDCT_CORE|Pituitary hypofunction|Hypopituitarism
C0020635|T047|SY|74728003|SNOMEDCT_CORE|Pituitary insufficiency|Hypopituitarism
C0020635|T047|IS|74728003|SNOMEDCT_CORE|Pituitary insufficiency, NOS|Hypopituitarism
C0020639|T047|PTGB|8900005|SNOMEDCT_CORE|Hypoproteinaemia|Hypoproteinemia
C0020639|T047|IS|8900005|SNOMEDCT_CORE|Hypoproteinaemia, NOS|Hypoproteinemia
C0020639|T047|PT|8900005|SNOMEDCT_CORE|Hypoproteinemia|Hypoproteinemia
C0020639|T047|FN|8900005|SNOMEDCT_CORE|Hypoproteinemia|Hypoproteinemia
C0020639|T047|IS|8900005|SNOMEDCT_CORE|Hypoproteinemia, NOS|Hypoproteinemia
C0020645|T033|PTGB|267447008|SNOMEDCT_CORE|Hypo-osmolality and or hyponatraemia|Hypo-osmolality and or hyponatremia
C0020645|T033|PT|267447008|SNOMEDCT_CORE|Hypo-osmolality and or hyponatremia|Hypo-osmolality and or hyponatremia
C0020645|T033|FN|267447008|SNOMEDCT_CORE|Hypo-osmolality and or hyponatremia|Hypo-osmolality and or hyponatremia
C0020649|T033|SY|45007003|SNOMEDCT_CORE|Arterial hypotension|Low blood pressure
C0020649|T033|IS|45007003|SNOMEDCT_CORE|Arterial hypotension, NOS|Low blood pressure
C0020649|T033|SY|45007003|SNOMEDCT_CORE|Hypopiesis|Low blood pressure
C0020649|T033|SY|45007003|SNOMEDCT_CORE|Hypotension|Low blood pressure
C0020649|T033|IS|45007003|SNOMEDCT_CORE|Hypotension, NOS|Low blood pressure
C0020649|T033|PT|45007003|SNOMEDCT_CORE|Low blood pressure|Low blood pressure
C0020649|T033|FN|45007003|SNOMEDCT_CORE|Low blood pressure|Low blood pressure
C0020651|T047|PT|28651003|SNOMEDCT_CORE|Orthostatic hypotension|Orthostatic hypotension
C0020651|T047|FN|28651003|SNOMEDCT_CORE|Orthostatic hypotension|Orthostatic hypotension
C0020651|T047|SY|28651003|SNOMEDCT_CORE|Postural hypotension|Orthostatic hypotension
C0020672|T033|SY|386689009|SNOMEDCT_CORE|Body temperature below normal|Hypothermia
C0020672|T033|SY|386689009|SNOMEDCT_CORE|Decreased body temperature|Hypothermia
C0020672|T033|PT|386689009|SNOMEDCT_CORE|Hypothermia|Hypothermia
C0020672|T033|FN|386689009|SNOMEDCT_CORE|Hypothermia|Hypothermia
C0020672|T033|SY|386689009|SNOMEDCT_CORE|State of hypothermia|Hypothermia
C0020672|T033|SY|386689009|SNOMEDCT_CORE|Temperature subnormal|Hypothermia
C0020676|T047|SY|40930008|SNOMEDCT_CORE|Hypothyroid|Hypothyroidism
C0020676|T047|PT|40930008|SNOMEDCT_CORE|Hypothyroidism|Hypothyroidism
C0020676|T047|FN|40930008|SNOMEDCT_CORE|Hypothyroidism|Hypothyroidism
C0020676|T047|IS|40930008|SNOMEDCT_CORE|Hypothyroidism, NOS|Hypothyroidism
C0020683|T046|PTGB|39419009|SNOMEDCT_CORE|Hypovolaemic shock|Hypovolemic shock
C0020683|T046|PT|39419009|SNOMEDCT_CORE|Hypovolemic shock|Hypovolemic shock
C0020683|T046|FN|39419009|SNOMEDCT_CORE|Hypovolemic shock|Hypovolemic shock
C0020683|T046|SY|39419009|SNOMEDCT_CORE|Low volume shock|Hypovolemic shock
C0020796|T048|SY|31216003|SNOMEDCT_CORE|Profound intellectual development disorder|Profound intellectual disability
C0020796|T048|FN|31216003|SNOMEDCT_CORE|Profound intellectual disability|Profound intellectual disability
C0020796|T048|PT|31216003|SNOMEDCT_CORE|Profound intellectual disability|Profound intellectual disability
C0020796|T048|SY|31216003|SNOMEDCT_CORE|Profound mental handicap|Profound intellectual disability
C0020877|T047|PT|52457000|SNOMEDCT_CORE|Ileitis|Ileitis
C0020877|T047|FN|52457000|SNOMEDCT_CORE|Ileitis|Ileitis
C0020877|T047|IS|52457000|SNOMEDCT_CORE|Ileitis, NOS|Ileitis
C0021051|T047|SY|234532001|SNOMEDCT_CORE|Immunodeficiency|Immunodeficiency disorder
C0021051|T047|SY|234532001|SNOMEDCT_CORE|Immunodeficiency disease|Immunodeficiency disorder
C0021051|T047|PT|234532001|SNOMEDCT_CORE|Immunodeficiency disorder|Immunodeficiency disorder
C0021051|T047|FN|234532001|SNOMEDCT_CORE|Immunodeficiency disorder|Immunodeficiency disorder
C0021092|T033|PT|18070006|SNOMEDCT_CORE|Impacted cerumen|Impacted cerumen
C0021092|T033|FN|18070006|SNOMEDCT_CORE|Impacted cerumen|Impacted cerumen
C0021092|T033|SY|18070006|SNOMEDCT_CORE|Impacted wax|Impacted cerumen
C0021099|T047|PT|48277006|SNOMEDCT_CORE|Impetigo|Impetigo
C0021099|T047|FN|48277006|SNOMEDCT_CORE|Impetigo|Impetigo
C0021099|T047|IS|48277006|SNOMEDCT_CORE|Impetigo, NOS|Impetigo
C0021122|T048|PT|66347000|SNOMEDCT_CORE|Impulse control disorder|Impulse control disorder
C0021122|T048|FN|66347000|SNOMEDCT_CORE|Impulse control disorder|Impulse control disorder
C0021122|T048|IS|66347000|SNOMEDCT_CORE|Impulse control disorder, NOS|Impulse control disorder
C0021141|T047|SY|55004003|SNOMEDCT_CORE|Schwartz-Bartter syndrome|Syndrome of inappropriate vasopressin secretion
C0021141|T047|IS|55004003|SNOMEDCT_CORE|Schwarz-Bartter syndrome|Syndrome of inappropriate vasopressin secretion
C0021141|T047|SY|55004003|SNOMEDCT_CORE|SIAD - Syndrome of inappropriate antidiuresis|Syndrome of inappropriate vasopressin secretion
C0021141|T047|SY|55004003|SNOMEDCT_CORE|SIADH|Syndrome of inappropriate vasopressin secretion
C0021141|T047|SY|55004003|SNOMEDCT_CORE|SIADH - Syndrome of inappropriate secretion of antidiuretic hormone|Syndrome of inappropriate vasopressin secretion
C0021141|T047|SY|55004003|SNOMEDCT_CORE|Syndrome of inappropriate ADH production|Syndrome of inappropriate vasopressin secretion
C0021141|T047|SY|55004003|SNOMEDCT_CORE|Syndrome of inappropriate antidiuresis|Syndrome of inappropriate vasopressin secretion
C0021141|T047|SY|55004003|SNOMEDCT_CORE|Syndrome of inappropriate antidiuretic hormone secretion|Syndrome of inappropriate vasopressin secretion
C0021141|T047|SY|55004003|SNOMEDCT_CORE|Syndrome of inappropriate secretion of antidiuretic hormone|Syndrome of inappropriate vasopressin secretion
C0021141|T047|PT|55004003|SNOMEDCT_CORE|Syndrome of inappropriate vasopressin secretion|Syndrome of inappropriate vasopressin secretion
C0021141|T047|FN|55004003|SNOMEDCT_CORE|Syndrome of inappropriate vasopressin secretion|Syndrome of inappropriate vasopressin secretion
C0021167|T047|PT|48340000|SNOMEDCT_CORE|Incontinence|Incontinence
C0021167|T047|FN|48340000|SNOMEDCT_CORE|Incontinence|Incontinence
C0021167|T047|IS|48340000|SNOMEDCT_CORE|Incontinence, NOS|Incontinence
C0021294|T033|PT|395507008|SNOMEDCT_CORE|Premature infant|Prematurity of infant
C0021294|T033|FN|395507008|SNOMEDCT_CORE|Premature infant|Prematurity of infant
C0021294|T033|PT|771299009|SNOMEDCT_CORE|Prematurity of infant|Prematurity of infant
C0021294|T033|FN|771299009|SNOMEDCT_CORE|Prematurity of infant|Prematurity of infant
C0021313|T047|FN|129128006|SNOMEDCT_CORE|Infectious disorder of kidney|Infectious disorder of kidney
C0021313|T047|PT|129128006|SNOMEDCT_CORE|Infectious disorder of kidney|Infectious disorder of kidney
C0021313|T047|SY|129128006|SNOMEDCT_CORE|Kidney infection|Infectious disorder of kidney
C0021313|T047|SY|129128006|SNOMEDCT_CORE|Renal infection|Infectious disorder of kidney
C0021345|T047|IS|271558008|SNOMEDCT_CORE|Gammaherpesviral mononucleosis|Infectious mononucleosis
C0021345|T047|SY|271558008|SNOMEDCT_CORE|GF - Glandular fever|Infectious mononucleosis
C0021345|T047|SY|271558008|SNOMEDCT_CORE|Glandular fever|Infectious mononucleosis
C0021345|T047|SY|271558008|SNOMEDCT_CORE|IM - Infectious mononucleosis|Infectious mononucleosis
C0021345|T047|SY|271558008|SNOMEDCT_CORE|IM - Infective mononucleosis|Infectious mononucleosis
C0021345|T047|PT|271558008|SNOMEDCT_CORE|Infectious mononucleosis|Infectious mononucleosis
C0021345|T047|FN|271558008|SNOMEDCT_CORE|Infectious mononucleosis|Infectious mononucleosis
C0021345|T047|SY|271558008|SNOMEDCT_CORE|Infective mononucleosis|Infectious mononucleosis
C0021345|T047|SY|271558008|SNOMEDCT_CORE|Monocytic angina|Infectious mononucleosis
C0021345|T047|SY|271558008|SNOMEDCT_CORE|Mononucleosis syndrome|Infectious mononucleosis
C0021345|T047|SY|271558008|SNOMEDCT_CORE|Pfeiffer's disease|Infectious mononucleosis
C0021355|T047|SY|86981007|SNOMEDCT_CORE|Infective OE|Infective otitis externa
C0021355|T047|PT|86981007|SNOMEDCT_CORE|Infective otitis externa|Infective otitis externa
C0021355|T047|FN|86981007|SNOMEDCT_CORE|Infective otitis externa|Infective otitis externa
C0021355|T047|IS|86981007|SNOMEDCT_CORE|Infective otitis externa, NOS|Infective otitis externa
C0021355|T047|IS|86981007|SNOMEDCT_CORE|Swimmer's ear|Infective otitis externa
C0021355|T047|SY|3135009|SNOMEDCT_CORE|Swimmer's ear|Infective otitis externa
C0021359|T046|SY|8619003|SNOMEDCT_CORE|Cannot achieve a pregnancy|Infertile
C0021359|T046|SY|8619003|SNOMEDCT_CORE|Difficulty conceiving|Infertile
C0021359|T046|PT|8619003|SNOMEDCT_CORE|Infertile|Infertile
C0021359|T046|FN|8619003|SNOMEDCT_CORE|Infertile|Infertile
C0021359|T046|IS|8619003|SNOMEDCT_CORE|Infertility|Infertile
C0021359|T046|IS|8619003|SNOMEDCT_CORE|Infertility, NOS|Infertile
C0021361|T046|PT|6738008|SNOMEDCT_CORE|Female infertility|Female infertility
C0021361|T046|FN|6738008|SNOMEDCT_CORE|Female infertility|Female infertility
C0021361|T046|IS|6738008|SNOMEDCT_CORE|Female infertility, NOS|Female infertility
C0021364|T047|PT|2904007|SNOMEDCT_CORE|Male infertility|Male infertility
C0021364|T047|FN|2904007|SNOMEDCT_CORE|Male infertility|Male infertility
C0021364|T047|OF|2904007|SNOMEDCT_CORE|Male infertility|Male infertility
C0021364|T047|IS|2904007|SNOMEDCT_CORE|Male infertility, NOS|Male infertility
C0021390|T047|SY|24526004|SNOMEDCT_CORE|IBD - Inflammatory bowel disease|Inflammatory bowel disease
C0021390|T047|PT|24526004|SNOMEDCT_CORE|Inflammatory bowel disease|Inflammatory bowel disease
C0021390|T047|FN|24526004|SNOMEDCT_CORE|Inflammatory bowel disease|Inflammatory bowel disease
C0021390|T047|IS|24526004|SNOMEDCT_CORE|Inflammatory bowel disease, NOS|Inflammatory bowel disease
C0021400|T047|SY|6142004|SNOMEDCT_CORE|Flu|Influenza
C0021400|T047|SY|6142004|SNOMEDCT_CORE|Grippe|Influenza
C0021400|T047|PT|6142004|SNOMEDCT_CORE|Influenza|Influenza
C0021400|T047|FN|6142004|SNOMEDCT_CORE|Influenza|Influenza
C0021400|T047|IS|6142004|SNOMEDCT_CORE|Influenza, NOS|Influenza
C0021564|T037|SY|276433004|SNOMEDCT_CORE|Insect bite|Insect bite - wound
C0021564|T037|PT|276433004|SNOMEDCT_CORE|Insect bite - wound|Insect bite - wound
C0021564|T037|FN|276433004|SNOMEDCT_CORE|Insect bite - wound|Insect bite - wound
C0021607|T048|PT|81608000|SNOMEDCT_CORE|Insomnia disorder related to known organic factor|Insomnia disorder related to known organic factor
C0021607|T048|FN|81608000|SNOMEDCT_CORE|Insomnia disorder related to known organic factor|Insomnia disorder related to known organic factor
C0021607|T048|SY|81608000|SNOMEDCT_CORE|Organic insomnia|Insomnia disorder related to known organic factor
C0021655|T046|PT|48606007|SNOMEDCT_CORE|Drug resistance to insulin|Drug resistance to insulin
C0021655|T046|FN|48606007|SNOMEDCT_CORE|Drug resistance to insulin|Drug resistance to insulin
C0021655|T046|IS|48606007|SNOMEDCT_CORE|Insulin resistance|Drug resistance to insulin
C0021775|T047|IS|63491006|SNOMEDCT_CORE|Charcot's syndrome|Intermittent claudication
C0021775|T047|SY|63491006|SNOMEDCT_CORE|Claudication|Intermittent claudication
C0021775|T047|SY|63491006|SNOMEDCT_CORE|IC - Intermittent claudication|Intermittent claudication
C0021775|T047|PT|63491006|SNOMEDCT_CORE|Intermittent claudication|Intermittent claudication
C0021775|T047|FN|63491006|SNOMEDCT_CORE|Intermittent claudication|Intermittent claudication
C0021775|T047|OF|63491006|SNOMEDCT_CORE|Intermittent claudication|Intermittent claudication
C0021775|T047|SY|63491006|SNOMEDCT_CORE|Myasthenia angiosclerotica|Intermittent claudication
C0021776|T048|PT|40987004|SNOMEDCT_CORE|Intermittent explosive disorder|Intermittent explosive disorder
C0021776|T048|FN|40987004|SNOMEDCT_CORE|Intermittent explosive disorder|Intermittent explosive disorder
C0021807|T047|SY|58759008|SNOMEDCT_CORE|Eczema intertrigo|Intertrigo
C0021807|T047|SY|58759008|SNOMEDCT_CORE|Erythema intertrigo|Intertrigo
C0021807|T047|PT|58759008|SNOMEDCT_CORE|Intertrigo|Intertrigo
C0021807|T047|FN|58759008|SNOMEDCT_CORE|Intertrigo|Intertrigo
C0021818|T047|SY|73589001|SNOMEDCT_CORE|Displacement of intervertebral disc|Displacement of intervertebral disc
C0021831|T047|IS|85919009|SNOMEDCT_CORE|Disease of intestine|Disorder of intestine
C0021831|T047|OF|85919009|SNOMEDCT_CORE|Disease of intestine|Disorder of intestine
C0021831|T047|IS|85919009|SNOMEDCT_CORE|Disease of intestine, NOS|Disorder of intestine
C0021831|T047|PT|85919009|SNOMEDCT_CORE|Disorder of intestine|Disorder of intestine
C0021831|T047|FN|85919009|SNOMEDCT_CORE|Disorder of intestine|Disorder of intestine
C0021831|T047|SY|85919009|SNOMEDCT_CORE|Enteropathy|Disorder of intestine
C0021831|T047|IS|85919009|SNOMEDCT_CORE|Enteropathy, NOS|Disorder of intestine
C0021831|T047|SY|85919009|SNOMEDCT_CORE|Intestinal disease|Disorder of intestine
C0021843|T047|SY|81060008|SNOMEDCT_CORE|Bowel obstruction|Intestinal obstruction
C0021843|T047|PT|81060008|SNOMEDCT_CORE|Intestinal obstruction|Intestinal obstruction
C0021843|T047|FN|81060008|SNOMEDCT_CORE|Intestinal obstruction|Intestinal obstruction
C0021843|T047|IS|81060008|SNOMEDCT_CORE|Intestinal obstruction, NOS|Intestinal obstruction
C0021843|T047|IS|81060008|SNOMEDCT_CORE|Intestinal occlusion|Intestinal obstruction
C0021843|T047|IS|81060008|SNOMEDCT_CORE|Intestinal occlusion, NOS|Intestinal obstruction
C0021843|T047|SY|81060008|SNOMEDCT_CORE|IO - Intestinal obstruction|Intestinal obstruction
C0021843|T047|SY|81060008|SNOMEDCT_CORE|Obstruction of intestine|Intestinal obstruction
C0021845|T047|SY|56905009|SNOMEDCT_CORE|Intestinal perforation|Perforation of intestine
C0021845|T047|PT|56905009|SNOMEDCT_CORE|Perforation of intestine|Perforation of intestine
C0021845|T047|FN|56905009|SNOMEDCT_CORE|Perforation of intestine|Perforation of intestine
C0021845|T047|IS|56905009|SNOMEDCT_CORE|Perforation of intestine, NOS|Perforation of intestine
C0021846|T190|SY|254588001|SNOMEDCT_CORE|Bowel polyp|Polyp of intestine
C0021846|T190|SY|254588001|SNOMEDCT_CORE|Intestinal polyp|Polyp of intestine
C0021846|T190|PT|254588001|SNOMEDCT_CORE|Polyp of intestine|Polyp of intestine
C0021846|T190|FN|254588001|SNOMEDCT_CORE|Polyp of intestine|Polyp of intestine
C0021847|T047|PT|235825006|SNOMEDCT_CORE|Pseudo-obstruction of intestine|Pseudo-obstruction of intestine
C0021847|T047|FN|235825006|SNOMEDCT_CORE|Pseudo-obstruction of intestine|Pseudo-obstruction of intestine
C0021933|T047|SY|49723003|SNOMEDCT_CORE|Intestinal intussusception|Intussusception of intestine
C0021933|T047|PT|49723003|SNOMEDCT_CORE|Intussusception of intestine|Intussusception of intestine
C0021933|T047|FN|49723003|SNOMEDCT_CORE|Intussusception of intestine|Intussusception of intestine
C0021933|T047|SY|49723003|SNOMEDCT_CORE|Intussusception of the intestine|Intussusception of intestine
C0021933|T047|SY|49723003|SNOMEDCT_CORE|Invagination of intestine|Intussusception of intestine
C0021933|T047|SY|49723003|SNOMEDCT_CORE|ISN - Intussusception|Intussusception of intestine
C0022073|T047|PT|77971008|SNOMEDCT_CORE|Iridocyclitis|Iridocyclitis
C0022073|T047|FN|77971008|SNOMEDCT_CORE|Iridocyclitis|Iridocyclitis
C0022073|T047|IS|77971008|SNOMEDCT_CORE|Iridocyclitis, NOS|Iridocyclitis
C0022081|T047|PT|65074000|SNOMEDCT_CORE|Iritis|Iritis
C0022081|T047|FN|65074000|SNOMEDCT_CORE|Iritis|Iritis
C0022081|T047|IS|65074000|SNOMEDCT_CORE|Iritis, NOS|Iritis
C0022104|T047|SY|10743008|SNOMEDCT_CORE|Adaptive colitis|Irritable bowel syndrome
C0022104|T047|SY|10743008|SNOMEDCT_CORE|Colon spasm|Irritable bowel syndrome
C0022104|T047|SY|10743008|SNOMEDCT_CORE|Functional bowel disease|Irritable bowel syndrome
C0022104|T047|SY|10743008|SNOMEDCT_CORE|IBS - Irritable bowel syndrome|Irritable bowel syndrome
C0022104|T047|SY|10743008|SNOMEDCT_CORE|IC - Irritable colon|Irritable bowel syndrome
C0022104|T047|SY|10743008|SNOMEDCT_CORE|Irritable bowel|Irritable bowel syndrome
C0022104|T047|PT|10743008|SNOMEDCT_CORE|Irritable bowel syndrome|Irritable bowel syndrome
C0022104|T047|FN|10743008|SNOMEDCT_CORE|Irritable bowel syndrome|Irritable bowel syndrome
C0022104|T047|SY|10743008|SNOMEDCT_CORE|Irritable colon|Irritable bowel syndrome
C0022104|T047|OF|10743008|SNOMEDCT_CORE|Irritable colon|Irritable bowel syndrome
C0022104|T047|SY|10743008|SNOMEDCT_CORE|Irritable colon syndrome|Irritable bowel syndrome
C0022104|T047|SY|10743008|SNOMEDCT_CORE|Membranous colitis|Irritable bowel syndrome
C0022104|T047|SY|10743008|SNOMEDCT_CORE|Mucous colitis|Irritable bowel syndrome
C0022104|T047|SY|10743008|SNOMEDCT_CORE|Nervous colitis|Irritable bowel syndrome
C0022104|T047|IS|10743008|SNOMEDCT_CORE|Psychogenic IBS|Irritable bowel syndrome
C0022104|T047|SY|10743008|SNOMEDCT_CORE|Spastic colitis|Irritable bowel syndrome
C0022104|T047|SY|10743008|SNOMEDCT_CORE|Spastic colon|Irritable bowel syndrome
C0022107|T033|PT|55929007|SNOMEDCT_CORE|Feeling irritable|Feeling irritable
C0022107|T033|FN|55929007|SNOMEDCT_CORE|Feeling irritable|Feeling irritable
C0022107|T033|SY|55929007|SNOMEDCT_CORE|Fussiness|Feeling irritable
C0022107|T033|SY|55929007|SNOMEDCT_CORE|Irritability|Feeling irritable
C0022107|T033|IS|55929007|SNOMEDCT_CORE|Irritable mood|Feeling irritable
C0022116|T046|PTGB|52674009|SNOMEDCT_CORE|Ischaemia|Ischemia
C0022116|T046|IS|52674009|SNOMEDCT_CORE|Ischaemia, NOS|Ischemia
C0022116|T046|PT|52674009|SNOMEDCT_CORE|Ischemia|Ischemia
C0022116|T046|FN|52674009|SNOMEDCT_CORE|Ischemia|Ischemia
C0022116|T046|IS|52674009|SNOMEDCT_CORE|Ischemia, NOS|Ischemia
C0022346|T184|SY|18165001|SNOMEDCT_CORE|Icteric|Jaundice
C0022346|T184|SY|18165001|SNOMEDCT_CORE|Icterus|Jaundice
C0022346|T184|IS|18165001|SNOMEDCT_CORE|Icterus, NOS|Jaundice
C0022346|T184|PT|18165001|SNOMEDCT_CORE|Jaundice|Jaundice
C0022346|T184|FN|18165001|SNOMEDCT_CORE|Jaundice|Jaundice
C0022346|T184|IS|18165001|SNOMEDCT_CORE|Jaundice, NOS|Jaundice
C0022346|T184|SY|18165001|SNOMEDCT_CORE|Jaundiced|Jaundice
C0022353|T047|IS|276549000|SNOMEDCT_CORE|Icterus neonatorum|Neonatal jaundice
C0022353|T047|SY|387712008|SNOMEDCT_CORE|Icterus neonatorum|Neonatal jaundice
C0022353|T047|PT|387712008|SNOMEDCT_CORE|Neonatal jaundice|Neonatal jaundice
C0022353|T047|FN|387712008|SNOMEDCT_CORE|Neonatal jaundice|Neonatal jaundice
C0022354|T047|PTGB|59848001|SNOMEDCT_CORE|Obstructive hyperbilirubinaemia|Obstructive hyperbilirubinemia
C0022354|T047|PT|59848001|SNOMEDCT_CORE|Obstructive hyperbilirubinemia|Obstructive hyperbilirubinemia
C0022354|T047|FN|59848001|SNOMEDCT_CORE|Obstructive hyperbilirubinemia|Obstructive hyperbilirubinemia
C0022354|T047|SY|59848001|SNOMEDCT_CORE|Obstructive jaundice|Obstructive hyperbilirubinemia
C0022361|T020|PT|43144004|SNOMEDCT_CORE|Cyst of jaw|Cyst of jaw
C0022361|T020|FN|43144004|SNOMEDCT_CORE|Cyst of jaw|Cyst of jaw
C0022361|T020|IS|43144004|SNOMEDCT_CORE|Cyst of jaw, NOS|Cyst of jaw
C0022408|T047|PT|399269003|SNOMEDCT_CORE|Arthropathy|Arthropathy
C0022408|T047|FN|399269003|SNOMEDCT_CORE|Arthropathy|Arthropathy
C0022408|T047|SY|399269003|SNOMEDCT_CORE|Arthrosis|Arthropathy
C0022408|T047|SY|399269003|SNOMEDCT_CORE|Disorder of joint|Arthropathy
C0022408|T047|SY|399269003|SNOMEDCT_CORE|Joint disease|Arthropathy
C0022408|T047|SY|399269003|SNOMEDCT_CORE|Joint disorder|Arthropathy
C0022548|T020|SY|33659008|SNOMEDCT_CORE|Cheloid|Keloid scar
C0022548|T020|SY|33659008|SNOMEDCT_CORE|Cheloid of skin|Keloid scar
C0022548|T020|SY|33659008|SNOMEDCT_CORE|Keloid|Keloid scar
C0022548|T020|SY|33659008|SNOMEDCT_CORE|Keloid cicatrix|Keloid scar
C0022548|T020|SY|33659008|SNOMEDCT_CORE|Keloid of skin|Keloid scar
C0022548|T020|PT|33659008|SNOMEDCT_CORE|Keloid scar|Keloid scar
C0022548|T020|FN|33659008|SNOMEDCT_CORE|Keloid scar|Keloid scar
C0022548|T020|IS|33659008|SNOMEDCT_CORE|Keloid scar of skin|Keloid scar
C0022568|T047|PT|5888003|SNOMEDCT_CORE|Keratitis|Keratitis
C0022568|T047|FN|5888003|SNOMEDCT_CORE|Keratitis|Keratitis
C0022568|T047|IS|5888003|SNOMEDCT_CORE|Keratitis, NOS|Keratitis
C0022570|T047|PT|29943008|SNOMEDCT_CORE|Herpes simplex dendritic keratitis|Herpes simplex dendritic keratitis
C0022570|T047|FN|29943008|SNOMEDCT_CORE|Herpes simplex dendritic keratitis|Herpes simplex dendritic keratitis
C0022570|T047|SY|29943008|SNOMEDCT_CORE|HSV dendritic keratitis|Herpes simplex dendritic keratitis
C0022573|T047|PT|88151007|SNOMEDCT_CORE|Keratoconjunctivitis|Keratoconjunctivitis
C0022573|T047|FN|88151007|SNOMEDCT_CORE|Keratoconjunctivitis|Keratoconjunctivitis
C0022573|T047|IS|88151007|SNOMEDCT_CORE|Keratoconjunctivitis, NOS|Keratoconjunctivitis
C0022573|T047|SY|88151007|SNOMEDCT_CORE|Superficial keratitis with conjunctivitis|Keratoconjunctivitis
C0022573|T047|IS|88151007|SNOMEDCT_CORE|Superficial keratitis with conjunctivitis, NOS|Keratoconjunctivitis
C0022575|T047|SY|302896008|SNOMEDCT_CORE|KCS - Keratoconjunctivitis sicca|Keratoconjunctivitis sicca
C0022575|T047|PT|302896008|SNOMEDCT_CORE|Keratoconjunctivitis sicca|Keratoconjunctivitis sicca
C0022575|T047|FN|302896008|SNOMEDCT_CORE|Keratoconjunctivitis sicca|Keratoconjunctivitis sicca
C0022578|T047|SY|65636009|SNOMEDCT_CORE|Cornea conical|Keratoconus
C0022578|T047|PT|65636009|SNOMEDCT_CORE|Keratoconus|Keratoconus
C0022578|T047|FN|65636009|SNOMEDCT_CORE|Keratoconus|Keratoconus
C0022578|T047|IS|65636009|SNOMEDCT_CORE|Keratoconus, NOS|Keratoconus
C0022593|T047|PT|254666005|SNOMEDCT_CORE|Keratosis|Keratosis
C0022593|T047|FN|254666005|SNOMEDCT_CORE|Keratosis|Keratosis
C0022595|T047|PT|48611009|SNOMEDCT_CORE|Darier disease|Darier disease
C0022595|T047|FN|48611009|SNOMEDCT_CORE|Darier disease|Darier disease
C0022595|T047|SY|48611009|SNOMEDCT_CORE|Darier-White disease|Darier disease
C0022595|T047|SY|48611009|SNOMEDCT_CORE|Darier's disease|Darier disease
C0022595|T047|SY|48611009|SNOMEDCT_CORE|Dyskeratosis follicularis|Darier disease
C0022595|T047|IS|48611009|SNOMEDCT_CORE|Follicular keratosis|Darier disease
C0022595|T047|OP|48611009|SNOMEDCT_CORE|Hereditary follicular keratosis|Darier disease
C0022595|T047|SY|48611009|SNOMEDCT_CORE|Keratosis follicularis|Darier disease
C0022595|T047|OF|48611009|SNOMEDCT_CORE|Keratosis follicularis|Darier disease
C0022595|T047|SY|48611009|SNOMEDCT_CORE|Psorospermosis|Darier disease
C0022595|T047|SY|48611009|SNOMEDCT_CORE|Psorospermosis follicularis vegetans|Darier disease
C0022602|T191|PT|201101007|SNOMEDCT_CORE|Actinic keratosis|Actinic keratosis
C0022602|T191|IS|46795000|SNOMEDCT_CORE|Actinic keratosis|Actinic keratosis
C0022602|T191|FN|201101007|SNOMEDCT_CORE|Actinic keratosis|Actinic keratosis
C0022602|T191|IS|46795000|SNOMEDCT_CORE|AK - Actinic keratosis|Actinic keratosis
C0022602|T191|SY|201101007|SNOMEDCT_CORE|AK - Actinic keratosis|Actinic keratosis
C0022602|T191|IS|46795000|SNOMEDCT_CORE|Atrophic keratosis|Actinic keratosis
C0022602|T191|SY|201101007|SNOMEDCT_CORE|Atrophic keratosis|Actinic keratosis
C0022602|T191|IS|46795000|SNOMEDCT_CORE|Hyperplastic keratosis|Actinic keratosis
C0022602|T191|SY|201101007|SNOMEDCT_CORE|Hyperplastic keratosis|Actinic keratosis
C0022602|T191|IS|201101007|SNOMEDCT_CORE|Senile hyperkeratosis|Actinic keratosis
C0022602|T191|IS|46795000|SNOMEDCT_CORE|Senile hyperkeratosis|Actinic keratosis
C0022602|T191|IS|46795000|SNOMEDCT_CORE|Senile keratoma|Actinic keratosis
C0022602|T191|SY|201101007|SNOMEDCT_CORE|Senile keratoma|Actinic keratosis
C0022602|T191|IS|201101007|SNOMEDCT_CORE|Senile keratosis|Actinic keratosis
C0022602|T191|IS|46795000|SNOMEDCT_CORE|Senile keratosis|Actinic keratosis
C0022602|T191|IS|46795000|SNOMEDCT_CORE|SK - Solar keratosis|Actinic keratosis
C0022602|T191|SY|201101007|SNOMEDCT_CORE|SK - Solar keratosis|Actinic keratosis
C0022602|T191|IS|46795000|SNOMEDCT_CORE|Solar keratosis|Actinic keratosis
C0022602|T191|OF|201101007|SNOMEDCT_CORE|Solar keratosis|Actinic keratosis
C0022602|T191|SY|201101007|SNOMEDCT_CORE|Solar keratosis|Actinic keratosis
C0022603|T191|IS|398838000|SNOMEDCT_CORE|Seborrheic keratosis|Seborrheic keratosis
C0022603|T191|IS|50563003|SNOMEDCT_CORE|Seborrheic wart|Seborrheic keratosis
C0022603|T191|IS|398838000|SNOMEDCT_CORE|Seborrhoeic keratosis|Seborrheic keratosis
C0022603|T191|IS|50563003|SNOMEDCT_CORE|Seborrhoeic wart|Seborrheic keratosis
C0022603|T191|IS|50563003|SNOMEDCT_CORE|Senile wart|Seborrheic keratosis
C0022650|T047|SY|95570007|SNOMEDCT_CORE|Calculus of kidney|Kidney stone
C0022650|T047|SY|95570007|SNOMEDCT_CORE|Kidney calculus|Kidney stone
C0022650|T047|PT|95570007|SNOMEDCT_CORE|Kidney stone|Kidney stone
C0022650|T047|FN|95570007|SNOMEDCT_CORE|Kidney stone|Kidney stone
C0022650|T047|SY|95570007|SNOMEDCT_CORE|Nephrolith|Kidney stone
C0022650|T047|SY|95570007|SNOMEDCT_CORE|Nephrolithiasis|Kidney stone
C0022650|T047|SY|95570007|SNOMEDCT_CORE|Renal calculus|Kidney stone
C0022650|T047|SY|95570007|SNOMEDCT_CORE|Renal stone|Kidney stone
C0022658|T047|SY|90708001|SNOMEDCT_CORE|Disease of kidney|Kidney disease
C0022658|T047|SY|90708001|SNOMEDCT_CORE|Disorder of kidney|Kidney disease
C0022658|T047|PT|90708001|SNOMEDCT_CORE|Kidney disease|Kidney disease
C0022658|T047|FN|90708001|SNOMEDCT_CORE|Kidney disease|Kidney disease
C0022658|T047|IS|90708001|SNOMEDCT_CORE|Kidney disease, NOS|Kidney disease
C0022658|T047|SY|90708001|SNOMEDCT_CORE|Nephropathy|Kidney disease
C0022658|T047|IS|90708001|SNOMEDCT_CORE|Nephropathy, NOS|Kidney disease
C0022658|T047|SY|90708001|SNOMEDCT_CORE|Renal disease|Kidney disease
C0022658|T047|IS|90708001|SNOMEDCT_CORE|Renal disease, NOS|Kidney disease
C0022658|T047|SY|90708001|SNOMEDCT_CORE|Renal disorder|Kidney disease
C0022658|T047|IS|90708001|SNOMEDCT_CORE|Renal disorder, NOS|Kidney disease
C0022660|T047|SY|14669001|SNOMEDCT_CORE|Acute renal failure|Acute renal failure syndrome
C0022660|T047|PT|14669001|SNOMEDCT_CORE|Acute renal failure syndrome|Acute renal failure syndrome
C0022660|T047|FN|14669001|SNOMEDCT_CORE|Acute renal failure syndrome|Acute renal failure syndrome
C0022660|T047|IS|14669001|SNOMEDCT_CORE|Acute renal failure syndrome, NOS|Acute renal failure syndrome
C0022660|T047|SY|14669001|SNOMEDCT_CORE|ARF - Acute renal failure|Acute renal failure syndrome
C0022661|T047|PT|90688005|SNOMEDCT_CORE|Chronic renal failure|Chronic renal failure
C0022661|T047|SY|90688005|SNOMEDCT_CORE|Chronic renal failure syndrome|Chronic renal failure
C0022661|T047|FN|90688005|SNOMEDCT_CORE|Chronic renal failure syndrome|Chronic renal failure
C0022661|T047|IS|90688005|SNOMEDCT_CORE|Chronic renal failure syndrome, NOS|Chronic renal failure
C0022661|T047|SY|90688005|SNOMEDCT_CORE|CRF - Chronic renal failure|Chronic renal failure
C0022661|T047|IS|46177005|SNOMEDCT_CORE|End stage chronc renal failure|Chronic renal failure
C0022661|T047|SY|46177005|SNOMEDCT_CORE|End stage chronic renal failure|Chronic renal failure
C0022661|T047|SY|46177005|SNOMEDCT_CORE|End stage kidney disease|Chronic renal failure
C0022661|T047|OP|46177005|SNOMEDCT_CORE|End stage renal disease|Chronic renal failure
C0022661|T047|OF|46177005|SNOMEDCT_CORE|End stage renal disease|Chronic renal failure
C0022661|T047|PT|46177005|SNOMEDCT_CORE|End-stage renal disease|Chronic renal failure
C0022661|T047|FN|46177005|SNOMEDCT_CORE|End-stage renal disease|Chronic renal failure
C0022661|T047|SY|46177005|SNOMEDCT_CORE|ESCRF - End stage chronic renal failure|Chronic renal failure
C0022661|T047|SY|46177005|SNOMEDCT_CORE|ESRD - End stage renal disease|Chronic renal failure
C0022661|T047|SY|46177005|SNOMEDCT_CORE|ESRF - End stage renal failure|Chronic renal failure
C0022665|T191|PT|126880001|SNOMEDCT_CORE|Neoplasm of kidney|Neoplasm of kidney
C0022665|T191|FN|126880001|SNOMEDCT_CORE|Neoplasm of kidney|Neoplasm of kidney
C0022665|T191|SY|126880001|SNOMEDCT_CORE|Renal tumor|Neoplasm of kidney
C0022665|T191|SYGB|126880001|SNOMEDCT_CORE|Renal tumour|Neoplasm of kidney
C0022665|T191|SY|126880001|SNOMEDCT_CORE|Tumor of kidney|Neoplasm of kidney
C0022665|T191|SYGB|126880001|SNOMEDCT_CORE|Tumour of kidney|Neoplasm of kidney
C0022680|T047|SY|82525005|SNOMEDCT_CORE|PCK - Polycystic kidney disease|PKD - Polycystic kidney disease
C0022680|T047|SY|82525005|SNOMEDCT_CORE|PKD - Polycystic kidney disease|PKD - Polycystic kidney disease
C0022680|T047|SY|82525005|SNOMEDCT_CORE|Polycystic kidney disease|PKD - Polycystic kidney disease
C0022681|T019|PT|236443009|SNOMEDCT_CORE|Medullary sponge kidney|Medullary sponge kidney
C0022681|T047|PT|236443009|SNOMEDCT_CORE|Medullary sponge kidney|Medullary sponge kidney
C0022681|T019|FN|236443009|SNOMEDCT_CORE|Medullary sponge kidney|Medullary sponge kidney
C0022681|T047|FN|236443009|SNOMEDCT_CORE|Medullary sponge kidney|Medullary sponge kidney
C0022739|T047|IS|721105004|SNOMEDCT_CORE|Angio-osteohypertrophy syndrome|Klippel Trenaunay syndrome
C0022739|T047|IS|721105004|SNOMEDCT_CORE|Angioosteohypertrophic syndrome|Klippel Trenaunay syndrome
C0022739|T047|OAS|59078009|SNOMEDCT_CORE|Cerebrofacial angiomatosis|Klippel Trenaunay syndrome
C0022739|T047|OAS|59078009|SNOMEDCT_CORE|Haemangiectatic hypertrophy|Klippel Trenaunay syndrome
C0022739|T047|OAS|59078009|SNOMEDCT_CORE|Hemangiectatic hypertrophy|Klippel Trenaunay syndrome
C0022739|T047|FN|721105004|SNOMEDCT_CORE|Klippel Trenaunay syndrome|Klippel Trenaunay syndrome
C0022739|T047|PT|721105004|SNOMEDCT_CORE|Klippel Trenaunay syndrome|Klippel Trenaunay syndrome
C0022739|T047|OAP|59078009|SNOMEDCT_CORE|Klippel-Trenaunay-Weber syndrome|Klippel Trenaunay syndrome
C0022739|T047|OAF|59078009|SNOMEDCT_CORE|Klippel-Trenaunay-Weber syndrome|Klippel Trenaunay syndrome
C0022744|T037|PT|125601008|SNOMEDCT_CORE|Injury of knee|Injury of knee
C0022744|T037|FN|125601008|SNOMEDCT_CORE|Injury of knee|Injury of knee
C0022744|T037|SY|125601008|SNOMEDCT_CORE|Knee injury|Injury of knee
C0022790|T191|SY|94455000|SNOMEDCT_CORE|Cancer metastatic to ovary|Secondary malignant neoplasm of ovary
C0022790|T191|SY|94455000|SNOMEDCT_CORE|Krukenburg tumor|Secondary malignant neoplasm of ovary
C0022790|T191|SYGB|94455000|SNOMEDCT_CORE|Krukenburg tumour|Secondary malignant neoplasm of ovary
C0022790|T191|SY|94455000|SNOMEDCT_CORE|Metastasis to ovary|Secondary malignant neoplasm of ovary
C0022790|T191|SY|94455000|SNOMEDCT_CORE|Metastatic malignant neoplasm to ovary|Secondary malignant neoplasm of ovary
C0022790|T191|SY|94455000|SNOMEDCT_CORE|Ovarian metastasis|Secondary malignant neoplasm of ovary
C0022790|T191|SY|94455000|SNOMEDCT_CORE|Secondary cancer of ovary|Secondary malignant neoplasm of ovary
C0022790|T191|PT|94455000|SNOMEDCT_CORE|Secondary malignant neoplasm of ovary|Secondary malignant neoplasm of ovary
C0022790|T191|FN|94455000|SNOMEDCT_CORE|Secondary malignant neoplasm of ovary|Secondary malignant neoplasm of ovary
C0022790|T191|SY|94455000|SNOMEDCT_CORE|Secondary tumor to ovary|Secondary malignant neoplasm of ovary
C0022790|T191|SYGB|94455000|SNOMEDCT_CORE|Secondary tumour to ovary|Secondary malignant neoplasm of ovary
C0022820|T190|PT|203638000|SNOMEDCT_CORE|Kyphoscoliosis and scoliosis|Kyphoscoliosis and scoliosis
C0022820|T190|FN|203638000|SNOMEDCT_CORE|Kyphoscoliosis and scoliosis|Kyphoscoliosis and scoliosis
C0022821|T190|SY|414564002|SNOMEDCT_CORE|Gibbosity|Kyphosis deformity of spine
C0022821|T190|SY|414564002|SNOMEDCT_CORE|Gibbus|Kyphosis deformity of spine
C0022821|T190|SY|414564002|SNOMEDCT_CORE|Humpback|Kyphosis deformity of spine
C0022821|T190|SY|414564002|SNOMEDCT_CORE|Hunchback|Kyphosis deformity of spine
C0022821|T190|SY|414564002|SNOMEDCT_CORE|Kyphosis|Kyphosis deformity of spine
C0022821|T190|PT|414564002|SNOMEDCT_CORE|Kyphosis deformity of spine|Kyphosis deformity of spine
C0022821|T190|FN|414564002|SNOMEDCT_CORE|Kyphosis deformity of spine|Kyphosis deformity of spine
C0022822|T020|SY|413428007|SNOMEDCT_CORE|Acquired hunchback|Acquired kyphosis
C0022822|T020|PT|413428007|SNOMEDCT_CORE|Acquired kyphosis|Acquired kyphosis
C0022822|T020|FN|413428007|SNOMEDCT_CORE|Acquired kyphosis|Acquired kyphosis
C0022876|T046|PT|6383007|SNOMEDCT_CORE|Premature labor|Premature labor
C0022876|T046|FN|6383007|SNOMEDCT_CORE|Premature labor|Premature labor
C0022876|T046|PTGB|6383007|SNOMEDCT_CORE|Premature labour|Premature labor
C0022876|T046|SY|6383007|SNOMEDCT_CORE|Premature onset of labor|Premature labor
C0022876|T046|SYGB|6383007|SNOMEDCT_CORE|Premature onset of labour|Premature labor
C0022876|T046|SY|6383007|SNOMEDCT_CORE|Preterm labor|Premature labor
C0022876|T046|SYGB|6383007|SNOMEDCT_CORE|Preterm labour|Premature labor
C0022890|T047|PT|20425006|SNOMEDCT_CORE|Labyrinthine disorder|Labyrinthine disorder
C0022890|T047|FN|20425006|SNOMEDCT_CORE|Labyrinthine disorder|Labyrinthine disorder
C0022890|T047|IS|20425006|SNOMEDCT_CORE|Labyrinthine disorder, NOS|Labyrinthine disorder
C0022893|T047|PT|23919004|SNOMEDCT_CORE|Labyrinthitis|Labyrinthitis
C0022893|T047|FN|23919004|SNOMEDCT_CORE|Labyrinthitis|Labyrinthitis
C0022893|T047|IS|23919004|SNOMEDCT_CORE|Labyrinthitis, NOS|Labyrinthitis
C0022906|T190|SY|416920000|SNOMEDCT_CORE|Canalicular obstruction|Obstruction of lacrimal canaliculus
C0022906|T190|SY|416920000|SNOMEDCT_CORE|Lacrimal canalicular obstruction|Obstruction of lacrimal canaliculus
C0022906|T190|PT|416920000|SNOMEDCT_CORE|Obstruction of lacrimal canaliculus|Obstruction of lacrimal canaliculus
C0022906|T190|FN|416920000|SNOMEDCT_CORE|Obstruction of lacrimal canaliculus|Obstruction of lacrimal canaliculus
C0022906|T190|SY|416920000|SNOMEDCT_CORE|Obstruction of lacrimal duct|Obstruction of lacrimal canaliculus
C0022951|T047|OAS|267425008|SNOMEDCT_CORE|Cow's milk enteropathy|LM - Lactose malabsorption
C0022951|T047|OAP|267425008|SNOMEDCT_CORE|Lactose intolerance|LM - Lactose malabsorption
C0022951|T047|OAF|267425008|SNOMEDCT_CORE|Lactose intolerance|LM - Lactose malabsorption
C0022951|T047|OAS|267425008|SNOMEDCT_CORE|Lactose malabsorption|LM - Lactose malabsorption
C0022951|T047|OAS|267425008|SNOMEDCT_CORE|LM - Lactose malabsorption|LM - Lactose malabsorption
C0023009|T047|PT|231543005|SNOMEDCT_CORE|Speech and language disorder|Speech and language disorder
C0023009|T047|FN|231543005|SNOMEDCT_CORE|Speech and language disorder|Speech and language disorder
C0023009|T047|SY|231543005|SNOMEDCT_CORE|Speech, language, communication disorder|Speech and language disorder
C0023014|T048|PT|280032002|SNOMEDCT_CORE|Developmental language disorder|Developmental language disorder
C0023014|T048|FN|280032002|SNOMEDCT_CORE|Developmental language disorder|Developmental language disorder
C0023014|T048|OAP|231535000|SNOMEDCT_CORE|Language development disorder|Developmental language disorder
C0023014|T048|OAF|231535000|SNOMEDCT_CORE|Language development disorder|Developmental language disorder
C0023051|T047|SY|60600009|SNOMEDCT_CORE|Disease of larynx|Disorder of the larynx
C0023051|T047|IS|60600009|SNOMEDCT_CORE|Disease of the larynx|Disorder of the larynx
C0023051|T047|OF|60600009|SNOMEDCT_CORE|Disease of the larynx|Disorder of the larynx
C0023051|T047|IS|60600009|SNOMEDCT_CORE|Disease of the larynx, NOS|Disorder of the larynx
C0023051|T047|SY|60600009|SNOMEDCT_CORE|Disorder of larynx|Disorder of the larynx
C0023051|T047|PT|60600009|SNOMEDCT_CORE|Disorder of the larynx|Disorder of the larynx
C0023051|T047|FN|60600009|SNOMEDCT_CORE|Disorder of the larynx|Disorder of the larynx
C0023055|T191|PT|126692004|SNOMEDCT_CORE|Neoplasm of larynx|Neoplasm of larynx
C0023055|T191|FN|126692004|SNOMEDCT_CORE|Neoplasm of larynx|Neoplasm of larynx
C0023055|T191|SY|126692004|SNOMEDCT_CORE|Tumor of larynx|Neoplasm of larynx
C0023055|T191|SYGB|126692004|SNOMEDCT_CORE|Tumour of larynx|Neoplasm of larynx
C0023066|T047|PT|53787002|SNOMEDCT_CORE|Laryngismus|Laryngismus
C0023066|T047|FN|53787002|SNOMEDCT_CORE|Laryngismus|Laryngismus
C0023066|T047|IS|53787002|SNOMEDCT_CORE|Laryngismus, NOS|Laryngismus
C0023067|T047|PT|45913009|SNOMEDCT_CORE|Laryngitis|Laryngitis
C0023067|T047|FN|45913009|SNOMEDCT_CORE|Laryngitis|Laryngitis
C0023067|T047|IS|45913009|SNOMEDCT_CORE|Laryngitis, NOS|Laryngitis
C0023176|T037|SY|38342005|SNOMEDCT_CORE|Lead - toxic effect|Toxic effect of lead compound
C0023176|T037|SY|38342005|SNOMEDCT_CORE|Lead compound poisoning|Toxic effect of lead compound
C0023176|T037|SY|38342005|SNOMEDCT_CORE|Lead poisoning|Toxic effect of lead compound
C0023176|T037|SY|38342005|SNOMEDCT_CORE|Plumbism|Toxic effect of lead compound
C0023176|T037|SY|38342005|SNOMEDCT_CORE|Saturnine poisoning|Toxic effect of lead compound
C0023176|T037|PT|38342005|SNOMEDCT_CORE|Toxic effect of lead compound|Toxic effect of lead compound
C0023176|T037|FN|38342005|SNOMEDCT_CORE|Toxic effect of lead compound|Toxic effect of lead compound
C0023176|T037|IS|38342005|SNOMEDCT_CORE|Toxic effect of lead compound, NOS|Toxic effect of lead compound
C0023186|T048|SY|1855002|SNOMEDCT_CORE|Academic skill disorder|Academic skill disorder
C0023186|T048|IS|1855002|SNOMEDCT_CORE|Academic skill disorder, NOS|Academic skill disorder
C0023186|T048|SY|1855002|SNOMEDCT_CORE|Learning disorder|Academic skill disorder
C0023186|T048|IS|1855002|SNOMEDCT_CORE|Learning disorder, NOS|Academic skill disorder
C0023211|T047|SY|63467002|SNOMEDCT_CORE|LBBB - Left bundle branch block|Left bundle branch block
C0023211|T047|PT|63467002|SNOMEDCT_CORE|Left bundle branch block|Left bundle branch block
C0023211|T047|FN|63467002|SNOMEDCT_CORE|Left bundle branch block|Left bundle branch block
C0023211|T047|IS|63467002|SNOMEDCT_CORE|Left bundle branch block, NOS|Left bundle branch block
C0023212|T047|PT|85232009|SNOMEDCT_CORE|Left heart failure|Left heart failure
C0023212|T047|FN|85232009|SNOMEDCT_CORE|Left heart failure|Left heart failure
C0023212|T047|SY|85232009|SNOMEDCT_CORE|Left ventricular failure|Left heart failure
C0023212|T047|SY|85232009|SNOMEDCT_CORE|Left-sided heart failure|Left heart failure
C0023212|T047|SY|85232009|SNOMEDCT_CORE|LVF - Left ventricular failure|Left heart failure
C0023218|T184|OAP|102550009|SNOMEDCT_CORE|Leg cramp|Leg cramps
C0023218|T184|OAF|102550009|SNOMEDCT_CORE|Leg cramp|Leg cramps
C0023218|T184|OAS|102550009|SNOMEDCT_CORE|Leg cramps|Leg cramps
C0023218|T184|IS|102550009|SNOMEDCT_CORE|Muscle cramps in leg|Leg cramps
C0023220|T037|PT|127279002|SNOMEDCT_CORE|Injury of lower extremity|Injury of lower extremity
C0023220|T037|FN|127279002|SNOMEDCT_CORE|Injury of lower extremity|Injury of lower extremity
C0023220|T037|SY|127279002|SNOMEDCT_CORE|Injury of lower limb|Injury of lower extremity
C0023220|T037|IS|127279002|SNOMEDCT_CORE|Leg injury|Injury of lower extremity
C0023221|T033|IS|45939007|SNOMEDCT_CORE|Leg length discrepancy|Leg length inequality
C0023221|T033|PT|45939007|SNOMEDCT_CORE|Leg length inequality|Leg length inequality
C0023221|T033|FN|45939007|SNOMEDCT_CORE|Leg length inequality|Leg length inequality
C0023221|T033|OF|45939007|SNOMEDCT_CORE|Leg length inequality|Leg length inequality
C0023221|T033|SY|45939007|SNOMEDCT_CORE|Lower limb length difference|Leg length inequality
C0023222|T184|IS|10601006|SNOMEDCT_CORE|Leg pain|Pain in lower limb
C0023222|T184|IS|10601006|SNOMEDCT_CORE|Leg pain, NOS|Pain in lower limb
C0023222|T184|PT|10601006|SNOMEDCT_CORE|Pain in lower limb|Pain in lower limb
C0023222|T184|FN|10601006|SNOMEDCT_CORE|Pain in lower limb|Pain in lower limb
C0023223|T047|SY|95344007|SNOMEDCT_CORE|Leg ulcer|Ulcer of lower extremity
C0023223|T047|OF|95344007|SNOMEDCT_CORE|Leg ulcer|Ulcer of lower extremity
C0023223|T047|IS|95344007|SNOMEDCT_CORE|Ulcer of leg|Ulcer of lower extremity
C0023223|T047|IS|95344007|SNOMEDCT_CORE|Ulcer of leg, NOS|Ulcer of lower extremity
C0023223|T047|PT|95344007|SNOMEDCT_CORE|Ulcer of lower extremity|Ulcer of lower extremity
C0023223|T047|FN|95344007|SNOMEDCT_CORE|Ulcer of lower extremity|Ulcer of lower extremity
C0023223|T047|SY|95344007|SNOMEDCT_CORE|Ulcer of lower limb|Ulcer of lower extremity
C0023234|T047|SY|111255008|SNOMEDCT_CORE|Legg-Calve-Perthes disease|Pseudocoxalgia
C0023234|T047|IS|111255008|SNOMEDCT_CORE|Perthe's disease|Pseudocoxalgia
C0023234|T047|IS|111255008|SNOMEDCT_CORE|Perthe's disease of hip|Pseudocoxalgia
C0023234|T047|SY|111255008|SNOMEDCT_CORE|Perthes disease - osteochondritis of the femoral head|Pseudocoxalgia
C0023234|T047|IS|111255008|SNOMEDCT_CORE|Perthes' disease - osteochondritis of the femoral head|Pseudocoxalgia
C0023234|T047|SY|111255008|SNOMEDCT_CORE|Pseudocoxalgia|Pseudocoxalgia
C0023269|T191|OF|51549004|SNOMEDCT_CORE|Leiomyomosarcoma, no subtype|Leiomyosarcoma
C0023269|T191|PT|443719001|SNOMEDCT_CORE|Leiomyosarcoma|Leiomyosarcoma
C0023269|T191|PT|51549004|SNOMEDCT_CORE|Leiomyosarcoma|Leiomyosarcoma
C0023269|T191|FN|443719001|SNOMEDCT_CORE|Leiomyosarcoma|Leiomyosarcoma
C0023269|T191|FN|51549004|SNOMEDCT_CORE|Leiomyosarcoma, no subtype|Leiomyosarcoma
C0023269|T191|SY|51549004|SNOMEDCT_CORE|Leiomyosarcoma, no subtype|Leiomyosarcoma
C0023269|T191|IS|51549004|SNOMEDCT_CORE|Leiomyosarcoma, NOS|Leiomyosarcoma
C0023269|T191|SY|51549004|SNOMEDCT_CORE|LMS - Leiomyosarcoma|Leiomyosarcoma
C0023316|T047|SY|65814009|SNOMEDCT_CORE|Partial dislocation of lens|Subluxation of lens
C0023316|T047|PT|65814009|SNOMEDCT_CORE|Subluxation of lens|Subluxation of lens
C0023316|T047|FN|65814009|SNOMEDCT_CORE|Subluxation of lens|Subluxation of lens
C0023321|T047|PT|402624000|SNOMEDCT_CORE|Lentiginosis|Lentiginosis
C0023321|T047|FN|402624000|SNOMEDCT_CORE|Lentiginosis|Lentiginosis
C0023321|T047|OAP|398744007|SNOMEDCT_CORE|Lentigo|Lentiginosis
C0023321|T047|OAF|398744007|SNOMEDCT_CORE|Lentigo|Lentiginosis
C0023380|T184|SY|214264003|SNOMEDCT_CORE|Lethargic|Lethargy
C0023380|T184|PT|214264003|SNOMEDCT_CORE|Lethargy|Lethargy
C0023380|T184|FN|214264003|SNOMEDCT_CORE|Lethargy|Lethargy
C0023418|T191|PTGB|93143009|SNOMEDCT_CORE|Leukaemia|Leukemia
C0023418|T191|SYGB|93143009|SNOMEDCT_CORE|Leukaemia, disease|Leukemia
C0023418|T191|IS|93143009|SNOMEDCT_CORE|Leukaemia, NOS, without mention of remission|Leukemia
C0023418|T191|PT|93143009|SNOMEDCT_CORE|Leukemia|Leukemia
C0023418|T191|FN|93143009|SNOMEDCT_CORE|Leukemia, disease|Leukemia
C0023418|T191|SY|93143009|SNOMEDCT_CORE|Leukemia, disease|Leukemia
C0023418|T191|IS|93143009|SNOMEDCT_CORE|Leukemia, NOS, without mention of remission|Leukemia
C0023434|T191|SYGB|92814006|SNOMEDCT_CORE|Chronic lymphoid leukaemia|Chronic lymphoid leukemia, disease
C0023434|T191|PTGB|92814006|SNOMEDCT_CORE|Chronic lymphoid leukaemia, disease|Chronic lymphoid leukemia, disease
C0023434|T191|SY|92814006|SNOMEDCT_CORE|Chronic lymphoid leukemia|Chronic lymphoid leukemia, disease
C0023434|T191|FN|92814006|SNOMEDCT_CORE|Chronic lymphoid leukemia, disease|Chronic lymphoid leukemia, disease
C0023434|T191|PT|92814006|SNOMEDCT_CORE|Chronic lymphoid leukemia, disease|Chronic lymphoid leukemia, disease
C0023434|T191|SYGB|92814006|SNOMEDCT_CORE|CLL - Chronic lymphocytic leukaemia|Chronic lymphoid leukemia, disease
C0023434|T191|SY|92814006|SNOMEDCT_CORE|CLL - Chronic lymphocytic leukemia|Chronic lymphoid leukemia, disease
C0023443|T191|SYGB|118613001|SNOMEDCT_CORE|Hairy cell leukaemia|Hairy cell leukemia
C0023443|T191|PTGB|118613001|SNOMEDCT_CORE|Hairy cell leukaemia|Hairy cell leukemia
C0023443|T191|SY|118613001|SNOMEDCT_CORE|Hairy cell leukemia|Hairy cell leukemia
C0023443|T191|PT|118613001|SNOMEDCT_CORE|Hairy cell leukemia|Hairy cell leukemia
C0023443|T191|FN|118613001|SNOMEDCT_CORE|Hairy cell leukemia|Hairy cell leukemia
C0023443|T191|SYGB|118613001|SNOMEDCT_CORE|HCL - Hairy cell leukaemia|Hairy cell leukemia
C0023443|T191|SY|118613001|SNOMEDCT_CORE|HCL - Hairy cell leukemia|Hairy cell leukemia
C0023443|T191|SYGB|118613001|SNOMEDCT_CORE|Leukaemic reticuloendotheliosis|Hairy cell leukemia
C0023443|T191|SY|118613001|SNOMEDCT_CORE|Leukemic reticuloendotheliosis|Hairy cell leukemia
C0023443|T191|SYGB|118613001|SNOMEDCT_CORE|LRE - Leukaemic reticuloendotheliosis|Hairy cell leukemia
C0023443|T191|SY|118613001|SNOMEDCT_CORE|LRE - Leukemic reticuloendotheliosis|Hairy cell leukemia
C0023449|T191|PTGB|91857003|SNOMEDCT_CORE|Acute lymphoid leukaemia|Acute lymphoid leukemia
C0023449|T191|SYGB|91857003|SNOMEDCT_CORE|Acute lymphoid leukaemia, disease|Acute lymphoid leukemia
C0023449|T191|PT|91857003|SNOMEDCT_CORE|Acute lymphoid leukemia|Acute lymphoid leukemia
C0023449|T191|FN|91857003|SNOMEDCT_CORE|Acute lymphoid leukemia, disease|Acute lymphoid leukemia
C0023449|T191|SY|91857003|SNOMEDCT_CORE|Acute lymphoid leukemia, disease|Acute lymphoid leukemia
C0023449|T191|SYGB|91857003|SNOMEDCT_CORE|ALL - Acute lymphoblastic leukaemia|Acute lymphoid leukemia
C0023449|T191|SY|91857003|SNOMEDCT_CORE|ALL - Acute lymphoblastic leukemia|Acute lymphoid leukemia
C0023467|T191|SYGB|91861009|SNOMEDCT_CORE|Acute myelocytic leukaemia|Acute myeloid leukemia, disease
C0023467|T191|SY|91861009|SNOMEDCT_CORE|Acute myelocytic leukemia|Acute myeloid leukemia, disease
C0023467|T191|SYGB|91861009|SNOMEDCT_CORE|Acute myeloid leukaemia|Acute myeloid leukemia, disease
C0023467|T191|PTGB|91861009|SNOMEDCT_CORE|Acute myeloid leukaemia, disease|Acute myeloid leukemia, disease
C0023467|T191|SY|91861009|SNOMEDCT_CORE|Acute myeloid leukemia|Acute myeloid leukemia, disease
C0023467|T191|FN|91861009|SNOMEDCT_CORE|Acute myeloid leukemia, disease|Acute myeloid leukemia, disease
C0023467|T191|PT|91861009|SNOMEDCT_CORE|Acute myeloid leukemia, disease|Acute myeloid leukemia, disease
C0023467|T191|SYGB|91861009|SNOMEDCT_CORE|AML - Acute myeloblastic leukaemia|Acute myeloid leukemia, disease
C0023467|T191|SY|91861009|SNOMEDCT_CORE|AML - Acute myeloblastic leukemia|Acute myeloid leukemia, disease
C0023467|T191|SYGB|91861009|SNOMEDCT_CORE|AML - Acute myeloid leukaemia|Acute myeloid leukemia, disease
C0023467|T191|SY|91861009|SNOMEDCT_CORE|AML - Acute myeloid leukemia|Acute myeloid leukemia, disease
C0023473|T191|SYGB|92818009|SNOMEDCT_CORE|CGL - Chronic granulocytic leukaemia|Chronic myeloid leukemia
C0023473|T191|SY|92818009|SNOMEDCT_CORE|CGL - Chronic granulocytic leukemia|Chronic myeloid leukemia
C0023473|T191|SYGB|92818009|SNOMEDCT_CORE|Chronic myelocytic leukaemia|Chronic myeloid leukemia
C0023473|T191|SY|92818009|SNOMEDCT_CORE|Chronic myelocytic leukemia|Chronic myeloid leukemia
C0023473|T191|PTGB|92818009|SNOMEDCT_CORE|Chronic myeloid leukaemia|Chronic myeloid leukemia
C0023473|T191|SYGB|92818009|SNOMEDCT_CORE|Chronic myeloid leukaemia, disease|Chronic myeloid leukemia
C0023473|T191|PT|92818009|SNOMEDCT_CORE|Chronic myeloid leukemia|Chronic myeloid leukemia
C0023473|T191|FN|92818009|SNOMEDCT_CORE|Chronic myeloid leukemia, disease|Chronic myeloid leukemia
C0023473|T191|SY|92818009|SNOMEDCT_CORE|Chronic myeloid leukemia, disease|Chronic myeloid leukemia
C0023473|T191|SYGB|92818009|SNOMEDCT_CORE|CML - Chronic myeloid leukaemia|Chronic myeloid leukemia
C0023473|T191|SY|92818009|SNOMEDCT_CORE|CML - Chronic myeloid leukemia|Chronic myeloid leukemia
C0023479|T191|SYGB|110005000|SNOMEDCT_CORE|Acute myelomonocytic leukaemia|Acute myelomonocytic leukemia, FAB M4
C0023479|T191|PTGB|110005000|SNOMEDCT_CORE|Acute myelomonocytic leukaemia, FAB M4|Acute myelomonocytic leukemia, FAB M4
C0023479|T191|SY|110005000|SNOMEDCT_CORE|Acute myelomonocytic leukemia|Acute myelomonocytic leukemia, FAB M4
C0023479|T191|PT|110005000|SNOMEDCT_CORE|Acute myelomonocytic leukemia, FAB M4|Acute myelomonocytic leukemia, FAB M4
C0023479|T191|FN|110005000|SNOMEDCT_CORE|Acute myelomonocytic leukemia, FAB M4|Acute myelomonocytic leukemia, FAB M4
C0023479|T191|SYGB|110005000|SNOMEDCT_CORE|AMML - Acute myelomonocytic leukaemia|Acute myelomonocytic leukemia, FAB M4
C0023479|T191|SY|110005000|SNOMEDCT_CORE|AMML - Acute myelomonocytic leukemia|Acute myelomonocytic leukemia, FAB M4
C0023479|T191|OF|110005000|SNOMEDCT_CORE|Disorder: Acute myelomonocytic leukemia, FAB M4|Acute myelomonocytic leukemia, FAB M4
C0023479|T191|SYGB|110005000|SNOMEDCT_CORE|M4 - Acute myelomonocytic leukaemia|Acute myelomonocytic leukemia, FAB M4
C0023479|T191|SY|110005000|SNOMEDCT_CORE|M4 - Acute myelomonocytic leukemia|Acute myelomonocytic leukemia, FAB M4
C0023480|T191|PTGB|127225006|SNOMEDCT_CORE|Chronic myelomonocytic leukaemia|Chronic myelomonocytic leukemia
C0023480|T191|IS|127225006|SNOMEDCT_CORE|Chronic myelomonocytic leukaemia|Chronic myelomonocytic leukemia
C0023480|T191|PT|127225006|SNOMEDCT_CORE|Chronic myelomonocytic leukemia|Chronic myelomonocytic leukemia
C0023480|T191|IS|127225006|SNOMEDCT_CORE|Chronic myelomonocytic leukemia|Chronic myelomonocytic leukemia
C0023480|T191|FN|127225006|SNOMEDCT_CORE|Chronic myelomonocytic leukemia|Chronic myelomonocytic leukemia
C0023487|T191|SYGB|110004001|SNOMEDCT_CORE|Acute promyelocytic leukaemia|Acute promyelocytic leukemia, FAB M3
C0023487|T191|PTGB|110004001|SNOMEDCT_CORE|Acute promyelocytic leukaemia, FAB M3|Acute promyelocytic leukemia, FAB M3
C0023487|T191|SY|110004001|SNOMEDCT_CORE|Acute promyelocytic leukemia|Acute promyelocytic leukemia, FAB M3
C0023487|T191|PT|110004001|SNOMEDCT_CORE|Acute promyelocytic leukemia, FAB M3|Acute promyelocytic leukemia, FAB M3
C0023487|T191|FN|110004001|SNOMEDCT_CORE|Acute promyelocytic leukemia, FAB M3|Acute promyelocytic leukemia, FAB M3
C0023487|T191|SYGB|110004001|SNOMEDCT_CORE|APL - Acute promyelocytic leukaemia|Acute promyelocytic leukemia, FAB M3
C0023487|T191|SY|110004001|SNOMEDCT_CORE|APL - Acute promyelocytic leukemia|Acute promyelocytic leukemia, FAB M3
C0023487|T191|SYGB|110004001|SNOMEDCT_CORE|APML - Acute promyelocytic leukaemia|Acute promyelocytic leukemia, FAB M3
C0023487|T191|SY|110004001|SNOMEDCT_CORE|APML - Acute promyelocytic leukemia|Acute promyelocytic leukemia, FAB M3
C0023487|T191|OF|110004001|SNOMEDCT_CORE|Disorder: Acute promyelocytic leukemia, FAB M3|Acute promyelocytic leukemia, FAB M3
C0023487|T191|SYGB|110004001|SNOMEDCT_CORE|M3 - Acute promyelocytic leukaemia|Acute promyelocytic leukemia, FAB M3
C0023487|T191|SY|110004001|SNOMEDCT_CORE|M3 - Acute promyelocytic leukemia|Acute promyelocytic leukemia, FAB M3
C0023494|T191|PTGB|277545003|SNOMEDCT_CORE|T-cell chronic lymphocytic leukaemia|T-cell chronic lymphocytic leukemia
C0023494|T191|PT|277545003|SNOMEDCT_CORE|T-cell chronic lymphocytic leukemia|T-cell chronic lymphocytic leukemia
C0023494|T191|FN|277545003|SNOMEDCT_CORE|T-cell chronic lymphocytic leukemia|T-cell chronic lymphocytic leukemia
C0023494|T191|SYGB|277545003|SNOMEDCT_CORE|TCLL - T-cell chronic lymphocytic leukaemia|T-cell chronic lymphocytic leukemia
C0023494|T191|SY|277545003|SNOMEDCT_CORE|TCLL - T-cell chronic lymphocytic leukemia|T-cell chronic lymphocytic leukemia
C0023510|T047|SY|54097007|SNOMEDCT_CORE|WBC diseases|White blood cell disorder
C0023510|T047|PT|54097007|SNOMEDCT_CORE|White blood cell disorder|White blood cell disorder
C0023510|T047|FN|54097007|SNOMEDCT_CORE|White blood cell disorder|White blood cell disorder
C0023510|T047|IS|54097007|SNOMEDCT_CORE|White blood cell disorder, NOS|White blood cell disorder
C0023518|T047|PTGB|111583006|SNOMEDCT_CORE|Leucocytosis|Leukocytosis
C0023518|T047|IS|111583006|SNOMEDCT_CORE|Leucocytosis, NOS|Leukocytosis
C0023518|T047|PT|111583006|SNOMEDCT_CORE|Leukocytosis|Leukocytosis
C0023518|T047|FN|111583006|SNOMEDCT_CORE|Leukocytosis|Leukocytosis
C0023518|T047|IS|111583006|SNOMEDCT_CORE|Leukocytosis, NOS|Leukocytosis
C0023530|T047|SYGB|84828003|SNOMEDCT_CORE|Leucocytopenia|Leukopenia
C0023530|T047|PTGB|84828003|SNOMEDCT_CORE|Leucopenia|Leukopenia
C0023530|T047|IS|84828003|SNOMEDCT_CORE|Leucopenia, NOS|Leukopenia
C0023530|T047|SY|84828003|SNOMEDCT_CORE|Leukocytopenia|Leukopenia
C0023530|T047|FN|84828003|SNOMEDCT_CORE|Leukopenia|Leukopenia
C0023530|T047|PT|84828003|SNOMEDCT_CORE|Leukopenia|Leukopenia
C0023530|T047|IS|84828003|SNOMEDCT_CORE|Leukopenia, NOS|Leukopenia
C0023531|T191|PTGB|274134003|SNOMEDCT_CORE|Leucoplakia|Leukoplakia
C0023531|T191|PT|274134003|SNOMEDCT_CORE|Leukoplakia|Leukoplakia
C0023531|T191|FN|274134003|SNOMEDCT_CORE|Leukoplakia|Leukoplakia
C0023532|T191|PTGB|414603003|SNOMEDCT_CORE|Leucoplakia of oral mucosa|Leukoplakia of oral mucosa
C0023532|T191|PT|414603003|SNOMEDCT_CORE|Leukoplakia of oral mucosa|Leukoplakia of oral mucosa
C0023532|T191|FN|414603003|SNOMEDCT_CORE|Leukoplakia of oral mucosa|Leukoplakia of oral mucosa
C0023646|T047|PT|4776004|SNOMEDCT_CORE|Lichen planus|Lichen planus
C0023646|T047|FN|4776004|SNOMEDCT_CORE|Lichen planus|Lichen planus
C0023646|T047|SY|4776004|SNOMEDCT_CORE|LP - Lichen planus|Lichen planus
C0023646|T047|SY|4776004|SNOMEDCT_CORE|Ruber planus|Lichen planus
C0023652|T047|SY|25674000|SNOMEDCT_CORE|Lichen sclerosus|Lichen sclerosus et atrophicus
C0023652|T047|PT|25674000|SNOMEDCT_CORE|Lichen sclerosus et atrophicus|Lichen sclerosus et atrophicus
C0023652|T047|FN|25674000|SNOMEDCT_CORE|Lichen sclerosus et atrophicus|Lichen sclerosus et atrophicus
C0023652|T047|IS|25674000|SNOMEDCT_CORE|Lichen sclerosus et atrophicus, NOS|Lichen sclerosus et atrophicus
C0023652|T047|SY|25674000|SNOMEDCT_CORE|White spot disease|Lichen sclerosus et atrophicus
C0023787|T047|SY|71325002|SNOMEDCT_CORE|Dystrophy of fatty tissue|Lipodystrophy
C0023787|T047|PT|71325002|SNOMEDCT_CORE|Lipodystrophy|Lipodystrophy
C0023787|T047|FN|71325002|SNOMEDCT_CORE|Lipodystrophy|Lipodystrophy
C0023787|T047|IS|71325002|SNOMEDCT_CORE|Lipodystrophy, NOS|Lipodystrophy
C0023798|T191|SY|93163002|SNOMEDCT_CORE|Lipoma|Lipoma
C0023798|T191|PT|93163002|SNOMEDCT_CORE|Lipoma|Lipoma
C0023798|T191|FN|93163002|SNOMEDCT_CORE|Lipoma|Lipoma
C0023798|T191|IS|93163002|SNOMEDCT_CORE|Lipoma of unspecified body site|Lipoma
C0023817|T047|SYGB|238086005|SNOMEDCT_CORE|Familial hyperlipoproteinaemia, type I|Familial lipoprotein lipase deficiency
C0023817|T047|SY|238086005|SNOMEDCT_CORE|Familial hyperlipoproteinemia, type I|Familial lipoprotein lipase deficiency
C0023817|T047|PT|238086005|SNOMEDCT_CORE|Familial lipoprotein lipase deficiency|Familial lipoprotein lipase deficiency
C0023817|T047|SYGB|238086005|SNOMEDCT_CORE|Fredrickson type I hyperlipoproteinaemia|Familial lipoprotein lipase deficiency
C0023817|T047|SY|238086005|SNOMEDCT_CORE|Fredrickson type I hyperlipoproteinemia|Familial lipoprotein lipase deficiency
C0023817|T047|FN|238086005|SNOMEDCT_CORE|Fredrickson type I hyperlipoproteinemia|Familial lipoprotein lipase deficiency
C0023827|T191|PT|254829001|SNOMEDCT_CORE|Liposarcoma|Liposarcoma
C0023827|T191|FN|254829001|SNOMEDCT_CORE|Liposarcoma|Liposarcoma
C0023882|T047|OAF|1178005|SNOMEDCT_CORE|Infantile spastic cerebral palsy|Infantile spastic cerebral palsy
C0023882|T047|OAP|1178005|SNOMEDCT_CORE|Infantile spastic cerebral palsy|Infantile spastic cerebral palsy
C0023882|T047|IS|1178005|SNOMEDCT_CORE|Little's disease|Infantile spastic cerebral palsy
C0023882|T047|IS|1178005|SNOMEDCT_CORE|Spastic infantile paralysis|Infantile spastic cerebral palsy
C0023885|T047|PT|27916005|SNOMEDCT_CORE|Abscess of liver|Abscess of liver
C0023885|T047|FN|27916005|SNOMEDCT_CORE|Abscess of liver|Abscess of liver
C0023885|T047|IS|27916005|SNOMEDCT_CORE|Abscess of liver, NOS|Abscess of liver
C0023885|T047|SY|27916005|SNOMEDCT_CORE|Hepatic abscess|Abscess of liver
C0023885|T047|IS|27916005|SNOMEDCT_CORE|Hepatic abscess, NOS|Abscess of liver
C0023890|T047|PT|19943007|SNOMEDCT_CORE|Cirrhosis of liver|Cirrhosis of liver
C0023890|T047|FN|19943007|SNOMEDCT_CORE|Cirrhosis of liver|Cirrhosis of liver
C0023890|T047|IS|19943007|SNOMEDCT_CORE|Cirrhosis of liver, NOS|Cirrhosis of liver
C0023890|T047|SY|19943007|SNOMEDCT_CORE|CL - Cirrhosis of liver|Cirrhosis of liver
C0023890|T047|SY|19943007|SNOMEDCT_CORE|Hepatic cirrhosis|Cirrhosis of liver
C0023890|T047|IS|19943007|SNOMEDCT_CORE|Hepatic cirrhosis, NOS|Cirrhosis of liver
C0023891|T047|PT|420054005|SNOMEDCT_CORE|Alcoholic cirrhosis|Alcoholic cirrhosis
C0023891|T047|FN|420054005|SNOMEDCT_CORE|Alcoholic cirrhosis|Alcoholic cirrhosis
C0023891|T047|SY|420054005|SNOMEDCT_CORE|Alcoholic cirrhosis of liver|Alcoholic cirrhosis
C0023891|T047|SY|420054005|SNOMEDCT_CORE|Alcoholic liver cirrhosis|Alcoholic cirrhosis
C0023892|T047|PT|1761006|SNOMEDCT_CORE|Biliary cirrhosis|Biliary cirrhosis
C0023892|T047|FN|1761006|SNOMEDCT_CORE|Biliary cirrhosis|Biliary cirrhosis
C0023892|T047|SY|1761006|SNOMEDCT_CORE|Cholangitic cirrhosis|Biliary cirrhosis
C0023892|T047|SY|1761006|SNOMEDCT_CORE|Cholestatic cirrhosis|Biliary cirrhosis
C0023895|T047|PT|235856003|SNOMEDCT_CORE|Disease of liver|Disease of liver
C0023895|T047|SY|235856003|SNOMEDCT_CORE|Disorder of liver|Disease of liver
C0023895|T047|FN|235856003|SNOMEDCT_CORE|Disorder of liver|Disease of liver
C0023895|T047|SY|235856003|SNOMEDCT_CORE|Hepatopathy|Disease of liver
C0023895|T047|SY|235856003|SNOMEDCT_CORE|LD - Liver disease|Disease of liver
C0023895|T047|SY|235856003|SNOMEDCT_CORE|Liver disease|Disease of liver
C0023896|T047|SY|41309000|SNOMEDCT_CORE|Alcoholic liver disease|ALD - Alcoholic liver disease
C0023896|T047|IS|41309000|SNOMEDCT_CORE|Alcoholic liver disease, NOS|ALD - Alcoholic liver disease
C0023896|T047|SY|41309000|SNOMEDCT_CORE|ALD - Alcoholic liver disease|ALD - Alcoholic liver disease
C0023903|T191|SY|126851005|SNOMEDCT_CORE|Hepatic tumor|Neoplasm of liver
C0023903|T191|SYGB|126851005|SNOMEDCT_CORE|Hepatic tumour|Neoplasm of liver
C0023903|T191|SY|126851005|SNOMEDCT_CORE|Hepatoma|Neoplasm of liver
C0023903|T191|PT|126851005|SNOMEDCT_CORE|Neoplasm of liver|Neoplasm of liver
C0023903|T191|FN|126851005|SNOMEDCT_CORE|Neoplasm of liver|Neoplasm of liver
C0023903|T191|SY|126851005|SNOMEDCT_CORE|Tumor of liver|Neoplasm of liver
C0023903|T191|SYGB|126851005|SNOMEDCT_CORE|Tumour of liver|Neoplasm of liver
C0024031|T184|SY|279039007|SNOMEDCT_CORE|LBP - Low back pain|Low back pain
C0024031|T184|PT|279039007|SNOMEDCT_CORE|Low back pain|Low back pain
C0024031|T184|FN|279039007|SNOMEDCT_CORE|Low back pain|Low back pain
C0024031|T184|OF|279039007|SNOMEDCT_CORE|Low back pain|Low back pain
C0024031|T184|SY|279039007|SNOMEDCT_CORE|Low back syndrome|Low back pain
C0024031|T184|SY|279039007|SNOMEDCT_CORE|Lumbago|Low back pain
C0024031|T184|SY|279039007|SNOMEDCT_CORE|Lumbalgia|Low back pain
C0024031|T184|SY|279039007|SNOMEDCT_CORE|Lumbar pain|Low back pain
C0024031|T184|SY|279039007|SNOMEDCT_CORE|Nonspecific pain in the lumbar region|Low back pain
C0024032|T033|SY|276610007|SNOMEDCT_CORE|Low birth weight|Low birth weight
C0024050|T046|SY|87763006|SNOMEDCT_CORE|Lower gastrointestinal bleeding|Lower gastrointestinal hemorrhage
C0024050|T046|PTGB|87763006|SNOMEDCT_CORE|Lower gastrointestinal haemorrhage|Lower gastrointestinal hemorrhage
C0024050|T046|PT|87763006|SNOMEDCT_CORE|Lower gastrointestinal hemorrhage|Lower gastrointestinal hemorrhage
C0024050|T046|FN|87763006|SNOMEDCT_CORE|Lower gastrointestinal hemorrhage|Lower gastrointestinal hemorrhage
C0024050|T046|SY|87763006|SNOMEDCT_CORE|Lower GI bleeding|Lower gastrointestinal hemorrhage
C0024050|T046|SYGB|87763006|SNOMEDCT_CORE|Lower GI haemorrhage|Lower gastrointestinal hemorrhage
C0024050|T046|SY|87763006|SNOMEDCT_CORE|Lower GI hemorrhage|Lower gastrointestinal hemorrhage
C0024050|T046|SYGB|87763006|SNOMEDCT_CORE|Lower GIT - gastrointestinal haemorrhage|Lower gastrointestinal hemorrhage
C0024050|T046|SY|87763006|SNOMEDCT_CORE|Lower GIT - gastrointestinal hemorrhage|Lower gastrointestinal hemorrhage
C0024103|T033|SY|89164003|SNOMEDCT_CORE|Breast irregular nodularity|Breast lump
C0024103|T033|PT|89164003|SNOMEDCT_CORE|Breast lump|Breast lump
C0024103|T033|FN|89164003|SNOMEDCT_CORE|Breast lump|Breast lump
C0024103|T033|SY|89164003|SNOMEDCT_CORE|Breast mass|Breast lump
C0024103|T033|IS|89164003|SNOMEDCT_CORE|Lump in breast|Breast lump
C0024103|T033|SY|89164003|SNOMEDCT_CORE|Lumpy breast|Breast lump
C0024103|T033|SY|89164003|SNOMEDCT_CORE|Lumpy breasts|Breast lump
C0024103|T033|SY|89164003|SNOMEDCT_CORE|Mass in breast|Breast lump
C0024110|T047|PT|73452002|SNOMEDCT_CORE|Abscess of lung|Abscess of lung
C0024110|T047|FN|73452002|SNOMEDCT_CORE|Abscess of lung|Abscess of lung
C0024115|T047|IS|19829001|SNOMEDCT_CORE|Disease of lung|Disorder of lung
C0024115|T047|OF|19829001|SNOMEDCT_CORE|Disease of lung|Disorder of lung
C0024115|T047|IS|19829001|SNOMEDCT_CORE|Disease of lung, NOS|Disorder of lung
C0024115|T047|PT|19829001|SNOMEDCT_CORE|Disorder of lung|Disorder of lung
C0024115|T047|FN|19829001|SNOMEDCT_CORE|Disorder of lung|Disorder of lung
C0024115|T047|SY|19829001|SNOMEDCT_CORE|Lung disorder|Disorder of lung
C0024115|T047|IS|19829001|SNOMEDCT_CORE|Lung disorder, NOS|Disorder of lung
C0024115|T047|SY|19829001|SNOMEDCT_CORE|Pulmonary disease|Disorder of lung
C0024115|T047|IS|19829001|SNOMEDCT_CORE|Pulmonary disease, NOS|Disorder of lung
C0024117|T047|SY|13645005|SNOMEDCT_CORE|CAFL - Chronic airflow limitation|Chronic obstructive lung disease
C0024117|T047|SY|13645005|SNOMEDCT_CORE|CAL - Chronic airflow limitation|Chronic obstructive lung disease
C0024117|T047|SY|13645005|SNOMEDCT_CORE|Chronic airflow limitation|Chronic obstructive lung disease
C0024117|T047|SY|13645005|SNOMEDCT_CORE|Chronic airway disease|Chronic obstructive lung disease
C0024117|T047|SY|13645005|SNOMEDCT_CORE|Chronic airway obstruction|Chronic obstructive lung disease
C0024117|T047|SY|13645005|SNOMEDCT_CORE|Chronic irreversible airway obstruction|Chronic obstructive lung disease
C0024117|T047|SY|13645005|SNOMEDCT_CORE|Chronic obstructive airway disease|Chronic obstructive lung disease
C0024117|T047|PT|13645005|SNOMEDCT_CORE|Chronic obstructive lung disease|Chronic obstructive lung disease
C0024117|T047|FN|13645005|SNOMEDCT_CORE|Chronic obstructive lung disease|Chronic obstructive lung disease
C0024117|T047|IS|13645005|SNOMEDCT_CORE|Chronic obstructive lung disease, NOS|Chronic obstructive lung disease
C0024117|T047|SY|13645005|SNOMEDCT_CORE|Chronic obstructive pulmonary disease|Chronic obstructive lung disease
C0024117|T047|SY|13645005|SNOMEDCT_CORE|COAD - Chronic obstructive airways disease|Chronic obstructive lung disease
C0024117|T047|IS|13645005|SNOMEDCT_CORE|COLD|Chronic obstructive lung disease
C0024117|T047|SY|13645005|SNOMEDCT_CORE|COLD - Chronic obstructive lung disease|Chronic obstructive lung disease
C0024117|T047|IS|13645005|SNOMEDCT_CORE|COPD|Chronic obstructive lung disease
C0024117|T047|SY|13645005|SNOMEDCT_CORE|COPD - Chronic obstructive pulmonary disease|Chronic obstructive lung disease
C0024121|T191|PT|126713003|SNOMEDCT_CORE|Neoplasm of lung|Neoplasm of lung
C0024121|T191|FN|126713003|SNOMEDCT_CORE|Neoplasm of lung|Neoplasm of lung
C0024121|T191|SY|126713003|SNOMEDCT_CORE|Tumor of lung|Neoplasm of lung
C0024121|T191|SYGB|126713003|SNOMEDCT_CORE|Tumour of lung|Neoplasm of lung
C0024131|T047|SY|10528009|SNOMEDCT_CORE|Lupus exedens|Lupus vulgaris
C0024131|T047|PT|10528009|SNOMEDCT_CORE|Lupus vulgaris|Lupus vulgaris
C0024131|T047|FN|10528009|SNOMEDCT_CORE|Lupus vulgaris|Lupus vulgaris
C0024131|T047|SY|10528009|SNOMEDCT_CORE|LV - Lupus vulgaris|Lupus vulgaris
C0024131|T047|SY|10528009|SNOMEDCT_CORE|Tuberculosis cutis luposa|Lupus vulgaris
C0024131|T047|SY|10528009|SNOMEDCT_CORE|Tuberculosis luposa cutis|Lupus vulgaris
C0024131|T047|SY|10528009|SNOMEDCT_CORE|Tuberculosis lupus exedens|Lupus vulgaris
C0024138|T047|PT|200938002|SNOMEDCT_CORE|Discoid lupus erythematosus|Discoid lupus erythematosus
C0024138|T047|FN|200938002|SNOMEDCT_CORE|Discoid lupus erythematosus|Discoid lupus erythematosus
C0024138|T047|SY|200938002|SNOMEDCT_CORE|DLE - Discoid lupus erythematosus|Discoid lupus erythematosus
C0024138|T047|SY|200938002|SNOMEDCT_CORE|LE - Discoid lupus erythematosus|Discoid lupus erythematosus
C0024141|T047|SY|55464009|SNOMEDCT_CORE|Disseminated lupus erythematosus|Systemic lupus erythematosus
C0024141|T047|IS|55464009|SNOMEDCT_CORE|SLE|Systemic lupus erythematosus
C0024141|T047|SY|55464009|SNOMEDCT_CORE|SLE - Systemic lupus erythematosus|Systemic lupus erythematosus
C0024141|T047|PT|55464009|SNOMEDCT_CORE|Systemic lupus erythematosus|Systemic lupus erythematosus
C0024141|T047|FN|55464009|SNOMEDCT_CORE|Systemic lupus erythematosus|Systemic lupus erythematosus
C0024143|T047|SY|68815009|SNOMEDCT_CORE|Lupus nephritis|SLE glomerulonephritis syndrome
C0024143|T047|IS|68815009|SNOMEDCT_CORE|Lupus nephritis, NOS|SLE glomerulonephritis syndrome
C0024143|T047|PT|68815009|SNOMEDCT_CORE|SLE glomerulonephritis syndrome|SLE glomerulonephritis syndrome
C0024143|T047|OF|68815009|SNOMEDCT_CORE|SLE glomerulonephritis syndrome|SLE glomerulonephritis syndrome
C0024143|T047|IS|68815009|SNOMEDCT_CORE|SLE glomerulonephritis syndrome, NOS|SLE glomerulonephritis syndrome
C0024143|T047|FN|68815009|SNOMEDCT_CORE|Systemic lupus erythematosus glomerulonephritis syndrome|SLE glomerulonephritis syndrome
C0024143|T047|SY|68815009|SNOMEDCT_CORE|Systemic lupus erythematosus glomerulonephritis syndrome|SLE glomerulonephritis syndrome
C0024198|T047|IS|23502006|SNOMEDCT_CORE|Infection by Borrelia burgdorferi|Lyme disease
C0024198|T047|SY|23502006|SNOMEDCT_CORE|Infection due to Borrelia burgdorferi sensu lato|Lyme disease
C0024198|T047|SY|23502006|SNOMEDCT_CORE|Lyme borreliosis|Lyme disease
C0024198|T047|PT|23502006|SNOMEDCT_CORE|Lyme disease|Lyme disease
C0024198|T047|FN|23502006|SNOMEDCT_CORE|Lyme disease|Lyme disease
C0024198|T047|SY|23502006|SNOMEDCT_CORE|Steere's disease|Lyme disease
C0024205|T047|SY|19471005|SNOMEDCT_CORE|Adenitis|Lymphadenitis
C0024205|T047|IS|19471005|SNOMEDCT_CORE|Adenitis, NOS|Lymphadenitis
C0024205|T047|SY|19471005|SNOMEDCT_CORE|Inflammation of lymph node|Lymphadenitis
C0024205|T047|PT|19471005|SNOMEDCT_CORE|Lymphadenitis|Lymphadenitis
C0024205|T047|FN|19471005|SNOMEDCT_CORE|Lymphadenitis|Lymphadenitis
C0024205|T047|IS|19471005|SNOMEDCT_CORE|Lymphadenitis, NOS|Lymphadenitis
C0024221|T191|PT|400178008|SNOMEDCT_CORE|Lymphangioma|Lymphangioma
C0024221|T191|FN|400178008|SNOMEDCT_CORE|Lymphangioma|Lymphangioma
C0024225|T047|SY|1415005|SNOMEDCT_CORE|Inflammation of lymphatics|Lymphangitis
C0024225|T047|PT|1415005|SNOMEDCT_CORE|Lymphangitis|Lymphangitis
C0024225|T047|FN|1415005|SNOMEDCT_CORE|Lymphangitis|Lymphangitis
C0024225|T047|IS|1415005|SNOMEDCT_CORE|Lymphangitis, NOS|Lymphangitis
C0024228|T047|FN|362971004|SNOMEDCT_CORE|Disorder of lymphatic system|Disorder of lymphatic system
C0024228|T047|PT|362971004|SNOMEDCT_CORE|Disorder of lymphatic system|Disorder of lymphatic system
C0024236|T046|SY|234097001|SNOMEDCT_CORE|Lymphatic edema|Lymphedema
C0024236|T046|SYGB|234097001|SNOMEDCT_CORE|Lymphatic oedema|Lymphedema
C0024236|T046|PT|234097001|SNOMEDCT_CORE|Lymphedema|Lymphedema
C0024236|T046|FN|234097001|SNOMEDCT_CORE|Lymphedema|Lymphedema
C0024236|T046|PTGB|234097001|SNOMEDCT_CORE|Lymphoedema|Lymphedema
C0024248|T047|PT|234109007|SNOMEDCT_CORE|Lymphocele|Lymphocele
C0024248|T047|FN|234109007|SNOMEDCT_CORE|Lymphocele|Lymphocele
C0024282|T047|PT|67023009|SNOMEDCT_CORE|Lymphocytosis|Lymphocytosis
C0024282|T047|FN|67023009|SNOMEDCT_CORE|Lymphocytosis|Lymphocytosis
C0024282|T047|IS|67023009|SNOMEDCT_CORE|Lymphocytosis, NOS|Lymphocytosis
C0024299|T191|SY|118600007|SNOMEDCT_CORE|Lymphoma|Malignant lymphoma
C0024299|T191|IS|118600007|SNOMEDCT_CORE|Lymphoma|Malignant lymphoma
C0024299|T191|PT|118600007|SNOMEDCT_CORE|Malignant lymphoma|Malignant lymphoma
C0024299|T191|OP|118600007|SNOMEDCT_CORE|Malignant lymphoma|Malignant lymphoma
C0024299|T191|FN|118600007|SNOMEDCT_CORE|Malignant lymphoma|Malignant lymphoma
C0024301|T191|PT|269476000|SNOMEDCT_CORE|Nodular lymphoma|Nodular lymphoma
C0024301|T191|FN|269476000|SNOMEDCT_CORE|Nodular lymphoma|Nodular lymphoma
C0024302|T191|PT|373168002|SNOMEDCT_CORE|Reticulosarcoma|Reticulosarcoma
C0024302|T191|FN|373168002|SNOMEDCT_CORE|Reticulosarcoma|Reticulosarcoma
C0024302|T191|SY|373168002|SNOMEDCT_CORE|Reticulum cell sarcoma|Reticulosarcoma
C0024305|T191|SY|118601006|SNOMEDCT_CORE|Malignant lymphoma, non-Hodgkin's type|Non-Hodgkin's lymphoma
C0024305|T191|SY|118601006|SNOMEDCT_CORE|NHL - Non-Hodgkin's lymphoma|Non-Hodgkin's lymphoma
C0024305|T191|SY|118601006|SNOMEDCT_CORE|Non-Hodgkin lymphoma|Non-Hodgkin's lymphoma
C0024305|T191|SY|118601006|SNOMEDCT_CORE|Non-Hodgkin's lymphoma|Non-Hodgkin's lymphoma
C0024305|T191|PT|118601006|SNOMEDCT_CORE|Non-Hodgkin's lymphoma|Non-Hodgkin's lymphoma
C0024305|T191|FN|118601006|SNOMEDCT_CORE|Non-Hodgkin's lymphoma|Non-Hodgkin's lymphoma
C0024305|T191|SY|118601006|SNOMEDCT_CORE|Non-Hodgkin's lymphoma - disorder|Non-Hodgkin's lymphoma
C0024312|T047|PT|48813009|SNOMEDCT_CORE|Lymphocytopenia|Lymphocytopenia
C0024312|T047|FN|48813009|SNOMEDCT_CORE|Lymphocytopenia|Lymphocytopenia
C0024312|T047|IS|48813009|SNOMEDCT_CORE|Lymphocytopenia, NOS|Lymphocytopenia
C0024312|T047|SY|48813009|SNOMEDCT_CORE|Lymphopenia|Lymphocytopenia
C0024314|T191|PT|277466009|SNOMEDCT_CORE|Lymphoproliferative disorder|Lymphoproliferative disorder
C0024314|T191|FN|277466009|SNOMEDCT_CORE|Lymphoproliferative disorder|Lymphoproliferative disorder
C0024419|T191|PTGB|190818004|SNOMEDCT_CORE|Waldenström macroglobulinaemia|Waldenström macroglobulinemia
C0024419|T191|PT|190818004|SNOMEDCT_CORE|Waldenström macroglobulinemia|Waldenström macroglobulinemia
C0024419|T191|FN|190818004|SNOMEDCT_CORE|Waldenström macroglobulinemia|Waldenström macroglobulinemia
C0024419|T191|SYGB|190818004|SNOMEDCT_CORE|Waldenstrom's macroglobulinaemia|Waldenström macroglobulinemia
C0024419|T191|SY|190818004|SNOMEDCT_CORE|Waldenstrom's macroglobulinemia|Waldenström macroglobulinemia
C0024419|T191|OF|190818004|SNOMEDCT_CORE|Waldenstrom's macroglobulinemia|Waldenström macroglobulinemia
C0024437|T047|FN|422338006|SNOMEDCT_CORE|Degenerative disorder of macula|Degenerative disorder of macula
C0024437|T047|PT|422338006|SNOMEDCT_CORE|Degenerative disorder of macula|Degenerative disorder of macula
C0024440|T047|SY|193387007|SNOMEDCT_CORE|CME - cystoid macular edema|Cystoid macular edema
C0024440|T047|IS|193387007|SNOMEDCT_CORE|CME - cystoid macular oedema|Cystoid macular edema
C0024440|T047|IS|193387007|SNOMEDCT_CORE|CMO - cystoid macular edema|Cystoid macular edema
C0024440|T047|SYGB|193387007|SNOMEDCT_CORE|CMO - cystoid macular oedema|Cystoid macular edema
C0024440|T047|PT|193387007|SNOMEDCT_CORE|Cystoid macular edema|Cystoid macular edema
C0024440|T047|FN|193387007|SNOMEDCT_CORE|Cystoid macular edema|Cystoid macular edema
C0024440|T047|PTGB|193387007|SNOMEDCT_CORE|Cystoid macular oedema|Cystoid macular edema
C0024441|T047|PT|232006002|SNOMEDCT_CORE|Macular hole|Macular hole
C0024441|T047|FN|232006002|SNOMEDCT_CORE|Macular hole|Macular hole
C0024517|T048|PT|36923009|SNOMEDCT_CORE|Major depression, single episode|Major depression, single episode
C0024517|T048|FN|36923009|SNOMEDCT_CORE|Major depression, single episode|Major depression, single episode
C0024517|T048|IS|36923009|SNOMEDCT_CORE|Major depression, single episode, NOS|Major depression, single episode
C0024517|T048|SY|36923009|SNOMEDCT_CORE|Major depressive disorder, single episode|Major depression, single episode
C0024517|T048|OAF|268620009|SNOMEDCT_CORE|Single major depressive episode|Major depression, single episode
C0024517|T048|OAP|268620009|SNOMEDCT_CORE|Single major depressive episode|Major depression, single episode
C0024523|T047|IS|32230006|SNOMEDCT_CORE|Intestinal malabsorption|Malabsorption syndrome
C0024523|T047|IS|32230006|SNOMEDCT_CORE|Intestinal malabsorption, NOS|Malabsorption syndrome
C0024523|T047|SY|32230006|SNOMEDCT_CORE|Malabsorption|Malabsorption syndrome
C0024523|T047|PT|32230006|SNOMEDCT_CORE|Malabsorption syndrome|Malabsorption syndrome
C0024523|T047|FN|32230006|SNOMEDCT_CORE|Malabsorption syndrome|Malabsorption syndrome
C0024523|T047|IS|32230006|SNOMEDCT_CORE|Malabsorption syndrome, NOS|Malabsorption syndrome
C0024523|T047|IS|32230006|SNOMEDCT_CORE|Malabsorption, NOS|Malabsorption syndrome
C0024528|T184|PT|271795006|SNOMEDCT_CORE|Malaise and fatigue|Malaise and fatigue
C0024528|T184|FN|271795006|SNOMEDCT_CORE|Malaise and fatigue|Malaise and fatigue
C0024530|T047|PT|61462000|SNOMEDCT_CORE|Malaria|Malaria
C0024530|T047|FN|61462000|SNOMEDCT_CORE|Malaria|Malaria
C0024530|T047|IS|61462000|SNOMEDCT_CORE|Malaria, NOS|Malaria
C0024530|T047|SY|61462000|SNOMEDCT_CORE|Paludism|Malaria
C0024530|T047|SY|61462000|SNOMEDCT_CORE|Plasmodiosis|Malaria
C0024586|T047|PT|35868009|SNOMEDCT_CORE|Carcinoid syndrome|Carcinoid syndrome
C0024586|T047|FN|35868009|SNOMEDCT_CORE|Carcinoid syndrome|Carcinoid syndrome
C0024586|T047|SY|35868009|SNOMEDCT_CORE|Excessive serotonin secretion|Carcinoid syndrome
C0024586|T047|SY|35868009|SNOMEDCT_CORE|Hormonal tumor|Carcinoid syndrome
C0024586|T047|SYGB|35868009|SNOMEDCT_CORE|Hormonal tumour|Carcinoid syndrome
C0024586|T047|SY|35868009|SNOMEDCT_CORE|Hormone secretion by carcinoid tumor|Carcinoid syndrome
C0024586|T047|SYGB|35868009|SNOMEDCT_CORE|Hormone secretion by carcinoid tumour|Carcinoid syndrome
C0024586|T047|IS|35868009|SNOMEDCT_CORE|Serotonin syndrome|Carcinoid syndrome
C0024588|T047|SY|78975002|SNOMEDCT_CORE|Accelerated essential hypertension|Malignant essential hypertension
C0024588|T047|PT|78975002|SNOMEDCT_CORE|Malignant essential hypertension|Malignant essential hypertension
C0024588|T047|FN|78975002|SNOMEDCT_CORE|Malignant essential hypertension|Malignant essential hypertension
C0024620|T191|SY|95214007|SNOMEDCT_CORE|Ca liver - primary|Primary malignant neoplasm of liver
C0024620|T191|IS|93870000|SNOMEDCT_CORE|Primary malignant neoplasm of liver|Primary malignant neoplasm of liver
C0024620|T191|PT|95214007|SNOMEDCT_CORE|Primary malignant neoplasm of liver|Primary malignant neoplasm of liver
C0024620|T191|FN|95214007|SNOMEDCT_CORE|Primary malignant neoplasm of liver|Primary malignant neoplasm of liver
C0024623|T191|SY|363349007|SNOMEDCT_CORE|CA - Cancer of stomach|Malignant tumor of stomach
C0024623|T191|SY|363349007|SNOMEDCT_CORE|Cancer of stomach|Malignant tumor of stomach
C0024623|T191|SY|363349007|SNOMEDCT_CORE|Gastric cancer|Malignant tumor of stomach
C0024623|T191|PT|363349007|SNOMEDCT_CORE|Malignant tumor of stomach|Malignant tumor of stomach
C0024623|T191|FN|363349007|SNOMEDCT_CORE|Malignant tumor of stomach|Malignant tumor of stomach
C0024623|T191|PTGB|363349007|SNOMEDCT_CORE|Malignant tumour of stomach|Malignant tumor of stomach
C0024633|T047|IS|35265002|SNOMEDCT_CORE|Gastresophageal laceration-hemorrhage syndrome|Mallory-Weiss syndrome
C0024633|T047|SY|35265002|SNOMEDCT_CORE|Gastro-esophageal laceration-hemorrhage syndrome|Mallory-Weiss syndrome
C0024633|T047|SYGB|35265002|SNOMEDCT_CORE|Gastro-oesophageal laceration-haemorrhage syndrome|Mallory-Weiss syndrome
C0024633|T047|SY|35265002|SNOMEDCT_CORE|Gastroesophageal laceration-hemorrhage syndrome|Mallory-Weiss syndrome
C0024633|T047|SYGB|35265002|SNOMEDCT_CORE|Gastrooesophageal laceration-hemorrhage syndrome|Mallory-Weiss syndrome
C0024633|T047|PT|35265002|SNOMEDCT_CORE|Mallory-Weiss syndrome|Mallory-Weiss syndrome
C0024633|T047|FN|35265002|SNOMEDCT_CORE|Mallory-Weiss syndrome|Mallory-Weiss syndrome
C0024636|T190|SY|47944004|SNOMEDCT_CORE|Malocclusion|Malocclusion of teeth
C0024636|T190|PT|47944004|SNOMEDCT_CORE|Malocclusion of teeth|Malocclusion of teeth
C0024636|T190|FN|47944004|SNOMEDCT_CORE|Malocclusion of teeth|Malocclusion of teeth
C0024636|T190|IS|47944004|SNOMEDCT_CORE|Malocclusion of teeth, NOS|Malocclusion of teeth
C0024636|T190|IS|47944004|SNOMEDCT_CORE|Malocclusion, NOS|Malocclusion of teeth
C0024692|T037|SY|263172003|SNOMEDCT_CORE|Fracture of lower jaw|Fracture of mandible
C0024692|T037|PT|263172003|SNOMEDCT_CORE|Fracture of mandible|Fracture of mandible
C0024692|T037|FN|263172003|SNOMEDCT_CORE|Fracture of mandible|Fracture of mandible
C0024713|T048|IS|68569003|SNOMEDCT_CORE|Bipolar I disorder, most recent episode manic|Manic bipolar I disorder
C0024713|T048|IS|68569003|SNOMEDCT_CORE|Manic bipolar disorder, NOS|Manic bipolar I disorder
C0024713|T048|PT|68569003|SNOMEDCT_CORE|Manic bipolar I disorder|Manic bipolar I disorder
C0024713|T048|FN|68569003|SNOMEDCT_CORE|Manic bipolar I disorder|Manic bipolar I disorder
C0024713|T048|IS|68569003|SNOMEDCT_CORE|Manic bipolar I disorder, NOS|Manic bipolar I disorder
C0024790|T047|SY|1963002|SNOMEDCT_CORE|Marchiafava-Micheli syndrome|Paroxysmal nocturnal hemoglobinuria
C0024790|T047|IS|1963002|SNOMEDCT_CORE|Paroxysmal noctural hemoglobinuria|Paroxysmal nocturnal hemoglobinuria
C0024790|T047|PTGB|1963002|SNOMEDCT_CORE|Paroxysmal nocturnal haemoglobinuria|Paroxysmal nocturnal hemoglobinuria
C0024790|T047|PT|1963002|SNOMEDCT_CORE|Paroxysmal nocturnal hemoglobinuria|Paroxysmal nocturnal hemoglobinuria
C0024790|T047|FN|1963002|SNOMEDCT_CORE|Paroxysmal nocturnal hemoglobinuria|Paroxysmal nocturnal hemoglobinuria
C0024790|T047|SY|1963002|SNOMEDCT_CORE|PNH|Paroxysmal nocturnal hemoglobinuria
C0024790|T047|SYGB|1963002|SNOMEDCT_CORE|PNH - Paroxysmal nocturnal haemoglobinuria|Paroxysmal nocturnal hemoglobinuria
C0024790|T047|SY|1963002|SNOMEDCT_CORE|PNH - Paroxysmal nocturnal hemoglobinuria|Paroxysmal nocturnal hemoglobinuria
C0024796|T047|SY|19346006|SNOMEDCT_CORE|Marfan syndrome|Marfan's syndrome
C0024796|T047|SY|19346006|SNOMEDCT_CORE|Marfan's disease|Marfan's syndrome
C0024796|T047|PT|19346006|SNOMEDCT_CORE|Marfan's syndrome|Marfan's syndrome
C0024796|T047|FN|19346006|SNOMEDCT_CORE|Marfan's syndrome|Marfan's syndrome
C0024894|T047|OAP|45198002|SNOMEDCT_CORE|Mastitis|Mastitis
C0024894|T047|OAF|45198002|SNOMEDCT_CORE|Mastitis|Mastitis
C0024894|T047|IS|45198002|SNOMEDCT_CORE|Mastitis, NOS|Mastitis
C0024902|T184|SY|53430007|SNOMEDCT_CORE|Breast pain|Pain of breast
C0024902|T184|SY|53430007|SNOMEDCT_CORE|Breast painful|Pain of breast
C0024902|T184|SY|53430007|SNOMEDCT_CORE|Mastalgia|Pain of breast
C0024902|T184|SY|53430007|SNOMEDCT_CORE|Mastodynia|Pain of breast
C0024902|T184|SY|53430007|SNOMEDCT_CORE|Pain in the breast|Pain of breast
C0024902|T184|PT|53430007|SNOMEDCT_CORE|Pain of breast|Pain of breast
C0024902|T184|FN|53430007|SNOMEDCT_CORE|Pain of breast|Pain of breast
C0024902|T184|SY|53430007|SNOMEDCT_CORE|Painful breasts|Pain of breast
C0024904|T047|PT|52404001|SNOMEDCT_CORE|Mastoiditis|Mastoiditis
C0024904|T047|FN|52404001|SNOMEDCT_CORE|Mastoiditis|Mastoiditis
C0024904|T047|IS|52404001|SNOMEDCT_CORE|Mastoiditis, NOS|Mastoiditis
C0025007|T047|PT|14189004|SNOMEDCT_CORE|Measles|Measles
C0025007|T047|FN|14189004|SNOMEDCT_CORE|Measles|Measles
C0025007|T047|SY|14189004|SNOMEDCT_CORE|Morbilli|Measles
C0025007|T047|SY|14189004|SNOMEDCT_CORE|Rubeola|Measles
C0025037|T019|SY|37373007|SNOMEDCT_CORE|MD - Meckel's diverticulum|Meckel's diverticulum
C0025037|T019|SY|37373007|SNOMEDCT_CORE|Meckel diverticulum|Meckel's diverticulum
C0025037|T019|PT|37373007|SNOMEDCT_CORE|Meckel's diverticulum|Meckel's diverticulum
C0025037|T019|FN|37373007|SNOMEDCT_CORE|Meckel's diverticulum|Meckel's diverticulum
C0025037|T019|SY|37373007|SNOMEDCT_CORE|Persistent intestinal end of vitelline duct|Meckel's diverticulum
C0025037|T019|SY|37373007|SNOMEDCT_CORE|Persistent omphalomesenteric duct|Meckel's diverticulum
C0025037|T019|SY|37373007|SNOMEDCT_CORE|Persistent vitelline duct|Meckel's diverticulum
C0025048|T047|SY|206292002|SNOMEDCT_CORE|MAS - Meconium aspiration syndrome|Meconium aspiration syndrome
C0025048|T047|PT|206292002|SNOMEDCT_CORE|Meconium aspiration syndrome|Meconium aspiration syndrome
C0025048|T047|FN|206292002|SNOMEDCT_CORE|Meconium aspiration syndrome|Meconium aspiration syndrome
C0025062|T047|PT|16838000|SNOMEDCT_CORE|Mediastinal emphysema|Mediastinal emphysema
C0025062|T047|FN|16838000|SNOMEDCT_CORE|Mediastinal emphysema|Mediastinal emphysema
C0025062|T047|SY|16838000|SNOMEDCT_CORE|Pneumomediastinum|Mediastinal emphysema
C0025063|T191|IS|94147001|SNOMEDCT_CORE|Tumor of mediastinum|Tumor of mediastinum
C0025063|T191|IS|94147001|SNOMEDCT_CORE|Tumour of mediastinum|Tumor of mediastinum
C0025149|T191|SY|83217000|SNOMEDCT_CORE|MDB - Medulloblastoma|Medulloblastoma
C0025149|T191|PT|443333004|SNOMEDCT_CORE|Medulloblastoma|Medulloblastoma
C0025149|T191|PT|83217000|SNOMEDCT_CORE|Medulloblastoma|Medulloblastoma
C0025149|T191|OF|83217000|SNOMEDCT_CORE|Medulloblastoma|Medulloblastoma
C0025149|T191|FN|443333004|SNOMEDCT_CORE|Medulloblastoma|Medulloblastoma
C0025149|T191|SY|83217000|SNOMEDCT_CORE|Medulloblastoma, no ICD-O subtype|Medulloblastoma
C0025149|T191|OF|83217000|SNOMEDCT_CORE|Medulloblastoma, no ICD-O subtype|Medulloblastoma
C0025149|T191|FN|83217000|SNOMEDCT_CORE|Medulloblastoma, no International Classification of Diseases for Oncology subtype|Medulloblastoma
C0025149|T191|SY|83217000|SNOMEDCT_CORE|Medulloblastoma, no International Classification of Diseases for Oncology subtype|Medulloblastoma
C0025149|T191|IS|83217000|SNOMEDCT_CORE|Medulloblastoma, NOS|Medulloblastoma
C0025183|T047|SY|230325003|SNOMEDCT_CORE|Blepharospasm - oromandibular dystonia|Meige syndrome
C0025183|T047|SY|230325003|SNOMEDCT_CORE|Brueghel syndrome|Meige syndrome
C0025183|T047|PT|230325003|SNOMEDCT_CORE|Meige syndrome|Meige syndrome
C0025183|T047|FN|230325003|SNOMEDCT_CORE|Meige syndrome|Meige syndrome
C0025193|T048|IS|35489007|SNOMEDCT_CORE|Melancholia|Melancholia
C0025193|T048|IS|35489007|SNOMEDCT_CORE|Melancholia, NOS|Melancholia
C0025202|T191|PT|372244006|SNOMEDCT_CORE|Malignant melanoma|Malignant melanoma
C0025202|T191|FN|372244006|SNOMEDCT_CORE|Malignant melanoma|Malignant melanoma
C0025202|T191|SY|372244006|SNOMEDCT_CORE|Melanosarcoma|Malignant melanoma
C0025218|T047|PT|36209000|SNOMEDCT_CORE|Chloasma|Chloasma
C0025218|T047|FN|36209000|SNOMEDCT_CORE|Chloasma|Chloasma
C0025218|T047|IS|36209000|SNOMEDCT_CORE|Chloasma, NOS|Chloasma
C0025218|T047|SY|36209000|SNOMEDCT_CORE|Melasma|Chloasma
C0025218|T047|IS|36209000|SNOMEDCT_CORE|Melasma, NOS|Chloasma
C0025222|T046|SY|2901004|SNOMEDCT_CORE|Altered blood in stool|Melena
C0025222|T046|SY|2901004|SNOMEDCT_CORE|Altered blood passed per rectum|Melena
C0025222|T046|SY|2901004|SNOMEDCT_CORE|Black, tarry stool|Melena
C0025222|T046|PTGB|2901004|SNOMEDCT_CORE|Melaena|Melena
C0025222|T046|PT|2901004|SNOMEDCT_CORE|Melena|Melena
C0025222|T046|FN|2901004|SNOMEDCT_CORE|Melena|Melena
C0025222|T046|SY|2901004|SNOMEDCT_CORE|Tarry stools|Melena
C0025267|T191|SY|30664006|SNOMEDCT_CORE|MEA, type 1|Multiple endocrine neoplasia, type 1
C0025267|T191|SY|30664006|SNOMEDCT_CORE|MEN 1 - Multiple endocrine neoplasia syndrome type 1|Multiple endocrine neoplasia, type 1
C0025267|T191|SY|30664006|SNOMEDCT_CORE|MEN 1 syndrome|Multiple endocrine neoplasia, type 1
C0025267|T191|SY|30664006|SNOMEDCT_CORE|MEN, type 1|Multiple endocrine neoplasia, type 1
C0025267|T191|SY|30664006|SNOMEDCT_CORE|Multiple endocrine adenomatosis, type 1|Multiple endocrine neoplasia, type 1
C0025267|T191|SY|30664006|SNOMEDCT_CORE|Multiple endocrine neoplasia syndrome type 1|Multiple endocrine neoplasia, type 1
C0025267|T191|PT|30664006|SNOMEDCT_CORE|Multiple endocrine neoplasia, type 1|Multiple endocrine neoplasia, type 1
C0025267|T191|FN|30664006|SNOMEDCT_CORE|Multiple endocrine neoplasia, type 1|Multiple endocrine neoplasia, type 1
C0025267|T191|SY|30664006|SNOMEDCT_CORE|Wermer syndrome|Multiple endocrine neoplasia, type 1
C0025281|T047|SY|13445001|SNOMEDCT_CORE|Auditory vertigo|Ménière's disease
C0025281|T047|SY|13445001|SNOMEDCT_CORE|Meniere disease|Ménière's disease
C0025281|T047|SY|13445001|SNOMEDCT_CORE|Meniere disorder|Ménière's disease
C0025281|T047|SY|13445001|SNOMEDCT_CORE|Meniere syndrome|Ménière's disease
C0025281|T047|PT|13445001|SNOMEDCT_CORE|Ménière's disease|Ménière's disease
C0025281|T047|FN|13445001|SNOMEDCT_CORE|Ménière's disease|Ménière's disease
C0025281|T047|IS|13445001|SNOMEDCT_CORE|Meniere's disease, NOS|Ménière's disease
C0025281|T047|SY|13445001|SNOMEDCT_CORE|Ménière's syndrome|Ménière's disease
C0025281|T047|IS|13445001|SNOMEDCT_CORE|Ménière's syndrome, NOS|Ménière's disease
C0025281|T047|SY|13445001|SNOMEDCT_CORE|Ménière's vertigo|Ménière's disease
C0025281|T047|IS|13445001|SNOMEDCT_CORE|Meniere's vertigo, NOS|Ménière's disease
C0025281|T047|SY|13445001|SNOMEDCT_CORE|Menieres disease|Ménière's disease
C0025281|T047|SY|13445001|SNOMEDCT_CORE|Otogenic vertigo|Ménière's disease
C0025289|T047|PT|7180009|SNOMEDCT_CORE|Meningitis|Meningitis
C0025289|T047|FN|7180009|SNOMEDCT_CORE|Meningitis|Meningitis
C0025289|T047|IS|7180009|SNOMEDCT_CORE|Meningitis, NOS|Meningitis
C0025290|T047|IS|58170007|SNOMEDCT_CORE|Aseptic meningitis|Aseptic meningitis
C0025297|T047|SY|58170007|SNOMEDCT_CORE|Abacterial meningitis|Viral meningitis
C0025297|T047|SY|58170007|SNOMEDCT_CORE|Aseptic meningitis, viral|Viral meningitis
C0025297|T047|SY|58170007|SNOMEDCT_CORE|Meningitis, viral|Viral meningitis
C0025297|T047|PT|58170007|SNOMEDCT_CORE|Viral meningitis|Viral meningitis
C0025297|T047|FN|58170007|SNOMEDCT_CORE|Viral meningitis|Viral meningitis
C0025297|T047|IS|58170007|SNOMEDCT_CORE|Viral meningitis NOS|Viral meningitis
C0025312|T019|PT|414667000|SNOMEDCT_CORE|Meningomyelocele|Meningomyelocele
C0025312|T019|FN|414667000|SNOMEDCT_CORE|Meningomyelocele|Meningomyelocele
C0025312|T019|SY|414667000|SNOMEDCT_CORE|Myelomeningocele|Meningomyelocele
C0025319|T047|PT|123756000|SNOMEDCT_CORE|Menopausal syndrome|Menopausal syndrome
C0025319|T047|FN|123756000|SNOMEDCT_CORE|Menopausal syndrome|Menopausal syndrome
C0025322|T047|PT|373717006|SNOMEDCT_CORE|Premature menopause|Premature menopause
C0025322|T047|FN|373717006|SNOMEDCT_CORE|Premature menopause|Premature menopause
C0025323|T046|SY|386692008|SNOMEDCT_CORE|Flooding during periods|Menorrhagia
C0025323|T046|SY|386692008|SNOMEDCT_CORE|Heavy menstrual bleeding|Menorrhagia
C0025323|T046|SY|386692008|SNOMEDCT_CORE|Heavy period|Menorrhagia
C0025323|T046|SY|386692008|SNOMEDCT_CORE|Heavy periods|Menorrhagia
C0025323|T046|SY|386692008|SNOMEDCT_CORE|Hypermenorrhea|Menorrhagia
C0025323|T046|SYGB|386692008|SNOMEDCT_CORE|Hypermenorrhoea|Menorrhagia
C0025323|T046|PT|386692008|SNOMEDCT_CORE|Menorrhagia|Menorrhagia
C0025323|T046|FN|386692008|SNOMEDCT_CORE|Menorrhagia|Menorrhagia
C0025323|T046|SY|386692008|SNOMEDCT_CORE|Profuse menstrual flow|Menorrhagia
C0025345|T046|SY|386804004|SNOMEDCT_CORE|Abnormal menstruation|Disorder of menstruation
C0025345|T046|PT|386804004|SNOMEDCT_CORE|Disorder of menstruation|Disorder of menstruation
C0025345|T046|FN|386804004|SNOMEDCT_CORE|Disorder of menstruation|Disorder of menstruation
C0025345|T046|SY|386804004|SNOMEDCT_CORE|Menstrual disorder|Disorder of menstruation
C0025345|T046|SY|386804004|SNOMEDCT_CORE|Period disorder|Disorder of menstruation
C0025362|T048|OAP|91138005|SNOMEDCT_CORE|Mental retardation|MR - Mental retardation
C0025362|T048|IS|1855002|SNOMEDCT_CORE|Mental retardation|MR - Mental retardation
C0025362|T048|OAF|91138005|SNOMEDCT_CORE|Mental retardation|MR - Mental retardation
C0025362|T048|IS|91138005|SNOMEDCT_CORE|Mental retardation, NOS|MR - Mental retardation
C0025362|T048|OAS|91138005|SNOMEDCT_CORE|MR - Mental retardation|MR - Mental retardation
C0025362|T048|IS|1855002|SNOMEDCT_CORE|MR - Mental retardation|MR - Mental retardation
C0025469|T047|PT|44897000|SNOMEDCT_CORE|Mesenteric lymphadenitis|Mesenteric lymphadenitis
C0025469|T047|FN|44897000|SNOMEDCT_CORE|Mesenteric lymphadenitis|Mesenteric lymphadenitis
C0025469|T047|IS|44897000|SNOMEDCT_CORE|Mesenteric lymphadenitis, NOS|Mesenteric lymphadenitis
C0025517|T047|SY|75934005|SNOMEDCT_CORE|MD - Metabolic disorders|Metabolic disease
C0025517|T047|PT|75934005|SNOMEDCT_CORE|Metabolic disease|Metabolic disease
C0025517|T047|FN|75934005|SNOMEDCT_CORE|Metabolic disease|Metabolic disease
C0025517|T047|IS|75934005|SNOMEDCT_CORE|Metabolic disease, NOS|Metabolic disease
C0025517|T047|SY|75934005|SNOMEDCT_CORE|Metabolic disorder|Metabolic disease
C0025517|T047|IS|75934005|SNOMEDCT_CORE|Metabolic disorder, NOS|Metabolic disease
C0025587|T184|PT|10085004|SNOMEDCT_CORE|Metatarsalgia|Metatarsalgia
C0025587|T184|FN|10085004|SNOMEDCT_CORE|Metatarsalgia|Metatarsalgia
C0025587|T184|SY|10085004|SNOMEDCT_CORE|Pain in ball of foot|Metatarsalgia
C0025874|T046|OAS|19155002|SNOMEDCT_CORE|DUB - Dysfunctional uterine bleeding|DUH - Dysfunctional uterine haemorrhage
C0025874|T046|OAS|19155002|SNOMEDCT_CORE|DUH - Dysfunctional uterine haemorrhage|DUH - Dysfunctional uterine haemorrhage
C0025874|T046|OAS|19155002|SNOMEDCT_CORE|DUH - Dysfunctional uterine hemorrhage|DUH - Dysfunctional uterine haemorrhage
C0025874|T046|OAP|19155002|SNOMEDCT_CORE|Dysfunctional uterine bleeding|DUH - Dysfunctional uterine haemorrhage
C0025874|T046|OAF|19155002|SNOMEDCT_CORE|Dysfunctional uterine bleeding|DUH - Dysfunctional uterine haemorrhage
C0025874|T046|OAS|19155002|SNOMEDCT_CORE|Dysfunctional uterine haemorrhage|DUH - Dysfunctional uterine haemorrhage
C0025874|T046|OAS|19155002|SNOMEDCT_CORE|Dysfunctional uterine hemorrhage|DUH - Dysfunctional uterine haemorrhage
C0025958|T019|SY|1829003|SNOMEDCT_CORE|Micrencephaly|Microcephalus
C0025958|T019|PT|1829003|SNOMEDCT_CORE|Microcephalus|Microcephalus
C0025958|T019|FN|1829003|SNOMEDCT_CORE|Microcephalus|Microcephalus
C0025958|T019|SY|1829003|SNOMEDCT_CORE|Microcephaly|Microcephalus
C0025958|T019|SY|1829003|SNOMEDCT_CORE|Nanocephaly|Microcephalus
C0026106|T048|SY|86765009|SNOMEDCT_CORE|Mild intellectual development disorder|Mild intellectual disability
C0026106|T048|FN|86765009|SNOMEDCT_CORE|Mild intellectual disability|Mild intellectual disability
C0026106|T048|PT|86765009|SNOMEDCT_CORE|Mild intellectual disability|Mild intellectual disability
C0026106|T048|SY|86765009|SNOMEDCT_CORE|Mild mental handicap|Mild intellectual disability
C0026106|T048|SY|86765009|SNOMEDCT_CORE|Mild mental retardation, IQ in range 50-70|Mild intellectual disability
C0026265|T047|SY|11851006|SNOMEDCT_CORE|Mitral valve disease|Mitral valve disorder
C0026265|T047|PT|11851006|SNOMEDCT_CORE|Mitral valve disorder|Mitral valve disorder
C0026265|T047|FN|11851006|SNOMEDCT_CORE|Mitral valve disorder|Mitral valve disorder
C0026265|T047|IS|11851006|SNOMEDCT_CORE|Mitral valve disorder, NOS|Mitral valve disorder
C0026265|T047|SY|11851006|SNOMEDCT_CORE|MVD - Mitral valve disease|Mitral valve disorder
C0026266|T046|SY|48724000|SNOMEDCT_CORE|MI - Mitral incompetence|Mitral valve regurgitation
C0026266|T046|SY|48724000|SNOMEDCT_CORE|Mitral insufficiency|Mitral valve regurgitation
C0026266|T046|SY|48724000|SNOMEDCT_CORE|Mitral regurgitation|Mitral valve regurgitation
C0026266|T046|IS|48724000|SNOMEDCT_CORE|Mitral regurgitation, NOS|Mitral valve regurgitation
C0026266|T046|SY|48724000|SNOMEDCT_CORE|Mitral valve incompetence|Mitral valve regurgitation
C0026266|T046|IS|48724000|SNOMEDCT_CORE|Mitral valve incompetence, NOS|Mitral valve regurgitation
C0026266|T046|SY|48724000|SNOMEDCT_CORE|Mitral valve insufficiency|Mitral valve regurgitation
C0026266|T046|IS|48724000|SNOMEDCT_CORE|Mitral valve insufficiency, NOS|Mitral valve regurgitation
C0026266|T046|PT|48724000|SNOMEDCT_CORE|Mitral valve regurgitation|Mitral valve regurgitation
C0026266|T046|FN|48724000|SNOMEDCT_CORE|Mitral valve regurgitation|Mitral valve regurgitation
C0026266|T046|IS|48724000|SNOMEDCT_CORE|Mitral valve regurgitation, NOS|Mitral valve regurgitation
C0026266|T046|SY|48724000|SNOMEDCT_CORE|MR - Mitral regurgitation|Mitral valve regurgitation
C0026267|T047|PT|409712001|SNOMEDCT_CORE|Mitral valve prolapse|Mitral valve prolapse
C0026267|T047|FN|409712001|SNOMEDCT_CORE|Mitral valve prolapse|Mitral valve prolapse
C0026267|T047|SY|409712001|SNOMEDCT_CORE|MVP - Mitral valve prolapse|Mitral valve prolapse
C0026269|T047|SY|79619009|SNOMEDCT_CORE|Mitral stenosis|Mitral valve stenosis
C0026269|T047|PT|79619009|SNOMEDCT_CORE|Mitral valve stenosis|Mitral valve stenosis
C0026269|T047|FN|79619009|SNOMEDCT_CORE|Mitral valve stenosis|Mitral valve stenosis
C0026269|T047|IS|79619009|SNOMEDCT_CORE|Mitral valve stenosis, NOS|Mitral valve stenosis
C0026269|T047|SY|79619009|SNOMEDCT_CORE|MS - Mitral stenosis|Mitral valve stenosis
C0026272|T047|SY|398049005|SNOMEDCT_CORE|MCTD - Mixed connective tissue disease|Mixed collagen vascular disease
C0026272|T047|PT|398049005|SNOMEDCT_CORE|Mixed collagen vascular disease|Mixed collagen vascular disease
C0026272|T047|FN|398049005|SNOMEDCT_CORE|Mixed collagen vascular disease|Mixed collagen vascular disease
C0026272|T047|SY|398049005|SNOMEDCT_CORE|Mixed connective tissue disease|Mixed collagen vascular disease
C0026272|T047|SY|398049005|SNOMEDCT_CORE|Sharp's syndrome|Mixed collagen vascular disease
C0026351|T048|SY|61152003|SNOMEDCT_CORE|Moderate intellectual development disorder|Moderate intellectual disability
C0026351|T048|PT|61152003|SNOMEDCT_CORE|Moderate intellectual disability|Moderate intellectual disability
C0026351|T048|FN|61152003|SNOMEDCT_CORE|Moderate intellectual disability|Moderate intellectual disability
C0026351|T048|SY|61152003|SNOMEDCT_CORE|Moderate mental handicap|Moderate intellectual disability
C0026393|T047|FN|40070004|SNOMEDCT_CORE|Infection caused by Molluscum contagiosum|Molluscum contagiosum infection
C0026393|T047|SY|40070004|SNOMEDCT_CORE|Infection caused by Molluscum contagiosum|Molluscum contagiosum infection
C0026393|T047|IS|40070004|SNOMEDCT_CORE|MC - Molluscum contagiosum|Molluscum contagiosum infection
C0026393|T047|IS|40070004|SNOMEDCT_CORE|Molluscum contagiosum|Molluscum contagiosum infection
C0026393|T047|PT|40070004|SNOMEDCT_CORE|Molluscum contagiosum infection|Molluscum contagiosum infection
C0026393|T047|OF|40070004|SNOMEDCT_CORE|Molluscum contagiosum infection|Molluscum contagiosum infection
C0026393|T047|IS|40070004|SNOMEDCT_CORE|Molluscum verrucosum|Molluscum contagiosum infection
C0026470|T191|SY|58648008|SNOMEDCT_CORE|Asymptomatic monoclonal gammopathy|Benign monoclonal gammopathy
C0026470|T191|PT|58648008|SNOMEDCT_CORE|Benign monoclonal gammopathy|Benign monoclonal gammopathy
C0026470|T191|FN|58648008|SNOMEDCT_CORE|Benign monoclonal gammopathy|Benign monoclonal gammopathy
C0026470|T191|SY|277577000|SNOMEDCT_CORE|MGUS - Monoclonal gammopathy of uncertain significance|Benign monoclonal gammopathy
C0026470|T191|PT|277577000|SNOMEDCT_CORE|Monoclonal gammopathy of uncertain significance|Benign monoclonal gammopathy
C0026470|T191|FN|277577000|SNOMEDCT_CORE|Monoclonal gammopathy of uncertain significance|Benign monoclonal gammopathy
C0026470|T191|SY|277577000|SNOMEDCT_CORE|Monoclonal gammopathy of undetermined significance|Benign monoclonal gammopathy
C0026471|T191|OAP|267440005|SNOMEDCT_CORE|Monoclonal paraproteinaemia|Monoclonal paraproteinaemia
C0026471|T191|OAP|267440005|SNOMEDCT_CORE|Monoclonal paraproteinemia|Monoclonal paraproteinemia
C0026471|T191|OAF|267440005|SNOMEDCT_CORE|Monoclonal paraproteinemia|Monoclonal paraproteinemia
C0026603|T047|PT|37031009|SNOMEDCT_CORE|Motion sickness|Motion sickness
C0026603|T047|OF|37031009|SNOMEDCT_CORE|Motion sickness|Motion sickness
C0026603|T047|FN|37031009|SNOMEDCT_CORE|Motion sickness|Motion sickness
C0026603|T047|IS|37031009|SNOMEDCT_CORE|Motion sickness, NOS|Motion sickness
C0026603|T047|SY|37031009|SNOMEDCT_CORE|Riders' vertigo|Motion sickness
C0026603|T047|SY|37031009|SNOMEDCT_CORE|Travel sickness|Motion sickness
C0026636|T047|PT|118938008|SNOMEDCT_CORE|Disease of mouth|Disease of mouth
C0026636|T047|OF|118938008|SNOMEDCT_CORE|Disease of mouth|Disease of mouth
C0026636|T047|SY|118938008|SNOMEDCT_CORE|Disorder of mouth|Disease of mouth
C0026636|T047|FN|118938008|SNOMEDCT_CORE|Disorder of mouth|Disease of mouth
C0026636|T047|SY|118938008|SNOMEDCT_CORE|Disorder of oral cavity|Disease of mouth
C0026636|T047|SY|118938008|SNOMEDCT_CORE|Mouth disorder|Disease of mouth
C0026644|T033|PT|278650002|SNOMEDCT_CORE|Edentulous|Edentulous
C0026644|T033|FN|278650002|SNOMEDCT_CORE|Edentulous|Edentulous
C0026644|T033|SY|278650002|SNOMEDCT_CORE|No natural teeth|Edentulous
C0026650|T047|PT|60342002|SNOMEDCT_CORE|Movement disorder|Movement disorder
C0026650|T047|FN|60342002|SNOMEDCT_CORE|Movement disorder|Movement disorder
C0026650|T047|IS|60342002|SNOMEDCT_CORE|Movement disorder, NOS|Movement disorder
C0026686|T047|PT|69825009|SNOMEDCT_CORE|Mucocele of salivary gland|Mucocele of salivary gland
C0026686|T047|FN|69825009|SNOMEDCT_CORE|Mucocele of salivary gland|Mucocele of salivary gland
C0026686|T047|SY|69825009|SNOMEDCT_CORE|Mucous retention cyst of salivary gland|Mucocele of salivary gland
C0026686|T047|SY|69825009|SNOMEDCT_CORE|Ptyalocele|Mucocele of salivary gland
C0026686|T047|SY|69825009|SNOMEDCT_CORE|Retention cyst of salivary gland|Mucocele of salivary gland
C0026686|T047|SY|69825009|SNOMEDCT_CORE|Salivary cyst|Mucocele of salivary gland
C0026686|T047|SY|69825009|SNOMEDCT_CORE|Sialocele|Mucocele of salivary gland
C0026691|T047|PT|75053002|SNOMEDCT_CORE|Acute febrile mucocutaneous lymph node syndrome|Acute febrile mucocutaneous lymph node syndrome
C0026691|T047|FN|75053002|SNOMEDCT_CORE|Acute febrile mucocutaneous lymph node syndrome|Acute febrile mucocutaneous lymph node syndrome
C0026691|T047|SY|75053002|SNOMEDCT_CORE|Kawasaki disease|Acute febrile mucocutaneous lymph node syndrome
C0026691|T047|SY|75053002|SNOMEDCT_CORE|Kawasaki syndrome|Acute febrile mucocutaneous lymph node syndrome
C0026691|T047|SY|75053002|SNOMEDCT_CORE|Kawasaki's disease|Acute febrile mucocutaneous lymph node syndrome
C0026691|T047|SY|75053002|SNOMEDCT_CORE|Kawasaki's syndrome|Acute febrile mucocutaneous lymph node syndrome
C0026691|T047|SY|75053002|SNOMEDCT_CORE|Kawasakis mucocutaneous lymph node syndrome|Acute febrile mucocutaneous lymph node syndrome
C0026691|T047|SY|75053002|SNOMEDCT_CORE|MCLS|Acute febrile mucocutaneous lymph node syndrome
C0026691|T047|SY|75053002|SNOMEDCT_CORE|MLNS|Acute febrile mucocutaneous lymph node syndrome
C0026691|T047|SY|75053002|SNOMEDCT_CORE|Mucocutaneous lymph node syndrome|Acute febrile mucocutaneous lymph node syndrome
C0026751|T033|IS|28079008|SNOMEDCT_CORE|Multiparity|Multiparous
C0026751|T033|PT|28079008|SNOMEDCT_CORE|Multiparous|Multiparous
C0026751|T033|FN|28079008|SNOMEDCT_CORE|Multiparous|Multiparous
C0026764|T191|SY|109989006|SNOMEDCT_CORE|Kahler's disease|Multiple myeloma
C0026764|T191|PT|109989006|SNOMEDCT_CORE|Multiple myeloma|Multiple myeloma
C0026764|T191|SY|109989006|SNOMEDCT_CORE|Multiple myeloma|Multiple myeloma
C0026764|T191|FN|109989006|SNOMEDCT_CORE|Multiple myeloma|Multiple myeloma
C0026764|T191|SY|109989006|SNOMEDCT_CORE|Myeloma|Multiple myeloma
C0026764|T191|SY|109989006|SNOMEDCT_CORE|Myelomatosis|Multiple myeloma
C0026764|T191|SY|109989006|SNOMEDCT_CORE|Plasmacytic myeloma|Multiple myeloma
C0026769|T047|SY|24700007|SNOMEDCT_CORE|Disseminated sclerosis|Multiple sclerosis
C0026769|T047|SY|24700007|SNOMEDCT_CORE|DS - Disseminated sclerosis|Multiple sclerosis
C0026769|T047|IS|24700007|SNOMEDCT_CORE|Generalised multiple sclerosis|Multiple sclerosis
C0026769|T047|IS|24700007|SNOMEDCT_CORE|Generalized multiple sclerosis|Multiple sclerosis
C0026769|T047|SY|24700007|SNOMEDCT_CORE|MS - Multiple sclerosis|Multiple sclerosis
C0026769|T047|PT|24700007|SNOMEDCT_CORE|Multiple sclerosis|Multiple sclerosis
C0026769|T047|FN|24700007|SNOMEDCT_CORE|Multiple sclerosis|Multiple sclerosis
C0026769|T047|IS|24700007|SNOMEDCT_CORE|Multiple sclerosis, NOS|Multiple sclerosis
C0026773|T048|SY|31611000|SNOMEDCT_CORE|Dissociative identity disorder|Multiple personality disorder
C0026773|T048|PT|31611000|SNOMEDCT_CORE|Multiple personality disorder|Multiple personality disorder
C0026773|T048|FN|31611000|SNOMEDCT_CORE|Multiple personality disorder|Multiple personality disorder
C0026780|T047|IS|36989005|SNOMEDCT_CORE|Epidemic parotitis|Mumps
C0026780|T047|IS|36989005|SNOMEDCT_CORE|Infectious parotitis|Mumps
C0026780|T047|PT|36989005|SNOMEDCT_CORE|Mumps|Mumps
C0026780|T047|FN|36989005|SNOMEDCT_CORE|Mumps|Mumps
C0026780|T047|IS|36989005|SNOMEDCT_CORE|Mumps, NOS|Mumps
C0026821|T184|PT|55300003|SNOMEDCT_CORE|Cramp|Cramp
C0026821|T184|FN|55300003|SNOMEDCT_CORE|Cramp|Cramp
C0026821|T184|SY|55300003|SNOMEDCT_CORE|Cramp in muscle|Cramp
C0026821|T184|IS|55300003|SNOMEDCT_CORE|Cramp in muscle, NOS|Cramp
C0026821|T184|IS|55300003|SNOMEDCT_CORE|Cramp, NOS|Cramp
C0026821|T184|SY|55300003|SNOMEDCT_CORE|Muscle cramp|Cramp
C0026821|T184|IS|55300003|SNOMEDCT_CORE|Muscle cramp, NOS|Cramp
C0026821|T184|SY|55300003|SNOMEDCT_CORE|Muscle cramps|Cramp
C0026827|T033|PT|398151007|SNOMEDCT_CORE|Decreased muscle tone|Decreased muscle tone
C0026827|T033|FN|398151007|SNOMEDCT_CORE|Decreased muscle tone|Decreased muscle tone
C0026838|T184|SY|221360009|SNOMEDCT_CORE|Muscle spasm - tone|Spasticity
C0026838|T184|SY|221360009|SNOMEDCT_CORE|Muscle spasticity|Spasticity
C0026838|T184|SY|221360009|SNOMEDCT_CORE|Muscular spasticity|Spasticity
C0026838|T184|PT|221360009|SNOMEDCT_CORE|Spasticity|Spasticity
C0026838|T184|FN|221360009|SNOMEDCT_CORE|Spasticity|Spasticity
C0026846|T046|SY|88092000|SNOMEDCT_CORE|Amyotrophia|Muscle atrophy
C0026846|T046|IS|88092000|SNOMEDCT_CORE|Amyotrophia, NOS|Muscle atrophy
C0026846|T046|SY|88092000|SNOMEDCT_CORE|Amyotrophy|Muscle atrophy
C0026846|T046|IS|88092000|SNOMEDCT_CORE|Amyotrophy, NOS|Muscle atrophy
C0026846|T046|PT|88092000|SNOMEDCT_CORE|Muscle atrophy|Muscle atrophy
C0026846|T046|FN|88092000|SNOMEDCT_CORE|Muscle atrophy|Muscle atrophy
C0026846|T046|IS|88092000|SNOMEDCT_CORE|Muscle atrophy, NOS|Muscle atrophy
C0026846|T046|SY|88092000|SNOMEDCT_CORE|Muscle thinning|Muscle atrophy
C0026846|T046|SY|88092000|SNOMEDCT_CORE|Muscle wasting|Muscle atrophy
C0026846|T046|SY|88092000|SNOMEDCT_CORE|Muscle wasting disorder|Muscle atrophy
C0026846|T046|IS|88092000|SNOMEDCT_CORE|Muscle wasting, NOS|Muscle atrophy
C0026846|T046|SY|88092000|SNOMEDCT_CORE|Muscular atrophy|Muscle atrophy
C0026846|T046|IS|88092000|SNOMEDCT_CORE|Muscular atrophy, NOS|Muscle atrophy
C0026848|T047|PT|129565002|SNOMEDCT_CORE|Disorder of muscle|Disorder of muscle
C0026848|T047|SY|129565002|SNOMEDCT_CORE|Disorder of skeletal AND/OR smooth muscle|Disorder of muscle
C0026848|T047|FN|129565002|SNOMEDCT_CORE|Disorder of skeletal AND/OR smooth muscle|Disorder of muscle
C0026848|T047|SY|129565002|SNOMEDCT_CORE|Myopathic disease|Disorder of muscle
C0026848|T047|SY|129565002|SNOMEDCT_CORE|Myopathy|Disorder of muscle
C0026850|T047|SY|73297009|SNOMEDCT_CORE|MD - Muscular dystrophy|Muscular dystrophy
C0026850|T047|PT|73297009|SNOMEDCT_CORE|Muscular dystrophy|Muscular dystrophy
C0026850|T047|FN|73297009|SNOMEDCT_CORE|Muscular dystrophy|Muscular dystrophy
C0026850|T047|IS|73297009|SNOMEDCT_CORE|Muscular dystrophy, NOS|Muscular dystrophy
C0026850|T047|SY|73297009|SNOMEDCT_CORE|PMD - Progressive muscular dystrophy|Muscular dystrophy
C0026850|T047|SY|73297009|SNOMEDCT_CORE|Progressive muscular dystrophy|Muscular dystrophy
C0026858|T033|PT|279069000|SNOMEDCT_CORE|Musculoskeletal pain|Musculoskeletal pain
C0026858|T033|FN|279069000|SNOMEDCT_CORE|Musculoskeletal pain|Musculoskeletal pain
C0026858|T033|SY|279069000|SNOMEDCT_CORE|Rheumatic pain|Musculoskeletal pain
C0026896|T047|SY|91637004|SNOMEDCT_CORE|Erb-Goldflam disease|Myasthenia gravis
C0026896|T047|SY|91637004|SNOMEDCT_CORE|MG - Myasthenia gravis|Myasthenia gravis
C0026896|T047|PT|91637004|SNOMEDCT_CORE|Myasthenia gravis|Myasthenia gravis
C0026896|T047|FN|91637004|SNOMEDCT_CORE|Myasthenia gravis|Myasthenia gravis
C0026896|T047|IS|91637004|SNOMEDCT_CORE|Myasthenia gravis, NOS|Myasthenia gravis
C0026916|T047|SY|373436002|SNOMEDCT_CORE|Infection caused by Mycobacterium intracellulare|Infection due to Mycobacterium intracellulare
C0026916|T047|FN|373436002|SNOMEDCT_CORE|Infection caused by Mycobacterium intracellulare|Infection due to Mycobacterium intracellulare
C0026916|T047|PT|373436002|SNOMEDCT_CORE|Infection due to Mycobacterium intracellulare|Infection due to Mycobacterium intracellulare
C0026916|T047|OF|373436002|SNOMEDCT_CORE|Infection due to Mycobacterium intracellulare|Infection due to Mycobacterium intracellulare
C0026918|T047|SY|88415009|SNOMEDCT_CORE|Infection due to mycobacteria|Mycobacteriosis
C0026918|T047|SY|88415009|SNOMEDCT_CORE|Mycobacterial disease|Mycobacteriosis
C0026918|T047|PT|88415009|SNOMEDCT_CORE|Mycobacteriosis|Mycobacteriosis
C0026918|T047|FN|88415009|SNOMEDCT_CORE|Mycobacteriosis|Mycobacteriosis
C0026918|T047|IS|88415009|SNOMEDCT_CORE|Mycobacteriosis, NOS|Mycobacteriosis
C0026919|T047|IS|88415009|SNOMEDCT_CORE|Atypical mycobacterial infection, NOS|Atypical mycobacterial infection, NOS
C0026946|T047|SY|3218000|SNOMEDCT_CORE|Disease caused by fungus|Mycosis
C0026946|T047|IS|3218000|SNOMEDCT_CORE|Disease caused by fungus, NOS|Mycosis
C0026946|T047|SY|3218000|SNOMEDCT_CORE|Fungal infection|Mycosis
C0026946|T047|IS|3218000|SNOMEDCT_CORE|Fungal infection, NOS|Mycosis
C0026946|T047|SY|3218000|SNOMEDCT_CORE|Fungal infectious disease|Mycosis
C0026946|T047|IS|3218000|SNOMEDCT_CORE|Fungal infectious disease, NOS|Mycosis
C0026946|T047|SY|3218000|SNOMEDCT_CORE|Fungus infection|Mycosis
C0026946|T047|IS|3218000|SNOMEDCT_CORE|Fungus infection, NOS|Mycosis
C0026946|T047|SY|3218000|SNOMEDCT_CORE|Mycoses|Mycosis
C0026946|T047|PT|3218000|SNOMEDCT_CORE|Mycosis|Mycosis
C0026946|T047|FN|3218000|SNOMEDCT_CORE|Mycosis|Mycosis
C0026946|T047|IS|3218000|SNOMEDCT_CORE|Mycosis, NOS|Mycosis
C0026946|T047|SY|3218000|SNOMEDCT_CORE|Mycotic disease|Mycosis
C0026948|T191|SY|118618005|SNOMEDCT_CORE|MF - Mycosis fungoides|Mycosis fungoides
C0026948|T191|SY|118618005|SNOMEDCT_CORE|Mycosis fungoides|Mycosis fungoides
C0026948|T191|PT|118618005|SNOMEDCT_CORE|Mycosis fungoides|Mycosis fungoides
C0026948|T191|FN|118618005|SNOMEDCT_CORE|Mycosis fungoides|Mycosis fungoides
C0026976|T047|SY|16631009|SNOMEDCT_CORE|Transverse myelitis|Transverse myelopathy syndrome
C0026976|T047|PT|16631009|SNOMEDCT_CORE|Transverse myelopathy syndrome|Transverse myelopathy syndrome
C0026976|T047|FN|16631009|SNOMEDCT_CORE|Transverse myelopathy syndrome|Transverse myelopathy syndrome
C0026987|T191|SY|52967002|SNOMEDCT_CORE|MF - Myelofibrosis|Myelofibrosis
C0026987|T191|PT|52967002|SNOMEDCT_CORE|Myelofibrosis|Myelofibrosis
C0026987|T191|FN|52967002|SNOMEDCT_CORE|Myelofibrosis|Myelofibrosis
C0026987|T191|IS|52967002|SNOMEDCT_CORE|Myelofibrosis, NOS|Myelofibrosis
C0026987|T191|SY|52967002|SNOMEDCT_CORE|Myelosclerosis|Myelofibrosis
C0027013|T047|PT|443230004|SNOMEDCT_CORE|Myeloid metaplasia|Myeloid metaplasia
C0027013|T047|PT|82513007|SNOMEDCT_CORE|Myeloid metaplasia|Myeloid metaplasia
C0027013|T047|FN|82513007|SNOMEDCT_CORE|Myeloid metaplasia|Myeloid metaplasia
C0027013|T047|FN|443230004|SNOMEDCT_CORE|Myeloid metaplasia|Myeloid metaplasia
C0027022|T191|PT|425333006|SNOMEDCT_CORE|Myeloproliferative disorder|Myeloproliferative disorder
C0027022|T191|FN|425333006|SNOMEDCT_CORE|Myeloproliferative disorder|Myeloproliferative disorder
C0027051|T047|SY|22298006|SNOMEDCT_CORE|Cardiac infarction|Myocardial infarction
C0027051|T047|IS|22298006|SNOMEDCT_CORE|Cardiac infarction, NOS|Myocardial infarction
C0027051|T047|SY|22298006|SNOMEDCT_CORE|Heart attack|Myocardial infarction
C0027051|T047|IS|22298006|SNOMEDCT_CORE|Heart attack, NOS|Myocardial infarction
C0027051|T047|SY|22298006|SNOMEDCT_CORE|Infarction of heart|Myocardial infarction
C0027051|T047|IS|22298006|SNOMEDCT_CORE|Infarction of heart, NOS|Myocardial infarction
C0027051|T047|SY|22298006|SNOMEDCT_CORE|MI - myocardial infarction|Myocardial infarction
C0027051|T047|IS|22298006|SNOMEDCT_CORE|MI - Myocardial infarction|Myocardial infarction
C0027051|T047|SY|22298006|SNOMEDCT_CORE|Myocardial infarct|Myocardial infarction
C0027051|T047|PT|22298006|SNOMEDCT_CORE|Myocardial infarction|Myocardial infarction
C0027051|T047|FN|22298006|SNOMEDCT_CORE|Myocardial infarction|Myocardial infarction
C0027051|T047|IS|22298006|SNOMEDCT_CORE|Myocardial infarction, NOS|Myocardial infarction
C0027059|T047|SY|50920009|SNOMEDCT_CORE|Myocardial inflammation|Myocarditis
C0027059|T047|PT|50920009|SNOMEDCT_CORE|Myocarditis|Myocarditis
C0027059|T047|FN|50920009|SNOMEDCT_CORE|Myocarditis|Myocarditis
C0027059|T047|IS|50920009|SNOMEDCT_CORE|Myocarditis, NOS|Myocarditis
C0027066|T184|SY|17450006|SNOMEDCT_CORE|Myoclonia|Myoclonus
C0027066|T184|PT|17450006|SNOMEDCT_CORE|Myoclonus|Myoclonus
C0027066|T184|FN|17450006|SNOMEDCT_CORE|Myoclonus|Myoclonus
C0027092|T047|PT|57190000|SNOMEDCT_CORE|Myopia|Myopia
C0027092|T047|FN|57190000|SNOMEDCT_CORE|Myopia|Myopia
C0027092|T047|SY|57190000|SNOMEDCT_CORE|Near sighted|Myopia
C0027092|T047|SY|57190000|SNOMEDCT_CORE|Nearsightedness|Myopia
C0027121|T047|SY|26889001|SNOMEDCT_CORE|Inflammatory disorder of muscle|Myositis
C0027121|T047|SY|26889001|SNOMEDCT_CORE|Inflammatory myopathy|Myositis
C0027121|T047|SY|26889001|SNOMEDCT_CORE|Muscle inflammation|Myositis
C0027121|T047|PT|26889001|SNOMEDCT_CORE|Myositis|Myositis
C0027121|T047|FN|26889001|SNOMEDCT_CORE|Myositis|Myositis
C0027121|T047|IS|26889001|SNOMEDCT_CORE|Myositis, NOS|Myositis
C0027126|T047|SY|77956009|SNOMEDCT_CORE|DM - Dystrophia myotonica|Steinert myotonic dystrophy syndrome
C0027126|T047|SY|77956009|SNOMEDCT_CORE|Dystrophia myotonica|Steinert myotonic dystrophy syndrome
C0027126|T047|SY|77956009|SNOMEDCT_CORE|Myotonia dystrophica|Steinert myotonic dystrophy syndrome
C0027126|T047|SY|77956009|SNOMEDCT_CORE|Myotonic dystrophy|Steinert myotonic dystrophy syndrome
C0027126|T047|PT|77956009|SNOMEDCT_CORE|Steinert myotonic dystrophy syndrome|Steinert myotonic dystrophy syndrome
C0027126|T047|FN|77956009|SNOMEDCT_CORE|Steinert myotonic dystrophy syndrome|Steinert myotonic dystrophy syndrome
C0027126|T047|SY|77956009|SNOMEDCT_CORE|Steinert syndrome|Steinert myotonic dystrophy syndrome
C0027343|T033|SY|400200009|SNOMEDCT_CORE|Embedded toenail|Ingrowing nail
C0027343|T033|SY|400200009|SNOMEDCT_CORE|IGTN - Ingrowing toenail|Ingrowing nail
C0027343|T033|PT|400097005|SNOMEDCT_CORE|Ingrowing nail|Ingrowing nail
C0027343|T033|FN|400097005|SNOMEDCT_CORE|Ingrowing nail|Ingrowing nail
C0027343|T033|PT|400200009|SNOMEDCT_CORE|Ingrowing toenail|Ingrowing nail
C0027343|T033|FN|400200009|SNOMEDCT_CORE|Ingrowing toenail|Ingrowing nail
C0027343|T033|SY|400097005|SNOMEDCT_CORE|Ingrown nail|Ingrowing nail
C0027343|T033|SY|400200009|SNOMEDCT_CORE|Ingrown toenail|Ingrowing nail
C0027343|T033|SY|400097005|SNOMEDCT_CORE|OC - Onychocryptosis|Ingrowing nail
C0027343|T033|SY|400097005|SNOMEDCT_CORE|Onychocryptosis|Ingrowing nail
C0027343|T033|SY|400097005|SNOMEDCT_CORE|Onyxis|Ingrowing nail
C0027343|T033|SY|400097005|SNOMEDCT_CORE|Unguis aduncus|Ingrowing nail
C0027343|T033|SY|400097005|SNOMEDCT_CORE|Unguis incarnatus|Ingrowing nail
C0027402|T048|PT|80711002|SNOMEDCT_CORE|Narcissistic personality disorder|Narcissistic personality disorder
C0027402|T048|FN|80711002|SNOMEDCT_CORE|Narcissistic personality disorder|Narcissistic personality disorder
C0027404|T047|SY|60380001|SNOMEDCT_CORE|Gelineau's syndrome|Narcolepsy
C0027404|T047|PT|60380001|SNOMEDCT_CORE|Narcolepsy|Narcolepsy
C0027404|T047|FN|60380001|SNOMEDCT_CORE|Narcolepsy|Narcolepsy
C0027404|T047|SY|60380001|SNOMEDCT_CORE|Narcoleptic syndrome|Narcolepsy
C0027404|T047|SY|60380001|SNOMEDCT_CORE|Paroxysmal sleep|Narcolepsy
C0027424|T184|SY|68235000|SNOMEDCT_CORE|Congested nose|Nasal congestion
C0027424|T184|FN|68235000|SNOMEDCT_CORE|Nasal congestion|Nasal congestion
C0027424|T184|PT|68235000|SNOMEDCT_CORE|Nasal congestion|Nasal congestion
C0027424|T184|SY|68235000|SNOMEDCT_CORE|Stuffed-up nose|Nasal congestion
C0027429|T033|SY|232209000|SNOMEDCT_CORE|Nasal airway obstruction|Nasal obstruction
C0027429|T033|PT|232209000|SNOMEDCT_CORE|Nasal obstruction|Nasal obstruction
C0027429|T033|FN|232209000|SNOMEDCT_CORE|Nasal obstruction|Nasal obstruction
C0027429|T033|SY|232209000|SNOMEDCT_CORE|Nasal obstruction present|Nasal obstruction
C0027429|T033|SY|232209000|SNOMEDCT_CORE|NO - Nasal obstruction|Nasal obstruction
C0027430|T047|OAP|52756005|SNOMEDCT_CORE|Nasal polyp|Polyp of nasal cavity
C0027430|T047|OAF|52756005|SNOMEDCT_CORE|Nasal polyp|Polyp of nasal cavity
C0027430|T047|OAS|52756005|SNOMEDCT_CORE|Nasal polyp - anterior|Polyp of nasal cavity
C0027430|T047|IS|52756005|SNOMEDCT_CORE|Nasal polyp, NOS|Polyp of nasal cavity
C0027430|T047|OAS|52756005|SNOMEDCT_CORE|Nasal polyposis|Polyp of nasal cavity
C0027430|T047|OAS|52756005|SNOMEDCT_CORE|Polyp in anterior nares|Polyp of nasal cavity
C0027430|T047|OAS|52756005|SNOMEDCT_CORE|Polyp of nasal cavity|Polyp of nasal cavity
C0027430|T047|PT|736500007|SNOMEDCT_CORE|Polyp of nasal cavity|Polyp of nasal cavity
C0027430|T047|FN|736500007|SNOMEDCT_CORE|Polyp of nasal cavity|Polyp of nasal cavity
C0027430|T047|IS|52756005|SNOMEDCT_CORE|Polyp of nasal cavity, NOS|Polyp of nasal cavity
C0027441|T047|PT|51476001|SNOMEDCT_CORE|Nasopharyngitis|Nasopharyngitis
C0027441|T047|FN|51476001|SNOMEDCT_CORE|Nasopharyngitis|Nasopharyngitis
C0027441|T047|IS|51476001|SNOMEDCT_CORE|Nasopharyngitis, NOS|Nasopharyngitis
C0027441|T047|SY|51476001|SNOMEDCT_CORE|Rhinopharyngitis|Nasopharyngitis
C0027441|T047|IS|51476001|SNOMEDCT_CORE|Rhinopharyngitis, NOS|Nasopharyngitis
C0027497|T184|PT|422587007|SNOMEDCT_CORE|Nausea|Nausea
C0027497|T184|FN|422587007|SNOMEDCT_CORE|Nausea|Nausea
C0027497|T184|SY|422587007|SNOMEDCT_CORE|Nauseated|Nausea
C0027497|T184|SY|422587007|SNOMEDCT_CORE|Nauseous|Nausea
C0027497|T184|SY|422587007|SNOMEDCT_CORE|Observation of nausea|Nausea
C0027498|T184|SY|16932000|SNOMEDCT_CORE|N&V - Nausea and vomiting|Nausea and vomiting
C0027498|T184|SY|16932000|SNOMEDCT_CORE|N+V - Nausea and vomiting|Nausea and vomiting
C0027498|T184|PT|16932000|SNOMEDCT_CORE|Nausea and vomiting|Nausea and vomiting
C0027498|T184|FN|16932000|SNOMEDCT_CORE|Nausea and vomiting|Nausea and vomiting
C0027531|T037|PT|90460009|SNOMEDCT_CORE|Injury of neck|Injury of neck
C0027531|T037|FN|90460009|SNOMEDCT_CORE|Injury of neck|Injury of neck
C0027531|T037|SY|90460009|SNOMEDCT_CORE|Neck injury|Injury of neck
C0027535|T037|IS|39848009|SNOMEDCT_CORE|Acute cervical sprain|Neck sprain
C0027535|T037|IS|39848009|SNOMEDCT_CORE|Cervical sprain|Neck sprain
C0027535|T037|SY|209557005|SNOMEDCT_CORE|Cervical sprain|Neck sprain
C0027535|T037|PT|209557005|SNOMEDCT_CORE|Neck sprain|Neck sprain
C0027535|T037|FN|209557005|SNOMEDCT_CORE|Neck sprain|Neck sprain
C0027543|T047|PT|397758007|SNOMEDCT_CORE|Avascular necrosis of bone|Avascular necrosis of bone
C0027543|T047|FN|397758007|SNOMEDCT_CORE|Avascular necrosis of bone|Avascular necrosis of bone
C0027543|T047|SY|397758007|SNOMEDCT_CORE|AVN - Avascular necrosis of bone|Avascular necrosis of bone
C0027609|T047|OAP|61628006|SNOMEDCT_CORE|Drug withdrawal syndrome in newborn|Drug withdrawal syndrome in newborn
C0027609|T047|OAF|61628006|SNOMEDCT_CORE|Drug withdrawal syndrome in newborn|Drug withdrawal syndrome in newborn
C0027609|T047|IS|61628006|SNOMEDCT_CORE|Neonatal drug withdrawal syndrome|Drug withdrawal syndrome in newborn
C0027609|T047|IS|61628006|SNOMEDCT_CORE|Newborn drug withdrawal syndrome|Drug withdrawal syndrome in newborn
C0027611|T047|FN|206345004|SNOMEDCT_CORE|Neonatal dacryocystitis and conjunctivitis|Neonatal dacryocystitis and conjunctivitis
C0027611|T047|PT|206345004|SNOMEDCT_CORE|Neonatal dacryocystitis and conjunctivitis|Neonatal dacryocystitis and conjunctivitis
C0027667|T191|SY|255052006|SNOMEDCT_CORE|CA - Cancer of unknown origin|Malignant tumor of unknown origin
C0027667|T191|SY|255052006|SNOMEDCT_CORE|Cancer - unknown origin|Malignant tumor of unknown origin
C0027667|T191|SY|255052006|SNOMEDCT_CORE|Malignant neoplasm of unknown origin|Malignant tumor of unknown origin
C0027667|T191|FN|255052006|SNOMEDCT_CORE|Malignant neoplasm of unknown origin|Malignant tumor of unknown origin
C0027667|T191|SY|255052006|SNOMEDCT_CORE|Malignant tumor - unknown primary|Malignant tumor of unknown origin
C0027667|T191|PT|255052006|SNOMEDCT_CORE|Malignant tumor of unknown origin|Malignant tumor of unknown origin
C0027667|T191|OF|255052006|SNOMEDCT_CORE|Malignant tumor of unknown origin|Malignant tumor of unknown origin
C0027667|T191|SYGB|255052006|SNOMEDCT_CORE|Malignant tumour - unknown primary|Malignant tumor of unknown origin
C0027667|T191|PTGB|255052006|SNOMEDCT_CORE|Malignant tumour of unknown origin|Malignant tumor of unknown origin
C0027667|T191|SY|255052006|SNOMEDCT_CORE|Metastasis - unknown primary|Malignant tumor of unknown origin
C0027667|T191|SY|255052006|SNOMEDCT_CORE|UKP - Malignant tumor - unknown primary|Malignant tumor of unknown origin
C0027667|T191|SYGB|255052006|SNOMEDCT_CORE|UKP - Malignant tumour - unknown primary|Malignant tumor of unknown origin
C0027697|T047|PT|52845002|SNOMEDCT_CORE|Nephritis|Nephritis
C0027697|T047|FN|52845002|SNOMEDCT_CORE|Nephritis|Nephritis
C0027697|T047|IS|52845002|SNOMEDCT_CORE|Nephritis, NOS|Nephritis
C0027707|T047|OAP|28689008|SNOMEDCT_CORE|Interstitial nephritis|Interstitial nephritis
C0027707|T047|OAF|28689008|SNOMEDCT_CORE|Interstitial nephritis|Interstitial nephritis
C0027707|T047|IS|28689008|SNOMEDCT_CORE|Interstitial nephritis, NOS|Interstitial nephritis, NOS
C0027708|T191|PT|302849000|SNOMEDCT_CORE|Nephroblastoma|Nephroblastoma
C0027708|T191|FN|302849000|SNOMEDCT_CORE|Nephroblastoma|Nephroblastoma
C0027708|T191|SY|302849000|SNOMEDCT_CORE|Nephroma|Nephroblastoma
C0027708|T191|IS|302849000|SNOMEDCT_CORE|Perlman syndrome|Nephroblastoma
C0027708|T191|SY|302849000|SNOMEDCT_CORE|Wilm's tumor|Nephroblastoma
C0027708|T191|SY|302849000|SNOMEDCT_CORE|Wilms tumor|Nephroblastoma
C0027708|T191|SYGB|302849000|SNOMEDCT_CORE|Wilms tumour|Nephroblastoma
C0027708|T191|IS|302849000|SNOMEDCT_CORE|Wilms' tumor|Nephroblastoma
C0027708|T191|IS|302849000|SNOMEDCT_CORE|Wilms' tumour|Nephroblastoma
C0027719|T047|SY|32916005|SNOMEDCT_CORE|Arteriosclerosis of kidney|Nephrosclerosis
C0027719|T047|SY|32916005|SNOMEDCT_CORE|Chronic arteriosclerotic nephritis|Nephrosclerosis
C0027719|T047|SY|32916005|SNOMEDCT_CORE|Interstitial arteriosclerotic nephritis|Nephrosclerosis
C0027719|T047|PT|32916005|SNOMEDCT_CORE|Nephrosclerosis|Nephrosclerosis
C0027719|T047|FN|32916005|SNOMEDCT_CORE|Nephrosclerosis|Nephrosclerosis
C0027719|T047|SY|32916005|SNOMEDCT_CORE|Renal arteriosclerosis|Nephrosclerosis
C0027719|T047|SY|32916005|SNOMEDCT_CORE|Renal sclerosis|Nephrosclerosis
C0027720|T047|SY|90708001|SNOMEDCT_CORE|Nephrosis|Nephrosis
C0027720|T047|IS|90708001|SNOMEDCT_CORE|Nephrosis, NOS|Nephrosis
C0027726|T047|PT|52254009|SNOMEDCT_CORE|Nephrotic syndrome|Nephrotic syndrome
C0027726|T047|FN|52254009|SNOMEDCT_CORE|Nephrotic syndrome|Nephrotic syndrome
C0027726|T047|IS|52254009|SNOMEDCT_CORE|Nephrotic syndrome, NOS|Nephrotic syndrome
C0027726|T047|SY|52254009|SNOMEDCT_CORE|NS - Nephrotic syndrome|Nephrotic syndrome
C0027796|T184|PT|16269008|SNOMEDCT_CORE|Neuralgia|Neuralgia
C0027796|T184|FN|16269008|SNOMEDCT_CORE|Neuralgia|Neuralgia
C0027796|T184|OF|16269008|SNOMEDCT_CORE|Neuralgia|Neuralgia
C0027796|T184|IS|16269008|SNOMEDCT_CORE|Neuralgia, NOS|Neuralgia
C0027804|T048|IS|78667006|SNOMEDCT_CORE|Nervous debility|Neurasthenia
C0027804|T048|IS|78667006|SNOMEDCT_CORE|Neurasthaenia|Neurasthenia
C0027804|T048|IS|78667006|SNOMEDCT_CORE|Neurasthaenic neurosis|Neurasthenia
C0027804|T048|IS|78667006|SNOMEDCT_CORE|Neurasthenia|Neurasthenia
C0027804|T048|IS|78667006|SNOMEDCT_CORE|Neurasthenic neurosis|Neurasthenia
C0027809|T191|SY|189948006|SNOMEDCT_CORE|Neurilemmoma|Schwannoma
C0027809|T191|OAP|404022001|SNOMEDCT_CORE|Neurilemmoma|Schwannoma
C0027809|T191|OAF|404022001|SNOMEDCT_CORE|Neurilemmoma|Schwannoma
C0027809|T191|OAS|404022001|SNOMEDCT_CORE|Neurilemoma|Schwannoma
C0027809|T191|PT|189948006|SNOMEDCT_CORE|Schwannoma|Schwannoma
C0027809|T191|OAS|404022001|SNOMEDCT_CORE|Schwannoma|Schwannoma
C0027809|T191|OF|189948006|SNOMEDCT_CORE|Schwannoma|Schwannoma
C0027809|T191|FN|189948006|SNOMEDCT_CORE|Schwannoma|Schwannoma
C0027813|T047|OAP|84299009|SNOMEDCT_CORE|Neuritis|Neuritis
C0027813|T047|SY|21018002|SNOMEDCT_CORE|Neuritis|Neuritis
C0027813|T047|OAF|84299009|SNOMEDCT_CORE|Neuritis|Neuritis
C0027813|T047|IS|84299009|SNOMEDCT_CORE|Neuritis, NOS|Neuritis
C0027813|T047|IS|84299009|SNOMEDCT_CORE|Peripheral neuritis, NOS|Neuritis
C0027819|T191|PT|432328008|SNOMEDCT_CORE|Neuroblastoma|Neuroblastoma
C0027819|T191|FN|432328008|SNOMEDCT_CORE|Neuroblastoma|Neuroblastoma
C0027822|T047|OAP|267854005|SNOMEDCT_CORE|Neurodermatitis|Neurodermatitis
C0027822|T047|OAF|267854005|SNOMEDCT_CORE|Neurodermatitis|Neurodermatitis
C0027830|T191|PT|404029005|SNOMEDCT_CORE|Neurofibroma|Neurofibroma
C0027830|T191|FN|404029005|SNOMEDCT_CORE|Neurofibroma|Neurofibroma
C0027831|T191|IS|92824003|SNOMEDCT_CORE|Clinical von Reclinghausen's disease|Neurofibromatosis type 1
C0027831|T191|SY|92824003|SNOMEDCT_CORE|Multiple non-ossifying fibromatosis|Neurofibromatosis type 1
C0027831|T191|SY|92824003|SNOMEDCT_CORE|Neurofibromatosis 1|Neurofibromatosis type 1
C0027831|T191|PT|92824003|SNOMEDCT_CORE|Neurofibromatosis type 1|Neurofibromatosis type 1
C0027831|T191|FN|92824003|SNOMEDCT_CORE|Neurofibromatosis type 1|Neurofibromatosis type 1
C0027831|T191|SY|92824003|SNOMEDCT_CORE|Neurofibromatosis, peripheral type|Neurofibromatosis type 1
C0027831|T191|OP|92824003|SNOMEDCT_CORE|Neurofibromatosis, type 1|Neurofibromatosis type 1
C0027831|T191|OF|92824003|SNOMEDCT_CORE|Neurofibromatosis, type 1|Neurofibromatosis type 1
C0027831|T191|IS|92824003|SNOMEDCT_CORE|NF1|Neurofibromatosis type 1
C0027831|T191|SY|92824003|SNOMEDCT_CORE|NF1 - Neurofibromatosis type 1|Neurofibromatosis type 1
C0027831|T191|SY|92824003|SNOMEDCT_CORE|Von Recklinghausen disease|Neurofibromatosis type 1
C0027832|T191|SY|92503002|SNOMEDCT_CORE|BANF - Bilateral acoustic neurofibromatosis|Neurofibromatosis type 2
C0027832|T191|SY|92503002|SNOMEDCT_CORE|Bilateral acoustic neurofibromatosis|Neurofibromatosis type 2
C0027832|T191|SY|92503002|SNOMEDCT_CORE|Familial acoustic neuroma|Neurofibromatosis type 2
C0027832|T191|SY|92503002|SNOMEDCT_CORE|Familial vestibular schwannoma|Neurofibromatosis type 2
C0027832|T191|PT|92503002|SNOMEDCT_CORE|Neurofibromatosis type 2|Neurofibromatosis type 2
C0027832|T191|FN|92503002|SNOMEDCT_CORE|Neurofibromatosis type 2|Neurofibromatosis type 2
C0027832|T191|SY|92503002|SNOMEDCT_CORE|Neurofibromatosis, central type|Neurofibromatosis type 2
C0027832|T191|OP|92503002|SNOMEDCT_CORE|Neurofibromatosis, type 2|Neurofibromatosis type 2
C0027832|T191|OF|92503002|SNOMEDCT_CORE|Neurofibromatosis, type 2|Neurofibromatosis type 2
C0027832|T191|SY|92503002|SNOMEDCT_CORE|NF2|Neurofibromatosis type 2
C0027858|T191|SY|25169009|SNOMEDCT_CORE|Neuroma|Neuroma
C0027858|T191|PT|443892003|SNOMEDCT_CORE|Neuroma|Neuroma
C0027858|T191|OF|25169009|SNOMEDCT_CORE|Neuroma|Neuroma
C0027858|T191|FN|443892003|SNOMEDCT_CORE|Neuroma|Neuroma
C0027858|T191|PT|25169009|SNOMEDCT_CORE|Neuroma, no ICD-O subtype|Neuroma
C0027858|T191|OF|25169009|SNOMEDCT_CORE|Neuroma, no ICD-O subtype|Neuroma
C0027858|T191|FN|25169009|SNOMEDCT_CORE|Neuroma, no International Classification of Diseases for Oncology subtype|Neuroma
C0027858|T191|SY|25169009|SNOMEDCT_CORE|Neuroma, no International Classification of Diseases for Oncology subtype|Neuroma
C0027858|T191|IS|25169009|SNOMEDCT_CORE|Neuroma, NOS|Neuroma
C0027859|T191|SY|126949007|SNOMEDCT_CORE|Acoustic neurilemmoma|Acoustic neuroma
C0027859|T191|SY|126949007|SNOMEDCT_CORE|Acoustic neurinoma|Acoustic neuroma
C0027859|T191|PT|126949007|SNOMEDCT_CORE|Acoustic neuroma|Acoustic neuroma
C0027859|T191|FN|126949007|SNOMEDCT_CORE|Acoustic neuroma|Acoustic neuroma
C0027859|T191|SY|126949007|SNOMEDCT_CORE|Acoustic schwannoma|Acoustic neuroma
C0027859|T191|SY|126949007|SNOMEDCT_CORE|AN - Acoustic neuroma|Acoustic neuroma
C0027859|T191|SY|126949007|SNOMEDCT_CORE|Vestibular schwannoma|Acoustic neuroma
C0027888|T047|SY|398100001|SNOMEDCT_CORE|CMT - Charcot-Marie-Tooth disease|Hereditary motor and sensory neuropathy
C0027888|T047|PT|398100001|SNOMEDCT_CORE|Hereditary motor and sensory neuropathy|Hereditary motor and sensory neuropathy
C0027888|T047|FN|398100001|SNOMEDCT_CORE|Hereditary motor and sensory neuropathy|Hereditary motor and sensory neuropathy
C0027888|T047|SY|398100001|SNOMEDCT_CORE|Hereditary sensorimotor neuropathy|Hereditary motor and sensory neuropathy
C0027888|T047|SY|398100001|SNOMEDCT_CORE|Hereditary sensory and motor neuropathy|Hereditary motor and sensory neuropathy
C0027888|T047|SY|398100001|SNOMEDCT_CORE|Hereditary sensory-motor neuropathy|Hereditary motor and sensory neuropathy
C0027888|T047|SY|398100001|SNOMEDCT_CORE|HMSN|Hereditary motor and sensory neuropathy
C0027888|T047|SY|398100001|SNOMEDCT_CORE|HMSN - Hereditary motor and sensory neuropathy|Hereditary motor and sensory neuropathy
C0027888|T047|SY|398100001|SNOMEDCT_CORE|HSMN|Hereditary motor and sensory neuropathy
C0027888|T047|SY|398100001|SNOMEDCT_CORE|HSMN - Hereditary sensory and motor neuropathy|Hereditary motor and sensory neuropathy
C0027927|T047|PT|26039008|SNOMEDCT_CORE|Neurosyphilis|Neurosyphilis
C0027927|T047|FN|26039008|SNOMEDCT_CORE|Neurosyphilis|Neurosyphilis
C0027927|T047|IS|26039008|SNOMEDCT_CORE|Neurosyphilis, NOS|Neurosyphilis
C0027927|T047|SY|26039008|SNOMEDCT_CORE|Syphilis of central nervous system|Neurosyphilis
C0027927|T047|IS|26039008|SNOMEDCT_CORE|Syphilis of central nervous system, NOS|Neurosyphilis
C0027947|T047|IS|303011007|SNOMEDCT_CORE|Neutropenia|Neutropenic disorder
C0027947|T047|PT|303011007|SNOMEDCT_CORE|Neutropenic disorder|Neutropenic disorder
C0027947|T047|FN|303011007|SNOMEDCT_CORE|Neutropenic disorder|Neutropenic disorder
C0027962|T191|PTGB|400096001|SNOMEDCT_CORE|Melanocytic naevus|Melanocytic nevus
C0027962|T191|PT|400096001|SNOMEDCT_CORE|Melanocytic nevus|Melanocytic nevus
C0027962|T191|FN|400096001|SNOMEDCT_CORE|Melanocytic nevus|Melanocytic nevus
C0027962|T191|SY|400096001|SNOMEDCT_CORE|Mole|Melanocytic nevus
C0028043|T048|PT|56294008|SNOMEDCT_CORE|Nicotine dependence|Nicotine dependence
C0028043|T048|FN|56294008|SNOMEDCT_CORE|Nicotine dependence|Nicotine dependence
C0028081|T184|PT|42984000|SNOMEDCT_CORE|Night sweats|Night sweats
C0028081|T184|FN|42984000|SNOMEDCT_CORE|Night sweats|Night sweats
C0028084|T184|PT|419145002|SNOMEDCT_CORE|Nightmares|Nightmares
C0028084|T184|FN|419145002|SNOMEDCT_CORE|Nightmares|Nightmares
C0028431|T020|SY|18283000|SNOMEDCT_CORE|Acquired anomaly of nose|Acquired deformity of nose
C0028431|T020|PT|18283000|SNOMEDCT_CORE|Acquired deformity of nose|Acquired deformity of nose
C0028431|T020|FN|18283000|SNOMEDCT_CORE|Acquired deformity of nose|Acquired deformity of nose
C0028431|T020|SY|18283000|SNOMEDCT_CORE|Acquired nasal deformity|Acquired deformity of nose
C0028643|T184|SY|44077006|SNOMEDCT_CORE|Deadness - numbness|Numbness
C0028643|T184|SY|44077006|SNOMEDCT_CORE|Loss of sensation|Numbness
C0028643|T184|PT|44077006|SNOMEDCT_CORE|Numbness|Numbness
C0028643|T184|FN|44077006|SNOMEDCT_CORE|Numbness|Numbness
C0028734|T047|OAF|6408001|SNOMEDCT_CORE|Finding of nocturia|Nocturia
C0028734|T047|OAS|6408001|SNOMEDCT_CORE|Finding of nocturia|Nocturia
C0028734|T047|IS|6408001|SNOMEDCT_CORE|Nocturia|Nocturia
C0028734|T047|OF|139394000|SNOMEDCT_CORE|Nocturia|Nocturia
C0028734|T047|PT|139394000|SNOMEDCT_CORE|Nocturia|Nocturia
C0028734|T047|FN|139394000|SNOMEDCT_CORE|Nocturia|Nocturia
C0028734|T047|OAP|6408001|SNOMEDCT_CORE|Nocturia - finding|Nocturia
C0028734|T047|OAS|6408001|SNOMEDCT_CORE|Nycturia|Nocturia
C0028738|T047|PT|563001|SNOMEDCT_CORE|Nystagmus|Nystagmus
C0028738|T047|FN|563001|SNOMEDCT_CORE|Nystagmus|Nystagmus
C0028738|T047|IS|563001|SNOMEDCT_CORE|Nystagmus, NOS|Nystagmus
C0028754|T047|PT|414916001|SNOMEDCT_CORE|Obesity|Obesity
C0028754|T047|FN|414916001|SNOMEDCT_CORE|Obesity|Obesity
C0028756|T047|PT|238136002|SNOMEDCT_CORE|Morbid obesity|Morbid obesity
C0028756|T047|FN|238136002|SNOMEDCT_CORE|Morbid obesity|Morbid obesity
C0028768|T048|SY|191736004|SNOMEDCT_CORE|Anancastic neurosis|Obsessive-compulsive disorder
C0028768|T048|SY|191736004|SNOMEDCT_CORE|Anankastic neurosis|Obsessive-compulsive disorder
C0028768|T048|SY|191736004|SNOMEDCT_CORE|Obsessive compulsive disorder|Obsessive-compulsive disorder
C0028768|T048|SY|191736004|SNOMEDCT_CORE|Obsessive compulsive neurosis|Obsessive-compulsive disorder
C0028768|T048|PT|191736004|SNOMEDCT_CORE|Obsessive-compulsive disorder|Obsessive-compulsive disorder
C0028768|T048|FN|191736004|SNOMEDCT_CORE|Obsessive-compulsive disorder|Obsessive-compulsive disorder
C0028768|T048|SY|191736004|SNOMEDCT_CORE|OCD - Obsessive-compulsive disorder|Obsessive-compulsive disorder
C0028797|T047|PT|115966001|SNOMEDCT_CORE|Occupational disorder|Occupational disorder
C0028797|T047|FN|115966001|SNOMEDCT_CORE|Occupational disorder|Occupational disorder
C0028840|T047|PT|4210003|SNOMEDCT_CORE|Ocular hypertension|Ocular hypertension
C0028840|T047|FN|4210003|SNOMEDCT_CORE|Ocular hypertension|Ocular hypertension
C0028840|T047|SY|4210003|SNOMEDCT_CORE|OH - Ocular hypertension|Ocular hypertension
C0028840|T047|SY|4210003|SNOMEDCT_CORE|OHT - Ocular hypertension|Ocular hypertension
C0028879|T047|PT|235110008|SNOMEDCT_CORE|Odontogenic cyst|Odontogenic cyst
C0028879|T047|FN|235110008|SNOMEDCT_CORE|Odontogenic cyst|Odontogenic cyst
C0028945|T191|SY|73348003|SNOMEDCT_CORE|Oligodendroglioma|Oligodendroglioma, no ICD-O subtype
C0028945|T191|OF|73348003|SNOMEDCT_CORE|Oligodendroglioma|Oligodendroglioma, no ICD-O subtype
C0028945|T191|PT|73348003|SNOMEDCT_CORE|Oligodendroglioma, no ICD-O subtype|Oligodendroglioma, no ICD-O subtype
C0028945|T191|OF|73348003|SNOMEDCT_CORE|Oligodendroglioma, no ICD-O subtype|Oligodendroglioma, no ICD-O subtype
C0028945|T191|FN|73348003|SNOMEDCT_CORE|Oligodendroglioma, no International Classification of Diseases for Oncology subtype|Oligodendroglioma, no ICD-O subtype
C0028945|T191|SY|73348003|SNOMEDCT_CORE|Oligodendroglioma, no International Classification of Diseases for Oncology subtype|Oligodendroglioma, no ICD-O subtype
C0028945|T191|IS|73348003|SNOMEDCT_CORE|Oligodendroglioma, NOS|Oligodendroglioma, no ICD-O subtype
C0028949|T046|IS|52073004|SNOMEDCT_CORE|Abnormal long menstrual cycle|Oligomenorrhea
C0028949|T046|SY|52073004|SNOMEDCT_CORE|Infrequent menstruation|Oligomenorrhea
C0028949|T046|OF|52073004|SNOMEDCT_CORE|Infrequent menstruation|Oligomenorrhea
C0028949|T046|SY|52073004|SNOMEDCT_CORE|Infrequent periods|Oligomenorrhea
C0028949|T046|PT|52073004|SNOMEDCT_CORE|Oligomenorrhea|Oligomenorrhea
C0028949|T046|FN|52073004|SNOMEDCT_CORE|Oligomenorrhea|Oligomenorrhea
C0028949|T046|PTGB|52073004|SNOMEDCT_CORE|Oligomenorrhoea|Oligomenorrhea
C0028949|T046|SY|52073004|SNOMEDCT_CORE|Relative amenorrhea|Oligomenorrhea
C0028949|T046|SYGB|52073004|SNOMEDCT_CORE|Relative amenorrhoea|Oligomenorrhea
C0029095|T048|PT|5602001|SNOMEDCT_CORE|Opioid abuse|Opioid abuse
C0029095|T048|FN|5602001|SNOMEDCT_CORE|Opioid abuse|Opioid abuse
C0029100|T048|PT|77721001|SNOMEDCT_CORE|Opioid intoxication|Opioid intoxication
C0029100|T048|FN|77721001|SNOMEDCT_CORE|Opioid intoxication|Opioid intoxication
C0029104|T048|SY|87132004|SNOMEDCT_CORE|Narcotic withdrawal|Opioid withdrawal
C0029104|T048|PT|87132004|SNOMEDCT_CORE|Opioid withdrawal|Opioid withdrawal
C0029104|T048|FN|87132004|SNOMEDCT_CORE|Opioid withdrawal|Opioid withdrawal
C0029121|T048|PT|18941000|SNOMEDCT_CORE|Oppositional defiant disorder|Oppositional defiant disorder
C0029121|T048|FN|18941000|SNOMEDCT_CORE|Oppositional defiant disorder|Oppositional defiant disorder
C0029124|T047|SY|76976005|SNOMEDCT_CORE|OA - Optic atrophy|Optic atrophy
C0029124|T047|PT|76976005|SNOMEDCT_CORE|Optic atrophy|Optic atrophy
C0029124|T047|FN|76976005|SNOMEDCT_CORE|Optic atrophy|Optic atrophy
C0029124|T047|IS|76976005|SNOMEDCT_CORE|Optic atrophy, NOS|Optic atrophy
C0029124|T047|SY|76976005|SNOMEDCT_CORE|Optic nerve atrophy|Optic atrophy
C0029128|T047|PT|33629003|SNOMEDCT_CORE|Drusen of optic disc|Drusen of optic disc
C0029128|T047|FN|33629003|SNOMEDCT_CORE|Drusen of optic disc|Drusen of optic disc
C0029128|T047|OF|33629003|SNOMEDCT_CORE|Drusen of optic disc|Drusen of optic disc
C0029128|T047|SY|33629003|SNOMEDCT_CORE|Hyaline bodies of optic disc|Drusen of optic disc
C0029128|T047|SY|33629003|SNOMEDCT_CORE|Optic disc drusen|Drusen of optic disc
C0029128|T047|SY|33629003|SNOMEDCT_CORE|Optic nerve head drusen|Drusen of optic disc
C0029132|T047|PT|77157004|SNOMEDCT_CORE|Disorder of optic nerve|Disorder of optic nerve
C0029132|T047|FN|77157004|SNOMEDCT_CORE|Disorder of optic nerve|Disorder of optic nerve
C0029132|T047|IS|77157004|SNOMEDCT_CORE|Disorder of optic nerve, NOS|Disorder of optic nerve
C0029132|T047|SY|77157004|SNOMEDCT_CORE|Optic neuropathy|Disorder of optic nerve
C0029134|T047|SY|66760008|SNOMEDCT_CORE|ON - Optic neuritis|Optic neuritis
C0029134|T047|PT|66760008|SNOMEDCT_CORE|Optic neuritis|Optic neuritis
C0029134|T047|FN|66760008|SNOMEDCT_CORE|Optic neuritis|Optic neuritis
C0029134|T047|IS|66760008|SNOMEDCT_CORE|Optic neuritis, NOS|Optic neuritis
C0029184|T037|PT|95851007|SNOMEDCT_CORE|Fracture of orbit|Fracture of orbit
C0029184|T037|FN|95851007|SNOMEDCT_CORE|Fracture of orbit|Fracture of orbit
C0029184|T037|IS|95851007|SNOMEDCT_CORE|Fracture of orbit, NOS|Fracture of orbit
C0029184|T037|IS|95851007|SNOMEDCT_CORE|Fracture of orbital bones|Fracture of orbit
C0029184|T037|IS|95851007|SNOMEDCT_CORE|Fracture of orbital bones, NOS|Fracture of orbit
C0029184|T037|SY|95851007|SNOMEDCT_CORE|Fracture of orbital fossa|Fracture of orbit
C0029184|T037|SY|95851007|SNOMEDCT_CORE|Orbital fracture|Fracture of orbit
C0029184|T037|IS|95851007|SNOMEDCT_CORE|Orbital fracture, NOS|Fracture of orbit
C0029191|T047|SY|274718005|SNOMEDCT_CORE|Inflammation of testis|Orchitis
C0029191|T047|SY|274718005|SNOMEDCT_CORE|Non-specific orchitis|Orchitis
C0029191|T047|PT|274718005|SNOMEDCT_CORE|Orchitis|Orchitis
C0029191|T047|FN|274718005|SNOMEDCT_CORE|Orchitis|Orchitis
C0029191|T047|IS|274718005|SNOMEDCT_CORE|Orchititis|Orchitis
C0029221|T047|SY|2776000|SNOMEDCT_CORE|OBS - Organic brain syndrome|Organic brain syndrome
C0029221|T047|SY|2776000|SNOMEDCT_CORE|Organic brain syndrome|Organic brain syndrome
C0029221|T047|IS|2776000|SNOMEDCT_CORE|Organic brain syndrome, NOS|Organic brain syndrome
C0029225|T048|PT|5510009|SNOMEDCT_CORE|Organic delusional disorder|Organic delusional disorder
C0029225|T048|FN|5510009|SNOMEDCT_CORE|Organic delusional disorder|Organic delusional disorder
C0029225|T048|IS|5510009|SNOMEDCT_CORE|Organic delusional disorder, NOS|Organic delusional disorder
C0029227|T048|PT|111479008|SNOMEDCT_CORE|Organic mental disorder|Organic mental disorder
C0029227|T048|FN|111479008|SNOMEDCT_CORE|Organic mental disorder|Organic mental disorder
C0029227|T048|IS|111479008|SNOMEDCT_CORE|Organic mental disorder, NOS|Organic mental disorder
C0029232|T048|SY|23645006|SNOMEDCT_CORE|Organic affective disorder|Organic mood disorder
C0029232|T048|PT|23645006|SNOMEDCT_CORE|Organic mood disorder|Organic mood disorder
C0029232|T048|FN|23645006|SNOMEDCT_CORE|Organic mood disorder|Organic mood disorder
C0029232|T048|IS|23645006|SNOMEDCT_CORE|Organic mood disorder, NOS|Organic mood disorder
C0029295|T191|PT|126809003|SNOMEDCT_CORE|Neoplasm of oropharynx|Neoplasm of oropharynx
C0029295|T191|FN|126809003|SNOMEDCT_CORE|Neoplasm of oropharynx|Neoplasm of oropharynx
C0029295|T191|SY|126809003|SNOMEDCT_CORE|Tumor of oropharynx|Neoplasm of oropharynx
C0029295|T191|SYGB|126809003|SNOMEDCT_CORE|Tumour of oropharynx|Neoplasm of oropharynx
C0029376|T047|SY|72047008|SNOMEDCT_CORE|Juvenile osteochondrosis of tibial tubercle|Osgood Schlatter disease
C0029376|T047|FN|72047008|SNOMEDCT_CORE|Juvenile osteochondrosis of tibial tubercle|Osgood Schlatter disease
C0029376|T047|PT|72047008|SNOMEDCT_CORE|Osgood Schlatter disease|Osgood Schlatter disease
C0029376|T047|SY|72047008|SNOMEDCT_CORE|Osgood Schlatters disease|Osgood Schlatter disease
C0029376|T047|SY|72047008|SNOMEDCT_CORE|Osgood-Schlatter's disease|Osgood Schlatter disease
C0029401|T047|PT|2089002|SNOMEDCT_CORE|Osteitis deformans|Osteitis deformans
C0029401|T047|FN|2089002|SNOMEDCT_CORE|Osteitis deformans|Osteitis deformans
C0029401|T047|SY|2089002|SNOMEDCT_CORE|Paget's disease of bone|Osteitis deformans
C0029401|T047|SY|2089002|SNOMEDCT_CORE|Pagets disease of bone|Osteitis deformans
C0029403|T047|IS|2089002|SNOMEDCT_CORE|Osteitis deformans without mention of bone tumor|Osteitis deformans without mention of bone tumor
C0029408|T047|SY|396275006|SNOMEDCT_CORE|Degenerative arthritis|Osteoarthritis
C0029408|T047|SY|396275006|SNOMEDCT_CORE|Degenerative arthropathy|Osteoarthritis
C0029408|T047|SY|396275006|SNOMEDCT_CORE|Degenerative joint disease|Osteoarthritis
C0029408|T047|IS|396275006|SNOMEDCT_CORE|Degenerative polyarthritis|Osteoarthritis
C0029408|T047|SY|396275006|SNOMEDCT_CORE|Hypertrophic arthritis|Osteoarthritis
C0029408|T047|SY|396275006|SNOMEDCT_CORE|Hypertrophic polyarthritis|Osteoarthritis
C0029408|T047|SY|396275006|SNOMEDCT_CORE|OA - Osteoarthritis|Osteoarthritis
C0029408|T047|SY|396275006|SNOMEDCT_CORE|OA - Osteoarthrosis|Osteoarthritis
C0029408|T047|PT|396275006|SNOMEDCT_CORE|Osteoarthritis|Osteoarthritis
C0029408|T047|FN|396275006|SNOMEDCT_CORE|Osteoarthritis|Osteoarthritis
C0029408|T047|SY|396275006|SNOMEDCT_CORE|Osteoarthrosis|Osteoarthritis
C0029410|T047|SY|239872002|SNOMEDCT_CORE|Degenerative joint disease of hip|Osteoarthritis of hip
C0029410|T047|SY|239872002|SNOMEDCT_CORE|OA - Osteoarthritis of hip|Osteoarthritis of hip
C0029410|T047|PT|239872002|SNOMEDCT_CORE|Osteoarthritis of hip|Osteoarthritis of hip
C0029410|T047|FN|239872002|SNOMEDCT_CORE|Osteoarthritis of hip|Osteoarthritis of hip
C0029421|T047|SY|82562007|SNOMEDCT_CORE|Idiopathic avascular necrosis|Osteochondritis dissecans
C0029421|T047|IS|82562007|SNOMEDCT_CORE|OCC|Osteochondritis dissecans
C0029421|T047|IS|82562007|SNOMEDCT_CORE|OCD|Osteochondritis dissecans
C0029421|T047|SY|82562007|SNOMEDCT_CORE|OCD - Osteochondritis dissecans|Osteochondritis dissecans
C0029421|T047|SY|82562007|SNOMEDCT_CORE|OD - Osteochondritis dissecans|Osteochondritis dissecans
C0029421|T047|PT|82562007|SNOMEDCT_CORE|Osteochondritis dissecans|Osteochondritis dissecans
C0029421|T047|FN|82562007|SNOMEDCT_CORE|Osteochondritis dissecans|Osteochondritis dissecans
C0029421|T047|IS|82562007|SNOMEDCT_CORE|Osteochondrosis dessicans|Osteochondritis dissecans
C0029421|T047|SY|82562007|SNOMEDCT_CORE|Osteochondrosis dissecans|Osteochondritis dissecans
C0029423|T191|SY|52299001|SNOMEDCT_CORE|Cartilaginous exostosis|Osteochondroma
C0029423|T191|SY|52299001|SNOMEDCT_CORE|Ecchondroma|Osteochondroma
C0029423|T191|SY|52299001|SNOMEDCT_CORE|Osteocartilaginous exostosis|Osteochondroma
C0029423|T191|PT|443093007|SNOMEDCT_CORE|Osteochondroma|Osteochondroma
C0029423|T191|PT|52299001|SNOMEDCT_CORE|Osteochondroma|Osteochondroma
C0029423|T191|FN|52299001|SNOMEDCT_CORE|Osteochondroma|Osteochondroma
C0029423|T191|FN|443093007|SNOMEDCT_CORE|Osteochondroma|Osteochondroma
C0029434|T047|SY|78314001|SNOMEDCT_CORE|Brittle bone disease|Osteogenesis imperfecta
C0029434|T047|SY|78314001|SNOMEDCT_CORE|Brittle bone syndrome|Osteogenesis imperfecta
C0029434|T047|SY|78314001|SNOMEDCT_CORE|Fragilitas ossium|Osteogenesis imperfecta
C0029434|T047|SY|78314001|SNOMEDCT_CORE|OI - Osteogenesis imperfecta|Osteogenesis imperfecta
C0029434|T047|PT|78314001|SNOMEDCT_CORE|Osteogenesis imperfecta|Osteogenesis imperfecta
C0029434|T047|FN|78314001|SNOMEDCT_CORE|Osteogenesis imperfecta|Osteogenesis imperfecta
C0029434|T047|IS|78314001|SNOMEDCT_CORE|Osteogenesis imperfecta, NOS|Osteogenesis imperfecta
C0029434|T047|SY|78314001|SNOMEDCT_CORE|Osteopsathyrosis|Osteogenesis imperfecta
C0029442|T047|SY|4598005|SNOMEDCT_CORE|OM - Osteomalacia|Osteomalacia
C0029442|T047|PT|4598005|SNOMEDCT_CORE|Osteomalacia|Osteomalacia
C0029442|T047|FN|4598005|SNOMEDCT_CORE|Osteomalacia|Osteomalacia
C0029443|T047|SY|60168000|SNOMEDCT_CORE|OM - Osteomyelitis|Osteomyelitis
C0029443|T047|PT|60168000|SNOMEDCT_CORE|Osteomyelitis|Osteomyelitis
C0029443|T047|FN|60168000|SNOMEDCT_CORE|Osteomyelitis|Osteomyelitis
C0029443|T047|IS|60168000|SNOMEDCT_CORE|Osteomyelitis, NOS|Osteomyelitis
C0029443|T047|SY|60168000|SNOMEDCT_CORE|OSTM - Osteomyelitis|Osteomyelitis
C0029443|T047|SY|60168000|SNOMEDCT_CORE|Pyogenic inflammation of bone|Osteomyelitis
C0029443|T047|IS|60168000|SNOMEDCT_CORE|Pyogenic inflammation of bone, NOS|Osteomyelitis
C0029445|T046|PT|240196003|SNOMEDCT_CORE|Bone necrosis|Bone necrosis
C0029445|T046|FN|240196003|SNOMEDCT_CORE|Bone necrosis|Bone necrosis
C0029445|T046|IS|398199007|SNOMEDCT_CORE|Osteonecrosis|Bone necrosis
C0029445|T046|SY|240196003|SNOMEDCT_CORE|Osteonecrosis|Bone necrosis
C0029453|T047|PT|312894000|SNOMEDCT_CORE|Osteopenia|Osteopenia
C0029453|T047|FN|312894000|SNOMEDCT_CORE|Osteopenia|Osteopenia
C0029454|T047|IS|367489004|SNOMEDCT_CORE|Albers-Sch?nberg disease|Marble bone disease
C0029454|T047|IS|367489004|SNOMEDCT_CORE|Albers-Scho@nberg syndrome|Marble bone disease
C0029454|T047|IS|367489004|SNOMEDCT_CORE|Albers-Schoenberg syndrome|Marble bone disease
C0029454|T047|IS|367489004|SNOMEDCT_CORE|Albers-Schönberg disease|Marble bone disease
C0029454|T047|IS|367489004|SNOMEDCT_CORE|Albers-Schonberg syndrome|Marble bone disease
C0029454|T047|SY|367489004|SNOMEDCT_CORE|Congenital osteopetrosis|Marble bone disease
C0029454|T047|IS|367489004|SNOMEDCT_CORE|Ivory bones|Marble bone disease
C0029454|T047|SY|367489004|SNOMEDCT_CORE|Marble bone disease|Marble bone disease
C0029454|T047|IS|367489004|SNOMEDCT_CORE|Osteopetrosis - congenita type|Marble bone disease
C0029454|T047|IS|367489004|SNOMEDCT_CORE|Osteopetrosis generalisata|Marble bone disease
C0029456|T047|IS|64859006|SNOMEDCT_CORE|OP - Osteoporosis|Osteoporosis
C0029456|T047|PT|64859006|SNOMEDCT_CORE|Osteoporosis|Osteoporosis
C0029456|T047|FN|64859006|SNOMEDCT_CORE|Osteoporosis|Osteoporosis
C0029456|T047|IS|64859006|SNOMEDCT_CORE|Osteoporosis, NOS|Osteoporosis
C0029458|T047|PT|102447009|SNOMEDCT_CORE|Postmenopausal osteoporosis|Postmenopausal osteoporosis
C0029458|T047|FN|102447009|SNOMEDCT_CORE|Postmenopausal osteoporosis|Postmenopausal osteoporosis
C0029459|T047|SY|18040001|SNOMEDCT_CORE|Age related osteoporosis|Senile osteoporosis
C0029459|T047|SY|18040001|SNOMEDCT_CORE|Involutional osteoporosis|Senile osteoporosis
C0029459|T047|PT|18040001|SNOMEDCT_CORE|Senile osteoporosis|Senile osteoporosis
C0029459|T047|FN|18040001|SNOMEDCT_CORE|Senile osteoporosis|Senile osteoporosis
C0029459|T047|SY|18040001|SNOMEDCT_CORE|Type II osteoporosis|Senile osteoporosis
C0029463|T191|SY|307576001|SNOMEDCT_CORE|Osteosarcoma|Osteosarcoma
C0029463|T191|SY|307576001|SNOMEDCT_CORE|Osteosarcoma - disorder|Osteosarcoma
C0029877|T047|SY|43275000|SNOMEDCT_CORE|Inflammatory disorder of ear|Otitis
C0029877|T047|PT|43275000|SNOMEDCT_CORE|Otitis|Otitis
C0029877|T047|FN|43275000|SNOMEDCT_CORE|Otitis|Otitis
C0029877|T047|IS|43275000|SNOMEDCT_CORE|Otitis, NOS|Otitis
C0029878|T047|SY|3135009|SNOMEDCT_CORE|Inflammation of ear canal|Otitis externa
C0029878|T047|SY|3135009|SNOMEDCT_CORE|OE - Otitis externa|Otitis externa
C0029878|T047|PT|3135009|SNOMEDCT_CORE|Otitis externa|Otitis externa
C0029878|T047|FN|3135009|SNOMEDCT_CORE|Otitis externa|Otitis externa
C0029878|T047|IS|3135009|SNOMEDCT_CORE|Otitis externa, NOS|Otitis externa
C0029882|T047|SY|65363002|SNOMEDCT_CORE|OM - Otitis media|Otitis media
C0029882|T047|PT|65363002|SNOMEDCT_CORE|Otitis media|Otitis media
C0029882|T047|FN|65363002|SNOMEDCT_CORE|Otitis media|Otitis media
C0029882|T047|IS|65363002|SNOMEDCT_CORE|Otitis media, NOS|Otitis media
C0029883|T047|SY|78868004|SNOMEDCT_CORE|Glue ear|Secretory otitis media
C0029883|T047|SY|78868004|SNOMEDCT_CORE|Glue ear - mucoid|Secretory otitis media
C0029883|T047|SY|78868004|SNOMEDCT_CORE|Mucoid otitis media|Secretory otitis media
C0029883|T047|SY|78868004|SNOMEDCT_CORE|OME - Otitis media with effusion|Secretory otitis media
C0029883|T047|SY|78868004|SNOMEDCT_CORE|Otitis media with effusion|Secretory otitis media
C0029883|T047|SY|78868004|SNOMEDCT_CORE|Otitis media with effusion - mucoid|Secretory otitis media
C0029883|T047|SY|78868004|SNOMEDCT_CORE|Secretory otitis media|Secretory otitis media
C0029883|T047|SY|78868004|SNOMEDCT_CORE|SOM - Secretory otitis media|Secretory otitis media
C0029883|T047|SY|78868004|SNOMEDCT_CORE|Transudative otitis media|Secretory otitis media
C0029888|T047|SY|38394007|SNOMEDCT_CORE|Otitis media with effusion - purulent|Otitis media with effusion - purulent
C0029899|T047|PT|11543004|SNOMEDCT_CORE|Otosclerosis|Otosclerosis
C0029899|T047|FN|11543004|SNOMEDCT_CORE|Otosclerosis|Otosclerosis
C0029899|T047|IS|11543004|SNOMEDCT_CORE|Otosclerosis, NOS|Otosclerosis
C0029899|T047|SY|11543004|SNOMEDCT_CORE|Otospongiosis|Otosclerosis
C0029899|T047|IS|11543004|SNOMEDCT_CORE|Otospongiosis, NOS|Otosclerosis
C0029927|T047|IS|79883001|SNOMEDCT_CORE|Benign retention cyst|Cyst of ovary
C0029927|T047|PT|79883001|SNOMEDCT_CORE|Cyst of ovary|Cyst of ovary
C0029927|T047|FN|79883001|SNOMEDCT_CORE|Cyst of ovary|Cyst of ovary
C0029927|T047|SY|79883001|SNOMEDCT_CORE|Ovarian cyst|Cyst of ovary
C0029927|T047|IS|79883001|SNOMEDCT_CORE|Ovarian cyst, NOS|Cyst of ovary
C0029927|T047|SY|79883001|SNOMEDCT_CORE|Ovarian cystic mass|Cyst of ovary
C0029927|T047|IS|79883001|SNOMEDCT_CORE|Ovarian retention cyst|Cyst of ovary
C0029927|T047|IS|79883001|SNOMEDCT_CORE|Ovarian retention cyst, NOS|Cyst of ovary
C0029928|T047|IS|5552004|SNOMEDCT_CORE|Disease of ovary|Disorder of ovary
C0029928|T047|OF|5552004|SNOMEDCT_CORE|Disease of ovary|Disorder of ovary
C0029928|T047|IS|5552004|SNOMEDCT_CORE|Disease of ovary, NOS|Disorder of ovary
C0029928|T047|PT|5552004|SNOMEDCT_CORE|Disorder of ovary|Disorder of ovary
C0029928|T047|FN|5552004|SNOMEDCT_CORE|Disorder of ovary|Disorder of ovary
C0029928|T047|SY|5552004|SNOMEDCT_CORE|Ovarian disorder|Disorder of ovary
C0029928|T047|IS|5552004|SNOMEDCT_CORE|Ovarian disorder, NOS|Disorder of ovary
C0029944|T037|PT|55680006|SNOMEDCT_CORE|Drug overdose|Drug overdose
C0029944|T037|FN|55680006|SNOMEDCT_CORE|Drug overdose|Drug overdose
C0029944|T037|IS|55680006|SNOMEDCT_CORE|Drug overdose, NOS|Drug overdose
C0029944|T037|SY|55680006|SNOMEDCT_CORE|OD - Overdose of drug|Drug overdose
C0029944|T037|SY|55680006|SNOMEDCT_CORE|Overdose|Drug overdose
C0029944|T037|IS|55680006|SNOMEDCT_CORE|Overdose, NOS|Drug overdose
C0030100|T047|SY|266162007|SNOMEDCT_CORE|Oxyuriasis|Oxyuriasis
C0030193|T184|SY|22253000|SNOMEDCT_CORE|Dolor|Pain
C0030193|T184|PT|22253000|SNOMEDCT_CORE|Pain|Pain
C0030193|T184|FN|22253000|SNOMEDCT_CORE|Pain|Pain
C0030193|T184|SY|22253000|SNOMEDCT_CORE|Pain observations|Pain
C0030193|T184|IS|22253000|SNOMEDCT_CORE|Pain, NOS|Pain
C0030193|T184|SY|22253000|SNOMEDCT_CORE|Painful|Pain
C0030193|T184|SY|22253000|SNOMEDCT_CORE|Part hurts|Pain
C0030196|T184|SY|90834002|SNOMEDCT_CORE|Limb pain|Pain in limb
C0030196|T184|IS|90834002|SNOMEDCT_CORE|Limb pain, NOS|Pain in limb
C0030196|T184|PT|90834002|SNOMEDCT_CORE|Pain in limb|Pain in limb
C0030196|T184|FN|90834002|SNOMEDCT_CORE|Pain in limb|Pain in limb
C0030201|T184|PT|213299007|SNOMEDCT_CORE|Postoperative pain|Postoperative pain
C0030201|T184|FN|213299007|SNOMEDCT_CORE|Postoperative pain|Postoperative pain
C0030252|T033|PT|80313002|SNOMEDCT_CORE|Palpitations|Palpitations
C0030252|T033|FN|80313002|SNOMEDCT_CORE|Palpitations|Palpitations
C0030283|T047|PT|31258000|SNOMEDCT_CORE|Cyst of pancreas|Cyst of pancreas
C0030283|T047|FN|31258000|SNOMEDCT_CORE|Cyst of pancreas|Cyst of pancreas
C0030283|T047|SY|31258000|SNOMEDCT_CORE|Pancreatic cyst|Cyst of pancreas
C0030286|T047|IS|3855007|SNOMEDCT_CORE|Disease of pancreas|Disorder of pancreas
C0030286|T047|OF|3855007|SNOMEDCT_CORE|Disease of pancreas|Disorder of pancreas
C0030286|T047|IS|3855007|SNOMEDCT_CORE|Disease of pancreas, NOS|Disorder of pancreas
C0030286|T047|PT|3855007|SNOMEDCT_CORE|Disorder of pancreas|Disorder of pancreas
C0030286|T047|FN|3855007|SNOMEDCT_CORE|Disorder of pancreas|Disorder of pancreas
C0030286|T047|IS|3855007|SNOMEDCT_CORE|Disorder of pancreas, NOS|Disorder of pancreas
C0030293|T047|PT|37992001|SNOMEDCT_CORE|Pancreatic insufficiency|Pancreatic insufficiency
C0030293|T047|FN|37992001|SNOMEDCT_CORE|Pancreatic insufficiency|Pancreatic insufficiency
C0030293|T047|IS|37992001|SNOMEDCT_CORE|Pancreatic insufficiency, NOS|Pancreatic insufficiency
C0030299|T047|SY|111374002|SNOMEDCT_CORE|Pancreatic pseudocyst|Pseudocyst of pancreas
C0030299|T047|PT|111374002|SNOMEDCT_CORE|Pseudocyst of pancreas|Pseudocyst of pancreas
C0030299|T047|FN|111374002|SNOMEDCT_CORE|Pseudocyst of pancreas|Pseudocyst of pancreas
C0030305|T047|SY|75694006|SNOMEDCT_CORE|Inflammation of pancreas|Pancreatitis
C0030305|T047|PT|75694006|SNOMEDCT_CORE|Pancreatitis|Pancreatitis
C0030305|T047|FN|75694006|SNOMEDCT_CORE|Pancreatitis|Pancreatitis
C0030305|T047|IS|75694006|SNOMEDCT_CORE|Pancreatitis, NOS|Pancreatitis
C0030312|T047|IS|127034005|SNOMEDCT_CORE|Bone marrow failure|Pancytopenia
C0030312|T047|PT|127034005|SNOMEDCT_CORE|Pancytopenia|Pancytopenia
C0030312|T047|FN|127034005|SNOMEDCT_CORE|Pancytopenia|Pancytopenia
C0030319|T048|SY|371631005|SNOMEDCT_CORE|Episodic paroxysmal anxiety disorder|Panic disorder
C0030319|T048|PT|371631005|SNOMEDCT_CORE|Panic disorder|Panic disorder
C0030319|T048|FN|371631005|SNOMEDCT_CORE|Panic disorder|Panic disorder
C0030326|T047|PT|22125009|SNOMEDCT_CORE|Panniculitis|Panniculitis
C0030326|T047|FN|22125009|SNOMEDCT_CORE|Panniculitis|Panniculitis
C0030326|T047|IS|22125009|SNOMEDCT_CORE|Panniculitis, NOS|Panniculitis
C0030353|T047|SY|423341008|SNOMEDCT_CORE|Edema of optic disc|Optic disc edema
C0030353|T047|FN|423341008|SNOMEDCT_CORE|Edema of optic disc|Optic disc edema
C0030353|T047|PT|423341008|SNOMEDCT_CORE|Optic disc edema|Optic disc edema
C0030353|T047|OF|423341008|SNOMEDCT_CORE|Optic disc edema|Optic disc edema
C0030353|T047|PTGB|423341008|SNOMEDCT_CORE|Optic disc oedema|Optic disc edema
C0030353|T047|SY|423341008|SNOMEDCT_CORE|Papilledema|Optic disc edema
C0030353|T047|SYGB|423341008|SNOMEDCT_CORE|Papilloedema|Optic disc edema
C0030389|T047|PT|12188008|SNOMEDCT_CORE|Parainfluenza|Parainfluenza
C0030389|T047|FN|12188008|SNOMEDCT_CORE|Parainfluenza|Parainfluenza
C0030389|T047|IS|12188008|SNOMEDCT_CORE|Parainfluenza, NOS|Parainfluenza
C0030421|T191|PT|302833002|SNOMEDCT_CORE|Paraganglioma|Paraganglioma
C0030421|T191|FN|302833002|SNOMEDCT_CORE|Paraganglioma|Paraganglioma
C0030446|T047|SY|55525008|SNOMEDCT_CORE|Adynamic ileus|Paralytic ileus
C0030446|T047|SY|55525008|SNOMEDCT_CORE|Paralysis of intestine|Paralytic ileus
C0030446|T047|PT|55525008|SNOMEDCT_CORE|Paralytic ileus|Paralytic ileus
C0030446|T047|FN|55525008|SNOMEDCT_CORE|Paralytic ileus|Paralytic ileus
C0030483|T047|PT|13758004|SNOMEDCT_CORE|Paraphimosis|Paraphimosis
C0030483|T047|FN|13758004|SNOMEDCT_CORE|Paraphimosis|Paraphimosis
C0030486|T047|SY|60389000|SNOMEDCT_CORE|Lower paraplegia|Paraplegia
C0030486|T047|SY|60389000|SNOMEDCT_CORE|Paralysis of both lower limbs|Paraplegia
C0030486|T047|PT|60389000|SNOMEDCT_CORE|Paraplegia|Paraplegia
C0030486|T047|FN|60389000|SNOMEDCT_CORE|Paraplegia|Paraplegia
C0030508|T047|PT|58690002|SNOMEDCT_CORE|Parasomnia|Parasomnia
C0030508|T047|SY|58690002|SNOMEDCT_CORE|Parasomnia|Parasomnia
C0030508|T047|FN|58690002|SNOMEDCT_CORE|Parasomnia|Parasomnia
C0030508|T047|IS|58690002|SNOMEDCT_CORE|Parasomnia, NOS|Parasomnia
C0030540|T033|PT|52184009|SNOMEDCT_CORE|Parent-child problem|Parent-child problem
C0030540|T033|FN|52184009|SNOMEDCT_CORE|Parent-child problem|Parent-child problem
C0030552|T047|IS|26544005|SNOMEDCT_CORE|Incomplete paralysis|Paresis
C0030552|T047|IS|26544005|SNOMEDCT_CORE|Paresis|Paresis
C0030552|T047|IS|26544005|SNOMEDCT_CORE|Paresis, NOS|Paresis
C0030554|T047|PTGB|91019004|SNOMEDCT_CORE|Paraesthesia|Paresthesia
C0030554|T047|SYGB|91019004|SNOMEDCT_CORE|Paraesthesia|Paresthesia
C0030554|T047|PT|91019004|SNOMEDCT_CORE|Paresthesia|Paresthesia
C0030554|T047|SY|91019004|SNOMEDCT_CORE|Paresthesia|Paresthesia
C0030554|T047|FN|91019004|SNOMEDCT_CORE|Paresthesia|Paresthesia
C0030567|T047|SY|49049000|SNOMEDCT_CORE|Idiopathic Parkinson's disease|Parkinson's disease
C0030567|T047|SY|49049000|SNOMEDCT_CORE|Idiopathic Parkinsonism|Parkinson's disease
C0030567|T047|IS|49049000|SNOMEDCT_CORE|Idiopathic parkinsonism|Parkinson's disease
C0030567|T047|SY|49049000|SNOMEDCT_CORE|Paralysis agitans|Parkinson's disease
C0030567|T047|SY|49049000|SNOMEDCT_CORE|Parkinson disease|Parkinson's disease
C0030567|T047|PT|49049000|SNOMEDCT_CORE|Parkinson's disease|Parkinson's disease
C0030567|T047|FN|49049000|SNOMEDCT_CORE|Parkinson's disease|Parkinson's disease
C0030567|T047|IS|49049000|SNOMEDCT_CORE|Parkinson's disease, NOS|Parkinson's disease
C0030567|T047|SY|49049000|SNOMEDCT_CORE|Parkinsons disease|Parkinson's disease
C0030567|T047|SY|49049000|SNOMEDCT_CORE|PD - Parkinson's disease|Parkinson's disease
C0030567|T047|SY|49049000|SNOMEDCT_CORE|Primary Parkinsonism|Parkinson's disease
C0030567|T047|IS|49049000|SNOMEDCT_CORE|Primary parkinsonism|Parkinson's disease
C0030567|T047|SY|49049000|SNOMEDCT_CORE|Shaking palsy|Parkinson's disease
C0030569|T047|SY|32798002|SNOMEDCT_CORE|Disorders presenting primarily with parkinsonism|Secondary parkinsonism
C0030569|T047|SY|230292008|SNOMEDCT_CORE|Secondary Parkinson disease|Secondary parkinsonism
C0030569|T047|SY|230292008|SNOMEDCT_CORE|Secondary Parkinson's disease|Secondary parkinsonism
C0030569|T047|PT|230292008|SNOMEDCT_CORE|Secondary parkinsonism|Secondary parkinsonism
C0030569|T047|FN|230292008|SNOMEDCT_CORE|Secondary parkinsonism|Secondary parkinsonism
C0030578|T047|PT|71906005|SNOMEDCT_CORE|Paronychia|Paronychia
C0030578|T047|FN|71906005|SNOMEDCT_CORE|Paronychia|Paronychia
C0030578|T047|SY|71906005|SNOMEDCT_CORE|Perionychia|Paronychia
C0030581|T191|PT|126788000|SNOMEDCT_CORE|Neoplasm of parotid gland|Neoplasm of parotid gland
C0030581|T191|FN|126788000|SNOMEDCT_CORE|Neoplasm of parotid gland|Neoplasm of parotid gland
C0030581|T191|SY|126788000|SNOMEDCT_CORE|Tumor of parotid gland|Neoplasm of parotid gland
C0030581|T191|SYGB|126788000|SNOMEDCT_CORE|Tumour of parotid gland|Neoplasm of parotid gland
C0030584|T047|SY|64233004|SNOMEDCT_CORE|Congenital cyst of fimbria of fallopian tube|Embryonic fimbrial cyst
C0030584|T047|FN|64233004|SNOMEDCT_CORE|Embryonic cyst of fimbria of fallopian tube|Embryonic fimbrial cyst
C0030584|T047|SY|64233004|SNOMEDCT_CORE|Embryonic cyst of fimbria of fallopian tube|Embryonic fimbrial cyst
C0030584|T047|PT|64233004|SNOMEDCT_CORE|Embryonic fimbrial cyst|Embryonic fimbrial cyst
C0030584|T047|OF|64233004|SNOMEDCT_CORE|Embryonic fimbrial cyst|Embryonic fimbrial cyst
C0030584|T047|IS|64233004|SNOMEDCT_CORE|Fimbrial cyst|Embryonic fimbrial cyst
C0030584|T047|IS|64233004|SNOMEDCT_CORE|Parovarian cyst|Embryonic fimbrial cyst
C0030587|T033|PT|195069001|SNOMEDCT_CORE|Atrial paroxysmal tachycardia|Atrial paroxysmal tachycardia
C0030587|T033|SY|195069001|SNOMEDCT_CORE|Paroxysmal atrial tachycardia|Atrial paroxysmal tachycardia
C0030587|T033|FN|195069001|SNOMEDCT_CORE|Paroxysmal atrial tachycardia|Atrial paroxysmal tachycardia
C0030587|T033|SY|195069001|SNOMEDCT_CORE|PAT|Atrial paroxysmal tachycardia
C0030587|T033|SY|195069001|SNOMEDCT_CORE|PAT - Paroxysmal atrial tachycardia|Atrial paroxysmal tachycardia
C0030590|T047|PT|67198005|SNOMEDCT_CORE|Paroxysmal supraventricular tachycardia|Paroxysmal supraventricular tachycardia
C0030590|T047|FN|67198005|SNOMEDCT_CORE|Paroxysmal supraventricular tachycardia|Paroxysmal supraventricular tachycardia
C0030591|T047|PT|66657009|SNOMEDCT_CORE|Paroxysmal ventricular tachycardia|Paroxysmal ventricular tachycardia
C0030591|T047|FN|66657009|SNOMEDCT_CORE|Paroxysmal ventricular tachycardia|Paroxysmal ventricular tachycardia
C0030593|T047|PT|45688009|SNOMEDCT_CORE|Pars planitis|Pars planitis
C0030593|T047|FN|45688009|SNOMEDCT_CORE|Pars planitis|Pars planitis
C0030593|T047|IS|45688009|SNOMEDCT_CORE|Posterior cyclitis|Pars planitis
C0030662|T048|PT|18085000|SNOMEDCT_CORE|Compulsive gambling|Compulsive gambling
C0030662|T048|FN|18085000|SNOMEDCT_CORE|Compulsive gambling|Compulsive gambling
C0030662|T048|SY|18085000|SNOMEDCT_CORE|Gambling disorder|Compulsive gambling
C0030662|T048|IS|18085000|SNOMEDCT_CORE|Pathological gambling|Compulsive gambling
C0030662|T048|SY|18085000|SNOMEDCT_CORE|Pathological gambling disorder|Compulsive gambling
C0030756|T047|PT|20848007|SNOMEDCT_CORE|Infestation by Pediculus|Infestation by Pediculus
C0030756|T047|OF|20848007|SNOMEDCT_CORE|Infestation by Pediculus|Infestation by Pediculus
C0030756|T047|IS|20848007|SNOMEDCT_CORE|Infestation by Pediculus, NOS|Infestation by Pediculus
C0030756|T047|FN|20848007|SNOMEDCT_CORE|Infestation caused by Pediculus|Infestation by Pediculus
C0030756|T047|SY|20848007|SNOMEDCT_CORE|Infestation caused by Pediculus|Infestation by Pediculus
C0030756|T047|IS|74949007|SNOMEDCT_CORE|Lice infestation|Infestation by Pediculus
C0030756|T047|IS|74949007|SNOMEDCT_CORE|Lice infestation, NOS|Infestation by Pediculus
C0030756|T047|IS|20848007|SNOMEDCT_CORE|Louse infestation|Infestation by Pediculus
C0030756|T047|SY|20848007|SNOMEDCT_CORE|Pediculosis|Infestation by Pediculus
C0030757|T047|SY|81000006|SNOMEDCT_CORE|Head lice|Pediculosis capitis
C0030757|T047|SY|81000006|SNOMEDCT_CORE|Head lice infestation|Pediculosis capitis
C0030757|T047|SY|81000006|SNOMEDCT_CORE|Head louse infestation|Pediculosis capitis
C0030757|T047|SY|81000006|SNOMEDCT_CORE|Lice infested hair|Pediculosis capitis
C0030757|T047|SY|81000006|SNOMEDCT_CORE|Lousy hair|Pediculosis capitis
C0030757|T047|SY|81000006|SNOMEDCT_CORE|Nit infested hair|Pediculosis capitis
C0030757|T047|SY|81000006|SNOMEDCT_CORE|Nits|Pediculosis capitis
C0030757|T047|PT|81000006|SNOMEDCT_CORE|Pediculosis capitis|Pediculosis capitis
C0030757|T047|FN|81000006|SNOMEDCT_CORE|Pediculosis capitis|Pediculosis capitis
C0030757|T047|SY|81000006|SNOMEDCT_CORE|Pediculus capitis infestation|Pediculosis capitis
C0030793|T191|PT|126644004|SNOMEDCT_CORE|Neoplasm of pelvis|Neoplasm of pelvis
C0030793|T191|FN|126644004|SNOMEDCT_CORE|Neoplasm of pelvis|Neoplasm of pelvis
C0030793|T191|SY|126644004|SNOMEDCT_CORE|Tumor of pelvis|Neoplasm of pelvis
C0030793|T191|SYGB|126644004|SNOMEDCT_CORE|Tumour of pelvis|Neoplasm of pelvis
C0030794|T184|PT|30473006|SNOMEDCT_CORE|Pain in pelvis|Pain in pelvis
C0030794|T184|FN|30473006|SNOMEDCT_CORE|Pain in pelvis|Pain in pelvis
C0030794|T184|IS|30473006|SNOMEDCT_CORE|Pelvic pain|Pain in pelvis
C0030794|T184|IS|30473006|SNOMEDCT_CORE|Pelvic pain, NOS|Pain in pelvis
C0030795|T190|OAS|11374003|SNOMEDCT_CORE|Relaxation of pelvis|Relaxation of pelvis
C0030804|T047|SY|34250006|SNOMEDCT_CORE|Benign mucosal pemphigoid|Benign mucous membrane pemphigoid
C0030804|T047|PT|34250006|SNOMEDCT_CORE|Benign mucous membrane pemphigoid|Benign mucous membrane pemphigoid
C0030804|T047|FN|34250006|SNOMEDCT_CORE|Benign mucous membrane pemphigoid|Benign mucous membrane pemphigoid
C0030804|T047|SY|34250006|SNOMEDCT_CORE|Cicatricial pemphigoid|Benign mucous membrane pemphigoid
C0030804|T047|SY|34250006|SNOMEDCT_CORE|Mucosynechia atrophic bullous dermatitis|Benign mucous membrane pemphigoid
C0030804|T047|SY|34250006|SNOMEDCT_CORE|Mucous membrane pemphigoid|Benign mucous membrane pemphigoid
C0030804|T047|SY|34250006|SNOMEDCT_CORE|Scarring pemphigoid|Benign mucous membrane pemphigoid
C0030805|T047|SY|77090002|SNOMEDCT_CORE|BP - Bullous pemphigoid|Bullous pemphigoid
C0030805|T047|PT|77090002|SNOMEDCT_CORE|Bullous pemphigoid|Bullous pemphigoid
C0030805|T047|FN|77090002|SNOMEDCT_CORE|Bullous pemphigoid|Bullous pemphigoid
C0030824|T047|PT|91936005|SNOMEDCT_CORE|Allergy to penicillin|Allergy to penicillin
C0030824|T047|FN|91936005|SNOMEDCT_CORE|Allergy to penicillin|Allergy to penicillin
C0030824|T047|OF|91936005|SNOMEDCT_CORE|Allergy to penicillin|Allergy to penicillin
C0030824|T047|SY|91936005|SNOMEDCT_CORE|Penicillin allergy|Allergy to penicillin
C0030848|T047|SY|1335005|SNOMEDCT_CORE|Fibrous cavernositis|Induratio penis plastica
C0030848|T047|PT|1335005|SNOMEDCT_CORE|Induratio penis plastica|Induratio penis plastica
C0030848|T047|FN|1335005|SNOMEDCT_CORE|Induratio penis plastica|Induratio penis plastica
C0030848|T047|SY|1335005|SNOMEDCT_CORE|Penile fibromatosis|Induratio penis plastica
C0030848|T047|SY|1335005|SNOMEDCT_CORE|Peyronie's disease|Induratio penis plastica
C0030848|T047|SY|1335005|SNOMEDCT_CORE|Peyronies disease|Induratio penis plastica
C0030848|T047|SY|1335005|SNOMEDCT_CORE|Plastic induration of penis|Induratio penis plastica
C0030920|T047|SY|13200003|SNOMEDCT_CORE|Gastroduodenal ulcer|Peptic ulcer
C0030920|T047|IS|13200003|SNOMEDCT_CORE|Gastroduodenal ulcer, NOS|Peptic ulcer
C0030920|T047|PT|13200003|SNOMEDCT_CORE|Peptic ulcer|Peptic ulcer
C0030920|T047|FN|13200003|SNOMEDCT_CORE|Peptic ulcer|Peptic ulcer
C0030920|T047|SY|13200003|SNOMEDCT_CORE|Peptic ulcer disease|Peptic ulcer
C0030920|T047|IS|13200003|SNOMEDCT_CORE|Peptic ulcer, NOS|Peptic ulcer
C0030920|T047|SY|13200003|SNOMEDCT_CORE|Peptic ulceration|Peptic ulcer
C0030920|T047|SY|13200003|SNOMEDCT_CORE|PU - Peptic ulcer|Peptic ulcer
C0030920|T047|SY|13200003|SNOMEDCT_CORE|PUD - Peptic ulcer disease|Peptic ulcer
C0030922|T046|SY|64121000|SNOMEDCT_CORE|Bleeding peptic ulcer|Peptic ulcer with hemorrhage
C0030922|T046|PTGB|64121000|SNOMEDCT_CORE|Peptic ulcer with haemorrhage|Peptic ulcer with hemorrhage
C0030922|T046|PT|64121000|SNOMEDCT_CORE|Peptic ulcer with hemorrhage|Peptic ulcer with hemorrhage
C0030922|T046|FN|64121000|SNOMEDCT_CORE|Peptic ulcer with hemorrhage|Peptic ulcer with hemorrhage
C0030922|T046|IS|64121000|SNOMEDCT_CORE|Peptic ulcer, NOS with hemorrhage|Peptic ulcer with hemorrhage
C0031019|T047|PT|82127005|SNOMEDCT_CORE|Perianal abscess|Perianal abscess
C0031019|T047|FN|82127005|SNOMEDCT_CORE|Perianal abscess|Perianal abscess
C0031022|T047|IS|49120005|SNOMEDCT_CORE|Chronic peri-aortitis|Chronic peri-aortitis
C0031024|T047|SY|196341005|SNOMEDCT_CORE|Apical abscess|Periapical abscess
C0031024|T047|SY|196341005|SNOMEDCT_CORE|Dentoalveolar abscess|Periapical abscess
C0031024|T047|PT|196341005|SNOMEDCT_CORE|Periapical abscess|Periapical abscess
C0031024|T047|FN|196341005|SNOMEDCT_CORE|Periapical abscess|Periapical abscess
C0031036|T047|SY|155441006|SNOMEDCT_CORE|PAN - Polyarteritis nodosa|Polyarteritis nodosa
C0031036|T047|SY|155441006|SNOMEDCT_CORE|Periarteritis nodosa|Polyarteritis nodosa
C0031036|T047|OF|155441006|SNOMEDCT_CORE|Polyarteritis nodosa|Polyarteritis nodosa
C0031036|T047|PT|155441006|SNOMEDCT_CORE|Polyarteritis nodosa|Polyarteritis nodosa
C0031036|T047|FN|155441006|SNOMEDCT_CORE|Polyarteritis nodosa|Polyarteritis nodosa
C0031039|T047|PT|373945007|SNOMEDCT_CORE|Pericardial effusion|Pericardial effusion
C0031039|T047|FN|373945007|SNOMEDCT_CORE|Pericardial effusion|Pericardial effusion
C0031046|T047|PT|3238004|SNOMEDCT_CORE|Pericarditis|Pericarditis
C0031046|T047|FN|3238004|SNOMEDCT_CORE|Pericarditis|Pericarditis
C0031046|T047|IS|3238004|SNOMEDCT_CORE|Pericarditis, NOS|Pericarditis
C0031048|T047|PT|85598007|SNOMEDCT_CORE|Constrictive pericarditis|Constrictive pericarditis
C0031048|T047|FN|85598007|SNOMEDCT_CORE|Constrictive pericarditis|Constrictive pericarditis
C0031055|T047|PT|22240003|SNOMEDCT_CORE|Pericoronitis|Pericoronitis
C0031055|T047|FN|22240003|SNOMEDCT_CORE|Pericoronitis|Pericoronitis
C0031090|T047|SY|2556008|SNOMEDCT_CORE|Disease of supporting structures of teeth|Periodontal disease
C0031090|T047|PT|2556008|SNOMEDCT_CORE|Periodontal disease|Periodontal disease
C0031090|T047|FN|2556008|SNOMEDCT_CORE|Periodontal disease|Periodontal disease
C0031090|T047|IS|2556008|SNOMEDCT_CORE|Periodontal disease, NOS|Periodontal disease
C0031099|T047|PT|41565005|SNOMEDCT_CORE|Periodontitis|Periodontitis
C0031099|T047|FN|41565005|SNOMEDCT_CORE|Periodontitis|Periodontitis
C0031099|T047|IS|41565005|SNOMEDCT_CORE|Periodontitis, NOS|Periodontitis
C0031121|T047|PT|25416002|SNOMEDCT_CORE|Peripheral neuralgia|Peripheral neuralgia
C0031121|T047|FN|25416002|SNOMEDCT_CORE|Peripheral neuralgia|Peripheral neuralgia
C0031121|T047|OF|25416002|SNOMEDCT_CORE|Peripheral neuralgia|Peripheral neuralgia
C0031144|T047|FN|78609007|SNOMEDCT_CORE|Chronic peritoneal effusion|Chronic peritoneal effusion
C0031144|T047|PT|78609007|SNOMEDCT_CORE|Chronic peritoneal effusion|Chronic peritoneal effusion
C0031154|T046|PT|48661000|SNOMEDCT_CORE|Peritonitis|Peritonitis
C0031154|T046|FN|48661000|SNOMEDCT_CORE|Peritonitis|Peritonitis
C0031154|T046|IS|48661000|SNOMEDCT_CORE|Peritonitis of undetermined cause|Peritonitis
C0031154|T046|IS|48661000|SNOMEDCT_CORE|Peritonitis, NOS|Peritonitis
C0031157|T047|SY|15033003|SNOMEDCT_CORE|Angina tonsillaris|Peritonsillar abscess
C0031157|T047|PT|15033003|SNOMEDCT_CORE|Peritonsillar abscess|Peritonsillar abscess
C0031157|T047|FN|15033003|SNOMEDCT_CORE|Peritonsillar abscess|Peritonsillar abscess
C0031157|T047|SY|15033003|SNOMEDCT_CORE|Quinsy|Peritonsillar abscess
C0031190|T047|PT|233815004|SNOMEDCT_CORE|Persistent pulmonary hypertension of the newborn|Persistent pulmonary hypertension of the newborn
C0031190|T047|FN|233815004|SNOMEDCT_CORE|Persistent pulmonary hypertension of the newborn|Persistent pulmonary hypertension of the newborn
C0031190|T047|SY|233815004|SNOMEDCT_CORE|PFC - Persistent fetal circulation|Persistent pulmonary hypertension of the newborn
C0031190|T047|SY|233815004|SNOMEDCT_CORE|PFC - Persistent foetal circulation|Persistent pulmonary hypertension of the newborn
C0031190|T047|SY|233815004|SNOMEDCT_CORE|PPHN - Persistent pulmonary hypertension in newborn|Persistent pulmonary hypertension of the newborn
C0031212|T048|PT|33449004|SNOMEDCT_CORE|Personality disorder|Personality disorder
C0031212|T048|FN|33449004|SNOMEDCT_CORE|Personality disorder|Personality disorder
C0031212|T048|IS|33449004|SNOMEDCT_CORE|Personality disorder, NOS|Personality disorder
C0031256|T047|PT|271813007|SNOMEDCT_CORE|Petechiae|Petechiae
C0031256|T047|OF|271813007|SNOMEDCT_CORE|Petechiae|Petechiae
C0031256|T047|FN|271813007|SNOMEDCT_CORE|Petechiae|Petechiae
C0031256|T047|IS|271813007|SNOMEDCT_CORE|Petechial eruption|Petechiae
C0031256|T047|IS|271813007|SNOMEDCT_CORE|Petechial rash|Petechiae
C0031315|T047|SY|193114000|SNOMEDCT_CORE|FLS - Phantom limb syndrome|Phantom limb
C0031315|T047|PT|193114000|SNOMEDCT_CORE|Phantom limb|Phantom limb
C0031315|T047|FN|193114000|SNOMEDCT_CORE|Phantom limb|Phantom limb
C0031315|T047|SY|193114000|SNOMEDCT_CORE|Phantom limb syndrome|Phantom limb
C0031315|T047|SY|193114000|SNOMEDCT_CORE|PLS - Phantom limb syndrome|Phantom limb
C0031350|T047|PT|405737000|SNOMEDCT_CORE|Pharyngitis|Pharyngitis
C0031350|T047|FN|405737000|SNOMEDCT_CORE|Pharyngitis|Pharyngitis
C0031538|T033|PT|198006006|SNOMEDCT_CORE|Tight foreskin|Tight foreskin
C0031538|T033|FN|198006006|SNOMEDCT_CORE|Tight foreskin|Tight foreskin
C0031538|T033|SY|198006006|SNOMEDCT_CORE|Tight prepuce|Tight foreskin
C0031542|T046|SY|61599003|SNOMEDCT_CORE|Inflammation of vein|Phlebitis
C0031542|T046|IS|61599003|SNOMEDCT_CORE|Inflammation of vein, NOS|Phlebitis
C0031542|T046|PT|61599003|SNOMEDCT_CORE|Phlebitis|Phlebitis
C0031542|T046|FN|61599003|SNOMEDCT_CORE|Phlebitis|Phlebitis
C0031542|T046|IS|61599003|SNOMEDCT_CORE|Phlebitis, NOS|Phlebitis
C0031572|T048|SY|25501002|SNOMEDCT_CORE|Social anxiety disorder|Social phobia
C0031572|T048|PT|25501002|SNOMEDCT_CORE|Social phobia|Social phobia
C0031572|T048|FN|25501002|SNOMEDCT_CORE|Social phobia|Social phobia
C0031572|T048|IS|25501002|SNOMEDCT_CORE|Social phobia, NOS|Social phobia
C0031707|T047|PT|87049008|SNOMEDCT_CORE|Disorder of phosphorus metabolism|Disorder of phosphorus metabolism
C0031707|T047|FN|87049008|SNOMEDCT_CORE|Disorder of phosphorus metabolism|Disorder of phosphorus metabolism
C0031707|T047|IS|87049008|SNOMEDCT_CORE|Disorder of phosphorus metabolism, NOS|Disorder of phosphorus metabolism
C0031707|T047|SY|87049008|SNOMEDCT_CORE|Phosphorus metabolism disorder|Disorder of phosphorus metabolism
C0031736|T047|SY|238525001|SNOMEDCT_CORE|PLE - Polymorphic light eruption|Polymorphous light eruption
C0031736|T047|SY|238525001|SNOMEDCT_CORE|Polymorphic light eruption|Polymorphous light eruption
C0031736|T047|FN|238525001|SNOMEDCT_CORE|Polymorphic light eruption|Polymorphous light eruption
C0031736|T047|SY|238525001|SNOMEDCT_CORE|Polymorphic photodermatitis|Polymorphous light eruption
C0031736|T047|PT|238525001|SNOMEDCT_CORE|Polymorphous light eruption|Polymorphous light eruption
C0031876|T047|SY|85598007|SNOMEDCT_CORE|Pick disease of heart|Pick syndrome of heart
C0031876|T047|SY|85598007|SNOMEDCT_CORE|Pick syndrome of heart|Pick syndrome of heart
C0031925|T047|IS|47639008|SNOMEDCT_CORE|Coccygeal sinus|Pilonidal cyst
C0031925|T047|SY|47639008|SNOMEDCT_CORE|Cyst - pilonidal|Pilonidal cyst
C0031925|T047|OF|47639008|SNOMEDCT_CORE|Cyst - pilonidal|Pilonidal cyst
C0031925|T047|SY|47639008|SNOMEDCT_CORE|Piliferous cyst|Pilonidal cyst
C0031925|T047|PT|47639008|SNOMEDCT_CORE|Pilonidal cyst|Pilonidal cyst
C0031925|T047|FN|47639008|SNOMEDCT_CORE|Pilonidal cyst|Pilonidal cyst
C0031925|T047|IS|47639008|SNOMEDCT_CORE|Pilonidal cyst, NOS|Pilonidal cyst
C0031925|T047|IS|47639008|SNOMEDCT_CORE|Pilonidal sinus|Pilonidal cyst
C0032000|T191|SY|254956000|SNOMEDCT_CORE|Adenoma of pituitary|Pituitary adenoma
C0032000|T191|PT|254956000|SNOMEDCT_CORE|Pituitary adenoma|Pituitary adenoma
C0032000|T191|FN|254956000|SNOMEDCT_CORE|Pituitary adenoma|Pituitary adenoma
C0032002|T047|IS|399244003|SNOMEDCT_CORE|Disease of pituitary gland|Disorder of pituitary gland
C0032002|T047|OF|399244003|SNOMEDCT_CORE|Disease of pituitary gland|Disorder of pituitary gland
C0032002|T047|SY|399244003|SNOMEDCT_CORE|Disorder of pituitary|Disorder of pituitary gland
C0032002|T047|PT|399244003|SNOMEDCT_CORE|Disorder of pituitary gland|Disorder of pituitary gland
C0032002|T047|FN|399244003|SNOMEDCT_CORE|Disorder of pituitary gland|Disorder of pituitary gland
C0032002|T047|SY|399244003|SNOMEDCT_CORE|Dyspituitarism|Disorder of pituitary gland
C0032002|T047|SY|399244003|SNOMEDCT_CORE|Pituitary disease|Disorder of pituitary gland
C0032019|T191|PT|127024001|SNOMEDCT_CORE|Neoplasm of pituitary gland|Neoplasm of pituitary gland
C0032019|T191|FN|127024001|SNOMEDCT_CORE|Neoplasm of pituitary gland|Neoplasm of pituitary gland
C0032019|T191|SY|127024001|SNOMEDCT_CORE|Pituitary tumor|Neoplasm of pituitary gland
C0032019|T191|SYGB|127024001|SNOMEDCT_CORE|Pituitary tumour|Neoplasm of pituitary gland
C0032019|T191|SY|127024001|SNOMEDCT_CORE|Tumor of pituitary gland|Neoplasm of pituitary gland
C0032019|T191|SYGB|127024001|SNOMEDCT_CORE|Tumour of pituitary gland|Neoplasm of pituitary gland
C0032024|T047|PT|34630004|SNOMEDCT_CORE|Pityriasis|Pityriasis
C0032024|T047|FN|34630004|SNOMEDCT_CORE|Pityriasis|Pityriasis
C0032024|T047|IS|34630004|SNOMEDCT_CORE|Pityriasis, NOS|Pityriasis
C0032026|T047|SY|77252004|SNOMEDCT_CORE|Pityriasis circinata et maculata|Pityriasis rosea
C0032026|T047|PT|77252004|SNOMEDCT_CORE|Pityriasis rosea|Pityriasis rosea
C0032026|T047|FN|77252004|SNOMEDCT_CORE|Pityriasis rosea|Pityriasis rosea
C0032026|T047|SY|77252004|SNOMEDCT_CORE|PR - Pityriasis rosea|Pityriasis rosea
C0032046|T046|PTGB|36813001|SNOMEDCT_CORE|Placenta praevia|Placenta previa
C0032046|T046|PT|36813001|SNOMEDCT_CORE|Placenta previa|Placenta previa
C0032046|T046|FN|36813001|SNOMEDCT_CORE|Placenta previa|Placenta previa
C0032046|T046|IS|36813001|SNOMEDCT_CORE|Placenta previa, NOS|Placenta previa
C0032046|T046|SYGB|36813001|SNOMEDCT_CORE|PP - Placenta praevia|Placenta previa
C0032046|T046|SY|36813001|SNOMEDCT_CORE|PP - Placenta previa|Placenta previa
C0032131|T191|PT|415112005|SNOMEDCT_CORE|Plasmacytoma|Plasmacytoma
C0032131|T191|FN|415112005|SNOMEDCT_CORE|Plasmacytoma|Plasmacytoma
C0032131|T191|SY|415112005|SNOMEDCT_CORE|Plasmacytoma - disorder|Plasmacytoma
C0032227|T047|FN|60046008|SNOMEDCT_CORE|Pleural effusion|Pleural effusion
C0032227|T047|PT|60046008|SNOMEDCT_CORE|Pleural effusion|Pleural effusion
C0032227|T047|IS|60046008|SNOMEDCT_CORE|Pleural effusion, NOS|Pleural effusion
C0032231|T047|PT|196075003|SNOMEDCT_CORE|Pleurisy|Pleurisy
C0032231|T047|FN|196075003|SNOMEDCT_CORE|Pleurisy|Pleurisy
C0032231|T047|SY|196075003|SNOMEDCT_CORE|Pleuritis|Pleurisy
C0032269|T047|SY|16814004|SNOMEDCT_CORE|Pneumococcal disease|Pneumococcal infectious disease
C0032269|T047|SY|16814004|SNOMEDCT_CORE|Pneumococcal infection|Pneumococcal infectious disease
C0032269|T047|IS|16814004|SNOMEDCT_CORE|Pneumococcal infection, NOS|Pneumococcal infectious disease
C0032269|T047|PT|16814004|SNOMEDCT_CORE|Pneumococcal infectious disease|Pneumococcal infectious disease
C0032269|T047|FN|16814004|SNOMEDCT_CORE|Pneumococcal infectious disease|Pneumococcal infectious disease
C0032269|T047|IS|16814004|SNOMEDCT_CORE|Pneumococcal infectious disease, NOS|Pneumococcal infectious disease
C0032273|T047|SY|40122008|SNOMEDCT_CORE|PK - Pneumoconiosis|Pneumoconiosis
C0032273|T047|PT|40122008|SNOMEDCT_CORE|Pneumoconiosis|Pneumoconiosis
C0032273|T047|FN|40122008|SNOMEDCT_CORE|Pneumoconiosis|Pneumoconiosis
C0032273|T047|IS|40122008|SNOMEDCT_CORE|Pneumoconiosis, NOS|Pneumoconiosis
C0032285|T047|PT|233604007|SNOMEDCT_CORE|Pneumonia|Pneumonia
C0032285|T047|FN|233604007|SNOMEDCT_CORE|Pneumonia|Pneumonia
C0032290|T047|PT|422588002|SNOMEDCT_CORE|Aspiration pneumonia|Aspiration pneumonia
C0032290|T047|FN|422588002|SNOMEDCT_CORE|Aspiration pneumonia|Aspiration pneumonia
C0032290|T047|SY|422588002|SNOMEDCT_CORE|Inhalation pneumonia|Aspiration pneumonia
C0032300|T047|PT|278516003|SNOMEDCT_CORE|Lobar pneumonia|Lobar pneumonia
C0032300|T047|FN|278516003|SNOMEDCT_CORE|Lobar pneumonia|Lobar pneumonia
C0032302|T047|SY|46970008|SNOMEDCT_CORE|Eaton's agent pneumonia|Mycoplasma pneumonia
C0032302|T047|IS|46970008|SNOMEDCT_CORE|Eatons agent pneumonia|Mycoplasma pneumonia
C0032302|T047|SY|46970008|SNOMEDCT_CORE|Endemic pneumonia|Mycoplasma pneumonia
C0032302|T047|SY|46970008|SNOMEDCT_CORE|Infection by PPLO|Mycoplasma pneumonia
C0032302|T047|PT|46970008|SNOMEDCT_CORE|Mycoplasma pneumonia|Mycoplasma pneumonia
C0032302|T047|OF|46970008|SNOMEDCT_CORE|Mycoplasma pneumonia|Mycoplasma pneumonia
C0032302|T047|SY|46970008|SNOMEDCT_CORE|Mycoplasma pneumoniae pneumonia|Mycoplasma pneumonia
C0032302|T047|SY|46970008|SNOMEDCT_CORE|Mycoplasmal pneumonia|Mycoplasma pneumonia
C0032302|T047|SY|46970008|SNOMEDCT_CORE|PAP caused by Mycoplasma pneumoniae|Mycoplasma pneumonia
C0032302|T047|SY|46970008|SNOMEDCT_CORE|PAP due to Mycoplasma pneumoniae|Mycoplasma pneumonia
C0032302|T047|FN|46970008|SNOMEDCT_CORE|Pneumonia caused by Mycoplasma pneumoniae|Mycoplasma pneumonia
C0032302|T047|SY|46970008|SNOMEDCT_CORE|Pneumonia caused by Mycoplasma pneumoniae|Mycoplasma pneumonia
C0032302|T047|SY|46970008|SNOMEDCT_CORE|Pneumonia caused by PPLO|Mycoplasma pneumonia
C0032302|T047|SY|46970008|SNOMEDCT_CORE|Pneumonia due to Mycoplasma pneumoniae|Mycoplasma pneumonia
C0032302|T047|OF|46970008|SNOMEDCT_CORE|Pneumonia due to Mycoplasma pneumoniae|Mycoplasma pneumonia
C0032302|T047|SY|46970008|SNOMEDCT_CORE|Pneumonia due to PPLO|Mycoplasma pneumonia
C0032302|T047|SY|46970008|SNOMEDCT_CORE|Primary atypical pneumonia caused by Mycoplasma pneumoniae|Mycoplasma pneumonia
C0032302|T047|SY|46970008|SNOMEDCT_CORE|Primary atypical pneumonia due to Mycoplasma pneumoniae|Mycoplasma pneumonia
C0032308|T047|PT|22754005|SNOMEDCT_CORE|Staphylococcal pneumonia|Staphylococcal pneumonia
C0032308|T047|FN|22754005|SNOMEDCT_CORE|Staphylococcal pneumonia|Staphylococcal pneumonia
C0032310|T047|PT|75570004|SNOMEDCT_CORE|Viral pneumonia|Viral pneumonia
C0032310|T047|FN|75570004|SNOMEDCT_CORE|Viral pneumonia|Viral pneumonia
C0032310|T047|IS|75570004|SNOMEDCT_CORE|Viral pneumonia, NOS|Viral pneumonia
C0032326|T047|PT|36118008|SNOMEDCT_CORE|Pneumothorax|Pneumothorax
C0032326|T047|FN|36118008|SNOMEDCT_CORE|Pneumothorax|Pneumothorax
C0032326|T047|IS|36118008|SNOMEDCT_CORE|Pneumothorax, NOS|Pneumothorax
C0032371|T047|PT|398102009|SNOMEDCT_CORE|Acute poliomyelitis|Acute poliomyelitis
C0032371|T047|FN|398102009|SNOMEDCT_CORE|Acute poliomyelitis|Acute poliomyelitis
C0032371|T047|SY|398102009|SNOMEDCT_CORE|PM - Poliomyelitis|Acute poliomyelitis
C0032371|T047|SY|398102009|SNOMEDCT_CORE|Polio|Acute poliomyelitis
C0032371|T047|SY|398102009|SNOMEDCT_CORE|Poliomyelitis|Acute poliomyelitis
C0032453|T047|SY|72275000|SNOMEDCT_CORE|Chronic polychondritis|Relapsing polychondritis
C0032453|T047|SY|72275000|SNOMEDCT_CORE|Meyenburg's disease|Relapsing polychondritis
C0032453|T047|PT|72275000|SNOMEDCT_CORE|Relapsing polychondritis|Relapsing polychondritis
C0032453|T047|FN|72275000|SNOMEDCT_CORE|Relapsing polychondritis|Relapsing polychondritis
C0032453|T047|SY|72275000|SNOMEDCT_CORE|Systemic chondromalacia|Relapsing polychondritis
C0032460|T047|OAS|69878008|SNOMEDCT_CORE|Cystic disease of ovaries|Polycystic ovary
C0032460|T047|OAS|69878008|SNOMEDCT_CORE|Multicystic ovaries|Polycystic ovary
C0032460|T047|OAS|69878008|SNOMEDCT_CORE|PCO - Polycystic ovaries|Polycystic ovary
C0032460|T047|OAS|69878008|SNOMEDCT_CORE|PCOD - Polycystic ovarian disease|Polycystic ovary
C0032460|T047|OAS|69878008|SNOMEDCT_CORE|PCOS - Polycystic ovarian syndrome|Polycystic ovary
C0032460|T047|SY|237055002|SNOMEDCT_CORE|PCOS- polycystic ovary syndrome|Polycystic ovary
C0032460|T047|OAS|69878008|SNOMEDCT_CORE|Polycystic ovarian disease|Polycystic ovary
C0032460|T047|OAS|69878008|SNOMEDCT_CORE|Polycystic ovarian syndrome|Polycystic ovary
C0032460|T047|OAP|69878008|SNOMEDCT_CORE|Polycystic ovaries|Polycystic ovary
C0032460|T047|OAF|69878008|SNOMEDCT_CORE|Polycystic ovaries|Polycystic ovary
C0032460|T047|PT|781067001|SNOMEDCT_CORE|Polycystic ovary|Polycystic ovary
C0032460|T047|FN|781067001|SNOMEDCT_CORE|Polycystic ovary|Polycystic ovary
C0032460|T047|OAS|69878008|SNOMEDCT_CORE|Polycystic ovary syndrome|Polycystic ovary
C0032460|T047|OF|237055002|SNOMEDCT_CORE|Polycystic ovary syndrome|Polycystic ovary
C0032460|T047|PT|237055002|SNOMEDCT_CORE|Polycystic ovary syndrome|Polycystic ovary
C0032460|T047|FN|237055002|SNOMEDCT_CORE|Polycystic ovary syndrome|Polycystic ovary
C0032460|T047|OAS|69878008|SNOMEDCT_CORE|Sclerocystic ovary syndrome|Polycystic ovary
C0032460|T047|OAS|69878008|SNOMEDCT_CORE|Stein-Leventhal syndrome|Polycystic ovary
C0032461|T047|SYGB|109992005|SNOMEDCT_CORE|Erythrocythaemia|Polycythemia
C0032461|T047|SY|109992005|SNOMEDCT_CORE|Erythrocythemia|Polycythemia
C0032461|T047|SYGB|127062003|SNOMEDCT_CORE|Polycythaemia|Polycythemia
C0032461|T047|IS|44865000|SNOMEDCT_CORE|Polycythaemia, NOS|Polycythemia
C0032461|T047|SY|127062003|SNOMEDCT_CORE|Polycythemia|Polycythemia
C0032461|T047|IS|44865000|SNOMEDCT_CORE|Polycythemia, NOS|Polycythemia
C0032463|T191|SY|109992005|SNOMEDCT_CORE|Osler-Vaquez syndrome|Polycythemia vera
C0032463|T191|SY|109992005|SNOMEDCT_CORE|Osler's disease|Polycythemia vera
C0032463|T191|SYGB|109992005|SNOMEDCT_CORE|Polycythaemia rubra vera|Polycythemia vera
C0032463|T191|SYGB|109992005|SNOMEDCT_CORE|Polycythaemia vera|Polycythemia vera
C0032463|T191|PTGB|109992005|SNOMEDCT_CORE|Polycythaemia vera|Polycythemia vera
C0032463|T191|SY|109992005|SNOMEDCT_CORE|Polycythemia rubra vera|Polycythemia vera
C0032463|T191|SY|109992005|SNOMEDCT_CORE|Polycythemia vera|Polycythemia vera
C0032463|T191|PT|109992005|SNOMEDCT_CORE|Polycythemia vera|Polycythemia vera
C0032463|T191|FN|109992005|SNOMEDCT_CORE|Polycythemia vera|Polycythemia vera
C0032463|T191|SYGB|109992005|SNOMEDCT_CORE|PPP - Primary proliferative polycythaemia|Polycythemia vera
C0032463|T191|SY|109992005|SNOMEDCT_CORE|PPP - Primary proliferative polycythemia|Polycythemia vera
C0032463|T191|SYGB|109992005|SNOMEDCT_CORE|Primary polycythaemia|Polycythemia vera
C0032463|T191|SYGB|109992005|SNOMEDCT_CORE|Primary proliferative polycythaemia|Polycythemia vera
C0032463|T191|SY|109992005|SNOMEDCT_CORE|Primary proliferative polycythemia|Polycythemia vera
C0032463|T191|SYGB|109992005|SNOMEDCT_CORE|PRV - Polycythaemia rubra vera|Polycythemia vera
C0032463|T191|SY|109992005|SNOMEDCT_CORE|PRV - Polycythemia rubra vera|Polycythemia vera
C0032463|T191|SY|109992005|SNOMEDCT_CORE|Vaquez's disease|Polycythemia vera
C0032533|T047|SY|65323003|SNOMEDCT_CORE|Forestier-Certonciny syndrome|Polymyalgia rheumatica
C0032533|T047|SY|65323003|SNOMEDCT_CORE|PMR - Polymyalgia rheumatica|Polymyalgia rheumatica
C0032533|T047|PT|65323003|SNOMEDCT_CORE|Polymyalgia rheumatica|Polymyalgia rheumatica
C0032533|T047|FN|65323003|SNOMEDCT_CORE|Polymyalgia rheumatica|Polymyalgia rheumatica
C0032533|T047|SY|65323003|SNOMEDCT_CORE|Senile arthritis|Polymyalgia rheumatica
C0032580|T191|SY|72900001|SNOMEDCT_CORE|Adenomatous polyposis|Familial multiple polyposis syndrome
C0032580|T191|SY|72900001|SNOMEDCT_CORE|Adenomatous polyposis coli|Familial multiple polyposis syndrome
C0032580|T191|SY|72900001|SNOMEDCT_CORE|APC - Adenomatous polyposis coli|Familial multiple polyposis syndrome
C0032580|T191|SY|72900001|SNOMEDCT_CORE|Familial adenomatous polyposis|Familial multiple polyposis syndrome
C0032580|T191|PT|72900001|SNOMEDCT_CORE|Familial multiple polyposis syndrome|Familial multiple polyposis syndrome
C0032580|T191|FN|72900001|SNOMEDCT_CORE|Familial multiple polyposis syndrome|Familial multiple polyposis syndrome
C0032580|T191|SY|72900001|SNOMEDCT_CORE|Familial polyposis coli|Familial multiple polyposis syndrome
C0032580|T191|SY|72900001|SNOMEDCT_CORE|FAP - Familial adenomatous polyposis|Familial multiple polyposis syndrome
C0032580|T191|SY|72900001|SNOMEDCT_CORE|FPC - Familial polyposis coli|Familial multiple polyposis syndrome
C0032580|T191|SY|72900001|SNOMEDCT_CORE|Polyposis coli|Familial multiple polyposis syndrome
C0032584|T190|PT|441456002|SNOMEDCT_CORE|Polyp|Polyp
C0032584|T190|FN|441456002|SNOMEDCT_CORE|Polyp|Polyp
C0032586|T047|PT|75572007|SNOMEDCT_CORE|Polyradiculopathy|Polyradiculopathy
C0032586|T047|FN|75572007|SNOMEDCT_CORE|Polyradiculopathy|Polyradiculopathy
C0032587|T047|PT|128078004|SNOMEDCT_CORE|Polyradiculoneuropathy|Polyradiculoneuropathy
C0032587|T047|FN|128078004|SNOMEDCT_CORE|Polyradiculoneuropathy|Polyradiculoneuropathy
C0032606|T048|PT|51339003|SNOMEDCT_CORE|Polysubstance dependence|Polysubstance dependence
C0032606|T048|FN|51339003|SNOMEDCT_CORE|Polysubstance dependence|Polysubstance dependence
C0032617|T184|IS|28442001|SNOMEDCT_CORE|Increased urine volume|Polyuria
C0032617|T184|SY|28442001|SNOMEDCT_CORE|Passes too much urine|Polyuria
C0032617|T184|PT|28442001|SNOMEDCT_CORE|Polyuria|Polyuria
C0032617|T184|FN|28442001|SNOMEDCT_CORE|Polyuria|Polyuria
C0032617|T184|IS|28442001|SNOMEDCT_CORE|Urine output high|Polyuria
C0032633|T047|OAS|402567004|SNOMEDCT_CORE|Cheiropodopompholyx|Vesicular eczema of hands and/or feet
C0032633|T047|OAS|402567004|SNOMEDCT_CORE|Dyshidria|Vesicular eczema of hands and/or feet
C0032633|T047|OAS|402567004|SNOMEDCT_CORE|Dyshidrotic dermatitis|Vesicular eczema of hands and/or feet
C0032633|T047|OAS|402567004|SNOMEDCT_CORE|Dyshidrotic eczema|Vesicular eczema of hands and/or feet
C0032633|T047|OAS|402567004|SNOMEDCT_CORE|Pompholyx|Vesicular eczema of hands and/or feet
C0032633|T047|OAS|402567004|SNOMEDCT_CORE|Pompholyx eczema|Vesicular eczema of hands and/or feet
C0032633|T047|OAS|402567004|SNOMEDCT_CORE|Vesicular eczema of hands and feet|Vesicular eczema of hands and/or feet
C0032633|T047|OAF|402567004|SNOMEDCT_CORE|Vesicular eczema of hands and/or feet|Vesicular eczema of hands and/or feet
C0032633|T047|OAP|402567004|SNOMEDCT_CORE|Vesicular eczema of hands and/or feet|Vesicular eczema of hands and/or feet
C0032650|T020|OAS|82675004|SNOMEDCT_CORE|Baker's cyst|Synovial cyst of knee
C0032650|T020|SY|240008008|SNOMEDCT_CORE|Baker's cyst of knee|Synovial cyst of knee
C0032650|T020|OAS|82675004|SNOMEDCT_CORE|Popliteal cyst|Synovial cyst of knee
C0032650|T020|SY|240008008|SNOMEDCT_CORE|Popliteal cyst|Synovial cyst of knee
C0032650|T020|PT|240008008|SNOMEDCT_CORE|Synovial cyst of knee|Synovial cyst of knee
C0032650|T020|FN|240008008|SNOMEDCT_CORE|Synovial cyst of knee|Synovial cyst of knee
C0032650|T020|OAP|82675004|SNOMEDCT_CORE|Synovial cyst of popliteal space|Synovial cyst of knee
C0032650|T020|SY|240008008|SNOMEDCT_CORE|Synovial cyst of popliteal space|Synovial cyst of knee
C0032650|T020|OAF|82675004|SNOMEDCT_CORE|Synovial cyst of popliteal space|Synovial cyst of knee
C0032763|T047|SY|80193009|SNOMEDCT_CORE|Jejunal syndrome|Postgastric surgery syndrome
C0032763|T047|SY|80193009|SNOMEDCT_CORE|Post-cibal syndrome|Postgastric surgery syndrome
C0032763|T047|SY|80193009|SNOMEDCT_CORE|Postgastrectomy syndrome|Postgastric surgery syndrome
C0032763|T047|PT|80193009|SNOMEDCT_CORE|Postgastric surgery syndrome|Postgastric surgery syndrome
C0032763|T047|FN|80193009|SNOMEDCT_CORE|Postgastric surgery syndrome|Postgastric surgery syndrome
C0032768|T047|SY|2177002|SNOMEDCT_CORE|PHN - Post-herpetic neuralgia|Postherpetic neuralgia
C0032768|T047|SY|2177002|SNOMEDCT_CORE|Post-zoster neuralgia|Postherpetic neuralgia
C0032768|T047|PT|2177002|SNOMEDCT_CORE|Postherpetic neuralgia|Postherpetic neuralgia
C0032768|T047|FN|2177002|SNOMEDCT_CORE|Postherpetic neuralgia|Postherpetic neuralgia
C0032776|T046|SY|76742009|SNOMEDCT_CORE|Bleeding after menopause|Postmenopausal bleeding
C0032776|T046|SY|76742009|SNOMEDCT_CORE|PMB - Postmenopausal bleeding|Postmenopausal bleeding
C0032776|T046|PT|76742009|SNOMEDCT_CORE|Postmenopausal bleeding|Postmenopausal bleeding
C0032776|T046|FN|76742009|SNOMEDCT_CORE|Postmenopausal bleeding|Postmenopausal bleeding
C0032781|T184|SY|75803007|SNOMEDCT_CORE|Discharge from back of nose|Posterior rhinorrhea
C0032781|T184|SY|75803007|SNOMEDCT_CORE|Discharge from nasopharynx|Posterior rhinorrhea
C0032781|T184|SY|75803007|SNOMEDCT_CORE|PND - Postnasal drip|Posterior rhinorrhea
C0032781|T184|PT|75803007|SNOMEDCT_CORE|Posterior rhinorrhea|Posterior rhinorrhea
C0032781|T184|FN|75803007|SNOMEDCT_CORE|Posterior rhinorrhea|Posterior rhinorrhea
C0032781|T184|PTGB|75803007|SNOMEDCT_CORE|Posterior rhinorrhoea|Posterior rhinorrhea
C0032781|T184|SY|75803007|SNOMEDCT_CORE|Postnasal catarrh|Posterior rhinorrhea
C0032781|T184|IS|75803007|SNOMEDCT_CORE|Postnasal discharge|Posterior rhinorrhea
C0032781|T184|SY|75803007|SNOMEDCT_CORE|Postnasal drip|Posterior rhinorrhea
C0032787|T046|PT|385486001|SNOMEDCT_CORE|Postoperative complication|Postoperative complication
C0032787|T046|FN|385486001|SNOMEDCT_CORE|Postoperative complication|Postoperative complication
C0032787|T046|SY|385486001|SNOMEDCT_CORE|Postoperative problem|Postoperative complication
C0032788|T046|SYGB|110265006|SNOMEDCT_CORE|Haemorrhage postprocedure|Postoperative hemorrhage
C0032788|T046|SY|110265006|SNOMEDCT_CORE|Hemorrhage postprocedure|Postoperative hemorrhage
C0032788|T046|SY|110265006|SNOMEDCT_CORE|Postoperative bleeding|Postoperative hemorrhage
C0032788|T046|PTGB|110265006|SNOMEDCT_CORE|Postoperative haemorrhage|Postoperative hemorrhage
C0032788|T046|PT|110265006|SNOMEDCT_CORE|Postoperative hemorrhage|Postoperative hemorrhage
C0032788|T046|FN|110265006|SNOMEDCT_CORE|Postoperative hemorrhage|Postoperative hemorrhage
C0032797|T046|SY|47821001|SNOMEDCT_CORE|Bleeding postpartum|Postpartum hemorrhage
C0032797|T046|SYGB|47821001|SNOMEDCT_CORE|Haemorrhage after delivery of fetus|Postpartum hemorrhage
C0032797|T046|SYGB|47821001|SNOMEDCT_CORE|Haemorrhage after delivery of foetus|Postpartum hemorrhage
C0032797|T046|SY|47821001|SNOMEDCT_CORE|Hemorrhage after delivery of fetus|Postpartum hemorrhage
C0032797|T046|IS|47821001|SNOMEDCT_CORE|Hemorrhage after delivery of fetus, NOS|Postpartum hemorrhage
C0032797|T046|PTGB|47821001|SNOMEDCT_CORE|Postpartum haemorrhage|Postpartum hemorrhage
C0032797|T046|PT|47821001|SNOMEDCT_CORE|Postpartum hemorrhage|Postpartum hemorrhage
C0032797|T046|FN|47821001|SNOMEDCT_CORE|Postpartum hemorrhage|Postpartum hemorrhage
C0032797|T046|IS|47821001|SNOMEDCT_CORE|Postpartum hemorrhage, NOS|Postpartum hemorrhage
C0032797|T046|SYGB|47821001|SNOMEDCT_CORE|PPH - Postpartum haemorrhage|Postpartum hemorrhage
C0032797|T046|SY|47821001|SNOMEDCT_CORE|PPH - Postpartum hemorrhage|Postpartum hemorrhage
C0032807|T047|SY|20427003|SNOMEDCT_CORE|Postphlebitic syndrome|Postthrombotic syndrome
C0032807|T047|FN|20427003|SNOMEDCT_CORE|Postphlebitic syndrome|Postthrombotic syndrome
C0032807|T047|PT|20427003|SNOMEDCT_CORE|Postthrombotic syndrome|Postthrombotic syndrome
C0032807|T047|IS|20427003|SNOMEDCT_CORE|Venous ulcer of leg syndrome|Postthrombotic syndrome
C0032816|T046|FN|54012000|SNOMEDCT_CORE|Posttraumatic headache|Posttraumatic headache
C0032816|T046|PT|54012000|SNOMEDCT_CORE|Posttraumatic headache|Posttraumatic headache
C0032827|T047|SY|43339004|SNOMEDCT_CORE|K deficiency|K deficiency
C0032827|T047|SY|43339004|SNOMEDCT_CORE|Potassium deficiency|K deficiency
C0032914|T046|IS|46764007|SNOMEDCT_CORE|EPH - Edema, proteinuria and hypertension of pregnancy|Pre-eclampsia
C0032914|T046|SY|398254007|SNOMEDCT_CORE|EPH - Edema, proteinuria and hypertension of pregnancy|Pre-eclampsia
C0032914|T046|IS|46764007|SNOMEDCT_CORE|EPH - Oedema, proteinuria and hypertension of pregnancy|Pre-eclampsia
C0032914|T046|SYGB|398254007|SNOMEDCT_CORE|EPH - Oedema, proteinuria and hypertension of pregnancy|Pre-eclampsia
C0032914|T046|IS|46764007|SNOMEDCT_CORE|PE - Pre-eclampsia|Pre-eclampsia
C0032914|T046|SY|398254007|SNOMEDCT_CORE|PE - Pre-eclampsia|Pre-eclampsia
C0032914|T046|IS|46764007|SNOMEDCT_CORE|PET - Pre-eclamptic toxaemia|Pre-eclampsia
C0032914|T046|SYGB|398254007|SNOMEDCT_CORE|PET - Pre-eclamptic toxaemia|Pre-eclampsia
C0032914|T046|IS|46764007|SNOMEDCT_CORE|PET - Pre-eclamptic toxemia|Pre-eclampsia
C0032914|T046|SY|398254007|SNOMEDCT_CORE|PET - Pre-eclamptic toxemia|Pre-eclampsia
C0032914|T046|IS|46764007|SNOMEDCT_CORE|Pre-eclampsia|Pre-eclampsia
C0032914|T046|PT|398254007|SNOMEDCT_CORE|Pre-eclampsia|Pre-eclampsia
C0032914|T046|FN|398254007|SNOMEDCT_CORE|Pre-eclampsia|Pre-eclampsia
C0032914|T046|IS|46764007|SNOMEDCT_CORE|Pre-eclamptic toxaemia|Pre-eclampsia
C0032914|T046|SYGB|398254007|SNOMEDCT_CORE|Pre-eclamptic toxaemia|Pre-eclampsia
C0032914|T046|IS|46764007|SNOMEDCT_CORE|Pre-eclamptic toxemia|Pre-eclampsia
C0032914|T046|SY|398254007|SNOMEDCT_CORE|Pre-eclamptic toxemia|Pre-eclampsia
C0032914|T046|SY|398254007|SNOMEDCT_CORE|Preeclampsia|Pre-eclampsia
C0032914|T046|IS|46764007|SNOMEDCT_CORE|Proteinuric hypertension of pregnancy|Pre-eclampsia
C0032914|T046|SY|398254007|SNOMEDCT_CORE|Proteinuric hypertension of pregnancy|Pre-eclampsia
C0032962|T046|OAP|198881004|SNOMEDCT_CORE|Pregnancy complications|Pregnancy complications
C0032962|T046|OAF|198881004|SNOMEDCT_CORE|Pregnancy complications|Pregnancy complications
C0032967|T033|PT|271903000|SNOMEDCT_CORE|H/O: pregnancy|H/O: pregnancy
C0032967|T033|IS|271903000|SNOMEDCT_CORE|History of - pregnancy|H/O: pregnancy
C0032967|T033|OF|271903000|SNOMEDCT_CORE|History of - pregnancy|H/O: pregnancy
C0032967|T033|SY|271903000|SNOMEDCT_CORE|History of pregnancy|H/O: pregnancy
C0032967|T033|FN|271903000|SNOMEDCT_CORE|History of pregnancy|H/O: pregnancy
C0032968|T033|PT|237240001|SNOMEDCT_CORE|Teenage pregnancy|Teenage pregnancy
C0032968|T033|FN|237240001|SNOMEDCT_CORE|Teenage pregnancy|Teenage pregnancy
C0032984|T046|PT|82661006|SNOMEDCT_CORE|Abdominal pregnancy|Abdominal pregnancy
C0032984|T046|FN|82661006|SNOMEDCT_CORE|Abdominal pregnancy|Abdominal pregnancy
C0032987|T046|PT|34801009|SNOMEDCT_CORE|Ectopic pregnancy|Ectopic pregnancy
C0032987|T046|FN|34801009|SNOMEDCT_CORE|Ectopic pregnancy|Ectopic pregnancy
C0032987|T046|IS|34801009|SNOMEDCT_CORE|Ectopic pregnancy, NOS|Ectopic pregnancy
C0032987|T046|SY|34801009|SNOMEDCT_CORE|EP - Ectopic pregnancy|Ectopic pregnancy
C0032989|T033|IS|16356006|SNOMEDCT_CORE|Multiple gestation|Multiple pregnancy
C0032989|T033|IS|16356006|SNOMEDCT_CORE|Multiple gestation, NOS|Multiple pregnancy
C0032989|T033|PT|16356006|SNOMEDCT_CORE|Multiple pregnancy|Multiple pregnancy
C0032989|T033|FN|16356006|SNOMEDCT_CORE|Multiple pregnancy|Multiple pregnancy
C0032989|T033|IS|16356006|SNOMEDCT_CORE|Multiple pregnancy, NOS|Multiple pregnancy
C0032992|T033|SY|169565003|SNOMEDCT_CORE|Planned pregnancy|Pregnant - planned
C0032992|T033|PT|169565003|SNOMEDCT_CORE|Pregnant - planned|Pregnant - planned
C0032992|T033|FN|169565003|SNOMEDCT_CORE|Pregnant - planned|Pregnant - planned
C0032993|T046|SY|90968009|SNOMEDCT_CORE|Post term pregnancy|Post-term pregnancy
C0032993|T046|SY|90968009|SNOMEDCT_CORE|Post-dates|Post-term pregnancy
C0032993|T046|PT|90968009|SNOMEDCT_CORE|Post-term pregnancy|Post-term pregnancy
C0032993|T046|IS|90968009|SNOMEDCT_CORE|Pregnancy beyond 42 weeks of gestation|Post-term pregnancy
C0032993|T046|SY|90968009|SNOMEDCT_CORE|Prolonged gestation|Post-term pregnancy
C0032993|T046|SY|90968009|SNOMEDCT_CORE|Prolonged pregnancy|Post-term pregnancy
C0032993|T046|FN|90968009|SNOMEDCT_CORE|Prolonged pregnancy|Post-term pregnancy
C0032994|T046|SY|79586000|SNOMEDCT_CORE|Fallopian pregnancy|Tubal pregnancy
C0032994|T046|SY|79586000|SNOMEDCT_CORE|Fallopian tube pregnancy|Tubal pregnancy
C0032994|T046|PT|79586000|SNOMEDCT_CORE|Tubal pregnancy|Tubal pregnancy
C0032994|T046|FN|79586000|SNOMEDCT_CORE|Tubal pregnancy|Tubal pregnancy
C0033036|T047|SY|284470004|SNOMEDCT_CORE|Atrial ectopic|Premature atrial contraction
C0033036|T047|SY|284470004|SNOMEDCT_CORE|Atrial extrasystoles|Premature atrial contraction
C0033036|T047|PT|287057009|SNOMEDCT_CORE|Atrial premature complex|Premature atrial contraction
C0033036|T047|FN|287057009|SNOMEDCT_CORE|Atrial premature complex|Premature atrial contraction
C0033036|T047|SY|284470004|SNOMEDCT_CORE|Atrial premature contractions|Premature atrial contraction
C0033036|T047|SYGB|287057009|SNOMEDCT_CORE|Atrial premature depolarisation|Premature atrial contraction
C0033036|T047|SY|287057009|SNOMEDCT_CORE|Atrial premature depolarization|Premature atrial contraction
C0033036|T047|SY|284470004|SNOMEDCT_CORE|Atrial premature systoles|Premature atrial contraction
C0033036|T047|SY|284470004|SNOMEDCT_CORE|PAC - Premature atrial contraction|Premature atrial contraction
C0033036|T047|PT|284470004|SNOMEDCT_CORE|Premature atrial contraction|Premature atrial contraction
C0033036|T047|FN|284470004|SNOMEDCT_CORE|Premature atrial contraction|Premature atrial contraction
C0033038|T048|SY|44001008|SNOMEDCT_CORE|Ejaculates too soon|Premature ejaculation
C0033038|T048|SY|44001008|SNOMEDCT_CORE|Ejaculatio praecox|Premature ejaculation
C0033038|T048|PT|44001008|SNOMEDCT_CORE|Premature ejaculation|Premature ejaculation
C0033038|T048|FN|44001008|SNOMEDCT_CORE|Premature ejaculation|Premature ejaculation
C0033038|T048|SY|44001008|SNOMEDCT_CORE|Premature orgasm - male|Premature ejaculation
C0033046|T047|SY|82639001|SNOMEDCT_CORE|Menstrual molimen|Premenstrual syndrome
C0033046|T047|SY|82639001|SNOMEDCT_CORE|PMS|Premenstrual syndrome
C0033046|T047|SY|82639001|SNOMEDCT_CORE|PMS - Premenstrual syndrome|Premenstrual syndrome
C0033046|T047|SY|82639001|SNOMEDCT_CORE|Premenstrual syndrome|Premenstrual syndrome
C0033074|T046|SY|49526009|SNOMEDCT_CORE|Age-related hearing loss|Presbycusis
C0033074|T046|SY|49526009|SNOMEDCT_CORE|Presbyacusia|Presbycusis
C0033074|T046|PT|49526009|SNOMEDCT_CORE|Presbycusis|Presbycusis
C0033074|T046|OF|49526009|SNOMEDCT_CORE|Presbycusis|Presbycusis
C0033074|T046|FN|49526009|SNOMEDCT_CORE|Presbycusis|Presbycusis
C0033074|T046|SY|49526009|SNOMEDCT_CORE|Senile deafness|Presbycusis
C0033075|T047|PT|41256004|SNOMEDCT_CORE|Presbyopia|Presbyopia
C0033075|T047|FN|41256004|SNOMEDCT_CORE|Presbyopia|Presbyopia
C0033119|T037|SY|312609001|SNOMEDCT_CORE|Puncture wound|Puncture wound - injury
C0033119|T037|PT|312609001|SNOMEDCT_CORE|Puncture wound - injury|Puncture wound - injury
C0033119|T037|FN|312609001|SNOMEDCT_CORE|Puncture wound - injury|Puncture wound - injury
C0033139|T047|PT|3972004|SNOMEDCT_CORE|Primary insomnia|Primary insomnia
C0033139|T047|FN|3972004|SNOMEDCT_CORE|Primary insomnia|Primary insomnia
C0033141|T047|IS|89461002|SNOMEDCT_CORE|Idiopathic cardiomyopathy|Primary cardiomyopathy
C0033141|T047|PT|89461002|SNOMEDCT_CORE|Primary cardiomyopathy|Primary cardiomyopathy
C0033141|T047|FN|89461002|SNOMEDCT_CORE|Primary cardiomyopathy|Primary cardiomyopathy
C0033141|T047|IS|89461002|SNOMEDCT_CORE|Primary idiopathic cardiomyopathy|Primary cardiomyopathy
C0033246|T047|PT|3951002|SNOMEDCT_CORE|Proctitis|Proctitis
C0033246|T047|FN|3951002|SNOMEDCT_CORE|Proctitis|Proctitis
C0033246|T047|IS|3951002|SNOMEDCT_CORE|Proctitis, NOS|Proctitis
C0033375|T191|SY|134209002|SNOMEDCT_CORE|Prolactin-secreting pituitary adenoma|Prolactinoma
C0033375|T191|PT|134209002|SNOMEDCT_CORE|Prolactinoma|Prolactinoma
C0033375|T191|OF|134209002|SNOMEDCT_CORE|Prolactinoma|Prolactinoma
C0033375|T191|FN|134209002|SNOMEDCT_CORE|Prolactinoma|Prolactinoma
C0033575|T047|IS|30281009|SNOMEDCT_CORE|Disease of prostate|Disorder of prostate
C0033575|T047|OF|30281009|SNOMEDCT_CORE|Disease of prostate|Disorder of prostate
C0033575|T047|IS|30281009|SNOMEDCT_CORE|Disease of prostate, NOS|Disorder of prostate
C0033575|T047|PT|30281009|SNOMEDCT_CORE|Disorder of prostate|Disorder of prostate
C0033575|T047|FN|30281009|SNOMEDCT_CORE|Disorder of prostate|Disorder of prostate
C0033575|T047|IS|30281009|SNOMEDCT_CORE|Disorder of prostate, NOS|Disorder of prostate
C0033575|T047|SY|30281009|SNOMEDCT_CORE|Prostate disease|Disorder of prostate
C0033575|T047|SY|30281009|SNOMEDCT_CORE|Prostatic disorder|Disorder of prostate
C0033575|T047|IS|30281009|SNOMEDCT_CORE|Prostatic disorder, NOS|Disorder of prostate
C0033578|T191|PT|126906006|SNOMEDCT_CORE|Neoplasm of prostate|Neoplasm of prostate
C0033578|T191|FN|126906006|SNOMEDCT_CORE|Neoplasm of prostate|Neoplasm of prostate
C0033578|T191|SY|126906006|SNOMEDCT_CORE|NGP - New growth of prostate|Neoplasm of prostate
C0033578|T191|SY|126906006|SNOMEDCT_CORE|Tumor of prostate|Neoplasm of prostate
C0033578|T191|SYGB|126906006|SNOMEDCT_CORE|Tumour of prostate|Neoplasm of prostate
C0033581|T047|SY|9713002|SNOMEDCT_CORE|Inflammation of prostate|Prostatitis
C0033581|T047|PT|9713002|SNOMEDCT_CORE|Prostatitis|Prostatitis
C0033581|T047|FN|9713002|SNOMEDCT_CORE|Prostatitis|Prostatitis
C0033581|T047|IS|9713002|SNOMEDCT_CORE|Prostatitis, NOS|Prostatitis
C0033677|T046|PT|238107002|SNOMEDCT_CORE|Deficiency of macronutrients|Deficiency of macronutrients
C0033677|T046|FN|238107002|SNOMEDCT_CORE|Deficiency of macronutrients|Deficiency of macronutrients
C0033677|T046|SY|238107002|SNOMEDCT_CORE|PCM - Protein-calorie malnutrition|Deficiency of macronutrients
C0033677|T046|SY|238107002|SNOMEDCT_CORE|PEM - Protein-energy malnutrition|Deficiency of macronutrients
C0033677|T046|SY|238107002|SNOMEDCT_CORE|Protein calorie malnutrition|Deficiency of macronutrients
C0033677|T046|SY|238107002|SNOMEDCT_CORE|Protein-calorie malnutrition|Deficiency of macronutrients
C0033677|T046|SY|238107002|SNOMEDCT_CORE|Protein-calorie undernutrition|Deficiency of macronutrients
C0033677|T046|SY|238107002|SNOMEDCT_CORE|Protein-energy malnutrition|Deficiency of macronutrients
C0033687|T033|SY|29738008|SNOMEDCT_CORE|Abnormal presence of protein in urine|Proteinuria
C0033687|T033|PT|29738008|SNOMEDCT_CORE|Proteinuria|Proteinuria
C0033687|T033|FN|29738008|SNOMEDCT_CORE|Proteinuria|Proteinuria
C0033687|T033|IS|29738008|SNOMEDCT_CORE|Proteinuria, NOS|Proteinuria
C0033771|T047|SY|64144002|SNOMEDCT_CORE|Itchy skin eruption|Pruritic rash
C0033771|T047|IS|64144002|SNOMEDCT_CORE|Itchy skin eruption, NOS|Pruritic rash
C0033771|T047|SY|64144002|SNOMEDCT_CORE|Prurigo|Pruritic rash
C0033771|T047|IS|64144002|SNOMEDCT_CORE|Prurigo, NOS|Pruritic rash
C0033771|T047|PT|64144002|SNOMEDCT_CORE|Pruritic rash|Pruritic rash
C0033771|T047|FN|64144002|SNOMEDCT_CORE|Pruritic rash|Pruritic rash
C0033771|T047|IS|64144002|SNOMEDCT_CORE|Pruritic rash, NOS|Pruritic rash
C0033774|T033|SY|418290006|SNOMEDCT_CORE|Itch|Itching
C0033774|T033|PT|418290006|SNOMEDCT_CORE|Itching|Itching
C0033774|T033|FN|418290006|SNOMEDCT_CORE|Itching|Itching
C0033774|T033|SY|418290006|SNOMEDCT_CORE|Itchy|Itching
C0033774|T033|SY|279333002|SNOMEDCT_CORE|Pruritic dermatitis|Itching
C0033774|T033|SY|279333002|SNOMEDCT_CORE|Pruritic disorder|Itching
C0033774|T033|FN|279333002|SNOMEDCT_CORE|Pruritic disorder|Itching
C0033774|T033|IS|279333002|SNOMEDCT_CORE|Pruritic disorders|Itching
C0033774|T033|OF|279333002|SNOMEDCT_CORE|Pruritic disorders|Itching
C0033774|T033|SY|279333002|SNOMEDCT_CORE|Pruritus - disorder|Itching
C0033774|T033|PT|279333002|SNOMEDCT_CORE|Pruritus of skin|Itching
C0033775|T184|SY|90446007|SNOMEDCT_CORE|Anal itch|Pruritus ani
C0033775|T184|SY|90446007|SNOMEDCT_CORE|Perianal itch|Pruritus ani
C0033775|T184|PT|90446007|SNOMEDCT_CORE|Pruritus ani|Pruritus ani
C0033775|T184|OF|90446007|SNOMEDCT_CORE|Pruritus ani|Pruritus ani
C0033775|T184|FN|90446007|SNOMEDCT_CORE|Pruritus ani|Pruritus ani
C0033777|T184|SY|267802000|SNOMEDCT_CORE|Genital pruritus|Pruritus of genital organs
C0033777|T184|PT|267802000|SNOMEDCT_CORE|Pruritus of genital organs|Pruritus of genital organs
C0033777|T184|FN|267802000|SNOMEDCT_CORE|Pruritus of genital organs|Pruritus of genital organs
C0033778|T184|SY|67882000|SNOMEDCT_CORE|Itching of vulva|Pruritus of vulva
C0033778|T184|PT|67882000|SNOMEDCT_CORE|Pruritus of vulva|Pruritus of vulva
C0033778|T184|FN|67882000|SNOMEDCT_CORE|Pruritus of vulva|Pruritus of vulva
C0033778|T184|SY|67882000|SNOMEDCT_CORE|Pruritus vulvae|Pruritus of vulva
C0033778|T184|SY|67882000|SNOMEDCT_CORE|Vulval itching|Pruritus of vulva
C0033802|T047|OAF|60782007|SNOMEDCT_CORE|Pseudogout|Pseudogout
C0033802|T047|IS|60782007|SNOMEDCT_CORE|Pseudogout, NOS|Pseudogout, NOS
C0033806|T047|SYGB|58976002|SNOMEDCT_CORE|Constitutional chronic hypocalcaemia|Pseudohypoparathyroidism
C0033806|T047|SY|58976002|SNOMEDCT_CORE|Constitutional chronic hypocalcemia|Pseudohypoparathyroidism
C0033806|T047|SY|58976002|SNOMEDCT_CORE|Familial pseudohypoparathyroidism|Pseudohypoparathyroidism
C0033806|T047|SY|58976002|SNOMEDCT_CORE|Parathyroid hormone resistant hypoparathyroidism|Pseudohypoparathyroidism
C0033806|T047|PT|58976002|SNOMEDCT_CORE|Pseudohypoparathyroidism|Pseudohypoparathyroidism
C0033806|T047|FN|58976002|SNOMEDCT_CORE|Pseudohypoparathyroidism|Pseudohypoparathyroidism
C0033806|T047|IS|58976002|SNOMEDCT_CORE|Pseudohypoparathyroidism, NOS|Pseudohypoparathyroidism
C0033817|T047|SY|63398001|SNOMEDCT_CORE|Bacterial infection caused by Pseudomonas|Bacterial infection due to Pseudomonas
C0033817|T047|FN|63398001|SNOMEDCT_CORE|Bacterial infection caused by Pseudomonas|Bacterial infection due to Pseudomonas
C0033817|T047|PT|63398001|SNOMEDCT_CORE|Bacterial infection due to Pseudomonas|Bacterial infection due to Pseudomonas
C0033817|T047|OF|63398001|SNOMEDCT_CORE|Bacterial infection due to Pseudomonas|Bacterial infection due to Pseudomonas
C0033817|T047|SY|63398001|SNOMEDCT_CORE|Pseudomonas infection|Bacterial infection due to Pseudomonas
C0033822|T191|PT|307601000|SNOMEDCT_CORE|Pseudomyxoma peritonei|Pseudomyxoma peritonei
C0033822|T191|FN|307601000|SNOMEDCT_CORE|Pseudomyxoma peritonei|Pseudomyxoma peritonei
C0033845|T047|PT|68267002|SNOMEDCT_CORE|Benign intracranial hypertension|Benign intracranial hypertension
C0033845|T047|FN|68267002|SNOMEDCT_CORE|Benign intracranial hypertension|Benign intracranial hypertension
C0033845|T047|SY|68267002|SNOMEDCT_CORE|BIH - Benign intracranial hypertension|Benign intracranial hypertension
C0033845|T047|SY|68267002|SNOMEDCT_CORE|Idiopathic intracranial hypertension|Benign intracranial hypertension
C0033845|T047|SY|68267002|SNOMEDCT_CORE|IIH - Idiopathic intracranial hypertension|Benign intracranial hypertension
C0033845|T047|SY|68267002|SNOMEDCT_CORE|Noninfective serous meningitis|Benign intracranial hypertension
C0033845|T047|SY|68267002|SNOMEDCT_CORE|Nonne's syndrome|Benign intracranial hypertension
C0033845|T047|SY|68267002|SNOMEDCT_CORE|Otitic hydrocephalus syndrome|Benign intracranial hypertension
C0033845|T047|SY|68267002|SNOMEDCT_CORE|Pseudotumor cerebri|Benign intracranial hypertension
C0033845|T047|SYGB|68267002|SNOMEDCT_CORE|Pseudotumour cerebri|Benign intracranial hypertension
C0033860|T047|PT|9014002|SNOMEDCT_CORE|Psoriasis|Psoriasis
C0033860|T047|FN|9014002|SNOMEDCT_CORE|Psoriasis|Psoriasis
C0033860|T047|IS|9014002|SNOMEDCT_CORE|Psoriasis, NOS|Psoriasis
C0033883|T048|PT|11387009|SNOMEDCT_CORE|Psychoactive substance-induced organic mental disorder|Psychoactive substance-induced organic mental disorder
C0033883|T048|FN|11387009|SNOMEDCT_CORE|Psychoactive substance-induced organic mental disorder|Psychoactive substance-induced organic mental disorder
C0033883|T048|IS|11387009|SNOMEDCT_CORE|Psychoactive substance-induced organic mental disorder, NOS|Psychoactive substance-induced organic mental disorder
C0033893|T047|SY|398057008|SNOMEDCT_CORE|Tension headache|Tension-type headache
C0033893|T047|PT|398057008|SNOMEDCT_CORE|Tension-type headache|Tension-type headache
C0033893|T047|FN|398057008|SNOMEDCT_CORE|Tension-type headache|Tension-type headache
C0033936|T048|SY|42344001|SNOMEDCT_CORE|Alcohol induced psychosis|Alcohol-induced psychosis
C0033936|T048|PT|42344001|SNOMEDCT_CORE|Alcohol-induced psychosis|Alcohol-induced psychosis
C0033936|T048|FN|42344001|SNOMEDCT_CORE|Alcohol-induced psychosis|Alcohol-induced psychosis
C0033936|T048|IS|42344001|SNOMEDCT_CORE|Alcohol-induced psychosis, NOS|Alcohol-induced psychosis
C0033936|T048|SY|42344001|SNOMEDCT_CORE|Alcoholic psychosis|Alcohol-induced psychosis
C0033936|T048|IS|42344001|SNOMEDCT_CORE|Alcoholic psychosis, NOS|Alcohol-induced psychosis
C0033975|T048|IS|69322001|SNOMEDCT_CORE|Atypical psychosis|Psychotic disorder
C0033975|T048|SY|69322001|SNOMEDCT_CORE|Psychosis|Psychotic disorder
C0033975|T048|IS|69322001|SNOMEDCT_CORE|Psychosis, NOS|Psychotic disorder
C0033975|T048|IS|69322001|SNOMEDCT_CORE|Psychotic|Psychotic disorder
C0033975|T048|PT|69322001|SNOMEDCT_CORE|Psychotic disorder|Psychotic disorder
C0033975|T048|FN|69322001|SNOMEDCT_CORE|Psychotic disorder|Psychotic disorder
C0033975|T048|IS|69322001|SNOMEDCT_CORE|Psychotic disorder, NOS|Psychotic disorder
C0034012|T046|PT|400003000|SNOMEDCT_CORE|Delayed puberty|Delayed puberty
C0034012|T046|FN|400003000|SNOMEDCT_CORE|Delayed puberty|Delayed puberty
C0034013|T047|PT|400179000|SNOMEDCT_CORE|Precocious puberty|Precocious puberty
C0034013|T047|FN|400179000|SNOMEDCT_CORE|Precocious puberty|Precocious puberty
C0034063|T046|PT|19242006|SNOMEDCT_CORE|Pulmonary edema|Pulmonary edema
C0034063|T046|FN|19242006|SNOMEDCT_CORE|Pulmonary edema|Pulmonary edema
C0034063|T046|IS|19242006|SNOMEDCT_CORE|Pulmonary edema, NOS|Pulmonary edema
C0034063|T046|PTGB|19242006|SNOMEDCT_CORE|Pulmonary oedema|Pulmonary edema
C0034065|T046|SY|59282003|SNOMEDCT_CORE|PE - Pulmonary embolism|Pulmonary embolism
C0034065|T046|PT|59282003|SNOMEDCT_CORE|Pulmonary embolism|Pulmonary embolism
C0034065|T046|FN|59282003|SNOMEDCT_CORE|Pulmonary embolism|Pulmonary embolism
C0034067|T047|SY|87433001|SNOMEDCT_CORE|Emphysema of lung|Pulmonary emphysema
C0034067|T047|IS|87433001|SNOMEDCT_CORE|Emphysema of lung, NOS|Pulmonary emphysema
C0034067|T047|PT|87433001|SNOMEDCT_CORE|Pulmonary emphysema|Pulmonary emphysema
C0034067|T047|FN|87433001|SNOMEDCT_CORE|Pulmonary emphysema|Pulmonary emphysema
C0034067|T047|IS|87433001|SNOMEDCT_CORE|Pulmonary emphysema, NOS|Pulmonary emphysema
C0034069|T047|SY|51615001|SNOMEDCT_CORE|Cirrhosis of lung|Fibrosis of lung
C0034069|T047|IS|51615001|SNOMEDCT_CORE|Cirrhosis of lung, NOS|Fibrosis of lung
C0034069|T047|PT|51615001|SNOMEDCT_CORE|Fibrosis of lung|Fibrosis of lung
C0034069|T047|FN|51615001|SNOMEDCT_CORE|Fibrosis of lung|Fibrosis of lung
C0034069|T047|IS|51615001|SNOMEDCT_CORE|Fibrosis of lung, NOS|Fibrosis of lung
C0034069|T047|SY|51615001|SNOMEDCT_CORE|Pulmonary fibrosis|Fibrosis of lung
C0034072|T047|PT|83291003|SNOMEDCT_CORE|Cor pulmonale|Cor pulmonale
C0034072|T047|FN|83291003|SNOMEDCT_CORE|Cor pulmonale|Cor pulmonale
C0034072|T047|SY|83291003|SNOMEDCT_CORE|Right heart failure due to disorder of lung|Cor pulmonale
C0034072|T047|SY|83291003|SNOMEDCT_CORE|Right heart failure due to pulmonary disease|Cor pulmonale
C0034088|T046|SY|91434003|SNOMEDCT_CORE|PR - Pulmonary regurgitation|Pulmonic valve regurgitation
C0034088|T046|SY|91434003|SNOMEDCT_CORE|Pulmonary valve incompetence|Pulmonic valve regurgitation
C0034088|T046|IS|91434003|SNOMEDCT_CORE|Pulmonary valve incompetence, NOS|Pulmonic valve regurgitation
C0034088|T046|SY|91434003|SNOMEDCT_CORE|Pulmonary valve insufficiency|Pulmonic valve regurgitation
C0034088|T046|IS|91434003|SNOMEDCT_CORE|Pulmonary valve insufficiency, NOS|Pulmonic valve regurgitation
C0034088|T046|SY|91434003|SNOMEDCT_CORE|Pulmonary valve regurgitation|Pulmonic valve regurgitation
C0034088|T046|SY|91434003|SNOMEDCT_CORE|Pulmonic insufficiency|Pulmonic valve regurgitation
C0034088|T046|SY|91434003|SNOMEDCT_CORE|Pulmonic regurgitation|Pulmonic valve regurgitation
C0034088|T046|IS|91434003|SNOMEDCT_CORE|Pulmonic regurgitation, NOS|Pulmonic valve regurgitation
C0034088|T046|SY|91434003|SNOMEDCT_CORE|Pulmonic valve incompetence|Pulmonic valve regurgitation
C0034088|T046|IS|91434003|SNOMEDCT_CORE|Pulmonic valve incompetence, NOS|Pulmonic valve regurgitation
C0034088|T046|SY|91434003|SNOMEDCT_CORE|Pulmonic valve insufficiency|Pulmonic valve regurgitation
C0034088|T046|IS|91434003|SNOMEDCT_CORE|Pulmonic valve insufficiency, NOS|Pulmonic valve regurgitation
C0034088|T046|PT|91434003|SNOMEDCT_CORE|Pulmonic valve regurgitation|Pulmonic valve regurgitation
C0034088|T046|FN|91434003|SNOMEDCT_CORE|Pulmonic valve regurgitation|Pulmonic valve regurgitation
C0034088|T046|IS|91434003|SNOMEDCT_CORE|Pulmonic valve regurgitation, NOS|Pulmonic valve regurgitation
C0034088|T046|SY|91434003|SNOMEDCT_CORE|PVR - Pulmonary regurgitation|Pulmonic valve regurgitation
C0034150|T047|PT|423902002|SNOMEDCT_CORE|Purpura|Purpura
C0034150|T047|FN|423902002|SNOMEDCT_CORE|Purpura|Purpura
C0034152|T047|SY|191306005|SNOMEDCT_CORE|Acute vascular purpura|Henoch-Schönlein purpura
C0034152|T047|SY|191306005|SNOMEDCT_CORE|Anaphylactoid purpura|Henoch-Schönlein purpura
C0034152|T047|SY|191306005|SNOMEDCT_CORE|Autoimmune purpura|Henoch-Schönlein purpura
C0034152|T047|IS|191306005|SNOMEDCT_CORE|Henoch-Schoenlein purpura|Henoch-Schönlein purpura
C0034152|T047|SY|191306005|SNOMEDCT_CORE|Henoch-Schoenlein vasculitis|Henoch-Schönlein purpura
C0034152|T047|SY|191306005|SNOMEDCT_CORE|Henoch-Schonlein purpura|Henoch-Schönlein purpura
C0034152|T047|PT|191306005|SNOMEDCT_CORE|Henoch-Schönlein purpura|Henoch-Schönlein purpura
C0034152|T047|FN|191306005|SNOMEDCT_CORE|Henoch-Schönlein purpura|Henoch-Schönlein purpura
C0034152|T047|OF|191306005|SNOMEDCT_CORE|Henoch-Schonlein purpura|Henoch-Schönlein purpura
C0034152|T047|SY|191306005|SNOMEDCT_CORE|Henoch's purpura|Henoch-Schönlein purpura
C0034152|T047|SY|191306005|SNOMEDCT_CORE|HSP - Henoch-Schonlein purpura|Henoch-Schönlein purpura
C0034152|T047|SY|191306005|SNOMEDCT_CORE|Spring fever|Henoch-Schönlein purpura
C0034155|T047|SY|78129009|SNOMEDCT_CORE|Moschcowitz syndrome|Thrombotic thrombocytopenic purpura
C0034155|T047|SY|78129009|SNOMEDCT_CORE|Moschowitz's syndrome|Thrombotic thrombocytopenic purpura
C0034155|T047|PT|78129009|SNOMEDCT_CORE|Thrombotic thrombocytopenic purpura|Thrombotic thrombocytopenic purpura
C0034155|T047|FN|78129009|SNOMEDCT_CORE|Thrombotic thrombocytopenic purpura|Thrombotic thrombocytopenic purpura
C0034155|T047|SY|78129009|SNOMEDCT_CORE|TTP|Thrombotic thrombocytopenic purpura
C0034155|T047|SY|78129009|SNOMEDCT_CORE|TTP - Thrombotic thrombocytopenic purpura|Thrombotic thrombocytopenic purpura
C0034186|T047|PT|45816000|SNOMEDCT_CORE|Pyelonephritis|Pyelonephritis
C0034186|T047|FN|45816000|SNOMEDCT_CORE|Pyelonephritis|Pyelonephritis
C0034186|T047|IS|45816000|SNOMEDCT_CORE|Pyelonephritis, NOS|Pyelonephritis
C0034194|T046|SY|367403001|SNOMEDCT_CORE|PS - Pyloric stenosis|Pyloric stenosis
C0034194|T046|PT|367403001|SNOMEDCT_CORE|Pyloric stenosis|Pyloric stenosis
C0034194|T046|FN|367403001|SNOMEDCT_CORE|Pyloric stenosis|Pyloric stenosis
C0034212|T047|SY|70759006|SNOMEDCT_CORE|Purulent dermatitis|Pyoderma
C0034212|T047|PT|70759006|SNOMEDCT_CORE|Pyoderma|Pyoderma
C0034212|T047|FN|70759006|SNOMEDCT_CORE|Pyoderma|Pyoderma
C0034212|T047|SY|70759006|SNOMEDCT_CORE|Pyodermia|Pyoderma
C0034212|T047|SY|70759006|SNOMEDCT_CORE|Pyogenic dermatitis|Pyoderma
C0034212|T047|SY|70759006|SNOMEDCT_CORE|Pyogenic infection of skin and subcutis|Pyoderma
C0034212|T047|SY|70759006|SNOMEDCT_CORE|Septic dermatitis|Pyoderma
C0034212|T047|SY|70759006|SNOMEDCT_CORE|Suppurative dermatitis|Pyoderma
C0034215|T047|PT|88981003|SNOMEDCT_CORE|Pyometra|Pyometra
C0034215|T047|FN|88981003|SNOMEDCT_CORE|Pyometra|Pyometra
C0034215|T047|SY|88981003|SNOMEDCT_CORE|Pyometrium|Pyometra
C0034216|T047|PT|48631008|SNOMEDCT_CORE|Pyonephrosis|Pyonephrosis
C0034216|T047|FN|48631008|SNOMEDCT_CORE|Pyonephrosis|Pyonephrosis
C0034220|T047|SY|397810006|SNOMEDCT_CORE|Pyosalpingitis|Pyosalpinx
C0034220|T047|PT|397810006|SNOMEDCT_CORE|Pyosalpinx|Pyosalpinx
C0034220|T047|FN|397810006|SNOMEDCT_CORE|Pyosalpinx|Pyosalpinx
C0034359|T033|PT|4800001|SNOMEDCT_CORE|Pyuria|Pyuria
C0034359|T033|FN|4800001|SNOMEDCT_CORE|Pyuria|Pyuria
C0034372|T047|SY|11538006|SNOMEDCT_CORE|Quadriplegia|Tetraplegia
C0034372|T047|FN|11538006|SNOMEDCT_CORE|Quadriplegia|Tetraplegia
C0034372|T047|PT|11538006|SNOMEDCT_CORE|Tetraplegia|Tetraplegia
C0034561|T037|FN|49084001|SNOMEDCT_CORE|Dermatitis caused by radiation|Radiation dermatitis
C0034561|T037|SY|49084001|SNOMEDCT_CORE|Dermatitis caused by radiation|Radiation dermatitis
C0034561|T037|PT|49084001|SNOMEDCT_CORE|Radiation dermatitis|Radiation dermatitis
C0034561|T037|OF|49084001|SNOMEDCT_CORE|Radiation dermatitis|Radiation dermatitis
C0034561|T037|IS|49084001|SNOMEDCT_CORE|Radiation dermatitis, NOS|Radiation dermatitis
C0034561|T037|SY|49084001|SNOMEDCT_CORE|Radiodermatitis|Radiation dermatitis
C0034561|T037|IS|49084001|SNOMEDCT_CORE|Radiodermatitis, NOS|Radiation dermatitis
C0034628|T037|PT|12676007|SNOMEDCT_CORE|Fracture of radius|Fracture of radius
C0034628|T037|FN|12676007|SNOMEDCT_CORE|Fracture of radius|Fracture of radius
C0034628|T037|IS|12676007|SNOMEDCT_CORE|Fracture of radius, NOS|Fracture of radius
C0034642|T033|IS|48409008|SNOMEDCT_CORE|Crepitant rales|Respiratory crackles
C0034642|T033|SY|48409008|SNOMEDCT_CORE|Rales|Respiratory crackles
C0034642|T033|PT|48409008|SNOMEDCT_CORE|Respiratory crackles|Respiratory crackles
C0034642|T033|FN|48409008|SNOMEDCT_CORE|Respiratory crackles|Respiratory crackles
C0034642|T033|SY|48409008|SNOMEDCT_CORE|Respiratory crepitations|Respiratory crackles
C0034734|T047|SY|195295006|SNOMEDCT_CORE|Raynaud disease|Raynaud's disease
C0034734|T047|PT|195295006|SNOMEDCT_CORE|Raynaud's disease|Raynaud's disease
C0034734|T047|FN|195295006|SNOMEDCT_CORE|Raynaud's disease|Raynaud's disease
C0034734|T047|SY|195295006|SNOMEDCT_CORE|Raynauds disease|Raynaud's disease
C0034735|T047|SY|266261006|SNOMEDCT_CORE|Paroxysmal digital cyanosis|Raynaud's phenomenon
C0034735|T047|SY|266261006|SNOMEDCT_CORE|Raynaud phenomenon|Raynaud's phenomenon
C0034735|T047|PT|266261006|SNOMEDCT_CORE|Raynaud's phenomenon|Raynaud's phenomenon
C0034735|T047|OF|266261006|SNOMEDCT_CORE|Raynaud's phenomenon|Raynaud's phenomenon
C0034735|T047|FN|266261006|SNOMEDCT_CORE|Raynaud's phenomenon|Raynaud's phenomenon
C0034885|T191|PT|126847008|SNOMEDCT_CORE|Neoplasm of rectum|Neoplasm of rectum
C0034885|T191|FN|126847008|SNOMEDCT_CORE|Neoplasm of rectum|Neoplasm of rectum
C0034885|T191|SY|126847008|SNOMEDCT_CORE|Tumor of rectum|Neoplasm of rectum
C0034885|T191|SYGB|126847008|SNOMEDCT_CORE|Tumour of rectum|Neoplasm of rectum
C0034886|T184|SY|77880009|SNOMEDCT_CORE|Pain in rectum|Rectal pain
C0034886|T184|SY|77880009|SNOMEDCT_CORE|Proctalgia|Rectal pain
C0034886|T184|PT|77880009|SNOMEDCT_CORE|Rectal pain|Rectal pain
C0034886|T184|FN|77880009|SNOMEDCT_CORE|Rectal pain|Rectal pain
C0034886|T184|SY|77880009|SNOMEDCT_CORE|Rectalgia|Rectal pain
C0034887|T191|SY|39772007|SNOMEDCT_CORE|Polyp of rectum|Rectal polyp
C0034887|T191|PT|39772007|SNOMEDCT_CORE|Rectal polyp|Rectal polyp
C0034887|T191|FN|39772007|SNOMEDCT_CORE|Rectal polyp|Rectal polyp
C0034888|T047|SY|57773001|SNOMEDCT_CORE|Procidentia of rectum|Rectal prolapse
C0034888|T047|SY|57773001|SNOMEDCT_CORE|Rectal mucosa prolapse|Rectal prolapse
C0034888|T047|PT|57773001|SNOMEDCT_CORE|Rectal prolapse|Rectal prolapse
C0034888|T047|FN|57773001|SNOMEDCT_CORE|Rectal prolapse|Rectal prolapse
C0034888|T047|SY|57773001|SNOMEDCT_CORE|RP - Rectal prolapse|Rectal prolapse
C0034895|T190|PT|65619001|SNOMEDCT_CORE|Rectovaginal fistula|Rectovaginal fistula
C0034895|T190|FN|65619001|SNOMEDCT_CORE|Rectovaginal fistula|Rectovaginal fistula
C0034895|T190|SY|65619001|SNOMEDCT_CORE|RVF - Rectovaginal fistula|Rectovaginal fistula
C0034902|T047|SY|50715003|SNOMEDCT_CORE|Primary red cell aplasia|Pure red cell aplasia
C0034902|T047|SYGB|50715003|SNOMEDCT_CORE|Pure red cell anaemia|Pure red cell aplasia
C0034902|T047|SY|50715003|SNOMEDCT_CORE|Pure red cell anemia|Pure red cell aplasia
C0034902|T047|IS|50715003|SNOMEDCT_CORE|Pure red cell anemia, NOS|Pure red cell aplasia
C0034902|T047|PT|50715003|SNOMEDCT_CORE|Pure red cell aplasia|Pure red cell aplasia
C0034902|T047|FN|50715003|SNOMEDCT_CORE|Pure red cell aplasia|Pure red cell aplasia
C0034902|T047|IS|50715003|SNOMEDCT_CORE|Pure red cell aplasia, NOS|Pure red cell aplasia
C0034902|T047|SY|50715003|SNOMEDCT_CORE|Red cell hypoplasia|Pure red cell aplasia
C0034919|T047|PT|266570005|SNOMEDCT_CORE|Redundant prepuce and phimosis|Redundant prepuce and phimosis
C0034919|T047|FN|266570005|SNOMEDCT_CORE|Redundant prepuce and phimosis|Redundant prepuce and phimosis
C0034919|T047|SY|266570005|SNOMEDCT_CORE|Redundant prepuce with phimosis|Redundant prepuce and phimosis
C0034931|T047|OAS|50642008|SNOMEDCT_CORE|Algodystrophy|Complex regional pain syndrome type I
C0034931|T047|OAF|50642008|SNOMEDCT_CORE|Algodystrophy|Complex regional pain syndrome type I
C0034931|T047|OAS|50642008|SNOMEDCT_CORE|Algoneurodystrophy|Complex regional pain syndrome type I
C0034931|T047|SY|734947007|SNOMEDCT_CORE|Complex regional pain syndrome type 1|Complex regional pain syndrome type I
C0034931|T047|OAS|50642008|SNOMEDCT_CORE|Complex regional pain syndrome type I|Complex regional pain syndrome type I
C0034931|T047|PT|734947007|SNOMEDCT_CORE|Complex regional pain syndrome type I|Complex regional pain syndrome type I
C0034931|T047|FN|734947007|SNOMEDCT_CORE|Complex regional pain syndrome type I|Complex regional pain syndrome type I
C0034931|T047|OAS|128079007|SNOMEDCT_CORE|Complex regional pain syndrome, type I|Complex regional pain syndrome type I
C0034931|T047|OAP|50642008|SNOMEDCT_CORE|Complex regional pain syndrome, type I|Complex regional pain syndrome type I
C0034931|T047|OAS|50642008|SNOMEDCT_CORE|CRPS - Complex regional pain syndrome type I|Complex regional pain syndrome type I
C0034931|T047|OAP|128079007|SNOMEDCT_CORE|Reflex sympathetic dystrophy|Complex regional pain syndrome type I
C0034931|T047|IS|50642008|SNOMEDCT_CORE|Reflex sympathetic dystrophy|Complex regional pain syndrome type I
C0034931|T047|SY|734947007|SNOMEDCT_CORE|Reflex sympathetic dystrophy|Complex regional pain syndrome type I
C0034931|T047|OAF|128079007|SNOMEDCT_CORE|Reflex sympathetic dystrophy|Complex regional pain syndrome type I
C0034931|T047|OAS|50642008|SNOMEDCT_CORE|RSD - Reflex sympathetic dystrophy|Complex regional pain syndrome type I
C0034931|T047|OAS|128079007|SNOMEDCT_CORE|Sudek's atrophy|Complex regional pain syndrome type I
C0034931|T047|OAS|50642008|SNOMEDCT_CORE|Sudek's atrophy|Complex regional pain syndrome type I
C0034951|T047|PT|39021009|SNOMEDCT_CORE|Disorder of refraction|Disorder of refraction
C0034951|T047|FN|39021009|SNOMEDCT_CORE|Disorder of refraction|Disorder of refraction
C0034951|T047|IS|39021009|SNOMEDCT_CORE|Disorder of refraction, NOS|Disorder of refraction
C0034951|T047|SY|39021009|SNOMEDCT_CORE|Refractive error|Disorder of refraction
C0034951|T047|IS|39021009|SNOMEDCT_CORE|Refractive error, NOS|Disorder of refraction
C0035067|T047|SY|302233006|SNOMEDCT_CORE|RAS - Renal artery stenosis|Renal artery stenosis
C0035067|T047|PT|302233006|SNOMEDCT_CORE|Renal artery stenosis|Renal artery stenosis
C0035067|T047|FN|302233006|SNOMEDCT_CORE|Renal artery stenosis|Renal artery stenosis
C0035078|T047|SY|42399005|SNOMEDCT_CORE|Renal failure|Renal failure syndrome
C0035078|T047|PT|42399005|SNOMEDCT_CORE|Renal failure syndrome|Renal failure syndrome
C0035078|T047|FN|42399005|SNOMEDCT_CORE|Renal failure syndrome|Renal failure syndrome
C0035078|T047|IS|42399005|SNOMEDCT_CORE|Renal failure syndrome, NOS|Renal failure syndrome
C0035078|T047|IS|42399005|SNOMEDCT_CORE|Renal insufficiency|Renal failure syndrome
C0035078|T047|IS|42399005|SNOMEDCT_CORE|Renal insufficiency syndrome|Renal failure syndrome
C0035078|T047|IS|42399005|SNOMEDCT_CORE|Renal insufficiency syndrome, NOS|Renal failure syndrome
C0035078|T047|SY|42399005|SNOMEDCT_CORE|RF - Renal failure|Renal failure syndrome
C0035086|T047|SY|16726004|SNOMEDCT_CORE|Renal bone disease|Renal osteodystrophy
C0035086|T047|PT|16726004|SNOMEDCT_CORE|Renal osteodystrophy|Renal osteodystrophy
C0035086|T047|FN|16726004|SNOMEDCT_CORE|Renal osteodystrophy|Renal osteodystrophy
C0035086|T047|SY|16726004|SNOMEDCT_CORE|ROD - Renal osteodystrophy|Renal osteodystrophy
C0035127|T047|PT|788465007|SNOMEDCT_CORE|Repetitive motion disorder|Repetitive motion disorder
C0035127|T047|FN|788465007|SNOMEDCT_CORE|Repetitive motion disorder|Repetitive motion disorder
C0035127|T047|OAP|4308002|SNOMEDCT_CORE|Repetitive strain injury|Repetitive motion disorder
C0035127|T047|SY|788465007|SNOMEDCT_CORE|Repetitive strain injury|Repetitive motion disorder
C0035127|T047|OAF|4308002|SNOMEDCT_CORE|Repetitive strain injury|Repetitive motion disorder
C0035127|T047|OAS|4308002|SNOMEDCT_CORE|Repetitive strain injury syndrome|Repetitive motion disorder
C0035127|T047|SY|788465007|SNOMEDCT_CORE|Repetitive strain injury syndrome|Repetitive motion disorder
C0035127|T047|IS|4308002|SNOMEDCT_CORE|Repetitive strain injury, NOS|Repetitive motion disorder
C0035127|T047|SY|788465007|SNOMEDCT_CORE|Repetitive stress injury|Repetitive motion disorder
C0035127|T047|IS|4308002|SNOMEDCT_CORE|RSI|Repetitive motion disorder
C0035127|T047|OAS|4308002|SNOMEDCT_CORE|RSI - Repetitive strain injury|Repetitive motion disorder
C0035127|T047|SY|788465007|SNOMEDCT_CORE|RSI - Repetitive strain injury|Repetitive motion disorder
C0035127|T047|OAS|4308002|SNOMEDCT_CORE|RSIS - Repetitive strain injury syndrome|Repetitive motion disorder
C0035127|T047|SY|788465007|SNOMEDCT_CORE|RSIS - Repetitive strain injury syndrome|Repetitive motion disorder
C0035204|T047|IS|50043002|SNOMEDCT_CORE|Disease of respiratory system|Disorder of respiratory system
C0035204|T047|OF|50043002|SNOMEDCT_CORE|Disease of respiratory system|Disorder of respiratory system
C0035204|T047|IS|50043002|SNOMEDCT_CORE|Disease of respiratory system, NOS|Disorder of respiratory system
C0035204|T047|PT|50043002|SNOMEDCT_CORE|Disorder of respiratory system|Disorder of respiratory system
C0035204|T047|FN|50043002|SNOMEDCT_CORE|Disorder of respiratory system|Disorder of respiratory system
C0035204|T047|SY|50043002|SNOMEDCT_CORE|Respiratory disease|Disorder of respiratory system
C0035204|T047|SY|50043002|SNOMEDCT_CORE|Respiratory disorder|Disorder of respiratory system
C0035204|T047|IS|50043002|SNOMEDCT_CORE|Respiratory disorder, NOS|Disorder of respiratory system
C0035204|T047|SY|50043002|SNOMEDCT_CORE|Respiratory system disease|Disorder of respiratory system
C0035220|T047|SY|46775006|SNOMEDCT_CORE|Cardiorespiratory distress syndrome of newborn|Respiratory distress syndrome in the newborn
C0035220|T047|SY|46775006|SNOMEDCT_CORE|Congenital alveolar dysplasia|Respiratory distress syndrome in the newborn
C0035220|T047|SY|46775006|SNOMEDCT_CORE|Idiopathic respiratory distress syndrome|Respiratory distress syndrome in the newborn
C0035220|T047|SY|46775006|SNOMEDCT_CORE|Idiopathic respiratory distress syndrome of newborn|Respiratory distress syndrome in the newborn
C0035220|T047|SY|46775006|SNOMEDCT_CORE|IRDS - Idiopathic respiratory distress syndrome|Respiratory distress syndrome in the newborn
C0035220|T047|SY|46775006|SNOMEDCT_CORE|IRDS of newborn|Respiratory distress syndrome in the newborn
C0035220|T047|SY|46775006|SNOMEDCT_CORE|Neonatal respiratory distress syndrome|Respiratory distress syndrome in the newborn
C0035220|T047|SY|46775006|SNOMEDCT_CORE|Pulmonary hypoperfusion syndrome of newborn|Respiratory distress syndrome in the newborn
C0035220|T047|SY|46775006|SNOMEDCT_CORE|RDS - Respiratory distress syndrome of newborn|Respiratory distress syndrome in the newborn
C0035220|T047|SY|46775006|SNOMEDCT_CORE|RDS of newborn|Respiratory distress syndrome in the newborn
C0035220|T047|SY|46775006|SNOMEDCT_CORE|Respiratory distress syndrome in neonate|Respiratory distress syndrome in the newborn
C0035220|T047|PT|46775006|SNOMEDCT_CORE|Respiratory distress syndrome in the newborn|Respiratory distress syndrome in the newborn
C0035220|T047|FN|46775006|SNOMEDCT_CORE|Respiratory distress syndrome in the newborn|Respiratory distress syndrome in the newborn
C0035220|T047|SY|46775006|SNOMEDCT_CORE|Respiratory distress syndrome of newborn|Respiratory distress syndrome in the newborn
C0035220|T047|SY|46775006|SNOMEDCT_CORE|Wet lung disease of newborn|Respiratory distress syndrome in the newborn
C0035222|T047|SY|67782005|SNOMEDCT_CORE|Acquired respiratory distress syndrome|Acute respiratory distress syndrome
C0035222|T047|PT|67782005|SNOMEDCT_CORE|Acute respiratory distress syndrome|Acute respiratory distress syndrome
C0035222|T047|FN|67782005|SNOMEDCT_CORE|Acute respiratory distress syndrome|Acute respiratory distress syndrome
C0035222|T047|SY|67782005|SNOMEDCT_CORE|Adult hyaline membrane disease|Acute respiratory distress syndrome
C0035222|T047|SY|67782005|SNOMEDCT_CORE|Adult respiratory distress syndrome|Acute respiratory distress syndrome
C0035222|T047|OF|67782005|SNOMEDCT_CORE|Adult respiratory distress syndrome|Acute respiratory distress syndrome
C0035222|T047|IS|67782005|SNOMEDCT_CORE|Adult respiratory distress syndrome, NOS|Acute respiratory distress syndrome
C0035222|T047|IS|67782005|SNOMEDCT_CORE|ARDS|Acute respiratory distress syndrome
C0035222|T047|SY|67782005|SNOMEDCT_CORE|ARDS - Adult respiratory distress syndrome|Acute respiratory distress syndrome
C0035222|T047|SY|67782005|SNOMEDCT_CORE|Congestive atelectasis|Acute respiratory distress syndrome
C0035222|T047|SY|67782005|SNOMEDCT_CORE|DaNang lung|Acute respiratory distress syndrome
C0035222|T047|SY|67782005|SNOMEDCT_CORE|Pulmonary capillary leak syndrome|Acute respiratory distress syndrome
C0035222|T047|SY|67782005|SNOMEDCT_CORE|Shock lung|Acute respiratory distress syndrome
C0035222|T047|SY|67782005|SNOMEDCT_CORE|Vietnam lung|Acute respiratory distress syndrome
C0035229|T046|PT|409623005|SNOMEDCT_CORE|Respiratory insufficiency|Respiratory insufficiency
C0035229|T046|FN|409623005|SNOMEDCT_CORE|Respiratory insufficiency|Respiratory insufficiency
C0035235|T047|PT|55735004|SNOMEDCT_CORE|Respiratory syncytial virus infection|Respiratory syncytial virus infection
C0035235|T047|FN|55735004|SNOMEDCT_CORE|Respiratory syncytial virus infection|Respiratory syncytial virus infection
C0035235|T047|IS|55735004|SNOMEDCT_CORE|Respiratory syncytial virus infection, NOS|Respiratory syncytial virus infection
C0035235|T047|SY|55735004|SNOMEDCT_CORE|RSV - Respiratory syncytial virus infection|Respiratory syncytial virus infection
C0035243|T047|PT|275498002|SNOMEDCT_CORE|Respiratory tract infection|Respiratory tract infection
C0035243|T047|FN|275498002|SNOMEDCT_CORE|Respiratory tract infection|Respiratory tract infection
C0035243|T047|SY|275498002|SNOMEDCT_CORE|RTI - Respiratory tract infection|Respiratory tract infection
C0035258|T047|IS|32914008|SNOMEDCT_CORE|Ekbom syndrome|Restless legs
C0035258|T047|PT|32914008|SNOMEDCT_CORE|Restless legs|Restless legs
C0035258|T047|FN|32914008|SNOMEDCT_CORE|Restless legs|Restless legs
C0035258|T047|SY|32914008|SNOMEDCT_CORE|Restless legs syndrome|Restless legs
C0035258|T047|SY|32914008|SNOMEDCT_CORE|Willis-Ekbom disease|Restless legs
C0035305|T047|SY|42059000|SNOMEDCT_CORE|Detached retina|Retinal detachment
C0035305|T047|SY|42059000|SNOMEDCT_CORE|RD - Retinal detachment|Retinal detachment
C0035305|T047|PT|42059000|SNOMEDCT_CORE|Retinal detachment|Retinal detachment
C0035305|T047|FN|42059000|SNOMEDCT_CORE|Retinal detachment|Retinal detachment
C0035305|T047|IS|42059000|SNOMEDCT_CORE|Retinal detachment, NOS|Retinal detachment
C0035305|T047|SY|42059000|SNOMEDCT_CORE|Sensory retinal detachment|Retinal detachment
C0035309|T047|SY|29555009|SNOMEDCT_CORE|Retinal disease|Retinal disorder
C0035309|T047|IS|29555009|SNOMEDCT_CORE|Retinal disease, NOS|Retinal disorder
C0035309|T047|PT|29555009|SNOMEDCT_CORE|Retinal disorder|Retinal disorder
C0035309|T047|FN|29555009|SNOMEDCT_CORE|Retinal disorder|Retinal disorder
C0035309|T047|IS|29555009|SNOMEDCT_CORE|Retinal disorder, NOS|Retinal disorder
C0035309|T047|OAP|399625000|SNOMEDCT_CORE|Retinopathy|Retinal disorder
C0035309|T047|SY|29555009|SNOMEDCT_CORE|Retinopathy|Retinal disorder
C0035309|T047|OAF|399625000|SNOMEDCT_CORE|Retinopathy|Retinal disorder
C0035312|T047|SY|247153005|SNOMEDCT_CORE|Colloid bodies in retina|Retinal drusen
C0035312|T047|PT|247153005|SNOMEDCT_CORE|Retinal drusen|Retinal drusen
C0035312|T047|FN|247153005|SNOMEDCT_CORE|Retinal drusen|Retinal drusen
C0035317|T047|PTGB|28998008|SNOMEDCT_CORE|Retinal haemorrhage|Retinal hemorrhage
C0035317|T047|SYGB|28998008|SNOMEDCT_CORE|Retinal haemorrhages|Retinal hemorrhage
C0035317|T047|PT|28998008|SNOMEDCT_CORE|Retinal hemorrhage|Retinal hemorrhage
C0035317|T047|FN|28998008|SNOMEDCT_CORE|Retinal hemorrhage|Retinal hemorrhage
C0035317|T047|OF|28998008|SNOMEDCT_CORE|Retinal hemorrhage|Retinal hemorrhage
C0035317|T047|IS|28998008|SNOMEDCT_CORE|Retinal hemorrhage, NOS|Retinal hemorrhage
C0035317|T047|SY|28998008|SNOMEDCT_CORE|Retinal hemorrhages|Retinal hemorrhage
C0035320|T046|SYGB|61267008|SNOMEDCT_CORE|Neovascularisation of retina|Retinal neovascularization
C0035320|T046|SY|61267008|SNOMEDCT_CORE|Neovascularization of retina|Retinal neovascularization
C0035320|T046|PTGB|61267008|SNOMEDCT_CORE|Retinal neovascularisation|Retinal neovascularization
C0035320|T046|PT|61267008|SNOMEDCT_CORE|Retinal neovascularization|Retinal neovascularization
C0035320|T046|FN|61267008|SNOMEDCT_CORE|Retinal neovascularization|Retinal neovascularization
C0035320|T046|IS|61267008|SNOMEDCT_CORE|Retinal neovascularization, NOS|Retinal neovascularization
C0035320|T046|SY|61267008|SNOMEDCT_CORE|Retinal vascular proliferation|Retinal neovascularization
C0035320|T046|SY|61267008|SNOMEDCT_CORE|Vasoproliferative retinopathy|Retinal neovascularization
C0035321|T047|SY|40024006|SNOMEDCT_CORE|Retinal break|Retinal tear
C0035321|T047|IS|40024006|SNOMEDCT_CORE|Retinal break, NOS|Retinal tear
C0035321|T047|IS|40024006|SNOMEDCT_CORE|Retinal tear|Retinal tear
C0035321|T047|PT|95690009|SNOMEDCT_CORE|Retinal tear|Retinal tear
C0035321|T047|FN|95690009|SNOMEDCT_CORE|Retinal tear|Retinal tear
C0035321|T047|IS|95690009|SNOMEDCT_CORE|Retinal tear, NOS|Retinal tear
C0035334|T047|PT|28835009|SNOMEDCT_CORE|Retinitis pigmentosa|Retinitis pigmentosa
C0035334|T047|FN|28835009|SNOMEDCT_CORE|Retinitis pigmentosa|Retinitis pigmentosa
C0035334|T047|SY|28835009|SNOMEDCT_CORE|RP - Retinitis pigmentosa|Retinitis pigmentosa
C0035344|T047|PT|415297005|SNOMEDCT_CORE|Retinopathy of prematurity|Retinopathy of prematurity
C0035344|T047|FN|415297005|SNOMEDCT_CORE|Retinopathy of prematurity|Retinopathy of prematurity
C0035344|T047|SY|415297005|SNOMEDCT_CORE|Retrolental fibroplasia|Retinopathy of prematurity
C0035344|T047|SY|415297005|SNOMEDCT_CORE|RLF - Retrolental fibroplasia|Retinopathy of prematurity
C0035344|T047|IS|415297005|SNOMEDCT_CORE|ROP|Retinopathy of prematurity
C0035344|T047|SY|415297005|SNOMEDCT_CORE|ROP - Retinopathy of prematurity|Retinopathy of prematurity
C0035344|T047|SY|415297005|SNOMEDCT_CORE|Terry's syndrome|Retinopathy of prematurity
C0035357|T046|IS|49120005|SNOMEDCT_CORE|Idiopathic retroperitoneal fibrosis|Retroperitoneal fibrosis
C0035357|T046|SY|49120005|SNOMEDCT_CORE|Ormond's disease|Retroperitoneal fibrosis
C0035357|T046|PT|49120005|SNOMEDCT_CORE|Retroperitoneal fibrosis|Retroperitoneal fibrosis
C0035357|T046|FN|49120005|SNOMEDCT_CORE|Retroperitoneal fibrosis|Retroperitoneal fibrosis
C0035357|T046|SY|49120005|SNOMEDCT_CORE|RPF - Retroperitoneal fibrosis|Retroperitoneal fibrosis
C0035357|T046|SY|49120005|SNOMEDCT_CORE|Sclerosing retroperitonitis|Retroperitoneal fibrosis
C0035358|T191|PT|126872008|SNOMEDCT_CORE|Neoplasm of retroperitoneum|Neoplasm of retroperitoneum
C0035358|T191|FN|126872008|SNOMEDCT_CORE|Neoplasm of retroperitoneum|Neoplasm of retroperitoneum
C0035358|T191|SY|126872008|SNOMEDCT_CORE|Neoplasm of the retroperitoneum|Neoplasm of retroperitoneum
C0035358|T191|OF|126872008|SNOMEDCT_CORE|Neoplasm of the retroperitoneum|Neoplasm of retroperitoneum
C0035358|T191|SY|126872008|SNOMEDCT_CORE|Tumor of retroperitoneum|Neoplasm of retroperitoneum
C0035358|T191|SYGB|126872008|SNOMEDCT_CORE|Tumour of retroperitoneum|Neoplasm of retroperitoneum
C0035410|T046|PT|240131006|SNOMEDCT_CORE|Rhabdomyolysis|Rhabdomyolysis
C0035410|T046|FN|240131006|SNOMEDCT_CORE|Rhabdomyolysis|Rhabdomyolysis
C0035412|T191|PT|302847003|SNOMEDCT_CORE|Rhabdomyosarcoma|Rhabdomyosarcoma
C0035412|T191|FN|302847003|SNOMEDCT_CORE|Rhabdomyosarcoma|Rhabdomyosarcoma
C0035412|T191|SY|302847003|SNOMEDCT_CORE|Rhabdosarcoma|Rhabdomyosarcoma
C0035436|T047|PT|58718002|SNOMEDCT_CORE|Rheumatic fever|Rheumatic fever
C0035436|T047|FN|58718002|SNOMEDCT_CORE|Rheumatic fever|Rheumatic fever
C0035436|T047|IS|58718002|SNOMEDCT_CORE|Rheumatic fever, NOS|Rheumatic fever
C0035436|T047|SY|58718002|SNOMEDCT_CORE|RhF - Rheumatic fever|Rheumatic fever
C0035439|T047|SY|23685000|SNOMEDCT_CORE|Rheumatic carditis|Rheumatic heart disease
C0035439|T047|IS|23685000|SNOMEDCT_CORE|Rheumatic carditis, NOS|Rheumatic heart disease
C0035439|T047|PT|23685000|SNOMEDCT_CORE|Rheumatic heart disease|Rheumatic heart disease
C0035439|T047|FN|23685000|SNOMEDCT_CORE|Rheumatic heart disease|Rheumatic heart disease
C0035439|T047|IS|23685000|SNOMEDCT_CORE|Rheumatic heart disease, NOS|Rheumatic heart disease
C0035439|T047|SY|23685000|SNOMEDCT_CORE|Rheumatic pancarditis|Rheumatic heart disease
C0035455|T047|PT|70076002|SNOMEDCT_CORE|Rhinitis|Rhinitis
C0035455|T047|FN|70076002|SNOMEDCT_CORE|Rhinitis|Rhinitis
C0035455|T047|IS|70076002|SNOMEDCT_CORE|Rhinitis, NOS|Rhinitis
C0035460|T047|PT|8229003|SNOMEDCT_CORE|Vasomotor rhinitis|Vasomotor rhinitis
C0035460|T047|FN|8229003|SNOMEDCT_CORE|Vasomotor rhinitis|Vasomotor rhinitis
C0035460|T047|IS|8229003|SNOMEDCT_CORE|Vasomotor rhinitis, NOS|Vasomotor rhinitis
C0035460|T047|SY|8229003|SNOMEDCT_CORE|VMR - Vasomotor rhinitis|Vasomotor rhinitis
C0035466|T047|SY|19877001|SNOMEDCT_CORE|Hypertrophic rosacea|Rhinophyma
C0035466|T047|PT|19877001|SNOMEDCT_CORE|Rhinophyma|Rhinophyma
C0035466|T047|FN|19877001|SNOMEDCT_CORE|Rhinophyma|Rhinophyma
C0035522|T037|PT|33737001|SNOMEDCT_CORE|Fracture of rib|Fracture of rib
C0035522|T037|FN|33737001|SNOMEDCT_CORE|Fracture of rib|Fracture of rib
C0035522|T037|IS|33737001|SNOMEDCT_CORE|Fracture of rib, NOS|Fracture of rib
C0035522|T037|SY|33737001|SNOMEDCT_CORE|Rib fracture|Fracture of rib
C0035579|T047|PT|41345002|SNOMEDCT_CORE|Rickets|Rickets
C0035579|T047|FN|41345002|SNOMEDCT_CORE|Rickets|Rickets
C0035579|T047|IS|41345002|SNOMEDCT_CORE|Rickets, NOS|Rickets
C0035854|T047|SY|398909004|SNOMEDCT_CORE|Acne erythematosa|Rosacea
C0035854|T047|SY|398909004|SNOMEDCT_CORE|Acne rosacea|Rosacea
C0035854|T047|PT|398909004|SNOMEDCT_CORE|Rosacea|Rosacea
C0035854|T047|FN|398909004|SNOMEDCT_CORE|Rosacea|Rosacea
C0036114|T037|PT|302229004|SNOMEDCT_CORE|Salmonella food poisoning|Salmonella food poisoning
C0036114|T037|FN|302229004|SNOMEDCT_CORE|Salmonella food poisoning|Salmonella food poisoning
C0036114|T037|IS|302229004|SNOMEDCT_CORE|Salmonella gastroenteritis|Salmonella food poisoning
C0036202|T047|SY|31541009|SNOMEDCT_CORE|Benign lymphogranulomatosis of Schaumann|Sarcoidosis
C0036202|T047|SY|31541009|SNOMEDCT_CORE|Besnier-Boeck-Schaumann syndrome|Sarcoidosis
C0036202|T047|SY|31541009|SNOMEDCT_CORE|Boeck's sarcoid|Sarcoidosis
C0036202|T047|SY|31541009|SNOMEDCT_CORE|Boeck's sarcoidosis|Sarcoidosis
C0036202|T047|IS|31541009|SNOMEDCT_CORE|Boecks sarcoidosis|Sarcoidosis
C0036202|T047|SY|31541009|SNOMEDCT_CORE|Darier-Roussy sarcoid|Sarcoidosis
C0036202|T047|SY|31541009|SNOMEDCT_CORE|Lupus pernio of Besnier|Sarcoidosis
C0036202|T047|SY|31541009|SNOMEDCT_CORE|Miliary lupoid of Boeck|Sarcoidosis
C0036202|T047|PT|31541009|SNOMEDCT_CORE|Sarcoidosis|Sarcoidosis
C0036202|T047|FN|31541009|SNOMEDCT_CORE|Sarcoidosis|Sarcoidosis
C0036202|T047|IS|31541009|SNOMEDCT_CORE|Sarcoidosis, NOS|Sarcoidosis
C0036205|T047|PT|24369008|SNOMEDCT_CORE|Pulmonary sarcoidosis|Pulmonary sarcoidosis
C0036205|T047|FN|24369008|SNOMEDCT_CORE|Pulmonary sarcoidosis|Pulmonary sarcoidosis
C0036205|T047|SY|24369008|SNOMEDCT_CORE|Sarcoidosis of lung|Pulmonary sarcoidosis
C0036220|T191|SY|109385007|SNOMEDCT_CORE|Kaposi sarcoma|Kaposi's sarcoma
C0036220|T191|SY|109385007|SNOMEDCT_CORE|Kaposi's sarcoma|Kaposi's sarcoma
C0036220|T191|PT|109385007|SNOMEDCT_CORE|Kaposi's sarcoma|Kaposi's sarcoma
C0036220|T191|FN|109385007|SNOMEDCT_CORE|Kaposi's sarcoma|Kaposi's sarcoma
C0036220|T191|SY|109385007|SNOMEDCT_CORE|KS - Kaposi's sarcoma|Kaposi's sarcoma
C0036262|T047|OF|128869009|SNOMEDCT_CORE|Infestation by Sarcoptes scabiei var hominis|Infestation by Sarcoptes scabiei var hominis
C0036262|T047|PT|128869009|SNOMEDCT_CORE|Infestation by Sarcoptes scabiei var hominis|Infestation by Sarcoptes scabiei var hominis
C0036262|T047|FN|128869009|SNOMEDCT_CORE|Infestation caused by Sarcoptes scabiei var hominis|Infestation by Sarcoptes scabiei var hominis
C0036262|T047|SY|128869009|SNOMEDCT_CORE|Infestation caused by Sarcoptes scabiei var hominis|Infestation by Sarcoptes scabiei var hominis
C0036262|T047|SY|128869009|SNOMEDCT_CORE|Sarcoptic itch|Infestation by Sarcoptes scabiei var hominis
C0036262|T047|SY|128869009|SNOMEDCT_CORE|Scabies|Infestation by Sarcoptes scabiei var hominis
C0036285|T047|SY|30242009|SNOMEDCT_CORE|Scarlatina|Scarlet fever
C0036285|T047|PT|30242009|SNOMEDCT_CORE|Scarlet fever|Scarlet fever
C0036285|T047|FN|30242009|SNOMEDCT_CORE|Scarlet fever|Scarlet fever
C0036337|T048|PT|68890003|SNOMEDCT_CORE|Schizoaffective disorder|Schizoaffective disorder
C0036337|T048|FN|68890003|SNOMEDCT_CORE|Schizoaffective disorder|Schizoaffective disorder
C0036337|T048|IS|68890003|SNOMEDCT_CORE|Schizoaffective disorder, NOS|Schizoaffective disorder
C0036341|T048|PT|58214004|SNOMEDCT_CORE|Schizophrenia|Schizophrenia
C0036341|T048|FN|58214004|SNOMEDCT_CORE|Schizophrenia|Schizophrenia
C0036341|T048|IS|58214004|SNOMEDCT_CORE|Schizophrenia, NOS|Schizophrenia
C0036347|T048|PTGB|35252006|SNOMEDCT_CORE|Disorganised schizophrenia|Disorganized schizophrenia
C0036347|T048|PT|35252006|SNOMEDCT_CORE|Disorganized schizophrenia|Disorganized schizophrenia
C0036347|T048|FN|35252006|SNOMEDCT_CORE|Disorganized schizophrenia|Disorganized schizophrenia
C0036347|T048|IS|35252006|SNOMEDCT_CORE|Disorganized schizophrenia, NOS|Disorganized schizophrenia
C0036347|T048|SY|35252006|SNOMEDCT_CORE|Hebephrenic schizophrenia|Disorganized schizophrenia
C0036349|T048|PT|64905009|SNOMEDCT_CORE|Paranoid schizophrenia|Paranoid schizophrenia
C0036349|T048|FN|64905009|SNOMEDCT_CORE|Paranoid schizophrenia|Paranoid schizophrenia
C0036349|T048|IS|64905009|SNOMEDCT_CORE|Paranoid schizophrenia, NOS|Paranoid schizophrenia
C0036349|T048|SY|64905009|SNOMEDCT_CORE|Paraphrenic schizophrenia|Paranoid schizophrenia
C0036351|T048|PT|26025008|SNOMEDCT_CORE|Residual schizophrenia|Residual schizophrenia
C0036351|T048|FN|26025008|SNOMEDCT_CORE|Residual schizophrenia|Residual schizophrenia
C0036351|T048|IS|26025008|SNOMEDCT_CORE|Residual schizophrenia, NOS|Residual schizophrenia
C0036351|T048|SY|26025008|SNOMEDCT_CORE|Restzustand|Residual schizophrenia
C0036396|T184|SY|23056005|SNOMEDCT_CORE|Neuralgia-neuritis of sciatic nerve|Sciatica
C0036396|T184|SY|23056005|SNOMEDCT_CORE|Sciatic neuralgia|Sciatica
C0036396|T184|PT|23056005|SNOMEDCT_CORE|Sciatica|Sciatica
C0036396|T184|FN|23056005|SNOMEDCT_CORE|Sciatica|Sciatica
C0036396|T184|SY|23056005|SNOMEDCT_CORE|Sciatica neuralgia|Sciatica
C0036416|T047|SY|78370002|SNOMEDCT_CORE|Inflammation of white of eye|Scleritis
C0036416|T047|PT|78370002|SNOMEDCT_CORE|Scleritis|Scleritis
C0036416|T047|FN|78370002|SNOMEDCT_CORE|Scleritis|Scleritis
C0036416|T047|IS|78370002|SNOMEDCT_CORE|Scleritis, NOS|Scleritis
C0036420|T047|SY|201048007|SNOMEDCT_CORE|Addison's keloid|Localized scleroderma
C0036420|T047|SY|201048007|SNOMEDCT_CORE|Circumscribed scleroderma|Localized scleroderma
C0036420|T047|SYGB|201048007|SNOMEDCT_CORE|Localised dermatosclerosis|Localized scleroderma
C0036420|T047|SYGB|201048007|SNOMEDCT_CORE|Localised morphoea|Localized scleroderma
C0036420|T047|PTGB|201048007|SNOMEDCT_CORE|Localised scleroderma|Localized scleroderma
C0036420|T047|SY|201048007|SNOMEDCT_CORE|Localized dermatosclerosis|Localized scleroderma
C0036420|T047|SY|201048007|SNOMEDCT_CORE|Localized morphea|Localized scleroderma
C0036420|T047|FN|201048007|SNOMEDCT_CORE|Localized morphea|Localized scleroderma
C0036420|T047|PT|201048007|SNOMEDCT_CORE|Localized scleroderma|Localized scleroderma
C0036420|T047|SY|201048007|SNOMEDCT_CORE|Morphea scleroderma|Localized scleroderma
C0036420|T047|SYGB|201048007|SNOMEDCT_CORE|Morphoea scleroderma|Localized scleroderma
C0036421|T047|IS|89155008|SNOMEDCT_CORE|Progressive systemic sclerosis|Systemic sclerosis
C0036421|T047|IS|89155008|SNOMEDCT_CORE|PSS - Progressive systemic sclerosis|Systemic sclerosis
C0036421|T047|SY|89155008|SNOMEDCT_CORE|Scleroderma syndrome|Systemic sclerosis
C0036421|T047|SY|89155008|SNOMEDCT_CORE|SS - Systemic sclerosis|Systemic sclerosis
C0036421|T047|SY|89155008|SNOMEDCT_CORE|Systemic scleroderma|Systemic sclerosis
C0036421|T047|PT|89155008|SNOMEDCT_CORE|Systemic sclerosis|Systemic sclerosis
C0036421|T047|FN|89155008|SNOMEDCT_CORE|Systemic sclerosis|Systemic sclerosis
C0036439|T047|SY|298382003|SNOMEDCT_CORE|Scoliosis|Scoliosis deformity of spine
C0036439|T047|PT|298382003|SNOMEDCT_CORE|Scoliosis deformity of spine|Scoliosis deformity of spine
C0036439|T047|OF|298382003|SNOMEDCT_CORE|Scoliosis deformity of spine|Scoliosis deformity of spine
C0036439|T047|FN|298382003|SNOMEDCT_CORE|Scoliosis deformity of spine|Scoliosis deformity of spine
C0036440|T190|IS|30611007|SNOMEDCT_CORE|Idiopathic scoliosis and kyphoscoliosis|Idiopathic scoliosis AND/OR kyphoscoliosis
C0036440|T190|FN|30611007|SNOMEDCT_CORE|Idiopathic scoliosis AND/OR kyphoscoliosis|Idiopathic scoliosis AND/OR kyphoscoliosis
C0036440|T190|PT|30611007|SNOMEDCT_CORE|Idiopathic scoliosis AND/OR kyphoscoliosis|Idiopathic scoliosis AND/OR kyphoscoliosis
C0036454|T033|IS|23388006|SNOMEDCT_CORE|Scotoma|Visual field scotoma
C0036454|T033|IS|23388006|SNOMEDCT_CORE|Scotoma, NOS|Visual field scotoma
C0036454|T033|PT|23388006|SNOMEDCT_CORE|Visual field scotoma|Visual field scotoma
C0036454|T033|FN|23388006|SNOMEDCT_CORE|Visual field scotoma|Visual field scotoma
C0036467|T047|PT|54084005|SNOMEDCT_CORE|Cervical tuberculous lymphadenitis|Cervical tuberculous lymphadenitis
C0036467|T047|FN|54084005|SNOMEDCT_CORE|Cervical tuberculous lymphadenitis|Cervical tuberculous lymphadenitis
C0036467|T047|SY|54084005|SNOMEDCT_CORE|Scrofula|Cervical tuberculous lymphadenitis
C0036467|T047|SY|54084005|SNOMEDCT_CORE|Tuberculosis of cervical lymph nodes|Cervical tuberculous lymphadenitis
C0036467|T047|SY|54084005|SNOMEDCT_CORE|Tuberculous cervical lymphadenitis|Cervical tuberculous lymphadenitis
C0036508|T047|SY|50563003|SNOMEDCT_CORE|SBD - Seborrheic dermatitis|Seborrheic dermatitis
C0036508|T047|SYGB|50563003|SNOMEDCT_CORE|SBD - Seborrhoeic dermatitis|Seborrheic dermatitis
C0036508|T047|PT|86708008|SNOMEDCT_CORE|Seborrhea|Seborrheic dermatitis
C0036508|T047|FN|86708008|SNOMEDCT_CORE|Seborrhea|Seborrheic dermatitis
C0036508|T047|IS|86708008|SNOMEDCT_CORE|Seborrhea, NOS|Seborrheic dermatitis
C0036508|T047|PT|50563003|SNOMEDCT_CORE|Seborrheic dermatitis|Seborrheic dermatitis
C0036508|T047|FN|50563003|SNOMEDCT_CORE|Seborrheic dermatitis|Seborrheic dermatitis
C0036508|T047|SY|50563003|SNOMEDCT_CORE|Seborrheic eczema|Seborrheic dermatitis
C0036508|T047|PTGB|86708008|SNOMEDCT_CORE|Seborrhoea|Seborrheic dermatitis
C0036508|T047|IS|86708008|SNOMEDCT_CORE|Seborrhoea, NOS|Seborrheic dermatitis
C0036508|T047|PTGB|50563003|SNOMEDCT_CORE|Seborrhoeic dermatitis|Seborrheic dermatitis
C0036508|T047|SYGB|50563003|SNOMEDCT_CORE|Seborrhoeic eczema|Seborrheic dermatitis
C0036529|T047|OAP|89600009|SNOMEDCT_CORE|Secondary cardiomyopathy|Secondary cardiomyopathy
C0036529|T047|OAF|89600009|SNOMEDCT_CORE|Secondary cardiomyopathy|Secondary cardiomyopathy
C0036529|T047|IS|89600009|SNOMEDCT_CORE|Secondary cardiomyopathy, NOS|Secondary cardiomyopathy, NOS
C0036550|T048|SY|64386003|SNOMEDCT_CORE|Sedative, hypnotic AND/OR anxiolytic abuse|Sedative, hypnotic AND/OR anxiolytic abuse
C0036550|T048|IS|64386003|SNOMEDCT_CORE|Sedative, hypnotic or anxiolytic abuse|Sedative, hypnotic AND/OR anxiolytic abuse
C0036572|T184|SY|91175000|SNOMEDCT_CORE|Convulsion|Seizure
C0036572|T184|IS|91175000|SNOMEDCT_CORE|Convulsion, NOS|Seizure
C0036572|T184|IS|91175000|SNOMEDCT_CORE|Convulsions|Seizure
C0036572|T184|SY|91175000|SNOMEDCT_CORE|Fit|Seizure
C0036572|T184|SY|91175000|SNOMEDCT_CORE|Fit - convulsion|Seizure
C0036572|T184|IS|91175000|SNOMEDCT_CORE|Fit, NOS|Seizure
C0036572|T184|IS|91175000|SNOMEDCT_CORE|Fits - convulsions|Seizure
C0036572|T184|SY|91175000|SNOMEDCT_CORE|Fitting|Seizure
C0036572|T184|PT|91175000|SNOMEDCT_CORE|Seizure|Seizure
C0036572|T184|FN|91175000|SNOMEDCT_CORE|Seizure|Seizure
C0036572|T184|IS|91175000|SNOMEDCT_CORE|Seizure, NOS|Seizure
C0036631|T191|PT|443675005|SNOMEDCT_CORE|Seminoma|Seminoma
C0036631|T191|PT|36741007|SNOMEDCT_CORE|Seminoma|Seminoma
C0036631|T191|OF|36741007|SNOMEDCT_CORE|Seminoma|Seminoma
C0036631|T191|FN|443675005|SNOMEDCT_CORE|Seminoma|Seminoma
C0036631|T191|OF|36741007|SNOMEDCT_CORE|Seminoma, no ICD-O subtype|Seminoma
C0036631|T191|SY|36741007|SNOMEDCT_CORE|Seminoma, no ICD-O subtype|Seminoma
C0036631|T191|SY|36741007|SNOMEDCT_CORE|Seminoma, no International Classification of Diseases for Oncology subtype|Seminoma
C0036631|T191|FN|36741007|SNOMEDCT_CORE|Seminoma, no International Classification of Diseases for Oncology subtype|Seminoma
C0036631|T191|IS|36741007|SNOMEDCT_CORE|Seminoma, NOS|Seminoma
C0036646|T020|OP|39450006|SNOMEDCT_CORE|Age-related cataract|Senile cataract
C0036646|T020|OF|39450006|SNOMEDCT_CORE|Age-related cataract|Senile cataract
C0036646|T020|SY|39450006|SNOMEDCT_CORE|Old-age related cataract|Senile cataract
C0036646|T020|PT|39450006|SNOMEDCT_CORE|Senile cataract|Senile cataract
C0036646|T020|FN|39450006|SNOMEDCT_CORE|Senile cataract|Senile cataract
C0036646|T020|IS|39450006|SNOMEDCT_CORE|Senile cataract, NOS|Senile cataract
C0036651|T047|SY|72100002|SNOMEDCT_CORE|Actinic lentigo|Solar lentigo
C0036651|T047|SY|72100002|SNOMEDCT_CORE|Liver spot|Solar lentigo
C0036651|T047|SY|72100002|SNOMEDCT_CORE|Senile lentigo|Solar lentigo
C0036651|T047|OF|72100002|SNOMEDCT_CORE|Senile lentigo|Solar lentigo
C0036651|T047|PT|72100002|SNOMEDCT_CORE|Solar lentigo|Solar lentigo
C0036651|T047|FN|72100002|SNOMEDCT_CORE|Solar lentigo|Solar lentigo
C0036685|T047|IS|53869006|SNOMEDCT_CORE|Gram negative sepsis|Gram negative sepsis
C0036685|T047|OAP|53869006|SNOMEDCT_CORE|Gram negative septicaemia|Gram negative septicaemia
C0036685|T047|OAP|53869006|SNOMEDCT_CORE|Gram negative septicemia|Gram negative septicemia
C0036685|T047|OAF|53869006|SNOMEDCT_CORE|Gram negative septicemia|Gram negative septicemia
C0036685|T047|OAS|53869006|SNOMEDCT_CORE|Gram-negative septicaemia|Gram-negative septicaemia
C0036685|T047|OAS|53869006|SNOMEDCT_CORE|Gram-negative septicemia|Gram-negative septicemia
C0036689|T047|SY|43878008|SNOMEDCT_CORE|Septic sore throat|Streptococcal sore throat
C0036689|T047|SY|43878008|SNOMEDCT_CORE|Strep throat|Streptococcal sore throat
C0036689|T047|SY|43878008|SNOMEDCT_CORE|Strept throat|Streptococcal sore throat
C0036689|T047|SY|43878008|SNOMEDCT_CORE|Streptococcal angina|Streptococcal sore throat
C0036689|T047|SY|43878008|SNOMEDCT_CORE|Streptococcal pharyngitis|Streptococcal sore throat
C0036689|T047|PT|43878008|SNOMEDCT_CORE|Streptococcal sore throat|Streptococcal sore throat
C0036689|T047|FN|43878008|SNOMEDCT_CORE|Streptococcal sore throat|Streptococcal sore throat
C0036690|T047|OAP|105592009|SNOMEDCT_CORE|Septicaemia|Septicemia
C0036690|T047|IS|91302008|SNOMEDCT_CORE|Septicaemia, NOS|Septicemia
C0036690|T047|OAP|105592009|SNOMEDCT_CORE|Septicemia|Septicemia
C0036690|T047|OAF|105592009|SNOMEDCT_CORE|Septicemia|Septicemia
C0036690|T047|IS|91302008|SNOMEDCT_CORE|Septicemia, NOS|Septicemia
C0036857|T048|SY|40700009|SNOMEDCT_CORE|Severe intellectual development disorder|Severe intellectual disability
C0036857|T048|PT|40700009|SNOMEDCT_CORE|Severe intellectual disability|Severe intellectual disability
C0036857|T048|FN|40700009|SNOMEDCT_CORE|Severe intellectual disability|Severe intellectual disability
C0036857|T048|SY|40700009|SNOMEDCT_CORE|Severe mental handicap|Severe intellectual disability
C0036916|T047|SY|8098009|SNOMEDCT_CORE|Disease with a predominantly sexual mode of transmission|Sexually transmitted infectious disease
C0036916|T047|SY|8098009|SNOMEDCT_CORE|Sexually transmissible disease|Sexually transmitted infectious disease
C0036916|T047|SY|8098009|SNOMEDCT_CORE|Sexually transmitted disease|Sexually transmitted infectious disease
C0036916|T047|IS|8098009|SNOMEDCT_CORE|Sexually transmitted disease, NOS|Sexually transmitted infectious disease
C0036916|T047|PT|8098009|SNOMEDCT_CORE|Sexually transmitted infectious disease|Sexually transmitted infectious disease
C0036916|T047|FN|8098009|SNOMEDCT_CORE|Sexually transmitted infectious disease|Sexually transmitted infectious disease
C0036916|T047|IS|8098009|SNOMEDCT_CORE|Sexually transmitted infectious disease, NOS|Sexually transmitted infectious disease
C0036916|T047|SY|8098009|SNOMEDCT_CORE|Statutory venereal disease|Sexually transmitted infectious disease
C0036916|T047|SY|8098009|SNOMEDCT_CORE|STD - sexually transmitted disease|Sexually transmitted infectious disease
C0036916|T047|IS|8098009|SNOMEDCT_CORE|STD - Sexually transmitted disease|Sexually transmitted infectious disease
C0036916|T047|SY|8098009|SNOMEDCT_CORE|STI - sexually transmitted infection|Sexually transmitted infectious disease
C0036916|T047|SY|8098009|SNOMEDCT_CORE|VD - venereal disease|Sexually transmitted infectious disease
C0036916|T047|IS|8098009|SNOMEDCT_CORE|VD - Venereal disease|Sexually transmitted infectious disease
C0036916|T047|SY|8098009|SNOMEDCT_CORE|Venereal disease|Sexually transmitted infectious disease
C0036916|T047|IS|8098009|SNOMEDCT_CORE|Venereal disease, NOS|Sexually transmitted infectious disease
C0036973|T033|SY|43724002|SNOMEDCT_CORE|Shivering|Shivering
C0036974|T046|SY|27942005|SNOMEDCT_CORE|Acute circulatory failure|Shock
C0036974|T046|SY|27942005|SNOMEDCT_CORE|Circulatory collapse|Shock
C0036974|T046|SY|27942005|SNOMEDCT_CORE|Peripheral circulatory failure|Shock
C0036974|T046|SY|27942005|SNOMEDCT_CORE|Peripheral vascular failure|Shock
C0036974|T046|SY|27942005|SNOMEDCT_CORE|Peripheral vascular shutdown|Shock
C0036974|T046|PT|27942005|SNOMEDCT_CORE|Shock|Shock
C0036974|T046|FN|27942005|SNOMEDCT_CORE|Shock|Shock
C0036974|T046|SY|27942005|SNOMEDCT_CORE|Shock - physiological|Shock
C0036974|T046|IS|27942005|SNOMEDCT_CORE|Shock, NOS|Shock
C0036980|T046|PT|89138009|SNOMEDCT_CORE|Cardiogenic shock|Cardiogenic shock
C0036980|T046|FN|89138009|SNOMEDCT_CORE|Cardiogenic shock|Cardiogenic shock
C0036983|T046|SY|76571007|SNOMEDCT_CORE|Sepsis-associated hypotension|Septic shock
C0036983|T046|PT|76571007|SNOMEDCT_CORE|Septic shock|Septic shock
C0036983|T046|FN|76571007|SNOMEDCT_CORE|Septic shock|Septic shock
C0036983|T046|SYGB|76571007|SNOMEDCT_CORE|Septicaemic shock|Septic shock
C0036983|T046|SY|76571007|SNOMEDCT_CORE|Septicemic shock|Septic shock
C0036992|T047|IS|26629001|SNOMEDCT_CORE|Acquired short bowel syndrome|Short bowel syndrome
C0036992|T047|IS|26629001|SNOMEDCT_CORE|Post-resection malabsorption|Short bowel syndrome
C0036992|T047|IS|26629001|SNOMEDCT_CORE|Postresectional malabsorption syndrome|Short bowel syndrome
C0036992|T047|SY|26629001|SNOMEDCT_CORE|SBS - Short bowel syndrome|Short bowel syndrome
C0036992|T047|SY|26629001|SNOMEDCT_CORE|SGS - Short gut syndrome|Short bowel syndrome
C0036992|T047|PT|26629001|SNOMEDCT_CORE|Short bowel syndrome|Short bowel syndrome
C0036992|T047|FN|26629001|SNOMEDCT_CORE|Short bowel syndrome|Short bowel syndrome
C0036992|T047|SY|26629001|SNOMEDCT_CORE|Short gut syndrome|Short bowel syndrome
C0036992|T047|SY|26629001|SNOMEDCT_CORE|Short intestine syndrome|Short bowel syndrome
C0037005|T037|SY|417076003|SNOMEDCT_CORE|Dislocation of glenohumeral joint|Dislocation of shoulder joint
C0037005|T037|SY|417076003|SNOMEDCT_CORE|Dislocation of shoulder|Dislocation of shoulder joint
C0037005|T037|PT|417076003|SNOMEDCT_CORE|Dislocation of shoulder joint|Dislocation of shoulder joint
C0037005|T037|FN|417076003|SNOMEDCT_CORE|Dislocation of shoulder joint|Dislocation of shoulder joint
C0037005|T037|SY|417076003|SNOMEDCT_CORE|Shoulder dislocation|Dislocation of shoulder joint
C0037011|T184|IS|45326000|SNOMEDCT_CORE|Pain in shoulder|Shoulder pain
C0037011|T184|PT|45326000|SNOMEDCT_CORE|Shoulder pain|Shoulder pain
C0037011|T184|FN|45326000|SNOMEDCT_CORE|Shoulder pain|Shoulder pain
C0037011|T184|SY|45326000|SNOMEDCT_CORE|Shoulder region pain|Shoulder pain
C0037023|T047|SY|42982001|SNOMEDCT_CORE|Sialadenitis|Sialoadenitis
C0037023|T047|IS|42982001|SNOMEDCT_CORE|Sialadenitis, NOS|Sialoadenitis
C0037023|T047|PT|42982001|SNOMEDCT_CORE|Sialoadenitis|Sialoadenitis
C0037023|T047|FN|42982001|SNOMEDCT_CORE|Sialoadenitis|Sialoadenitis
C0037023|T047|IS|42982001|SNOMEDCT_CORE|Sialoadenitis, NOS|Sialoadenitis
C0037052|T047|PT|36083008|SNOMEDCT_CORE|Sick sinus syndrome|Sick sinus syndrome
C0037052|T047|FN|36083008|SNOMEDCT_CORE|Sick sinus syndrome|Sick sinus syndrome
C0037054|T047|SY|16402000|SNOMEDCT_CORE|AS - Sickle cell trait|Sickle cell trait
C0037054|T047|SY|16402000|SNOMEDCT_CORE|Drepanocytosis|Sickle cell trait
C0037054|T047|SYGB|16402000|SNOMEDCT_CORE|Haemoglobin A-S genotype|Sickle cell trait
C0037054|T047|SYGB|16402000|SNOMEDCT_CORE|Haemoglobin S trait|Sickle cell trait
C0037054|T047|SYGB|16402000|SNOMEDCT_CORE|Haemoglobin S-A disorder|Sickle cell trait
C0037054|T047|SY|16402000|SNOMEDCT_CORE|Hemoglobin A-S genotype|Sickle cell trait
C0037054|T047|SY|16402000|SNOMEDCT_CORE|Hemoglobin S trait|Sickle cell trait
C0037054|T047|SY|16402000|SNOMEDCT_CORE|Hemoglobin S-A disorder|Sickle cell trait
C0037054|T047|SY|16402000|SNOMEDCT_CORE|Heterozygous for Hb S|Sickle cell trait
C0037054|T047|SYGB|16402000|SNOMEDCT_CORE|Heterozygous haemoglobin S|Sickle cell trait
C0037054|T047|SY|16402000|SNOMEDCT_CORE|Heterozygous hemoglobin S|Sickle cell trait
C0037054|T047|SY|16402000|SNOMEDCT_CORE|RBC's - sickle cells present|Sickle cell trait
C0037054|T047|PT|16402000|SNOMEDCT_CORE|Sickle cell trait|Sickle cell trait
C0037054|T047|FN|16402000|SNOMEDCT_CORE|Sickle cell trait|Sickle cell trait
C0037054|T047|SY|16402000|SNOMEDCT_CORE|Sickle cells present|Sickle cell trait
C0037116|T047|SY|805002|SNOMEDCT_CORE|Nodular silicosis|Pneumoconiosis due to silica
C0037116|T047|SY|805002|SNOMEDCT_CORE|Pneumoconiosis caused by silica|Pneumoconiosis due to silica
C0037116|T047|FN|805002|SNOMEDCT_CORE|Pneumoconiosis caused by silica|Pneumoconiosis due to silica
C0037116|T047|PT|805002|SNOMEDCT_CORE|Pneumoconiosis due to silica|Pneumoconiosis due to silica
C0037116|T047|OF|805002|SNOMEDCT_CORE|Pneumoconiosis due to silica|Pneumoconiosis due to silica
C0037116|T047|IS|805002|SNOMEDCT_CORE|Pneumoconiosis due to silica, NOS|Pneumoconiosis due to silica
C0037116|T047|SY|805002|SNOMEDCT_CORE|Silicatosis|Pneumoconiosis due to silica
C0037116|T047|SY|805002|SNOMEDCT_CORE|Silicosis|Pneumoconiosis due to silica
C0037116|T047|IS|805002|SNOMEDCT_CORE|Silicosis, NOS|Pneumoconiosis due to silica
C0037195|T033|PT|4969004|SNOMEDCT_CORE|Sinus headache|Sinus headache
C0037195|T033|FN|4969004|SNOMEDCT_CORE|Sinus headache|Sinus headache
C0037199|T047|PT|36971009|SNOMEDCT_CORE|Sinusitis|Sinusitis
C0037199|T047|FN|36971009|SNOMEDCT_CORE|Sinusitis|Sinusitis
C0037199|T047|IS|36971009|SNOMEDCT_CORE|Sinusitis, NOS|Sinusitis
C0037268|T019|PT|199879009|SNOMEDCT_CORE|Congenital anomaly of skin|Congenital anomaly of skin
C0037268|T019|FN|199879009|SNOMEDCT_CORE|Congenital anomaly of skin|Congenital anomaly of skin
C0037268|T019|IS|199879009|SNOMEDCT_CORE|Congenital anomaly of skin, NOS|Congenital anomaly of skin
C0037268|T019|SY|199879009|SNOMEDCT_CORE|Congenital cutaneous anomaly|Congenital anomaly of skin
C0037268|T019|IS|199879009|SNOMEDCT_CORE|Congenital cutaneous anomaly, NOS|Congenital anomaly of skin
C0037268|T019|SY|199879009|SNOMEDCT_CORE|Congenital malformation of the skin|Congenital anomaly of skin
C0037268|T019|SY|199879009|SNOMEDCT_CORE|Congenital skin anomalies|Congenital anomaly of skin
C0037274|T047|SY|95320005|SNOMEDCT_CORE|Dermatological disease|Disorder of skin
C0037274|T047|SY|95320005|SNOMEDCT_CORE|Dermatological disorder|Disorder of skin
C0037274|T047|SY|95320005|SNOMEDCT_CORE|Dermatopathy|Disorder of skin
C0037274|T047|SY|95320005|SNOMEDCT_CORE|Dermatosis|Disorder of skin
C0037274|T047|IS|95320005|SNOMEDCT_CORE|Dermatosis, NOS|Disorder of skin
C0037274|T047|IS|80659006|SNOMEDCT_CORE|Dermatosis, NOS|Disorder of skin
C0037274|T047|IS|95320005|SNOMEDCT_CORE|Disease of skin|Disorder of skin
C0037274|T047|OF|95320005|SNOMEDCT_CORE|Disease of skin|Disorder of skin
C0037274|T047|IS|95320005|SNOMEDCT_CORE|Disease of skin, NOS|Disorder of skin
C0037274|T047|PT|95320005|SNOMEDCT_CORE|Disorder of skin|Disorder of skin
C0037274|T047|FN|95320005|SNOMEDCT_CORE|Disorder of skin|Disorder of skin
C0037274|T047|SY|95320005|SNOMEDCT_CORE|Skin disease|Disorder of skin
C0037274|T047|SY|95320005|SNOMEDCT_CORE|Skin disorder|Disorder of skin
C0037274|T047|IS|95320005|SNOMEDCT_CORE|Skin disorder, NOS|Disorder of skin
C0037277|T047|IS|199879009|SNOMEDCT_CORE|Genodermatosis, NOS|Genodermatosis, NOS
C0037278|T047|PT|108365000|SNOMEDCT_CORE|Infection of skin|Infection of skin
C0037278|T047|FN|108365000|SNOMEDCT_CORE|Infection of skin|Infection of skin
C0037284|T047|PT|95324001|SNOMEDCT_CORE|Skin lesion|Skin lesion
C0037284|T047|FN|95324001|SNOMEDCT_CORE|Skin lesion|Skin lesion
C0037284|T047|IS|95324001|SNOMEDCT_CORE|Skin lesion, NOS|Skin lesion
C0037286|T191|SY|126488004|SNOMEDCT_CORE|Cutaneous tumor|Neoplasm of skin
C0037286|T191|SYGB|126488004|SNOMEDCT_CORE|Cutaneous tumour|Neoplasm of skin
C0037286|T191|PT|126488004|SNOMEDCT_CORE|Neoplasm of skin|Neoplasm of skin
C0037286|T191|FN|126488004|SNOMEDCT_CORE|Neoplasm of skin|Neoplasm of skin
C0037286|T191|SY|126488004|SNOMEDCT_CORE|Skin tumor|Neoplasm of skin
C0037286|T191|SYGB|126488004|SNOMEDCT_CORE|Skin tumour|Neoplasm of skin
C0037286|T191|SY|126488004|SNOMEDCT_CORE|Tumor of skin|Neoplasm of skin
C0037286|T191|SYGB|126488004|SNOMEDCT_CORE|Tumour of skin|Neoplasm of skin
C0037287|T046|SY|95319004|SNOMEDCT_CORE|Cutaneous nodule|Skin nodule
C0037287|T046|SY|95319004|SNOMEDCT_CORE|Nodule of skin|Skin nodule
C0037287|T046|PT|95319004|SNOMEDCT_CORE|Skin nodule|Skin nodule
C0037287|T046|FN|95319004|SNOMEDCT_CORE|Skin nodule|Skin nodule
C0037287|T046|OF|95319004|SNOMEDCT_CORE|Skin nodule|Skin nodule
C0037293|T191|SY|201091002|SNOMEDCT_CORE|Achrochordon|Skin tag
C0037293|T191|PT|201091002|SNOMEDCT_CORE|Skin tag|Skin tag
C0037293|T191|FN|201091002|SNOMEDCT_CORE|Skin tag|Skin tag
C0037293|T191|SY|201091002|SNOMEDCT_CORE|SKT - Skin tag|Skin tag
C0037293|T191|SY|201091002|SNOMEDCT_CORE|Soft fibroma|Skin tag
C0037293|T191|SY|201091002|SNOMEDCT_CORE|Soft papilloma|Skin tag
C0037299|T047|SY|46742003|SNOMEDCT_CORE|Cutaneous ulcer|Skin ulcer
C0037299|T047|PT|46742003|SNOMEDCT_CORE|Skin ulcer|Skin ulcer
C0037299|T047|FN|46742003|SNOMEDCT_CORE|Skin ulcer|Skin ulcer
C0037299|T047|IS|46742003|SNOMEDCT_CORE|Ulcer of skin|Skin ulcer
C0037299|T047|IS|46742003|SNOMEDCT_CORE|Ulcer of skin, NOS|Skin ulcer
C0037301|T033|SY|247434009|SNOMEDCT_CORE|Rugosity of skin|Wrinkled skin
C0037301|T033|PT|247434009|SNOMEDCT_CORE|Wrinkled skin|Wrinkled skin
C0037301|T033|FN|247434009|SNOMEDCT_CORE|Wrinkled skin|Wrinkled skin
C0037304|T037|PT|71642004|SNOMEDCT_CORE|Fracture of skull|Fracture of skull
C0037304|T037|FN|71642004|SNOMEDCT_CORE|Fracture of skull|Fracture of skull
C0037304|T037|IS|71642004|SNOMEDCT_CORE|Fracture of skull, NOS|Fracture of skull
C0037304|T037|SY|71642004|SNOMEDCT_CORE|Fractured skull|Fracture of skull
C0037315|T047|SY|73430006|SNOMEDCT_CORE|SAS - Sleep apnea syndrome|Sleep apnea
C0037315|T047|SYGB|73430006|SNOMEDCT_CORE|SAS - Sleep apnoea syndrome|Sleep apnea
C0037315|T047|PT|73430006|SNOMEDCT_CORE|Sleep apnea|Sleep apnea
C0037315|T047|OF|73430006|SNOMEDCT_CORE|Sleep apnea|Sleep apnea
C0037315|T047|FN|73430006|SNOMEDCT_CORE|Sleep apnea|Sleep apnea
C0037315|T047|SY|73430006|SNOMEDCT_CORE|Sleep apnea syndrome|Sleep apnea
C0037315|T047|IS|73430006|SNOMEDCT_CORE|Sleep apnea, NOS|Sleep apnea
C0037315|T047|PTGB|73430006|SNOMEDCT_CORE|Sleep apnoea|Sleep apnea
C0037315|T047|SYGB|73430006|SNOMEDCT_CORE|Sleep apnoea syndrome|Sleep apnea
C0037315|T047|SY|73430006|SNOMEDCT_CORE|Sleep hypopnea|Sleep apnea
C0037315|T047|SYGB|73430006|SNOMEDCT_CORE|Sleep hypopnoea|Sleep apnea
C0037317|T184|PT|53888004|SNOMEDCT_CORE|Disturbance in sleep behavior|Disturbance in sleep behavior
C0037317|T184|FN|53888004|SNOMEDCT_CORE|Disturbance in sleep behavior|Disturbance in sleep behavior
C0037317|T184|IS|53888004|SNOMEDCT_CORE|Disturbance in sleep behavior, NOS|Disturbance in sleep behavior
C0037317|T184|PTGB|53888004|SNOMEDCT_CORE|Disturbance in sleep behaviour|Disturbance in sleep behavior
C0037320|T048|SY|89675003|SNOMEDCT_CORE|Night terrors|Sleep terror disorder
C0037320|T048|PT|89675003|SNOMEDCT_CORE|Sleep terror disorder|Sleep terror disorder
C0037320|T048|FN|89675003|SNOMEDCT_CORE|Sleep terror disorder|Sleep terror disorder
C0037320|T048|SY|89675003|SNOMEDCT_CORE|Sleep terrors|Sleep terror disorder
C0037367|T037|PT|426936004|SNOMEDCT_CORE|Smoke inhalation injury|Smoke inhalation injury
C0037367|T037|FN|426936004|SNOMEDCT_CORE|Smoke inhalation injury|Smoke inhalation injury
C0037384|T184|SY|72863001|SNOMEDCT_CORE|Finding of snoring|Snoring
C0037384|T184|SY|72863001|SNOMEDCT_CORE|Observation of snoring|Snoring
C0037384|T184|SY|72863001|SNOMEDCT_CORE|Snores|Snoring
C0037384|T184|PT|72863001|SNOMEDCT_CORE|Snoring|Snoring
C0037384|T184|FN|72863001|SNOMEDCT_CORE|Snoring|Snoring
C0037578|T037|PT|282026002|SNOMEDCT_CORE|Soft tissue injury|Soft tissue injury
C0037578|T037|FN|282026002|SNOMEDCT_CORE|Soft tissue injury|Soft tissue injury
C0037578|T037|SY|282026002|SNOMEDCT_CORE|STI - Soft tissue injury|Soft tissue injury
C0037580|T047|PT|298349001|SNOMEDCT_CORE|Soft tissue swelling|Soft tissue swelling
C0037580|T047|FN|298349001|SNOMEDCT_CORE|Soft tissue swelling|Soft tissue swelling
C0037672|T047|SY|80495009|SNOMEDCT_CORE|Sleep walking|Sleep walking disorder
C0037672|T047|PT|80495009|SNOMEDCT_CORE|Sleep walking disorder|Sleep walking disorder
C0037672|T047|FN|80495009|SNOMEDCT_CORE|Sleep walking disorder|Sleep walking disorder
C0037672|T047|SY|80495009|SNOMEDCT_CORE|Sleepwalking|Sleep walking disorder
C0037672|T047|SY|80495009|SNOMEDCT_CORE|Sleepwalking disorder|Sleep walking disorder
C0037672|T047|SY|80495009|SNOMEDCT_CORE|Somnambulism|Sleep walking disorder
C0037672|T047|IS|80495009|SNOMEDCT_CORE|Somnanbulism|Sleep walking disorder
C0037763|T184|PT|45352006|SNOMEDCT_CORE|Spasm|Spasm
C0037763|T184|FN|45352006|SNOMEDCT_CORE|Spasm|Spasm
C0037763|T184|IS|45352006|SNOMEDCT_CORE|Spasm, NOS|Spasm
C0037771|T184|PT|312444006|SNOMEDCT_CORE|Spastic paraparesis|Spastic paraparesis
C0037771|T184|FN|312444006|SNOMEDCT_CORE|Spastic paraparesis|Spastic paraparesis
C0037856|T047|PT|49198006|SNOMEDCT_CORE|Torsion of spermatic cord|Torsion of spermatic cord
C0037856|T047|FN|49198006|SNOMEDCT_CORE|Torsion of spermatic cord|Torsion of spermatic cord
C0037859|T047|PT|49263001|SNOMEDCT_CORE|Spermatocele|Spermatocele
C0037859|T047|FN|49263001|SNOMEDCT_CORE|Spermatocele|Spermatocele
C0037926|T047|SY|71286001|SNOMEDCT_CORE|Compression of spinal cord|Spinal cord compression
C0037926|T047|IS|71286001|SNOMEDCT_CORE|Cord compression, NOS|Spinal cord compression
C0037926|T047|SY|71286001|SNOMEDCT_CORE|SCC - Spinal cord compression|Spinal cord compression
C0037926|T047|PT|71286001|SNOMEDCT_CORE|Spinal cord compression|Spinal cord compression
C0037926|T047|FN|71286001|SNOMEDCT_CORE|Spinal cord compression|Spinal cord compression
C0037926|T047|IS|71286001|SNOMEDCT_CORE|Spinal cord compression, NOS|Spinal cord compression
C0037928|T047|IS|48522003|SNOMEDCT_CORE|Disease of spinal cord|Spinal cord disease
C0037928|T047|IS|48522003|SNOMEDCT_CORE|Disease of spinal cord, NOS|Spinal cord disease
C0037928|T047|SY|48522003|SNOMEDCT_CORE|MP - Myelopathy|Spinal cord disease
C0037928|T047|SY|48522003|SNOMEDCT_CORE|Myelopathy|Spinal cord disease
C0037928|T047|OF|48522003|SNOMEDCT_CORE|Myelopathy|Spinal cord disease
C0037928|T047|IS|48522003|SNOMEDCT_CORE|Myelopathy, NOS|Spinal cord disease
C0037928|T047|SY|48522003|SNOMEDCT_CORE|Neurologic myelopathy|Spinal cord disease
C0037928|T047|PT|48522003|SNOMEDCT_CORE|Spinal cord disease|Spinal cord disease
C0037928|T047|SY|48522003|SNOMEDCT_CORE|Spinal cord disorder|Spinal cord disease
C0037928|T047|FN|48522003|SNOMEDCT_CORE|Spinal cord disorder|Spinal cord disease
C0037929|T037|SY|90584004|SNOMEDCT_CORE|SCI - Spinal cord injury|Spinal cord injury
C0037929|T037|PT|90584004|SNOMEDCT_CORE|Spinal cord injury|Spinal cord injury
C0037929|T037|FN|90584004|SNOMEDCT_CORE|Spinal cord injury|Spinal cord injury
C0037929|T037|IS|90584004|SNOMEDCT_CORE|Spinal cord injury, NOS|Spinal cord injury
C0037929|T037|SY|90584004|SNOMEDCT_CORE|Spinal cord syndrome|Spinal cord injury
C0037944|T020|PT|76107001|SNOMEDCT_CORE|Spinal stenosis|Spinal stenosis
C0037944|T020|FN|76107001|SNOMEDCT_CORE|Spinal stenosis|Spinal stenosis
C0037944|T020|IS|76107001|SNOMEDCT_CORE|Spinal stenosis, NOS|Spinal stenosis
C0037944|T020|SY|76107001|SNOMEDCT_CORE|SS - Spinal stenosis|Spinal stenosis
C0037997|T047|SY|58381000|SNOMEDCT_CORE|Dyssplenism|Dyssplenism
C0038002|T033|SY|16294009|SNOMEDCT_CORE|Enlargement of spleen|Splenomegaly
C0038002|T033|IS|16294009|SNOMEDCT_CORE|Enlargement of spleen, NOS|Splenomegaly
C0038002|T033|SY|16294009|SNOMEDCT_CORE|Large spleen|Splenomegaly
C0038002|T033|PT|16294009|SNOMEDCT_CORE|Splenomegaly|Splenomegaly
C0038002|T033|FN|16294009|SNOMEDCT_CORE|Splenomegaly|Splenomegaly
C0038002|T033|IS|16294009|SNOMEDCT_CORE|Splenomegaly, NOS|Splenomegaly
C0038002|T033|IS|16294009|SNOMEDCT_CORE|Unspecified splenomegaly|Splenomegaly
C0038013|T047|PT|9631008|SNOMEDCT_CORE|Ankylosing spondylitis|Ankylosing spondylitis
C0038013|T047|FN|9631008|SNOMEDCT_CORE|Ankylosing spondylitis|Ankylosing spondylitis
C0038013|T047|IS|9631008|SNOMEDCT_CORE|Ankylosing spondylitis, NOS|Ankylosing spondylitis
C0038013|T047|SY|9631008|SNOMEDCT_CORE|AS - Ankylosing spondylitis|Ankylosing spondylitis
C0038013|T047|SY|9631008|SNOMEDCT_CORE|Bekhterev's disease|Ankylosing spondylitis
C0038013|T047|SY|9631008|SNOMEDCT_CORE|Idiopathic ankylosing spondylitis|Ankylosing spondylitis
C0038013|T047|IS|9631008|SNOMEDCT_CORE|Marie Strumpell spondylitis|Ankylosing spondylitis
C0038013|T047|SY|9631008|SNOMEDCT_CORE|Marie Strümpell spondylitis|Ankylosing spondylitis
C0038013|T047|SY|9631008|SNOMEDCT_CORE|Marie-Strumpell spondylitis|Ankylosing spondylitis
C0038013|T047|IS|9631008|SNOMEDCT_CORE|Rheumatoid arthritis of spine|Ankylosing spondylitis
C0038013|T047|IS|9631008|SNOMEDCT_CORE|Rheumatoid arthritis of spine, NOS|Ankylosing spondylitis
C0038013|T047|IS|9631008|SNOMEDCT_CORE|Rheumatoid spondylitis|Ankylosing spondylitis
C0038016|T047|SY|274152003|SNOMEDCT_CORE|SPL - Spondylolisthesis|Spondylolisthesis
C0038016|T047|PT|274152003|SNOMEDCT_CORE|Spondylolisthesis|Spondylolisthesis
C0038016|T047|FN|274152003|SNOMEDCT_CORE|Spondylolisthesis|Spondylolisthesis
C0038017|T019|PT|13236000|SNOMEDCT_CORE|Congenital spondylolisthesis|Congenital spondylolisthesis
C0038017|T019|FN|13236000|SNOMEDCT_CORE|Congenital spondylolisthesis|Congenital spondylolisthesis
C0038019|T047|PT|8847002|SNOMEDCT_CORE|Spondylosis|Spondylosis
C0038019|T047|FN|8847002|SNOMEDCT_CORE|Spondylosis|Spondylosis
C0038019|T047|IS|8847002|SNOMEDCT_CORE|Spondylosis, NOS|Spondylosis
C0038020|T047|SY|9631008|SNOMEDCT_CORE|Spondylosis deformans|Spondylosis deformans
C0038045|T037|PT|384709000|SNOMEDCT_CORE|Sprain|Sprain
C0038045|T037|FN|384709000|SNOMEDCT_CORE|Sprain|Sprain
C0038160|T047|SY|56038003|SNOMEDCT_CORE|Staphylococcal infection|Staphylococcal infectious disease
C0038160|T047|IS|56038003|SNOMEDCT_CORE|Staphylococcal infection, NOS|Staphylococcal infectious disease
C0038160|T047|PT|56038003|SNOMEDCT_CORE|Staphylococcal infectious disease|Staphylococcal infectious disease
C0038160|T047|FN|56038003|SNOMEDCT_CORE|Staphylococcal infectious disease|Staphylococcal infectious disease
C0038160|T047|IS|56038003|SNOMEDCT_CORE|Staphylococcal infectious disease, NOS|Staphylococcal infectious disease
C0038160|T047|SY|56038003|SNOMEDCT_CORE|Staphylococcosis|Staphylococcal infectious disease
C0038218|T047|OAS|57546000|SNOMEDCT_CORE|Acute severe asthma|Acute severe exacerbation of asthma
C0038218|T047|FN|708090002|SNOMEDCT_CORE|Acute severe exacerbation of asthma|Acute severe exacerbation of asthma
C0038218|T047|PT|708090002|SNOMEDCT_CORE|Acute severe exacerbation of asthma|Acute severe exacerbation of asthma
C0038218|T047|OAP|57546000|SNOMEDCT_CORE|Asthma with status asthmaticus|Acute severe exacerbation of asthma
C0038218|T047|OAF|57546000|SNOMEDCT_CORE|Asthma with status asthmaticus|Acute severe exacerbation of asthma
C0038218|T047|OAS|57546000|SNOMEDCT_CORE|Status asthmaticus|Acute severe exacerbation of asthma
C0038218|T047|OP|708090002|SNOMEDCT_CORE|Status asthmaticus|Acute severe exacerbation of asthma
C0038220|T047|IS|13973009|SNOMEDCT_CORE|Status epilepticus|Status epilepticus
C0038238|T033|PT|66187002|SNOMEDCT_CORE|Fatty stool|Fatty stool
C0038238|T033|FN|66187002|SNOMEDCT_CORE|Fatty stool|Fatty stool
C0038238|T033|SY|66187002|SNOMEDCT_CORE|Steatorrhea|Fatty stool
C0038238|T033|IS|66187002|SNOMEDCT_CORE|Steatorrhea, NOS|Fatty stool
C0038238|T033|SYGB|66187002|SNOMEDCT_CORE|Steatorrhoea|Fatty stool
C0038238|T033|IS|66187002|SNOMEDCT_CORE|Steatorrhoea, NOS|Fatty stool
C0038325|T047|IS|73442001|SNOMEDCT_CORE|Bullous erythema multiforme|Stevens-Johnson syndrome
C0038325|T047|IS|73442001|SNOMEDCT_CORE|Ectodermosis erosiva pluriorificialis|Stevens-Johnson syndrome
C0038325|T047|IS|73442001|SNOMEDCT_CORE|Erythema multiforme bullosum|Stevens-Johnson syndrome
C0038325|T047|IS|73442001|SNOMEDCT_CORE|Erythema multiforme exudativum|Stevens-Johnson syndrome
C0038325|T047|IS|73442001|SNOMEDCT_CORE|Erythema multiforme major|Stevens-Johnson syndrome
C0038325|T047|SY|73442001|SNOMEDCT_CORE|Stevens Johnson syndrome|Stevens-Johnson syndrome
C0038325|T047|PT|73442001|SNOMEDCT_CORE|Stevens-Johnson syndrome|Stevens-Johnson syndrome
C0038325|T047|FN|73442001|SNOMEDCT_CORE|Stevens-Johnson syndrome|Stevens-Johnson syndrome
C0038354|T047|IS|29384001|SNOMEDCT_CORE|Disease of stomach|Disorder of stomach
C0038354|T047|OF|29384001|SNOMEDCT_CORE|Disease of stomach|Disorder of stomach
C0038354|T047|IS|29384001|SNOMEDCT_CORE|Disease of stomach, NOS|Disorder of stomach
C0038354|T047|PT|29384001|SNOMEDCT_CORE|Disorder of stomach|Disorder of stomach
C0038354|T047|FN|29384001|SNOMEDCT_CORE|Disorder of stomach|Disorder of stomach
C0038354|T047|SY|29384001|SNOMEDCT_CORE|Gastropathy|Disorder of stomach
C0038356|T191|PT|126824007|SNOMEDCT_CORE|Neoplasm of stomach|Neoplasm of stomach
C0038356|T191|FN|126824007|SNOMEDCT_CORE|Neoplasm of stomach|Neoplasm of stomach
C0038356|T191|SY|126824007|SNOMEDCT_CORE|Tumor of stomach|Neoplasm of stomach
C0038356|T191|SYGB|126824007|SNOMEDCT_CORE|Tumour of stomach|Neoplasm of stomach
C0038358|T047|SY|397825006|SNOMEDCT_CORE|Gastric peptic ulcer|Gastric ulcer
C0038358|T047|PT|397825006|SNOMEDCT_CORE|Gastric ulcer|Gastric ulcer
C0038358|T047|FN|397825006|SNOMEDCT_CORE|Gastric ulcer|Gastric ulcer
C0038358|T047|SY|397825006|SNOMEDCT_CORE|Gastric ulceration|Gastric ulcer
C0038358|T047|SY|397825006|SNOMEDCT_CORE|GU - Gastric ulcer|Gastric ulcer
C0038358|T047|SY|397825006|SNOMEDCT_CORE|Peptic ulcer of stomach|Gastric ulcer
C0038358|T047|SY|397825006|SNOMEDCT_CORE|Stomach ulcer|Gastric ulcer
C0038362|T047|SY|61170000|SNOMEDCT_CORE|Inflammation of mouth|Stomatitis
C0038362|T047|SY|61170000|SNOMEDCT_CORE|Inflammatory condition of oral mucous membrane|Stomatitis
C0038362|T047|SY|61170000|SNOMEDCT_CORE|Oral mucositis|Stomatitis
C0038362|T047|IS|95361005|SNOMEDCT_CORE|Stomatitis|Stomatitis
C0038362|T047|PT|61170000|SNOMEDCT_CORE|Stomatitis|Stomatitis
C0038362|T047|FN|61170000|SNOMEDCT_CORE|Stomatitis|Stomatitis
C0038362|T047|IS|61170000|SNOMEDCT_CORE|Stomatitis, NOS|Stomatitis
C0038363|T047|SY|426965005|SNOMEDCT_CORE|Aphthous stomatitis|Aphthous ulcer of mouth
C0038363|T047|IS|426965005|SNOMEDCT_CORE|Aphthous ulcer|Aphthous ulcer of mouth
C0038363|T047|FN|426965005|SNOMEDCT_CORE|Aphthous ulcer of mouth|Aphthous ulcer of mouth
C0038363|T047|PT|426965005|SNOMEDCT_CORE|Aphthous ulcer of mouth|Aphthous ulcer of mouth
C0038363|T047|IS|426965005|SNOMEDCT_CORE|Aphthous ulceration|Aphthous ulcer of mouth
C0038363|T047|SY|426965005|SNOMEDCT_CORE|Canker sore|Aphthous ulcer of mouth
C0038363|T047|SY|426965005|SNOMEDCT_CORE|Oral aphthae|Aphthous ulcer of mouth
C0038366|T047|SY|57920007|SNOMEDCT_CORE|Herpes stomatitis|Herpes stomatitis
C0038379|T047|SY|22066006|SNOMEDCT_CORE|Disorder of binocular eye movements|Strabismus
C0038379|T047|IS|22066006|SNOMEDCT_CORE|Heterotropia, NOS|Strabismus
C0038379|T047|SY|22066006|SNOMEDCT_CORE|Ocular dissociation|Strabismus
C0038379|T047|SY|22066006|SNOMEDCT_CORE|Squint|Strabismus
C0038379|T047|IS|22066006|SNOMEDCT_CORE|Squint, NOS|Strabismus
C0038379|T047|PT|22066006|SNOMEDCT_CORE|Strabismus|Strabismus
C0038379|T047|FN|22066006|SNOMEDCT_CORE|Strabismus|Strabismus
C0038379|T047|IS|22066006|SNOMEDCT_CORE|Strabismus, NOS|Strabismus
C0038435|T033|IS|73595000|SNOMEDCT_CORE|Pressure, NOS|Stress
C0038435|T033|SY|73595000|SNOMEDCT_CORE|State of stress|Stress
C0038435|T033|PT|73595000|SNOMEDCT_CORE|Stress|Stress
C0038435|T033|FN|73595000|SNOMEDCT_CORE|Stress|Stress
C0038435|T033|IS|73595000|SNOMEDCT_CORE|Stress, NOS|Stress
C0038436|T048|SY|47505003|SNOMEDCT_CORE|Post-traumatic stress disorder|Posttraumatic stress disorder
C0038436|T048|SY|47505003|SNOMEDCT_CORE|Post-traumatic stress syndrome|Posttraumatic stress disorder
C0038436|T048|FN|47505003|SNOMEDCT_CORE|Posttraumatic stress disorder|Posttraumatic stress disorder
C0038436|T048|PT|47505003|SNOMEDCT_CORE|Posttraumatic stress disorder|Posttraumatic stress disorder
C0038436|T048|IS|47505003|SNOMEDCT_CORE|Posttraumatic stress disorder, NOS|Posttraumatic stress disorder
C0038436|T048|SY|47505003|SNOMEDCT_CORE|PTSD - Post-traumatic stress disorder|Posttraumatic stress disorder
C0038436|T048|SY|47505003|SNOMEDCT_CORE|Traumatic neurosis|Posttraumatic stress disorder
C0038437|T047|PT|60241006|SNOMEDCT_CORE|Female stress incontinence|Female stress incontinence
C0038437|T047|SY|60241006|SNOMEDCT_CORE|Female urinary stress incontinence|Female stress incontinence
C0038437|T047|FN|60241006|SNOMEDCT_CORE|Female urinary stress incontinence|Female stress incontinence
C0038443|T048|SY|73595000|SNOMEDCT_CORE|Psychological stress|Psychological stress
C0038450|T184|PT|70407001|SNOMEDCT_CORE|Stridor|Stridor
C0038450|T184|FN|70407001|SNOMEDCT_CORE|Stridor|Stridor
C0038450|T184|SY|70407001|SNOMEDCT_CORE|Stridulous breathing|Stridor
C0038454|T047|PT|230690007|SNOMEDCT_CORE|Cerebrovascular accident|Cerebrovascular accident
C0038454|T047|FN|230690007|SNOMEDCT_CORE|Cerebrovascular accident|Cerebrovascular accident
C0038454|T047|SY|230690007|SNOMEDCT_CORE|CVA - Cerebrovascular accident|Cerebrovascular accident
C0038454|T047|SY|230690007|SNOMEDCT_CORE|Stroke|Cerebrovascular accident
C0038506|T048|SY|39423001|SNOMEDCT_CORE|Dysphemia|Stuttering
C0038506|T048|IS|39423001|SNOMEDCT_CORE|dysphemia|Stuttering
C0038506|T048|SY|39423001|SNOMEDCT_CORE|Non-fluent speech|Stuttering
C0038506|T048|SYGB|39423001|SNOMEDCT_CORE|Stammer|Stuttering
C0038506|T048|PTGB|39423001|SNOMEDCT_CORE|Stammering|Stuttering
C0038506|T048|OF|39423001|SNOMEDCT_CORE|Stammering|Stuttering
C0038506|T048|SY|39423001|SNOMEDCT_CORE|Stutter|Stuttering
C0038506|T048|PT|39423001|SNOMEDCT_CORE|Stuttering|Stuttering
C0038506|T048|FN|39423001|SNOMEDCT_CORE|Stuttering|Stuttering
C0038525|T047|SYGB|21454007|SNOMEDCT_CORE|SAH - Subarachnoid haemorrhage|Subarachnoid hemorrhage
C0038525|T047|SY|21454007|SNOMEDCT_CORE|SAH - Subarachnoid hemorrhage|Subarachnoid hemorrhage
C0038525|T047|PTGB|21454007|SNOMEDCT_CORE|Subarachnoid haemorrhage|Subarachnoid hemorrhage
C0038525|T047|PT|21454007|SNOMEDCT_CORE|Subarachnoid hemorrhage|Subarachnoid hemorrhage
C0038525|T047|OF|21454007|SNOMEDCT_CORE|Subarachnoid hemorrhage|Subarachnoid hemorrhage
C0038525|T047|SYGB|21454007|SNOMEDCT_CORE|Subarachnoid intracranial haemorrhage|Subarachnoid hemorrhage
C0038525|T047|SY|21454007|SNOMEDCT_CORE|Subarachnoid intracranial hemorrhage|Subarachnoid hemorrhage
C0038525|T047|FN|21454007|SNOMEDCT_CORE|Subarachnoid intracranial hemorrhage|Subarachnoid hemorrhage
C0038531|T047|PT|15258001|SNOMEDCT_CORE|Subclavian steal syndrome|Subclavian steal syndrome
C0038531|T047|FN|15258001|SNOMEDCT_CORE|Subclavian steal syndrome|Subclavian steal syndrome
C0038534|T046|SY|78768009|SNOMEDCT_CORE|Subconjunctival bleed|Subconjunctival hemorrhage
C0038534|T046|PTGB|78768009|SNOMEDCT_CORE|Subconjunctival haemorrhage|Subconjunctival hemorrhage
C0038534|T046|PT|78768009|SNOMEDCT_CORE|Subconjunctival hemorrhage|Subconjunctival hemorrhage
C0038534|T046|FN|78768009|SNOMEDCT_CORE|Subconjunctival hemorrhage|Subconjunctival hemorrhage
C0038558|T191|OAP|254464000|SNOMEDCT_CORE|Tumor of submandibular gland|Tumor of submandibular gland
C0038558|T191|OAF|254464000|SNOMEDCT_CORE|Tumor of submandibular gland|Tumor of submandibular gland
C0038558|T191|OAP|254464000|SNOMEDCT_CORE|Tumour of submandibular gland|Tumour of submandibular gland
C0038580|T048|SY|2403008|SNOMEDCT_CORE|Substance dependence|Substance dependence
C0038580|T048|IS|2403008|SNOMEDCT_CORE|Substance dependence, NOS|Substance dependence
C0038661|T033|PT|44301001|SNOMEDCT_CORE|Suicide|Suicide
C0038661|T033|OF|44301001|SNOMEDCT_CORE|Suicide|Suicide
C0038661|T033|FN|44301001|SNOMEDCT_CORE|Suicide|Suicide
C0038661|T033|IS|44301001|SNOMEDCT_CORE|Suicide, NOS|Suicide
C0038663|T037|PT|82313006|SNOMEDCT_CORE|Suicide attempt|Suicide attempt
C0038663|T037|OF|82313006|SNOMEDCT_CORE|Suicide attempt|Suicide attempt
C0038663|T037|FN|82313006|SNOMEDCT_CORE|Suicide attempt|Suicide attempt
C0038663|T037|IS|82313006|SNOMEDCT_CORE|Suicide attempt, NOS|Suicide attempt
C0038814|T037|IS|23346002|SNOMEDCT_CORE|Erythema solare|Sunburn
C0038814|T037|IS|23346002|SNOMEDCT_CORE|Solar erythema|Sunburn
C0038814|T037|OAP|23346002|SNOMEDCT_CORE|Sunburn|Sunburn
C0038814|T037|OAF|23346002|SNOMEDCT_CORE|Sunburn|Sunburn
C0038833|T047|IS|63363004|SNOMEDCT_CORE|Superior vena cava obstruction|Superior vena cava syndrome
C0038833|T047|PT|63363004|SNOMEDCT_CORE|Superior vena cava syndrome|Superior vena cava syndrome
C0038833|T047|FN|63363004|SNOMEDCT_CORE|Superior vena cava syndrome|Superior vena cava syndrome
C0038833|T047|IS|63363004|SNOMEDCT_CORE|SVC - Superior vena cava obstruction|Superior vena cava syndrome
C0038833|T047|IS|63363004|SNOMEDCT_CORE|SVCO - Superior vena cava obstruction|Superior vena cava syndrome
C0038868|T047|IS|28978003|SNOMEDCT_CORE|Progressive supranuclear palsy|Progressive supranuclear palsy
C0038868|T047|IS|28978003|SNOMEDCT_CORE|PSP - Progressive supranuclear palsy|Progressive supranuclear palsy
C0038940|T046|SY|22247000|SNOMEDCT_CORE|Dehiscence of operation wound|Dehiscence of surgical wound
C0038940|T046|PT|22247000|SNOMEDCT_CORE|Dehiscence of surgical wound|Dehiscence of surgical wound
C0038940|T046|FN|22247000|SNOMEDCT_CORE|Dehiscence of surgical wound|Dehiscence of surgical wound
C0038940|T046|IS|22247000|SNOMEDCT_CORE|Disruption of operation wound|Dehiscence of surgical wound
C0038940|T046|SY|22247000|SNOMEDCT_CORE|Operation wound dehiscence|Dehiscence of surgical wound
C0038940|T046|SY|22247000|SNOMEDCT_CORE|Operation wound disruption|Dehiscence of surgical wound
C0038940|T046|OF|22247000|SNOMEDCT_CORE|Operation wound disruption|Dehiscence of surgical wound
C0038940|T046|SY|22247000|SNOMEDCT_CORE|Operation wound rupture|Dehiscence of surgical wound
C0038940|T046|IS|22247000|SNOMEDCT_CORE|Postoperative wound breakdown|Dehiscence of surgical wound
C0038940|T046|SY|22247000|SNOMEDCT_CORE|Rupture of operation wound|Dehiscence of surgical wound
C0038940|T046|SY|22247000|SNOMEDCT_CORE|Wound breakdown|Dehiscence of surgical wound
C0038941|T046|SY|58126003|SNOMEDCT_CORE|Infected surgical wound|Postoperative wound infection
C0038941|T046|PT|58126003|SNOMEDCT_CORE|Postoperative wound infection|Postoperative wound infection
C0038941|T046|FN|58126003|SNOMEDCT_CORE|Postoperative wound infection|Postoperative wound infection
C0038967|T046|PT|66962008|SNOMEDCT_CORE|Suture granuloma|Suture granuloma
C0038967|T046|FN|66962008|SNOMEDCT_CORE|Suture granuloma|Suture granuloma
C0038990|T033|PT|415690000|SNOMEDCT_CORE|Sweating|Sweating
C0038990|T033|FN|415690000|SNOMEDCT_CORE|Sweating|Sweating
C0038990|T033|SY|415690000|SNOMEDCT_CORE|Sweats|Sweating
C0038999|T033|SY|65124004|SNOMEDCT_CORE|Bulge|Swelling
C0038999|T033|IS|65124004|SNOMEDCT_CORE|Bulge, NOS|Swelling
C0038999|T033|SY|65124004|SNOMEDCT_CORE|Observation of swelling|Swelling
C0038999|T033|SY|65124004|SNOMEDCT_CORE|Part of body puffy|Swelling
C0038999|T033|SY|65124004|SNOMEDCT_CORE|Part of body swollen|Swelling
C0038999|T033|PT|65124004|SNOMEDCT_CORE|Swelling|Swelling
C0038999|T033|FN|65124004|SNOMEDCT_CORE|Swelling|Swelling
C0038999|T033|IS|65124004|SNOMEDCT_CORE|Swelling, NOS|Swelling
C0038999|T033|SY|65124004|SNOMEDCT_CORE|Tumefaction|Swelling
C0038999|T033|SY|65124004|SNOMEDCT_CORE|Tumescence|Swelling
C0039070|T184|SY|271594007|SNOMEDCT_CORE|Blackout|Syncope
C0039070|T184|SY|271594007|SNOMEDCT_CORE|Faint|Syncope
C0039070|T184|SY|271594007|SNOMEDCT_CORE|Fainting|Syncope
C0039070|T184|PT|271594007|SNOMEDCT_CORE|Syncope|Syncope
C0039070|T184|FN|271594007|SNOMEDCT_CORE|Syncope|Syncope
C0039070|T184|PT|309585006|SNOMEDCT_CORE|Syncope and collapse|Syncope
C0039070|T184|FN|309585006|SNOMEDCT_CORE|Syncope and collapse|Syncope
C0039070|T184|SY|271594007|SNOMEDCT_CORE|Syncope attack|Syncope
C0039101|T191|SY|302851001|SNOMEDCT_CORE|Malignant synovioma|Synovial sarcoma
C0039101|T191|PT|302851001|SNOMEDCT_CORE|Synovial sarcoma|Synovial sarcoma
C0039101|T191|FN|302851001|SNOMEDCT_CORE|Synovial sarcoma|Synovial sarcoma
C0039103|T047|PT|416209007|SNOMEDCT_CORE|Synovitis|Synovitis
C0039103|T047|FN|416209007|SNOMEDCT_CORE|Synovitis|Synovitis
C0039104|T047|PT|202900007|SNOMEDCT_CORE|Synovitis and tenosynovitis|Synovitis and tenosynovitis
C0039104|T047|FN|202900007|SNOMEDCT_CORE|Synovitis and tenosynovitis|Synovitis and tenosynovitis
C0039128|T047|SY|76272004|SNOMEDCT_CORE|Infection by Treponema pallidum|Syphilis
C0039128|T047|SY|76272004|SNOMEDCT_CORE|Lues|Syphilis
C0039128|T047|SY|76272004|SNOMEDCT_CORE|Luetic disease|Syphilis
C0039128|T047|PT|76272004|SNOMEDCT_CORE|Syphilis|Syphilis
C0039128|T047|FN|76272004|SNOMEDCT_CORE|Syphilis|Syphilis
C0039128|T047|IS|76272004|SNOMEDCT_CORE|Syphilis, NOS|Syphilis
C0039128|T047|IS|76272004|SNOMEDCT_CORE|Syphilis, stage unspecified|Syphilis
C0039131|T047|PT|35742006|SNOMEDCT_CORE|Congenital syphilis|Congenital syphilis
C0039131|T047|FN|35742006|SNOMEDCT_CORE|Congenital syphilis|Congenital syphilis
C0039131|T047|IS|35742006|SNOMEDCT_CORE|Congenital syphilis, NOS|Congenital syphilis
C0039133|T047|PT|444150000|SNOMEDCT_CORE|Latent syphilis|Latent syphilis
C0039133|T047|FN|444150000|SNOMEDCT_CORE|Latent syphilis|Latent syphilis
C0039144|T047|SY|111496009|SNOMEDCT_CORE|Myelosyringosis|Syringomyelia
C0039144|T047|PT|111496009|SNOMEDCT_CORE|Syringomyelia|Syringomyelia
C0039144|T047|FN|111496009|SNOMEDCT_CORE|Syringomyelia|Syringomyelia
C0039144|T047|SYGB|111496009|SNOMEDCT_CORE|Syringomyelia-anaesthesia syndrome|Syringomyelia
C0039144|T047|SY|111496009|SNOMEDCT_CORE|Syringomyelia-anesthesia syndrome|Syringomyelia
C0039231|T033|IS|6285003|SNOMEDCT_CORE|Heart rate fast|Tachycardia
C0039231|T033|SY|3424008|SNOMEDCT_CORE|Heart rate fast|Tachycardia
C0039231|T033|IS|6285003|SNOMEDCT_CORE|Increased heart rate|Tachycardia
C0039231|T033|SY|3424008|SNOMEDCT_CORE|Increased heart rate|Tachycardia
C0039231|T033|IS|6285003|SNOMEDCT_CORE|Rapid heart beat|Tachycardia
C0039231|T033|SY|3424008|SNOMEDCT_CORE|Rapid heart beat|Tachycardia
C0039231|T033|IS|6285003|SNOMEDCT_CORE|Tachycardia|Tachycardia
C0039231|T033|PT|3424008|SNOMEDCT_CORE|Tachycardia|Tachycardia
C0039231|T033|FN|3424008|SNOMEDCT_CORE|Tachycardia|Tachycardia
C0039231|T033|IS|3424008|SNOMEDCT_CORE|Tachycardia, NOS|Tachycardia
C0039232|T047|FN|251166008|SNOMEDCT_CORE|Atrioventricular nodal re-entry tachycardia|AV nodal re-entry tachycardia
C0039232|T047|SY|251166008|SNOMEDCT_CORE|Atrioventricular nodal re-entry tachycardia|AV nodal re-entry tachycardia
C0039232|T047|PT|251166008|SNOMEDCT_CORE|AV nodal re-entry tachycardia|AV nodal re-entry tachycardia
C0039232|T047|OF|251166008|SNOMEDCT_CORE|AV nodal re-entry tachycardia|AV nodal re-entry tachycardia
C0039236|T047|SY|12026006|SNOMEDCT_CORE|Bouveret-Hoffmann syndrome|Paroxysmal tachycardia
C0039236|T047|SY|12026006|SNOMEDCT_CORE|Essential paroxysmal tachycardia|Paroxysmal tachycardia
C0039236|T047|PT|12026006|SNOMEDCT_CORE|Paroxysmal tachycardia|Paroxysmal tachycardia
C0039236|T047|FN|12026006|SNOMEDCT_CORE|Paroxysmal tachycardia|Paroxysmal tachycardia
C0039236|T047|IS|12026006|SNOMEDCT_CORE|Paroxysmal tachycardia, NOS|Paroxysmal tachycardia
C0039236|T047|SY|12026006|SNOMEDCT_CORE|PT - Paroxysmal tachycardia|Paroxysmal tachycardia
C0039239|T047|PT|11092001|SNOMEDCT_CORE|Sinus tachycardia|Sinus tachycardia
C0039239|T047|FN|11092001|SNOMEDCT_CORE|Sinus tachycardia|Sinus tachycardia
C0039240|T047|PT|6456007|SNOMEDCT_CORE|Supraventricular tachycardia|Supraventricular tachycardia
C0039240|T047|FN|6456007|SNOMEDCT_CORE|Supraventricular tachycardia|Supraventricular tachycardia
C0039240|T047|IS|6456007|SNOMEDCT_CORE|Supraventricular tachycardia, NOS|Supraventricular tachycardia
C0039240|T047|SY|6456007|SNOMEDCT_CORE|SVT - Supraventricular tachycardia|Supraventricular tachycardia
C0039263|T047|SY|359789008|SNOMEDCT_CORE|Acquired aortoarteritis|Takayasu's disease
C0039263|T047|SY|359789008|SNOMEDCT_CORE|Aortic arch arteritis|Takayasu's disease
C0039263|T047|SY|359789008|SNOMEDCT_CORE|Atypical coarctation|Takayasu's disease
C0039263|T047|SY|359789008|SNOMEDCT_CORE|Idiopathic medial aortopathy AND arteriopathy|Takayasu's disease
C0039263|T047|SY|359789008|SNOMEDCT_CORE|Martorell syndrome|Takayasu's disease
C0039263|T047|IS|359789008|SNOMEDCT_CORE|Middle aortic syndrome|Takayasu's disease
C0039263|T047|SY|359789008|SNOMEDCT_CORE|Nonspecific aortoarteritis|Takayasu's disease
C0039263|T047|SY|359789008|SNOMEDCT_CORE|Nonspecific arteritis|Takayasu's disease
C0039263|T047|SY|359789008|SNOMEDCT_CORE|Occlusive thromboarteriopathy|Takayasu's disease
C0039263|T047|SY|359789008|SNOMEDCT_CORE|Primary arteritis|Takayasu's disease
C0039263|T047|SY|359789008|SNOMEDCT_CORE|Pulseless disease|Takayasu's disease
C0039263|T047|SY|359789008|SNOMEDCT_CORE|Raeder-Harbitz syndrome|Takayasu's disease
C0039263|T047|SY|359789008|SNOMEDCT_CORE|Reverse coarctation|Takayasu's disease
C0039263|T047|SY|359789008|SNOMEDCT_CORE|Sclerosing aortitis AND arteritis|Takayasu's disease
C0039263|T047|SY|359789008|SNOMEDCT_CORE|Takayasu disease|Takayasu's disease
C0039263|T047|SY|359789008|SNOMEDCT_CORE|Takayasu's arteriopathy|Takayasu's disease
C0039263|T047|SY|359789008|SNOMEDCT_CORE|Takayasu's arteritis|Takayasu's disease
C0039263|T047|PT|359789008|SNOMEDCT_CORE|Takayasu's disease|Takayasu's disease
C0039263|T047|FN|359789008|SNOMEDCT_CORE|Takayasu's disease|Takayasu's disease
C0039263|T047|SY|359789008|SNOMEDCT_CORE|Young female arteritis|Takayasu's disease
C0039292|T047|SYGB|15346004|SNOMEDCT_CORE|Analphalipoproteinaemia|Analphalipoproteinemia
C0039292|T047|SY|15346004|SNOMEDCT_CORE|Analphalipoproteinemia|Analphalipoproteinemia
C0039292|T047|SYGB|15346004|SNOMEDCT_CORE|Analphaliproteinaemia|Analphalipoproteinemia
C0039292|T047|SY|15346004|SNOMEDCT_CORE|Analphaliproteinemia|Analphalipoproteinemia
C0039292|T047|SY|15346004|SNOMEDCT_CORE|Cholesterol thesaurismosis|Analphalipoproteinemia
C0039292|T047|IS|15346004|SNOMEDCT_CORE|Tangier disease|Analphalipoproteinemia
C0039319|T047|PT|47374004|SNOMEDCT_CORE|Tarsal tunnel syndrome|Tarsal tunnel syndrome
C0039319|T047|SY|47374004|SNOMEDCT_CORE|Tarsal tunnel syndrome|Tarsal tunnel syndrome
C0039319|T047|FN|47374004|SNOMEDCT_CORE|Tarsal tunnel syndrome|Tarsal tunnel syndrome
C0039319|T047|SY|47374004|SNOMEDCT_CORE|TTS - Tarsal tunnel syndrome|Tarsal tunnel syndrome
C0039338|T047|PT|399993004|SNOMEDCT_CORE|Disorder of taste|Disorder of taste
C0039338|T047|FN|399993004|SNOMEDCT_CORE|Disorder of taste|Disorder of taste
C0039437|T033|PT|8004003|SNOMEDCT_CORE|Teething syndrome|Teething syndrome
C0039437|T033|FN|8004003|SNOMEDCT_CORE|Teething syndrome|Teething syndrome
C0039437|T033|OF|8004003|SNOMEDCT_CORE|Teething syndrome|Teething syndrome
C0039445|T047|SYGB|21877004|SNOMEDCT_CORE|Hereditary haemorrhagic telangiectasia|Osler hemorrhagic telangiectasia syndrome
C0039445|T047|SY|21877004|SNOMEDCT_CORE|Hereditary hemorrhagic telangiectasia|Osler hemorrhagic telangiectasia syndrome
C0039445|T047|SYGB|21877004|SNOMEDCT_CORE|HHT - Hereditary haemorrhagic telangiectasia|Osler hemorrhagic telangiectasia syndrome
C0039445|T047|SY|21877004|SNOMEDCT_CORE|HHT - Hereditary hemorrhagic telangiectasia|Osler hemorrhagic telangiectasia syndrome
C0039445|T047|PTGB|21877004|SNOMEDCT_CORE|Osler haemorrhagic telangiectasia syndrome|Osler hemorrhagic telangiectasia syndrome
C0039445|T047|PT|21877004|SNOMEDCT_CORE|Osler hemorrhagic telangiectasia syndrome|Osler hemorrhagic telangiectasia syndrome
C0039445|T047|FN|21877004|SNOMEDCT_CORE|Osler hemorrhagic telangiectasia syndrome|Osler hemorrhagic telangiectasia syndrome
C0039445|T047|SY|21877004|SNOMEDCT_CORE|Osler-Rendu-Weber disease|Osler hemorrhagic telangiectasia syndrome
C0039445|T047|SY|21877004|SNOMEDCT_CORE|Osler-Rendu-Weber syndrome|Osler hemorrhagic telangiectasia syndrome
C0039445|T047|SY|21877004|SNOMEDCT_CORE|Osler-Weber-Rendu disease|Osler hemorrhagic telangiectasia syndrome
C0039445|T047|SY|21877004|SNOMEDCT_CORE|Osler's disease|Osler hemorrhagic telangiectasia syndrome
C0039445|T047|IS|21877004|SNOMEDCT_CORE|Synonym deleted refer to DC-F4801|Osler hemorrhagic telangiectasia syndrome
C0039446|T033|SY|247479008|SNOMEDCT_CORE|Hyphenwebs|Telangiectasia disorder
C0039446|T033|OAP|276328002|SNOMEDCT_CORE|Telangiectasia|Telangiectasia disorder
C0039446|T033|OAF|276328002|SNOMEDCT_CORE|Telangiectasia|Telangiectasia disorder
C0039446|T033|PT|247479008|SNOMEDCT_CORE|Telangiectasia disorder|Telangiectasia disorder
C0039446|T033|FN|247479008|SNOMEDCT_CORE|Telangiectasia disorder|Telangiectasia disorder
C0039446|T033|SY|247479008|SNOMEDCT_CORE|Thread veins|Telangiectasia disorder
C0039483|T047|OAP|414341000|SNOMEDCT_CORE|Giant cell arteritis|Horton's disease
C0039483|T047|OAF|414341000|SNOMEDCT_CORE|Giant cell arteritis|Horton's disease
C0039483|T047|SY|400130008|SNOMEDCT_CORE|Horton's disease|Horton's disease
C0039494|T047|PT|41888000|SNOMEDCT_CORE|Temporomandibular joint disorder|Temporomandibular joint disorder
C0039494|T047|FN|41888000|SNOMEDCT_CORE|Temporomandibular joint disorder|Temporomandibular joint disorder
C0039494|T047|IS|41888000|SNOMEDCT_CORE|Temporomandibular joint disorder, NOS|Temporomandibular joint disorder
C0039494|T047|SY|41888000|SNOMEDCT_CORE|TMJ - Temporomandibular joint disorder|Temporomandibular joint disorder
C0039496|T047|SY|386207004|SNOMEDCT_CORE|Costen's complex|Temporomandibular joint-pain-dysfunction syndrome
C0039496|T047|SY|386207004|SNOMEDCT_CORE|Costen's syndrome|Temporomandibular joint-pain-dysfunction syndrome
C0039496|T047|SY|386207004|SNOMEDCT_CORE|Mandibular dysfunction|Temporomandibular joint-pain-dysfunction syndrome
C0039496|T047|SY|386207004|SNOMEDCT_CORE|Myofascial pain - dysfunction syndrome of TMJ|Temporomandibular joint-pain-dysfunction syndrome
C0039496|T047|SY|386207004|SNOMEDCT_CORE|Snapping jaw|Temporomandibular joint-pain-dysfunction syndrome
C0039496|T047|SY|386207004|SNOMEDCT_CORE|Temporomandibular joint pain dysfunction syndrome|Temporomandibular joint-pain-dysfunction syndrome
C0039496|T047|SY|41888000|SNOMEDCT_CORE|Temporomandibular joint syndrome|Temporomandibular joint-pain-dysfunction syndrome
C0039496|T047|IS|41888000|SNOMEDCT_CORE|Temporomandibular joint syndrome, NOS|Temporomandibular joint-pain-dysfunction syndrome
C0039496|T047|PT|386207004|SNOMEDCT_CORE|Temporomandibular joint-pain-dysfunction syndrome|Temporomandibular joint-pain-dysfunction syndrome
C0039496|T047|FN|386207004|SNOMEDCT_CORE|Temporomandibular joint-pain-dysfunction syndrome|Temporomandibular joint-pain-dysfunction syndrome
C0039496|T047|SY|386207004|SNOMEDCT_CORE|TMJ syndrome|Temporomandibular joint-pain-dysfunction syndrome
C0039496|T047|SY|386207004|SNOMEDCT_CORE|TMJPDS - Temporomandibular joint pain dysfunction syndrome|Temporomandibular joint-pain-dysfunction syndrome
C0039503|T047|SY|34840004|SNOMEDCT_CORE|Inflammatory disorder of tendon|Tendinitis
C0039503|T047|PT|34840004|SNOMEDCT_CORE|Tendinitis|Tendinitis
C0039503|T047|FN|34840004|SNOMEDCT_CORE|Tendinitis|Tendinitis
C0039503|T047|IS|34840004|SNOMEDCT_CORE|Tendinitis, NOS|Tendinitis
C0039503|T047|SY|34840004|SNOMEDCT_CORE|Tendonitis|Tendinitis
C0039503|T047|IS|34840004|SNOMEDCT_CORE|Tendonitis, NOS|Tendinitis
C0039516|T047|PT|202855006|SNOMEDCT_CORE|Lateral epicondylitis|Lateral epicondylitis
C0039516|T047|FN|202855006|SNOMEDCT_CORE|Lateral epicondylitis|Lateral epicondylitis
C0039516|T047|SY|202855006|SNOMEDCT_CORE|Lateral epicondylitis of elbow|Lateral epicondylitis
C0039516|T047|IS|202855006|SNOMEDCT_CORE|Tennis elbow|Lateral epicondylitis
C0039520|T047|SY|67801009|SNOMEDCT_CORE|Inflammation of tendon sheath|Tenosynovitis
C0039520|T047|SY|67801009|SNOMEDCT_CORE|Tendinous synovitis|Tenosynovitis
C0039520|T047|SY|67801009|SNOMEDCT_CORE|Tendovaginitis|Tenosynovitis
C0039520|T047|SY|67801009|SNOMEDCT_CORE|Tenontolemmitis|Tenosynovitis
C0039520|T047|PT|67801009|SNOMEDCT_CORE|Tenosynovitis|Tenosynovitis
C0039520|T047|FN|67801009|SNOMEDCT_CORE|Tenosynovitis|Tenosynovitis
C0039520|T047|IS|67801009|SNOMEDCT_CORE|Tenosynovitis, NOS|Tenosynovitis
C0039520|T047|SY|67801009|SNOMEDCT_CORE|Tenovaginitis|Tenosynovitis
C0039520|T047|IS|67801009|SNOMEDCT_CORE|Vaginal synovitis|Tenosynovitis
C0039591|T184|SY|63901009|SNOMEDCT_CORE|Orchialgia|Pain in testicle
C0039591|T184|IS|63901009|SNOMEDCT_CORE|Orchialgia, NOS|Pain in testicle
C0039591|T184|SY|63901009|SNOMEDCT_CORE|Orchidalgia|Pain in testicle
C0039591|T184|IS|63901009|SNOMEDCT_CORE|Orchidalgia, NOS|Pain in testicle
C0039591|T184|SY|63901009|SNOMEDCT_CORE|Orchidodynia|Pain in testicle
C0039591|T184|IS|63901009|SNOMEDCT_CORE|Orchidodynia, NOS|Pain in testicle
C0039591|T184|PT|63901009|SNOMEDCT_CORE|Pain in testicle|Pain in testicle
C0039591|T184|FN|63901009|SNOMEDCT_CORE|Pain in testicle|Pain in testicle
C0039591|T184|SY|63901009|SNOMEDCT_CORE|Pain in testis|Pain in testicle
C0039591|T184|SY|63901009|SNOMEDCT_CORE|Pain of testes|Pain in testicle
C0039591|T184|IS|63901009|SNOMEDCT_CORE|Testicular pain|Pain in testicle
C0039591|T184|IS|63901009|SNOMEDCT_CORE|Testicular pain, NOS|Pain in testicle
C0039614|T047|IS|76902006|SNOMEDCT_CORE|Infection due to Clostridium tetani|Tetanus
C0039614|T047|PT|76902006|SNOMEDCT_CORE|Tetanus|Tetanus
C0039614|T047|FN|76902006|SNOMEDCT_CORE|Tetanus|Tetanus
C0039685|T019|SY|86299006|SNOMEDCT_CORE|Fallot's tetralogy|Tetralogy of Fallot
C0039685|T019|SY|86299006|SNOMEDCT_CORE|Subpulmonic stenosis, ventricular septal defect, overriding aorta, AND right ventricular hypertrophy|Tetralogy of Fallot
C0039685|T019|IS|86299006|SNOMEDCT_CORE|Subpulmonic stenosis, ventricular septal defect, overriding aorta, and right ventricular hypertrophy|Tetralogy of Fallot
C0039685|T019|PT|86299006|SNOMEDCT_CORE|Tetralogy of Fallot|Tetralogy of Fallot
C0039685|T019|FN|86299006|SNOMEDCT_CORE|Tetralogy of Fallot|Tetralogy of Fallot
C0039685|T019|SY|86299006|SNOMEDCT_CORE|TOF - Tetralogy of Fallot|Tetralogy of Fallot
C0039730|T047|SY|40108008|SNOMEDCT_CORE|Hereditary leptocytosis|Thalassemia
C0039730|T047|PTGB|40108008|SNOMEDCT_CORE|Thalassaemia|Thalassemia
C0039730|T047|PT|40108008|SNOMEDCT_CORE|Thalassemia|Thalassemia
C0039730|T047|FN|40108008|SNOMEDCT_CORE|Thalassemia|Thalassemia
C0039730|T047|IS|40108008|SNOMEDCT_CORE|Thalassemia, NOS|Thalassemia
C0039841|T047|SY|399357009|SNOMEDCT_CORE|Aneurin deficiency|Thiamine deficiency
C0039841|T047|SY|399357009|SNOMEDCT_CORE|Thiamin deficiency|Thiamine deficiency
C0039841|T047|OF|399357009|SNOMEDCT_CORE|Thiamin deficiency|Thiamine deficiency
C0039841|T047|PT|399357009|SNOMEDCT_CORE|Thiamine deficiency|Thiamine deficiency
C0039841|T047|FN|399357009|SNOMEDCT_CORE|Thiamine deficiency|Thiamine deficiency
C0039841|T047|SY|399357009|SNOMEDCT_CORE|Vitamin B1 deficiency|Thiamine deficiency
C0039980|T037|PT|262525000|SNOMEDCT_CORE|Chest injury|Chest injury
C0039980|T037|FN|262525000|SNOMEDCT_CORE|Chest injury|Chest injury
C0039984|T047|PT|128210009|SNOMEDCT_CORE|Thoracic outlet syndrome|Thoracic outlet syndrome
C0039984|T047|FN|128210009|SNOMEDCT_CORE|Thoracic outlet syndrome|Thoracic outlet syndrome
C0039984|T047|SY|128210009|SNOMEDCT_CORE|TOS - Thoracic outlet syndrome|Thoracic outlet syndrome
C0040028|T047|PTGB|109994006|SNOMEDCT_CORE|Essential thrombocythaemia|Essential thrombocythemia
C0040028|T047|IS|109994006|SNOMEDCT_CORE|Essential thrombocythaemia|Essential thrombocythemia
C0040028|T047|OP|109994006|SNOMEDCT_CORE|Essential thrombocythaemia|Essential thrombocythemia
C0040028|T047|IS|109994006|SNOMEDCT_CORE|Essential thrombocythemia|Essential thrombocythemia
C0040028|T047|FN|109994006|SNOMEDCT_CORE|Essential thrombocythemia|Essential thrombocythemia
C0040028|T047|PT|109994006|SNOMEDCT_CORE|Essential thrombocythemia|Essential thrombocythemia
C0040028|T047|SY|109994006|SNOMEDCT_CORE|Essential thrombocythemia|Essential thrombocythemia
C0040028|T047|SY|109994006|SNOMEDCT_CORE|Essential thrombocytosis|Essential thrombocythemia
C0040028|T047|SYGB|109994006|SNOMEDCT_CORE|Idiopathic thrombocythaemia|Essential thrombocythemia
C0040028|T047|IS|109994006|SNOMEDCT_CORE|Idiopathic thrombocythaemia|Essential thrombocythemia
C0040028|T047|SY|109994006|SNOMEDCT_CORE|Idiopathic thrombocythemia|Essential thrombocythemia
C0040028|T047|IS|109994006|SNOMEDCT_CORE|Idiopathic thrombocythemia|Essential thrombocythemia
C0040034|T047|SY|302215000|SNOMEDCT_CORE|Thrombocytopenia|Thrombocytopenic disorder
C0040034|T047|PT|302215000|SNOMEDCT_CORE|Thrombocytopenic disorder|Thrombocytopenic disorder
C0040034|T047|FN|302215000|SNOMEDCT_CORE|Thrombocytopenic disorder|Thrombocytopenic disorder
C0040046|T046|PT|64156001|SNOMEDCT_CORE|Thrombophlebitis|Thrombophlebitis
C0040046|T046|FN|64156001|SNOMEDCT_CORE|Thrombophlebitis|Thrombophlebitis
C0040046|T046|IS|64156001|SNOMEDCT_CORE|Thrombophlebitis, NOS|Thrombophlebitis
C0040100|T191|PT|444231005|SNOMEDCT_CORE|Thymoma|Thymoma
C0040100|T191|PT|128856005|SNOMEDCT_CORE|Thymoma|Thymoma
C0040100|T191|OF|128856005|SNOMEDCT_CORE|Thymoma|Thymoma
C0040100|T191|FN|444231005|SNOMEDCT_CORE|Thymoma|Thymoma
C0040100|T191|OF|128856005|SNOMEDCT_CORE|Thymoma, no ICD-O subtype|Thymoma
C0040100|T191|SY|128856005|SNOMEDCT_CORE|Thymoma, no ICD-O subtype|Thymoma
C0040100|T191|SY|128856005|SNOMEDCT_CORE|Thymoma, no International Classification of Diseases for Oncology subtype|Thymoma
C0040100|T191|FN|128856005|SNOMEDCT_CORE|Thymoma, no International Classification of Diseases for Oncology subtype|Thymoma
C0040124|T019|IS|39462005|SNOMEDCT_CORE|Thryroglossal duct cyst|Thyroglossal duct cyst
C0040124|T019|SY|39462005|SNOMEDCT_CORE|Thyroglossal cyst|Thyroglossal duct cyst
C0040124|T019|PT|39462005|SNOMEDCT_CORE|Thyroglossal duct cyst|Thyroglossal duct cyst
C0040124|T019|FN|39462005|SNOMEDCT_CORE|Thyroglossal duct cyst|Thyroglossal duct cyst
C0040128|T047|IS|14304000|SNOMEDCT_CORE|Disease of thyroid gland|Disorder of thyroid gland
C0040128|T047|OF|14304000|SNOMEDCT_CORE|Disease of thyroid gland|Disorder of thyroid gland
C0040128|T047|IS|14304000|SNOMEDCT_CORE|Disease of thyroid gland, NOS|Disorder of thyroid gland
C0040128|T047|PT|14304000|SNOMEDCT_CORE|Disorder of thyroid gland|Disorder of thyroid gland
C0040128|T047|FN|14304000|SNOMEDCT_CORE|Disorder of thyroid gland|Disorder of thyroid gland
C0040128|T047|IS|14304000|SNOMEDCT_CORE|Disorder of thyroid gland, NOS|Disorder of thyroid gland
C0040128|T047|SY|14304000|SNOMEDCT_CORE|Thyroid disease|Disorder of thyroid gland
C0040128|T047|SY|14304000|SNOMEDCT_CORE|Thyroid disorder|Disorder of thyroid gland
C0040128|T047|IS|14304000|SNOMEDCT_CORE|Thyroid disorder, NOS|Disorder of thyroid gland
C0040136|T191|FN|127018007|SNOMEDCT_CORE|Neoplasm of thyroid gland|Neoplasm of thyroid gland
C0040136|T191|PT|127018007|SNOMEDCT_CORE|Neoplasm of thyroid gland|Neoplasm of thyroid gland
C0040136|T191|SY|127018007|SNOMEDCT_CORE|Thyroid tumor|Neoplasm of thyroid gland
C0040136|T191|SYGB|127018007|SNOMEDCT_CORE|Thyroid tumour|Neoplasm of thyroid gland
C0040136|T191|SY|127018007|SNOMEDCT_CORE|Tumor of thyroid gland|Neoplasm of thyroid gland
C0040136|T191|SYGB|127018007|SNOMEDCT_CORE|Tumour of thyroid gland|Neoplasm of thyroid gland
C0040137|T191|PT|237495005|SNOMEDCT_CORE|Thyroid nodule|Thyroid nodule
C0040137|T191|FN|237495005|SNOMEDCT_CORE|Thyroid nodule|Thyroid nodule
C0040147|T047|PT|82119001|SNOMEDCT_CORE|Thyroiditis|Thyroiditis
C0040147|T047|FN|82119001|SNOMEDCT_CORE|Thyroiditis|Thyroiditis
C0040147|T047|IS|82119001|SNOMEDCT_CORE|Thyroiditis, NOS|Thyroiditis
C0040156|T047|PT|90739004|SNOMEDCT_CORE|Thyrotoxicosis|Thyrotoxicosis
C0040156|T047|FN|90739004|SNOMEDCT_CORE|Thyrotoxicosis|Thyrotoxicosis
C0040156|T047|IS|90739004|SNOMEDCT_CORE|Thyrotoxicosis, NOS|Thyrotoxicosis
C0040185|T037|PT|31978002|SNOMEDCT_CORE|Fracture of tibia|Fracture of tibia
C0040185|T037|FN|31978002|SNOMEDCT_CORE|Fracture of tibia|Fracture of tibia
C0040185|T037|IS|31978002|SNOMEDCT_CORE|Fracture of tibia, NOS|Fracture of tibia
C0040188|T048|PT|568005|SNOMEDCT_CORE|Tic disorder|Tic disorder
C0040188|T048|FN|568005|SNOMEDCT_CORE|Tic disorder|Tic disorder
C0040188|T048|IS|568005|SNOMEDCT_CORE|Tic disorder, NOS|Tic disorder
C0040213|T047|PT|64109004|SNOMEDCT_CORE|Costal chondritis|Tietze's disease
C0040213|T047|FN|64109004|SNOMEDCT_CORE|Costal chondritis|Tietze's disease
C0040213|T047|OF|64109004|SNOMEDCT_CORE|Costalchondritis|Tietze's disease
C0040213|T047|IS|64109004|SNOMEDCT_CORE|Costalchondritis|Tietze's disease
C0040213|T047|IS|64109004|SNOMEDCT_CORE|Costalchondritis, NOS|Tietze's disease
C0040213|T047|SY|30128009|SNOMEDCT_CORE|Costochondral junction syndrome|Tietze's disease
C0040213|T047|SY|64109004|SNOMEDCT_CORE|Costochondritis|Tietze's disease
C0040213|T047|IS|64109004|SNOMEDCT_CORE|Costochondritis, NOS|Tietze's disease
C0040213|T047|SY|30128009|SNOMEDCT_CORE|Cyriax's syndrome|Tietze's disease
C0040213|T047|SY|30128009|SNOMEDCT_CORE|Peristernal perichondritis|Tietze's disease
C0040213|T047|SY|30128009|SNOMEDCT_CORE|Slipping rib syndrome|Tietze's disease
C0040213|T047|SY|30128009|SNOMEDCT_CORE|Tietze disease|Tietze's disease
C0040213|T047|PT|30128009|SNOMEDCT_CORE|Tietze's disease|Tietze's disease
C0040213|T047|FN|30128009|SNOMEDCT_CORE|Tietze's disease|Tietze's disease
C0040213|T047|SY|30128009|SNOMEDCT_CORE|Tietze's syndrome|Tietze's disease
C0040247|T047|SY|47382004|SNOMEDCT_CORE|Microsporic tinea|Tinea
C0040247|T047|IS|47382004|SNOMEDCT_CORE|Microsporic tinea, NOS|Tinea
C0040247|T047|SY|47382004|SNOMEDCT_CORE|Ringworm|Tinea
C0040247|T047|IS|47382004|SNOMEDCT_CORE|Ringworm, NOS|Tinea
C0040247|T047|SY|47382004|SNOMEDCT_CORE|Tinea|Tinea
C0040247|T047|IS|47382004|SNOMEDCT_CORE|Tinea, NOS|Tinea
C0040250|T047|SY|5441008|SNOMEDCT_CORE|Black dot ringworm|Tinea capitis
C0040250|T047|SY|5441008|SNOMEDCT_CORE|Dermatophytosis of scalp|Tinea capitis
C0040250|T047|SY|5441008|SNOMEDCT_CORE|Ringworm of the scalp|Tinea capitis
C0040250|T047|PT|5441008|SNOMEDCT_CORE|Tinea capitis|Tinea capitis
C0040250|T047|FN|5441008|SNOMEDCT_CORE|Tinea capitis|Tinea capitis
C0040250|T047|SY|5441008|SNOMEDCT_CORE|Tinea of scalp|Tinea capitis
C0040252|T047|SY|84849002|SNOMEDCT_CORE|Body tinea|Tinea corporis
C0040252|T047|SY|84849002|SNOMEDCT_CORE|Herpes circinatus|Tinea corporis
C0040252|T047|SY|84849002|SNOMEDCT_CORE|Tinea circinata|Tinea corporis
C0040252|T047|SY|84849002|SNOMEDCT_CORE|Tinea circinatus|Tinea corporis
C0040252|T047|FN|84849002|SNOMEDCT_CORE|Tinea corporis|Tinea corporis
C0040252|T047|PT|84849002|SNOMEDCT_CORE|Tinea corporis|Tinea corporis
C0040259|T047|SY|6020002|SNOMEDCT_CORE|Athlete's foot|Tinea pedis
C0040259|T047|SY|6020002|SNOMEDCT_CORE|Dermatophytosis of foot|Tinea pedis
C0040259|T047|SY|6020002|SNOMEDCT_CORE|Epidermophytosis pedis|Tinea pedis
C0040259|T047|SY|6020002|SNOMEDCT_CORE|Ringworm of foot|Tinea pedis
C0040259|T047|PT|6020002|SNOMEDCT_CORE|Tinea pedis|Tinea pedis
C0040259|T047|FN|6020002|SNOMEDCT_CORE|Tinea pedis|Tinea pedis
C0040259|T047|SY|6020002|SNOMEDCT_CORE|TP - Tinea pedis|Tinea pedis
C0040261|T047|SY|414941008|SNOMEDCT_CORE|Fungal infection of nail|Onychomycosis
C0040261|T047|PT|414941008|SNOMEDCT_CORE|Onychomycosis|Onychomycosis
C0040261|T047|FN|414941008|SNOMEDCT_CORE|Onychomycosis|Onychomycosis
C0040261|T047|SY|414941008|SNOMEDCT_CORE|Ringworm of nail|Onychomycosis
C0040261|T047|IS|414941008|SNOMEDCT_CORE|Tinea unguium|Onychomycosis
C0040262|T047|PT|56454009|SNOMEDCT_CORE|Pityriasis versicolor|Pityriasis versicolor
C0040262|T047|FN|56454009|SNOMEDCT_CORE|Pityriasis versicolor|Pityriasis versicolor
C0040262|T047|SY|56454009|SNOMEDCT_CORE|PV - Pityriasis versicolor|Pityriasis versicolor
C0040262|T047|SY|56454009|SNOMEDCT_CORE|Tinea flava|Pityriasis versicolor
C0040262|T047|SY|56454009|SNOMEDCT_CORE|Tinea versicolor|Pityriasis versicolor
C0040262|T047|SY|56454009|SNOMEDCT_CORE|Tinea versicolor due to Malassezia furfur|Pityriasis versicolor
C0040262|T047|SY|56454009|SNOMEDCT_CORE|Tinea versicolor due to Pityrosporum furfur|Pityriasis versicolor
C0040262|T047|SY|56454009|SNOMEDCT_CORE|TV - Tinea versicolor|Pityriasis versicolor
C0040264|T047|SY|60862001|SNOMEDCT_CORE|Noise in ears|Tinnitus
C0040264|T047|SY|60862001|SNOMEDCT_CORE|Ringing in ears|Tinnitus
C0040264|T047|PT|60862001|SNOMEDCT_CORE|Tinnitus|Tinnitus
C0040264|T047|FN|60862001|SNOMEDCT_CORE|Tinnitus|Tinnitus
C0040264|T047|IS|60862001|SNOMEDCT_CORE|Tinnitus, NOS|Tinnitus
C0040332|T048|SY|89765005|SNOMEDCT_CORE|Compulsive tobacco user syndrome|Tobacco dependence syndrome
C0040332|T048|SY|89765005|SNOMEDCT_CORE|Tobacco dependence|Tobacco dependence syndrome
C0040332|T048|PT|89765005|SNOMEDCT_CORE|Tobacco dependence syndrome|Tobacco dependence syndrome
C0040332|T048|FN|89765005|SNOMEDCT_CORE|Tobacco dependence syndrome|Tobacco dependence syndrome
C0040336|T048|SY|89765005|SNOMEDCT_CORE|Tobacco abuse|Tobacco abuse
C0040425|T047|PT|90176007|SNOMEDCT_CORE|Tonsillitis|Tonsillitis
C0040425|T047|FN|90176007|SNOMEDCT_CORE|Tonsillitis|Tonsillitis
C0040425|T047|IS|90176007|SNOMEDCT_CORE|Tonsillitis, NOS|Tonsillitis
C0040433|T033|PT|12351004|SNOMEDCT_CORE|Crowding of teeth|Crowding of teeth
C0040433|T033|FN|12351004|SNOMEDCT_CORE|Crowding of teeth|Crowding of teeth
C0040433|T033|SY|12351004|SNOMEDCT_CORE|Imbrication of teeth|Crowding of teeth
C0040435|T047|SY|234947003|SNOMEDCT_CORE|Disease of teeth|Tooth disorder
C0040435|T047|SY|234947003|SNOMEDCT_CORE|Tooth disease|Tooth disorder
C0040435|T047|PT|234947003|SNOMEDCT_CORE|Tooth disorder|Tooth disorder
C0040435|T047|FN|234947003|SNOMEDCT_CORE|Tooth disorder|Tooth disorder
C0040441|T037|SY|36202009|SNOMEDCT_CORE|Broken teeth|Fracture of tooth
C0040441|T037|SY|36202009|SNOMEDCT_CORE|Broken tooth|Fracture of tooth
C0040441|T037|SY|36202009|SNOMEDCT_CORE|BT - Broken tooth|Fracture of tooth
C0040441|T037|SY|36202009|SNOMEDCT_CORE|Chipped tooth|Fracture of tooth
C0040441|T037|PT|36202009|SNOMEDCT_CORE|Fracture of tooth|Fracture of tooth
C0040441|T037|FN|36202009|SNOMEDCT_CORE|Fracture of tooth|Fracture of tooth
C0040441|T037|SY|36202009|SNOMEDCT_CORE|Fractured tooth|Fracture of tooth
C0040441|T037|SY|36202009|SNOMEDCT_CORE|Tooth fracture|Fracture of tooth
C0040456|T047|SY|235104008|SNOMEDCT_CORE|Impacted teeth|Impacted tooth
C0040456|T047|PT|235104008|SNOMEDCT_CORE|Impacted tooth|Impacted tooth
C0040456|T047|FN|235104008|SNOMEDCT_CORE|Impacted tooth|Impacted tooth
C0040456|T047|SY|235104008|SNOMEDCT_CORE|Impacted tooth - disorder|Impacted tooth
C0040457|T033|IS|367534004|SNOMEDCT_CORE|Supernumerary teeth|Supernumerary tooth
C0040457|T033|OF|367534004|SNOMEDCT_CORE|Supernumerary teeth|Supernumerary tooth
C0040457|T033|PT|367534004|SNOMEDCT_CORE|Supernumerary tooth|Supernumerary tooth
C0040457|T033|FN|367534004|SNOMEDCT_CORE|Supernumerary tooth|Supernumerary tooth
C0040457|T033|SY|367534004|SNOMEDCT_CORE|Supplemental tooth|Supernumerary tooth
C0040460|T184|SY|27355003|SNOMEDCT_CORE|Dentagra|Toothache
C0040460|T184|SY|27355003|SNOMEDCT_CORE|Dentalgia|Toothache
C0040460|T184|SY|27355003|SNOMEDCT_CORE|Odontalgia|Toothache
C0040460|T184|SY|27355003|SNOMEDCT_CORE|Pain in tooth|Toothache
C0040460|T184|PT|27355003|SNOMEDCT_CORE|Toothache|Toothache
C0040460|T184|FN|27355003|SNOMEDCT_CORE|Toothache|Toothache
C0040485|T184|SY|70070008|SNOMEDCT_CORE|Contracture of neck|Torticollis
C0040485|T184|IS|70070008|SNOMEDCT_CORE|Contracture of neck, NOS|Torticollis
C0040485|T184|PT|70070008|SNOMEDCT_CORE|Torticollis|Torticollis
C0040485|T184|FN|70070008|SNOMEDCT_CORE|Torticollis|Torticollis
C0040485|T184|IS|70070008|SNOMEDCT_CORE|Torticollis, NOS|Torticollis
C0040485|T184|SY|70070008|SNOMEDCT_CORE|Wry neck|Torticollis
C0040517|T047|SY|5158005|SNOMEDCT_CORE|Combined vocal and multiple motor tic disorder|Gilles de la Tourette's syndrome
C0040517|T047|SY|5158005|SNOMEDCT_CORE|Gilles de la Tourette syndrome|Gilles de la Tourette's syndrome
C0040517|T047|PT|5158005|SNOMEDCT_CORE|Gilles de la Tourette's syndrome|Gilles de la Tourette's syndrome
C0040517|T047|FN|5158005|SNOMEDCT_CORE|Gilles de la Tourette's syndrome|Gilles de la Tourette's syndrome
C0040517|T047|SY|5158005|SNOMEDCT_CORE|Gilles de la Tourettes syndrome|Gilles de la Tourette's syndrome
C0040517|T047|SY|5158005|SNOMEDCT_CORE|Tourette's disorder|Gilles de la Tourette's syndrome
C0040517|T047|SY|5158005|SNOMEDCT_CORE|Tourette's syndrome|Gilles de la Tourette's syndrome
C0040583|T047|PT|11296007|SNOMEDCT_CORE|Stenosis of trachea|Stenosis of trachea
C0040583|T047|FN|11296007|SNOMEDCT_CORE|Stenosis of trachea|Stenosis of trachea
C0040583|T047|SY|11296007|SNOMEDCT_CORE|Tracheal stenosis|Stenosis of trachea
C0040583|T047|IS|11296007|SNOMEDCT_CORE|Tracheal stricture|Stenosis of trachea
C0040701|T048|SY|17226007|SNOMEDCT_CORE|Adjustment reaction|Adjustment reaction
C0040701|T048|IS|17226007|SNOMEDCT_CORE|Adjustment reaction, NOS|Adjustment reaction
C0040761|T019|SY|26146002|SNOMEDCT_CORE|Classical transposition of great vessels|Complete transposition of great vessels
C0040761|T019|SY|26146002|SNOMEDCT_CORE|Complete TGA|Complete transposition of great vessels
C0040761|T019|IS|26146002|SNOMEDCT_CORE|Complete transposition of great arteries|Complete transposition of great vessels
C0040761|T019|PT|26146002|SNOMEDCT_CORE|Complete transposition of great vessels|Complete transposition of great vessels
C0040761|T019|FN|26146002|SNOMEDCT_CORE|Complete transposition of great vessels|Complete transposition of great vessels
C0040761|T019|SY|26146002|SNOMEDCT_CORE|Total great vessel transposition|Complete transposition of great vessels
C0040761|T019|SY|26146002|SNOMEDCT_CORE|Transposition of the great arteries|Complete transposition of great vessels
C0040822|T184|SY|26079004|SNOMEDCT_CORE|Has a tremor|Tremor
C0040822|T184|SY|26079004|SNOMEDCT_CORE|Shakes|Tremor
C0040822|T184|SY|26079004|SNOMEDCT_CORE|Shaking|Tremor
C0040822|T184|SY|26079004|SNOMEDCT_CORE|Shaking all over|Tremor
C0040822|T184|SY|26079004|SNOMEDCT_CORE|The shakes|Tremor
C0040822|T184|PT|26079004|SNOMEDCT_CORE|Tremor|Tremor
C0040822|T184|FN|26079004|SNOMEDCT_CORE|Tremor|Tremor
C0040822|T184|IS|26079004|SNOMEDCT_CORE|Tremor, NOS|Tremor
C0040843|T047|SY|76272004|SNOMEDCT_CORE|Treponemal disease|Treponemal disease
C0040843|T047|SY|76272004|SNOMEDCT_CORE|Treponemal infection|Treponemal disease
C0040921|T047|PT|56335008|SNOMEDCT_CORE|Infection by Trichomonas|Infection by Trichomonas
C0040921|T047|OF|56335008|SNOMEDCT_CORE|Infection by Trichomonas|Infection by Trichomonas
C0040921|T047|IS|56335008|SNOMEDCT_CORE|Infection by Trichomonas, NOS|Infection by Trichomonas
C0040921|T047|FN|56335008|SNOMEDCT_CORE|Infection caused by Trichomonas|Infection by Trichomonas
C0040921|T047|SY|56335008|SNOMEDCT_CORE|Infection caused by Trichomonas|Infection by Trichomonas
C0040921|T047|SY|56335008|SNOMEDCT_CORE|Trichomonas infection|Infection by Trichomonas
C0040921|T047|SY|56335008|SNOMEDCT_CORE|Trichomoniasis|Infection by Trichomonas
C0040921|T047|SY|56335008|SNOMEDCT_CORE|Trichomonosis|Infection by Trichomonas
C0040923|T047|SY|276877003|SNOMEDCT_CORE|Trichomonal fluor vaginalis|Trichomonal vaginitis
C0040923|T047|SY|276877003|SNOMEDCT_CORE|Trichomonal leukorrhea vaginalis|Trichomonal vaginitis
C0040923|T047|SYGB|276877003|SNOMEDCT_CORE|Trichomonal leukorrhoea vaginalis|Trichomonal vaginitis
C0040923|T047|PT|276877003|SNOMEDCT_CORE|Trichomonal vaginitis|Trichomonal vaginitis
C0040923|T047|FN|276877003|SNOMEDCT_CORE|Trichomonal vaginitis|Trichomonal vaginitis
C0040923|T047|SY|276877003|SNOMEDCT_CORE|Vaginal trichomoniasis|Trichomonal vaginitis
C0040953|T048|SY|17155009|SNOMEDCT_CORE|Hair plucking|Trichotillomania
C0040953|T048|SY|17155009|SNOMEDCT_CORE|Trichologia|Trichotillomania
C0040953|T048|PT|17155009|SNOMEDCT_CORE|Trichotillomania|Trichotillomania
C0040953|T048|FN|17155009|SNOMEDCT_CORE|Trichotillomania|Trichotillomania
C0040961|T047|SY|111287006|SNOMEDCT_CORE|TI - Tricuspid incompetence|Tricuspid valve regurgitation
C0040961|T047|SY|111287006|SNOMEDCT_CORE|TR - Tricuspid regurgitation|Tricuspid valve regurgitation
C0040961|T047|SY|111287006|SNOMEDCT_CORE|Tricuspid insufficiency|Tricuspid valve regurgitation
C0040961|T047|SY|111287006|SNOMEDCT_CORE|Tricuspid regurgitation|Tricuspid valve regurgitation
C0040961|T047|IS|111287006|SNOMEDCT_CORE|Tricuspid regurgitation, NOS|Tricuspid valve regurgitation
C0040961|T047|SY|111287006|SNOMEDCT_CORE|Tricuspid valve incompetence|Tricuspid valve regurgitation
C0040961|T047|IS|111287006|SNOMEDCT_CORE|Tricuspid valve incompetence, NOS|Tricuspid valve regurgitation
C0040961|T047|SY|111287006|SNOMEDCT_CORE|Tricuspid valve insufficiency|Tricuspid valve regurgitation
C0040961|T047|IS|111287006|SNOMEDCT_CORE|Tricuspid valve insufficiency, NOS|Tricuspid valve regurgitation
C0040961|T047|PT|111287006|SNOMEDCT_CORE|Tricuspid valve regurgitation|Tricuspid valve regurgitation
C0040961|T047|FN|111287006|SNOMEDCT_CORE|Tricuspid valve regurgitation|Tricuspid valve regurgitation
C0040961|T047|IS|111287006|SNOMEDCT_CORE|Tricuspid valve regurgitation, NOS|Tricuspid valve regurgitation
C0040997|T047|SY|31681005|SNOMEDCT_CORE|Fothergill's neuralgia|Trigeminal neuralgia
C0040997|T047|SY|31681005|SNOMEDCT_CORE|Tic douloureux|Trigeminal neuralgia
C0040997|T047|SY|31681005|SNOMEDCT_CORE|TN - Trigeminal neuralgia|Trigeminal neuralgia
C0040997|T047|SY|31681005|SNOMEDCT_CORE|Trifacial neuralgia|Trigeminal neuralgia
C0040997|T047|PT|31681005|SNOMEDCT_CORE|Trigeminal neuralgia|Trigeminal neuralgia
C0040997|T047|FN|31681005|SNOMEDCT_CORE|Trigeminal neuralgia|Trigeminal neuralgia
C0040997|T047|IS|31681005|SNOMEDCT_CORE|Trigeminal neuralgia, NOS|Trigeminal neuralgia
C0041296|T047|IS|56717001|SNOMEDCT_CORE|Infection due to Mycobacterium tuberculosis|Tuberculosis
C0041296|T047|IS|56717001|SNOMEDCT_CORE|MTB - Mycobacterium tuberculosis infection|Tuberculosis
C0041296|T047|IS|56717001|SNOMEDCT_CORE|Mycobacterium tuberculosis infection|Tuberculosis
C0041296|T047|SY|56717001|SNOMEDCT_CORE|TB - Tuberculosis|Tuberculosis
C0041296|T047|PT|56717001|SNOMEDCT_CORE|Tuberculosis|Tuberculosis
C0041296|T047|FN|56717001|SNOMEDCT_CORE|Tuberculosis|Tuberculosis
C0041296|T047|IS|56717001|SNOMEDCT_CORE|Tuberculosis, NOS|Tuberculosis
C0041316|T047|SY|10893003|SNOMEDCT_CORE|Tuberculosis of lymph node|Tuberculous adenitis
C0041316|T047|PT|10893003|SNOMEDCT_CORE|Tuberculous adenitis|Tuberculous adenitis
C0041316|T047|FN|10893003|SNOMEDCT_CORE|Tuberculous adenitis|Tuberculous adenitis
C0041316|T047|IS|10893003|SNOMEDCT_CORE|Tuberculous adenitis, NOS|Tuberculous adenitis
C0041316|T047|SY|10893003|SNOMEDCT_CORE|Tuberculous lymphadenopathy|Tuberculous adenitis
C0041318|T047|SY|58437007|SNOMEDCT_CORE|TB - Tuberculous meningitis|Tuberculosis of meninges
C0041318|T047|SY|58437007|SNOMEDCT_CORE|TBM - Tuberculous meningitis|Tuberculosis of meninges
C0041318|T047|PT|58437007|SNOMEDCT_CORE|Tuberculosis of meninges|Tuberculosis of meninges
C0041318|T047|FN|58437007|SNOMEDCT_CORE|Tuberculosis of meninges|Tuberculosis of meninges
C0041318|T047|SY|58437007|SNOMEDCT_CORE|Tuberculous meningitis|Tuberculosis of meninges
C0041321|T047|PT|47604008|SNOMEDCT_CORE|Miliary tuberculosis|Miliary tuberculosis
C0041321|T047|FN|47604008|SNOMEDCT_CORE|Miliary tuberculosis|Miliary tuberculosis
C0041321|T047|IS|47604008|SNOMEDCT_CORE|Miliary tuberculosis, NOS|Miliary tuberculosis
C0041321|T047|SY|47604008|SNOMEDCT_CORE|MTB - Miliary tuberculosis|Miliary tuberculosis
C0041326|T047|PT|186182003|SNOMEDCT_CORE|Tuberculosis of pleura|Tuberculosis of pleura
C0041326|T047|FN|186182003|SNOMEDCT_CORE|Tuberculosis of pleura|Tuberculosis of pleura
C0041326|T047|SY|186182003|SNOMEDCT_CORE|Tuberculous pleurisy|Tuberculosis of pleura
C0041326|T047|SY|186182003|SNOMEDCT_CORE|Tuberculous pleuritis|Tuberculosis of pleura
C0041327|T047|SY|154283005|SNOMEDCT_CORE|PTB - Pulmonary tuberculosis|Pulmonary tuberculosis
C0041327|T047|OF|154283005|SNOMEDCT_CORE|Pulmonary tuberculosis|Pulmonary tuberculosis
C0041327|T047|PT|154283005|SNOMEDCT_CORE|Pulmonary tuberculosis|Pulmonary tuberculosis
C0041327|T047|FN|154283005|SNOMEDCT_CORE|Pulmonary tuberculosis|Pulmonary tuberculosis
C0041327|T047|SY|154283005|SNOMEDCT_CORE|TB - Pulmonary tuberculosis|Pulmonary tuberculosis
C0041330|T047|SY|35984006|SNOMEDCT_CORE|Pott's disease|Tuberculosis of vertebral column
C0041330|T047|PT|35984006|SNOMEDCT_CORE|Tuberculosis of vertebral column|Tuberculosis of vertebral column
C0041330|T047|FN|35984006|SNOMEDCT_CORE|Tuberculosis of vertebral column|Tuberculosis of vertebral column
C0041330|T047|SY|35984006|SNOMEDCT_CORE|Tuberculosis of vertebral column - Pott's|Tuberculosis of vertebral column
C0041330|T047|SY|35984006|SNOMEDCT_CORE|Tuberculous spondylitis|Tuberculosis of vertebral column
C0041341|T191|SY|7199000|SNOMEDCT_CORE|Adenoma sebaceum syndrome|Tuberous sclerosis syndrome
C0041341|T191|SY|7199000|SNOMEDCT_CORE|Bourneville's disease|Tuberous sclerosis syndrome
C0041341|T191|SY|7199000|SNOMEDCT_CORE|Epiloia|Tuberous sclerosis syndrome
C0041341|T191|SY|7199000|SNOMEDCT_CORE|TS - Tuberous sclerosis|Tuberous sclerosis syndrome
C0041341|T191|SY|7199000|SNOMEDCT_CORE|Tuberous sclerosis|Tuberous sclerosis syndrome
C0041341|T191|PT|7199000|SNOMEDCT_CORE|Tuberous sclerosis syndrome|Tuberous sclerosis syndrome
C0041341|T191|FN|7199000|SNOMEDCT_CORE|Tuberous sclerosis syndrome|Tuberous sclerosis syndrome
C0041343|T047|SY|58949002|SNOMEDCT_CORE|Tubo ovarian abscess|Tubo-ovarian abscess
C0041343|T047|PT|58949002|SNOMEDCT_CORE|Tubo-ovarian abscess|Tubo-ovarian abscess
C0041343|T047|FN|58949002|SNOMEDCT_CORE|Tubo-ovarian abscess|Tubo-ovarian abscess
C0041349|T047|SY|428255004|SNOMEDCT_CORE|Interstitial nephritis|Tubulointerstitial nephritis
C0041349|T047|OAS|28689008|SNOMEDCT_CORE|Renal tubulo-interstitial disease|Tubulointerstitial nephritis
C0041349|T047|SY|428255004|SNOMEDCT_CORE|Renal tubulo-interstitial disease|Tubulointerstitial nephritis
C0041349|T047|OAS|28689008|SNOMEDCT_CORE|T.I.N.|Tubulointerstitial nephritis
C0041349|T047|IS|28689008|SNOMEDCT_CORE|T.I.N., NOS|Tubulointerstitial nephritis
C0041349|T047|SY|428255004|SNOMEDCT_CORE|Tubulo-interstitial nephritis|Tubulointerstitial nephritis
C0041349|T047|PT|428255004|SNOMEDCT_CORE|Tubulointerstitial nephritis|Tubulointerstitial nephritis
C0041349|T047|FN|428255004|SNOMEDCT_CORE|Tubulointerstitial nephritis|Tubulointerstitial nephritis
C0041349|T047|OAS|28689008|SNOMEDCT_CORE|Tubulointerstitial nephropathy|Tubulointerstitial nephritis
C0041349|T047|SY|428255004|SNOMEDCT_CORE|Tubulointerstitial nephropathy|Tubulointerstitial nephritis
C0041349|T047|IS|28689008|SNOMEDCT_CORE|Tubulointerstitial nephropathy, NOS|Tubulointerstitial nephritis
C0041408|T047|IS|38804009|SNOMEDCT_CORE|45, X syndrome|Turner syndrome
C0041408|T047|IS|38804009|SNOMEDCT_CORE|45X0 - Turner's syndrome|Turner syndrome
C0041408|T047|IS|38804009|SNOMEDCT_CORE|Karyotype 45, X|Turner syndrome
C0041408|T047|SY|38804009|SNOMEDCT_CORE|Pterygolymphangiectasia syndrome|Turner syndrome
C0041408|T047|SY|38804009|SNOMEDCT_CORE|TS - Turner's syndrome|Turner syndrome
C0041408|T047|PT|38804009|SNOMEDCT_CORE|Turner syndrome|Turner syndrome
C0041408|T047|FN|38804009|SNOMEDCT_CORE|Turner syndrome|Turner syndrome
C0041408|T047|IS|38804009|SNOMEDCT_CORE|Turner syndrome, NOS|Turner syndrome
C0041408|T047|SY|38804009|SNOMEDCT_CORE|Turner's syndrome|Turner syndrome
C0041408|T047|IS|38804009|SNOMEDCT_CORE|X0 - Turner's syndrome|Turner syndrome
C0041408|T047|IS|38804009|SNOMEDCT_CORE|XO syndrome|Turner syndrome
C0041466|T047|SY|4834000|SNOMEDCT_CORE|Infection by Salmonella Typhi|Typhoid fever
C0041466|T047|IS|4834000|SNOMEDCT_CORE|Infection by Salmonella typhi|Typhoid fever
C0041466|T047|PT|4834000|SNOMEDCT_CORE|Typhoid fever|Typhoid fever
C0041466|T047|FN|4834000|SNOMEDCT_CORE|Typhoid fever|Typhoid fever
C0041601|T037|PT|54556006|SNOMEDCT_CORE|Fracture of ulna|Fracture of ulna
C0041601|T037|FN|54556006|SNOMEDCT_CORE|Fracture of ulna|Fracture of ulna
C0041601|T037|IS|54556006|SNOMEDCT_CORE|Fracture of ulna, NOS|Fracture of ulna
C0041657|T033|SY|418107008|SNOMEDCT_CORE|Mental status, unconsciousness|Unconscious
C0041657|T033|PT|418107008|SNOMEDCT_CORE|Unconscious|Unconscious
C0041657|T033|FN|418107008|SNOMEDCT_CORE|Unconscious|Unconscious
C0041657|T033|SY|418107008|SNOMEDCT_CORE|Unconsciousness|Unconscious
C0041667|T033|SY|248342006|SNOMEDCT_CORE|Low body weight|Underweight
C0041667|T033|SY|248342006|SNOMEDCT_CORE|Patient underweight|Underweight
C0041667|T033|PT|248342006|SNOMEDCT_CORE|Underweight|Underweight
C0041667|T033|FN|248342006|SNOMEDCT_CORE|Underweight|Underweight
C0041674|T033|SY|73438004|SNOMEDCT_CORE|Out of work|Unemployed
C0041674|T033|SY|73438004|SNOMEDCT_CORE|U/E - Unemployed|Unemployed
C0041674|T033|SY|73438004|SNOMEDCT_CORE|UE - Unemployed|Unemployed
C0041674|T033|PT|73438004|SNOMEDCT_CORE|Unemployed|Unemployed
C0041674|T033|FN|73438004|SNOMEDCT_CORE|Unemployed|Unemployed
C0041674|T033|IS|73438004|SNOMEDCT_CORE|Unemployment|Unemployed
C0041674|T033|SY|73438004|SNOMEDCT_CORE|Without employment|Unemployed
C0041747|T033|SY|83074005|SNOMEDCT_CORE|Accidental pregnancy|Unplanned pregnancy
C0041747|T033|IS|83074005|SNOMEDCT_CORE|Unintended pregnancy|Unplanned pregnancy
C0041747|T033|PT|83074005|SNOMEDCT_CORE|Unplanned pregnancy|Unplanned pregnancy
C0041747|T033|FN|83074005|SNOMEDCT_CORE|Unplanned pregnancy|Unplanned pregnancy
C0041755|T046|SY|62014003|SNOMEDCT_CORE|ADR - Adverse drug reaction|Adverse reaction to drug
C0041755|T046|SY|62014003|SNOMEDCT_CORE|Adverse drug effect|Adverse reaction to drug
C0041755|T046|IS|62014003|SNOMEDCT_CORE|Adverse drug effect, NOS|Adverse reaction to drug
C0041755|T046|SY|62014003|SNOMEDCT_CORE|Adverse drug reaction|Adverse reaction to drug
C0041755|T046|IS|62014003|SNOMEDCT_CORE|Adverse drug reaction, NOS|Adverse reaction to drug
C0041755|T046|SY|62014003|SNOMEDCT_CORE|Adverse reaction caused by drug|Adverse reaction to drug
C0041755|T046|FN|62014003|SNOMEDCT_CORE|Adverse reaction caused by drug|Adverse reaction to drug
C0041755|T046|PT|62014003|SNOMEDCT_CORE|Adverse reaction to drug|Adverse reaction to drug
C0041755|T046|OF|62014003|SNOMEDCT_CORE|Adverse reaction to drug|Adverse reaction to drug
C0041755|T046|SY|62014003|SNOMEDCT_CORE|Adverse reaction to medication|Adverse reaction to drug
C0041755|T046|SY|62014003|SNOMEDCT_CORE|Drug reaction|Adverse reaction to drug
C0041755|T046|IS|62014003|SNOMEDCT_CORE|Drug reaction, NOS|Adverse reaction to drug
C0041782|T047|PTGB|267513007|SNOMEDCT_CORE|Deficiency anaemias|Deficiency anemias
C0041782|T047|PT|267513007|SNOMEDCT_CORE|Deficiency anemias|Deficiency anemias
C0041782|T047|FN|267513007|SNOMEDCT_CORE|Deficiency anemias|Deficiency anemias
C0041785|T047|SY|81573002|SNOMEDCT_CORE|Diffuse disease of connective tissue|Diffuse disease of connective tissue
C0041785|T047|IS|81573002|SNOMEDCT_CORE|Diffuse disease of connective tissue, NOS|Diffuse disease of connective tissue
C0041834|T047|PT|247441003|SNOMEDCT_CORE|Erythema|Erythema
C0041834|T047|FN|247441003|SNOMEDCT_CORE|Erythema|Erythema
C0041834|T047|SY|247441003|SNOMEDCT_CORE|Erythema - observation|Erythema
C0041834|T047|IS|247441003|SNOMEDCT_CORE|Injection|Erythema
C0041834|T047|IS|247441003|SNOMEDCT_CORE|Red skin|Erythema
C0041844|T020|PTGB|82985000|SNOMEDCT_CORE|Haemorrhoids without complication|Hemorrhoids without complication
C0041844|T020|PT|82985000|SNOMEDCT_CORE|Hemorrhoids without complication|Hemorrhoids without complication
C0041844|T020|FN|82985000|SNOMEDCT_CORE|Hemorrhoids without complication|Hemorrhoids without complication
C0041909|T046|PT|37372002|SNOMEDCT_CORE|Upper gastrointestinal bleeding|Upper gastrointestinal bleeding
C0041909|T046|SYGB|37372002|SNOMEDCT_CORE|Upper gastrointestinal haemorrhage|Upper gastrointestinal bleeding
C0041909|T046|SY|37372002|SNOMEDCT_CORE|Upper gastrointestinal hemorrhage|Upper gastrointestinal bleeding
C0041909|T046|FN|37372002|SNOMEDCT_CORE|Upper gastrointestinal hemorrhage|Upper gastrointestinal bleeding
C0041909|T046|SYGB|37372002|SNOMEDCT_CORE|Upper GI - gastrointestinal haemorrhage|Upper gastrointestinal bleeding
C0041909|T046|SY|37372002|SNOMEDCT_CORE|Upper GI - gastrointestinal hemorrhage|Upper gastrointestinal bleeding
C0041909|T046|SY|37372002|SNOMEDCT_CORE|Upper GI bleeding|Upper gastrointestinal bleeding
C0041909|T046|SYGB|37372002|SNOMEDCT_CORE|Upper GI haemorrhage|Upper gastrointestinal bleeding
C0041909|T046|SY|37372002|SNOMEDCT_CORE|Upper GI hemorrhage|Upper gastrointestinal bleeding
C0041912|T047|PT|54150009|SNOMEDCT_CORE|Upper respiratory infection|Upper respiratory infection
C0041912|T047|FN|54150009|SNOMEDCT_CORE|Upper respiratory infection|Upper respiratory infection
C0041912|T047|IS|54150009|SNOMEDCT_CORE|Upper respiratory infection, NOS|Upper respiratory infection
C0041912|T047|SY|54150009|SNOMEDCT_CORE|Upper respiratory tract infection|Upper respiratory infection
C0041912|T047|SY|54150009|SNOMEDCT_CORE|URI - Upper respiratory infection|Upper respiratory infection
C0041912|T047|SY|54150009|SNOMEDCT_CORE|URTI - Infection of the upper respiratory tract|Upper respiratory infection
C0041948|T047|PTGB|44730006|SNOMEDCT_CORE|Uraemia|Uremia
C0041948|T047|IS|44730006|SNOMEDCT_CORE|Uraemia, NOS|Uremia
C0041948|T047|PT|44730006|SNOMEDCT_CORE|Uremia|Uremia
C0041948|T047|FN|44730006|SNOMEDCT_CORE|Uremia|Uremia
C0041948|T047|IS|44730006|SNOMEDCT_CORE|Uremia, NOS|Uremia
C0041952|T047|SY|31054009|SNOMEDCT_CORE|Calculus of ureter|Ureteric stone
C0041952|T047|SY|31054009|SNOMEDCT_CORE|Ureteral calculus|Ureteric stone
C0041952|T047|SY|31054009|SNOMEDCT_CORE|Ureteral stone|Ureteric stone
C0041952|T047|SY|31054009|SNOMEDCT_CORE|Ureteric calculus|Ureteric stone
C0041952|T047|PT|31054009|SNOMEDCT_CORE|Ureteric stone|Ureteric stone
C0041952|T047|FN|31054009|SNOMEDCT_CORE|Ureteric stone|Ureteric stone
C0041952|T047|SY|31054009|SNOMEDCT_CORE|Ureterolithiasis|Ureteric stone
C0041956|T047|IS|20018005|SNOMEDCT_CORE|Obstruction of ureter|Occlusion of ureter
C0041956|T047|PT|20018005|SNOMEDCT_CORE|Occlusion of ureter|Occlusion of ureter
C0041956|T047|FN|20018005|SNOMEDCT_CORE|Occlusion of ureter|Occlusion of ureter
C0041956|T047|IS|20018005|SNOMEDCT_CORE|Occlusion of ureter, NOS|Occlusion of ureter
C0041956|T047|IS|20018005|SNOMEDCT_CORE|Ureteral obstruction|Occlusion of ureter
C0041956|T047|IS|20018005|SNOMEDCT_CORE|Ureteric obstruction|Occlusion of ureter
C0041956|T047|IS|20018005|SNOMEDCT_CORE|Ureteric obstruction, NOS|Occlusion of ureter
C0041959|T047|SY|111405003|SNOMEDCT_CORE|Inflammation of ureter|Ureteritis
C0041959|T047|PT|111405003|SNOMEDCT_CORE|Ureteritis|Ureteritis
C0041959|T047|FN|111405003|SNOMEDCT_CORE|Ureteritis|Ureteritis
C0041959|T047|IS|111405003|SNOMEDCT_CORE|Ureteritis, NOS|Ureteritis
C0041970|T190|PT|14981000|SNOMEDCT_CORE|Urethral fistula|Urethral fistula
C0041970|T190|FN|14981000|SNOMEDCT_CORE|Urethral fistula|Urethral fistula
C0041970|T190|IS|14981000|SNOMEDCT_CORE|Urethral fistula, NOS|Urethral fistula
C0041976|T047|SY|31822004|SNOMEDCT_CORE|Inflammation of urethra|Urethritis
C0041976|T047|PT|31822004|SNOMEDCT_CORE|Urethritis|Urethritis
C0041976|T047|FN|31822004|SNOMEDCT_CORE|Urethritis|Urethritis
C0042023|T033|IS|162116003|SNOMEDCT_CORE|FOM - Frequency of micturition|Increased frequency of urination
C0042023|T033|IS|162116003|SNOMEDCT_CORE|Frequency of micturition|Increased frequency of urination
C0042023|T033|IS|162116003|SNOMEDCT_CORE|Frequency of urination|Increased frequency of urination
C0042023|T033|SY|162116003|SNOMEDCT_CORE|Increased frequency of micturition|Increased frequency of urination
C0042023|T033|PT|162116003|SNOMEDCT_CORE|Increased frequency of urination|Increased frequency of urination
C0042023|T033|FN|162116003|SNOMEDCT_CORE|Increased frequency of urination|Increased frequency of urination
C0042023|T033|SY|162116003|SNOMEDCT_CORE|Passes water too often|Increased frequency of urination
C0042023|T033|SY|162116003|SNOMEDCT_CORE|Pollakisuria|Increased frequency of urination
C0042023|T033|SY|162116003|SNOMEDCT_CORE|Pollakiuria|Increased frequency of urination
C0042023|T033|SY|162116003|SNOMEDCT_CORE|Urinary frequency|Increased frequency of urination
C0042024|T046|SY|165232002|SNOMEDCT_CORE|Absence of bladder continence|Urinary incontinence
C0042024|T046|SY|165232002|SNOMEDCT_CORE|Bladder incontinence|Urinary incontinence
C0042024|T046|SY|165232002|SNOMEDCT_CORE|Bladder: incontinent|Urinary incontinence
C0042024|T046|OF|165232002|SNOMEDCT_CORE|Bladder: incontinent|Urinary incontinence
C0042024|T046|SY|165232002|SNOMEDCT_CORE|Incontinence of urine|Urinary incontinence
C0042024|T046|SY|165232002|SNOMEDCT_CORE|Involuntary urination|Urinary incontinence
C0042024|T046|SY|165232002|SNOMEDCT_CORE|Lack of bladder control|Urinary incontinence
C0042024|T046|SY|165232002|SNOMEDCT_CORE|Leaking of urine|Urinary incontinence
C0042024|T046|SY|165232002|SNOMEDCT_CORE|Loss of bladder control|Urinary incontinence
C0042024|T046|SY|165232002|SNOMEDCT_CORE|UI - Urinary incontinence|Urinary incontinence
C0042024|T046|SY|165232002|SNOMEDCT_CORE|Unable to control bladder|Urinary incontinence
C0042024|T046|SY|165232002|SNOMEDCT_CORE|Unable to hold fluids|Urinary incontinence
C0042024|T046|SY|165232002|SNOMEDCT_CORE|Unable to hold urine|Urinary incontinence
C0042024|T046|SY|165232002|SNOMEDCT_CORE|Unable to prevent bladder emptying|Urinary incontinence
C0042024|T046|FN|165232002|SNOMEDCT_CORE|Urinary incontinence|Urinary incontinence
C0042024|T046|PT|165232002|SNOMEDCT_CORE|Urinary incontinence|Urinary incontinence
C0042024|T046|SY|165232002|SNOMEDCT_CORE|Urine incontinence|Urinary incontinence
C0042024|T046|SY|165232002|SNOMEDCT_CORE|Weak bladder|Urinary incontinence
C0042025|T047|PT|22220005|SNOMEDCT_CORE|Genuine stress incontinence|Genuine stress incontinence
C0042025|T047|FN|22220005|SNOMEDCT_CORE|Genuine stress incontinence|Genuine stress incontinence
C0042025|T047|SY|22220005|SNOMEDCT_CORE|GSI - Genuine stress incontinence|Genuine stress incontinence
C0042025|T047|SY|22220005|SNOMEDCT_CORE|Incontinence when straining|Genuine stress incontinence
C0042025|T047|SY|22220005|SNOMEDCT_CORE|SI - Stress incontinence|Genuine stress incontinence
C0042025|T047|SY|22220005|SNOMEDCT_CORE|Stress bladder incontinence|Genuine stress incontinence
C0042025|T047|IS|22220005|SNOMEDCT_CORE|Stress incontinence|Genuine stress incontinence
C0042025|T047|SY|22220005|SNOMEDCT_CORE|Stress urinary incontinence|Genuine stress incontinence
C0042025|T047|SY|22220005|SNOMEDCT_CORE|Urinary stress incontinence|Genuine stress incontinence
C0042029|T047|SY|68566005|SNOMEDCT_CORE|Urinary tract infection|Urinary tract infectious disease
C0042029|T047|IS|68566005|SNOMEDCT_CORE|Urinary tract infection, NOS|Urinary tract infectious disease
C0042029|T047|PT|68566005|SNOMEDCT_CORE|Urinary tract infectious disease|Urinary tract infectious disease
C0042029|T047|FN|68566005|SNOMEDCT_CORE|Urinary tract infectious disease|Urinary tract infectious disease
C0042029|T047|IS|68566005|SNOMEDCT_CORE|Urinary tract infectious disease, NOS|Urinary tract infectious disease
C0042029|T047|SY|68566005|SNOMEDCT_CORE|UTI - Urinary tract infection|Urinary tract infectious disease
C0042109|T047|PT|126485001|SNOMEDCT_CORE|Urticaria|Urticaria
C0042109|T047|FN|126485001|SNOMEDCT_CORE|Urticaria|Urticaria
C0042131|T047|IS|12337004|SNOMEDCT_CORE|Disease of uterus|Disorder of uterus
C0042131|T047|OF|12337004|SNOMEDCT_CORE|Disease of uterus|Disorder of uterus
C0042131|T047|IS|12337004|SNOMEDCT_CORE|Disease of uterus, NOS|Disorder of uterus
C0042131|T047|PT|12337004|SNOMEDCT_CORE|Disorder of uterus|Disorder of uterus
C0042131|T047|FN|12337004|SNOMEDCT_CORE|Disorder of uterus|Disorder of uterus
C0042131|T047|SY|12337004|SNOMEDCT_CORE|Uterine disease|Disorder of uterus
C0042131|T047|IS|12337004|SNOMEDCT_CORE|Uterine disease, NOS|Disorder of uterus
C0042131|T047|SY|12337004|SNOMEDCT_CORE|Uterine disorder|Disorder of uterus
C0042131|T047|IS|12337004|SNOMEDCT_CORE|Uterine disorder, NOS|Disorder of uterus
C0042133|T191|SY|95315005|SNOMEDCT_CORE|Fibroid uterus|Uterine leiomyoma
C0042133|T191|SY|95315005|SNOMEDCT_CORE|Fibroids|Uterine leiomyoma
C0042133|T191|SY|95315005|SNOMEDCT_CORE|Leiomyoma of body of uterus|Uterine leiomyoma
C0042133|T191|SY|95315005|SNOMEDCT_CORE|Leiomyoma of uterus|Uterine leiomyoma
C0042133|T191|SY|95315005|SNOMEDCT_CORE|Uterine fibroid|Uterine leiomyoma
C0042133|T191|SY|95315005|SNOMEDCT_CORE|Uterine fibroids|Uterine leiomyoma
C0042133|T191|PT|95315005|SNOMEDCT_CORE|Uterine leiomyoma|Uterine leiomyoma
C0042133|T191|FN|95315005|SNOMEDCT_CORE|Uterine leiomyoma|Uterine leiomyoma
C0042133|T191|SY|95315005|SNOMEDCT_CORE|Uterine leiomyoma - fibroids|Uterine leiomyoma
C0042133|T191|IS|95315005|SNOMEDCT_CORE|Uterine leiomyoma, NOS|Uterine leiomyoma
C0042134|T046|SYGB|38280009|SNOMEDCT_CORE|Haemorrhage in uterus|Uterine hemorrhage
C0042134|T046|SY|38280009|SNOMEDCT_CORE|Hemorrhage in uterus|Uterine hemorrhage
C0042134|T046|SYGB|38280009|SNOMEDCT_CORE|Uterine haemorrhage|Uterine hemorrhage
C0042134|T046|SY|38280009|SNOMEDCT_CORE|Uterine hemorrhage|Uterine hemorrhage
C0042140|T190|SY|24976005|SNOMEDCT_CORE|Descens uteri|Uterine prolapse
C0042140|T190|SY|24976005|SNOMEDCT_CORE|Descensus uteri|Uterine prolapse
C0042140|T190|SY|24976005|SNOMEDCT_CORE|Prolapse of uterus|Uterine prolapse
C0042140|T190|SY|24976005|SNOMEDCT_CORE|Prolapsed uterus|Uterine prolapse
C0042140|T190|SY|24976005|SNOMEDCT_CORE|Uterine hernia|Uterine prolapse
C0042140|T190|PT|24976005|SNOMEDCT_CORE|Uterine prolapse|Uterine prolapse
C0042140|T190|FN|24976005|SNOMEDCT_CORE|Uterine prolapse|Uterine prolapse
C0042140|T190|IS|24976005|SNOMEDCT_CORE|Uterine prolapse, NOS|Uterine prolapse
C0042164|T047|SY|128473001|SNOMEDCT_CORE|Intraocular inflammation|Uveitis
C0042164|T047|PT|128473001|SNOMEDCT_CORE|Uveitis|Uveitis
C0042164|T047|FN|128473001|SNOMEDCT_CORE|Uveitis|Uveitis
C0042165|T047|IS|77971008|SNOMEDCT_CORE|Anterior uveitis|Anterior uveitis
C0042165|T047|IS|77971008|SNOMEDCT_CORE|Anterior uveitis, NOS|Anterior uveitis
C0042167|T047|PT|43363007|SNOMEDCT_CORE|Posterior uveitis|Posterior uveitis
C0042167|T047|FN|43363007|SNOMEDCT_CORE|Posterior uveitis|Posterior uveitis
C0042167|T047|IS|43363007|SNOMEDCT_CORE|Posterior uveitis, NOS|Posterior uveitis
C0042171|T047|IS|31541009|SNOMEDCT_CORE|Uveoparotid fever|Uveoparotid fever
C0042237|T191|SY|363445000|SNOMEDCT_CORE|Cancer of vagina|Malignant tumor of vagina
C0042237|T191|PT|363445000|SNOMEDCT_CORE|Malignant tumor of vagina|Malignant tumor of vagina
C0042237|T191|FN|363445000|SNOMEDCT_CORE|Malignant tumor of vagina|Malignant tumor of vagina
C0042237|T191|PTGB|363445000|SNOMEDCT_CORE|Malignant tumour of vagina|Malignant tumor of vagina
C0042256|T184|SY|34363003|SNOMEDCT_CORE|Itching of vagina|Pruritus of vagina
C0042256|T184|PT|34363003|SNOMEDCT_CORE|Pruritus of vagina|Pruritus of vagina
C0042256|T184|FN|34363003|SNOMEDCT_CORE|Pruritus of vagina|Pruritus of vagina
C0042267|T047|SY|30800001|SNOMEDCT_CORE|Inflammation of vagina|Vaginitis
C0042267|T047|PT|30800001|SNOMEDCT_CORE|Vaginitis|Vaginitis
C0042267|T047|FN|30800001|SNOMEDCT_CORE|Vaginitis|Vaginitis
C0042267|T047|IS|30800001|SNOMEDCT_CORE|Vaginitis, NOS|Vaginitis
C0042331|T047|PT|193030005|SNOMEDCT_CORE|Migraine variants|Migraine variants
C0042331|T047|FN|193030005|SNOMEDCT_CORE|Migraine variants|Migraine variants
C0042341|T047|SY|51070004|SNOMEDCT_CORE|Scrotal varices|Varicocele
C0042341|T047|PT|51070004|SNOMEDCT_CORE|Varicocele|Varicocele
C0042341|T047|FN|51070004|SNOMEDCT_CORE|Varicocele|Varicocele
C0042344|T047|OAP|371032004|SNOMEDCT_CORE|Stasis ulcer|Stasis ulcer
C0042344|T047|OAF|371032004|SNOMEDCT_CORE|Stasis ulcer|Stasis ulcer
C0042344|T047|OAS|371032004|SNOMEDCT_CORE|Venous stasis ulcer|Stasis ulcer
C0042344|T047|OAS|371032004|SNOMEDCT_CORE|Venous ulcer|Stasis ulcer
C0042345|T047|OAP|276504003|SNOMEDCT_CORE|Varices|Venous varices
C0042345|T047|SY|128060009|SNOMEDCT_CORE|Varices|Venous varices
C0042345|T047|OAF|276504003|SNOMEDCT_CORE|Varices|Venous varices
C0042345|T047|SY|128060009|SNOMEDCT_CORE|Varicose veins|Venous varices
C0042345|T047|OAS|276504003|SNOMEDCT_CORE|Varicosities|Venous varices
C0042345|T047|SY|128060009|SNOMEDCT_CORE|Varicosities|Venous varices
C0042345|T047|PT|128060009|SNOMEDCT_CORE|Venous varices|Venous varices
C0042345|T047|FN|128060009|SNOMEDCT_CORE|Venous varices|Venous varices
C0042345|T047|OAS|276504003|SNOMEDCT_CORE|VV - Varicose veins|Venous varices
C0042345|T047|OAS|276504003|SNOMEDCT_CORE|VVs - Varicose veins|Venous varices
C0042373|T047|SY|27550009|SNOMEDCT_CORE|Angiopathy|Vascular disorder
C0042373|T047|IS|27550009|SNOMEDCT_CORE|Angiopathy, NOS|Vascular disorder
C0042373|T047|SY|27550009|SNOMEDCT_CORE|Disorder of blood vessel|Vascular disorder
C0042373|T047|FN|27550009|SNOMEDCT_CORE|Disorder of blood vessel|Vascular disorder
C0042373|T047|SY|27550009|SNOMEDCT_CORE|Vascular disease|Vascular disorder
C0042373|T047|OF|27550009|SNOMEDCT_CORE|Vascular disease|Vascular disorder
C0042373|T047|IS|27550009|SNOMEDCT_CORE|Vascular disease, NOS|Vascular disorder
C0042373|T047|PT|27550009|SNOMEDCT_CORE|Vascular disorder|Vascular disorder
C0042373|T047|IS|27550009|SNOMEDCT_CORE|Vascular disorder, NOS|Vascular disorder
C0042376|T047|PT|128187005|SNOMEDCT_CORE|Vascular headache|Vascular headache
C0042376|T047|FN|128187005|SNOMEDCT_CORE|Vascular headache|Vascular headache
C0042384|T047|SY|31996006|SNOMEDCT_CORE|Angiitis|Vasculitis
C0042384|T047|IS|31996006|SNOMEDCT_CORE|Angiitis, NOS|Vasculitis
C0042384|T047|PT|31996006|SNOMEDCT_CORE|Vasculitis|Vasculitis
C0042384|T047|FN|31996006|SNOMEDCT_CORE|Vasculitis|Vasculitis
C0042384|T047|IS|31996006|SNOMEDCT_CORE|Vasculitis, NOS|Vasculitis
C0042420|T047|OAS|398652001|SNOMEDCT_CORE|Gower's syndrome|Vasovagal syncope
C0042420|T047|SY|398665005|SNOMEDCT_CORE|Gower's syndrome|Vasovagal syncope
C0042420|T047|SY|398665005|SNOMEDCT_CORE|Neurally-mediated syncope|Vasovagal syncope
C0042420|T047|OAS|398652001|SNOMEDCT_CORE|Vagal attack|Vasovagal syncope
C0042420|T047|SY|398665005|SNOMEDCT_CORE|Vaso vagal episode|Vasovagal syncope
C0042420|T047|SY|398665005|SNOMEDCT_CORE|Vasodepressor syncope|Vasovagal syncope
C0042420|T047|OAP|398652001|SNOMEDCT_CORE|Vasovagal attack|Vasovagal syncope
C0042420|T047|SY|398665005|SNOMEDCT_CORE|Vasovagal attack|Vasovagal syncope
C0042420|T047|OAF|398652001|SNOMEDCT_CORE|Vasovagal attack|Vasovagal syncope
C0042420|T047|PT|398665005|SNOMEDCT_CORE|Vasovagal syncope|Vasovagal syncope
C0042420|T047|OF|398665005|SNOMEDCT_CORE|Vasovagal syncope|Vasovagal syncope
C0042420|T047|FN|398665005|SNOMEDCT_CORE|Vasovagal syncope|Vasovagal syncope
C0042485|T047|PT|20696009|SNOMEDCT_CORE|Peripheral venous insufficiency|Peripheral venous insufficiency
C0042485|T047|FN|20696009|SNOMEDCT_CORE|Peripheral venous insufficiency|Peripheral venous insufficiency
C0042485|T047|IS|20696009|SNOMEDCT_CORE|Peripheral venous insufficiency, NOS|Peripheral venous insufficiency
C0042487|T046|PT|111293003|SNOMEDCT_CORE|Venous thrombosis|Venous thrombosis
C0042487|T046|FN|111293003|SNOMEDCT_CORE|Venous thrombosis|Venous thrombosis
C0042487|T046|IS|111293003|SNOMEDCT_CORE|Venous thrombosis, NOS|Venous thrombosis
C0042510|T047|SY|71908006|SNOMEDCT_CORE|Cardiac arrest - ventricular fibrillation|Ventricular fibrillation
C0042510|T047|PT|71908006|SNOMEDCT_CORE|Ventricular fibrillation|Ventricular fibrillation
C0042510|T047|FN|71908006|SNOMEDCT_CORE|Ventricular fibrillation|Ventricular fibrillation
C0042510|T047|SY|71908006|SNOMEDCT_CORE|VF - Ventricular fibrillation|Ventricular fibrillation
C0042514|T047|IS|25569003|SNOMEDCT_CORE|Ventricular tachyarrhythmia|Ventricular tachycardia
C0042514|T047|PT|25569003|SNOMEDCT_CORE|Ventricular tachycardia|Ventricular tachycardia
C0042514|T047|FN|25569003|SNOMEDCT_CORE|Ventricular tachycardia|Ventricular tachycardia
C0042514|T047|IS|25569003|SNOMEDCT_CORE|Ventricular tachycardia, NOS|Ventricular tachycardia
C0042514|T047|SY|25569003|SNOMEDCT_CORE|VT - Ventricular tachycardia|Ventricular tachycardia
C0042548|T047|SY|63440008|SNOMEDCT_CORE|Plantar wart|Verruca plantaris
C0042548|T047|SY|63440008|SNOMEDCT_CORE|Verruca pedis|Verruca plantaris
C0042548|T047|PT|63440008|SNOMEDCT_CORE|Verruca plantaris|Verruca plantaris
C0042548|T047|FN|63440008|SNOMEDCT_CORE|Verruca plantaris|Verruca plantaris
C0042548|T047|SY|63440008|SNOMEDCT_CORE|VP - Verrucae pedis|Verruca plantaris
C0042568|T047|SY|64009001|SNOMEDCT_CORE|Vertebrobasilar arterial insufficiency|Vertebrobasilar insufficiency
C0042568|T047|SY|64009001|SNOMEDCT_CORE|Vertebrobasilar insufficiency|Vertebrobasilar insufficiency
C0042571|T184|SY|399153001|SNOMEDCT_CORE|Rotary vertigo|Vertigo
C0042571|T184|SY|399153001|SNOMEDCT_CORE|Rotatory vertigo|Vertigo
C0042571|T184|PT|399153001|SNOMEDCT_CORE|Vertigo|Vertigo
C0042571|T184|SY|399153001|SNOMEDCT_CORE|Vertigo|Vertigo
C0042571|T184|FN|399153001|SNOMEDCT_CORE|Vertigo|Vertigo
C0042580|T047|SY|197811007|SNOMEDCT_CORE|Ureteric reflux|Vesicoureteric reflux
C0042580|T047|SY|197811007|SNOMEDCT_CORE|Vesicoureteral reflux|Vesicoureteric reflux
C0042580|T047|PT|197811007|SNOMEDCT_CORE|Vesicoureteric reflux|Vesicoureteric reflux
C0042580|T047|FN|197811007|SNOMEDCT_CORE|Vesicoureteric reflux|Vesicoureteric reflux
C0042580|T047|SY|197811007|SNOMEDCT_CORE|VUR - Vesicoureteric reflux|Vesicoureteric reflux
C0042582|T047|PT|89405008|SNOMEDCT_CORE|Vesicovaginal fistula|Vesicovaginal fistula
C0042582|T047|FN|89405008|SNOMEDCT_CORE|Vesicovaginal fistula|Vesicovaginal fistula
C0042582|T047|SY|89405008|SNOMEDCT_CORE|VVF - Vesicovaginal fistula|Vesicovaginal fistula
C0042594|T047|SY|20425006|SNOMEDCT_CORE|Vestibular disorder|Vestibular disorder
C0042594|T047|IS|20425006|SNOMEDCT_CORE|Vestibular disorder, NOS|Vestibular disorder
C0042708|T047|PT|78420004|SNOMEDCT_CORE|Viral enteritis|Viral enteritis
C0042708|T047|FN|78420004|SNOMEDCT_CORE|Viral enteritis|Viral enteritis
C0042708|T047|IS|78420004|SNOMEDCT_CORE|Viral enteritis, NOS|Viral enteritis
C0042740|T047|SY|445939008|SNOMEDCT_CORE|Nonspecific syndrome suggestive of viral illness|Viral syndrome
C0042740|T047|FN|445939008|SNOMEDCT_CORE|Nonspecific syndrome suggestive of viral illness|Viral syndrome
C0042740|T047|PT|445939008|SNOMEDCT_CORE|Viral syndrome|Viral syndrome
C0042749|T047|PTGB|2528003|SNOMEDCT_CORE|Viraemia|Viremia
C0042749|T047|IS|2528003|SNOMEDCT_CORE|Viral sepsis|Viremia
C0042749|T047|PT|2528003|SNOMEDCT_CORE|Viremia|Viremia
C0042749|T047|OF|2528003|SNOMEDCT_CORE|Viremia|Viremia
C0042749|T047|FN|2528003|SNOMEDCT_CORE|Viremia|Viremia
C0042749|T047|IS|2528003|SNOMEDCT_CORE|Viremia, NOS|Viremia
C0042769|T047|SY|34014006|SNOMEDCT_CORE|Disease caused by virus|Viral disease
C0042769|T047|IS|34014006|SNOMEDCT_CORE|Disease caused by virus, NOS|Viral disease
C0042769|T047|SY|34014006|SNOMEDCT_CORE|Disease due to virus|Viral disease
C0042769|T047|PT|34014006|SNOMEDCT_CORE|Viral disease|Viral disease
C0042769|T047|FN|34014006|SNOMEDCT_CORE|Viral disease|Viral disease
C0042769|T047|IS|34014006|SNOMEDCT_CORE|Viral disease, NOS|Viral disease
C0042769|T047|SY|34014006|SNOMEDCT_CORE|Viral illness|Viral disease
C0042769|T047|IS|34014006|SNOMEDCT_CORE|Viral illness, NOS|Viral disease
C0042769|T047|SY|34014006|SNOMEDCT_CORE|Viral infection|Viral disease
C0042769|T047|IS|34014006|SNOMEDCT_CORE|Viral infection, NOS|Viral disease
C0042769|T047|SY|34014006|SNOMEDCT_CORE|Viral infectious disease|Viral disease
C0042769|T047|IS|34014006|SNOMEDCT_CORE|Viral infectious disease, NOS|Viral disease
C0042790|T033|PT|95677002|SNOMEDCT_CORE|Disorder of vision|Disorder of vision
C0042790|T033|FN|95677002|SNOMEDCT_CORE|Disorder of vision|Disorder of vision
C0042790|T033|IS|95677002|SNOMEDCT_CORE|Disorder of vision, NOS|Disorder of vision
C0042790|T033|SY|95677002|SNOMEDCT_CORE|Vision disorder|Disorder of vision
C0042790|T033|IS|95677002|SNOMEDCT_CORE|Vision disorder, NOS|Disorder of vision
C0042790|T033|IS|7973008|SNOMEDCT_CORE|Visual disorder|Disorder of vision
C0042798|T047|IS|7973008|SNOMEDCT_CORE|Low vision|LV - Low vision
C0042798|T047|IS|7973008|SNOMEDCT_CORE|LV - Low vision|LV - Low vision
C0042847|T047|PT|190634004|SNOMEDCT_CORE|Cobalamin deficiency|Cobalamin deficiency
C0042847|T047|FN|190634004|SNOMEDCT_CORE|Cobalamin deficiency|Cobalamin deficiency
C0042847|T047|MTH_SY|190634004|SNOMEDCT_CORE|Deficiency of vitamin B<sub>12</sub>|Cobalamin deficiency
C0042847|T047|SY|190634004|SNOMEDCT_CORE|Deficiency of vitamin B>12<|Cobalamin deficiency
C0042847|T047|MTH_SY|190634004|SNOMEDCT_CORE|Deficiency of vitamin B12|Cobalamin deficiency
C0042847|T047|SY|190634004|SNOMEDCT_CORE|Vitamin B12 deficiency|Cobalamin deficiency
C0042850|T047|SY|47903000|SNOMEDCT_CORE|Deficiency of vitamin B|Vitamin B-complex deficiency
C0042850|T047|PT|47903000|SNOMEDCT_CORE|Vitamin B deficiency|Vitamin B-complex deficiency
C0042850|T047|FN|47903000|SNOMEDCT_CORE|Vitamin B deficiency|Vitamin B-complex deficiency
C0042850|T047|IS|47903000|SNOMEDCT_CORE|Vitamin B deficiency, NOS|Vitamin B-complex deficiency
C0042850|T047|IS|47903000|SNOMEDCT_CORE|Vitamin B-complex deficiency|Vitamin B-complex deficiency
C0042850|T047|PT|190631007|SNOMEDCT_CORE|Vitamin B-complex deficiency|Vitamin B-complex deficiency
C0042850|T047|FN|190631007|SNOMEDCT_CORE|Vitamin B-complex deficiency|Vitamin B-complex deficiency
C0042850|T047|IS|47903000|SNOMEDCT_CORE|Vitamin B-complex deficiency, NOS|Vitamin B-complex deficiency
C0042870|T047|SY|34713006|SNOMEDCT_CORE|Avitaminosis D|Vitamin D deficiency
C0042870|T047|IS|34713006|SNOMEDCT_CORE|Avitaminosis D, NOS|Vitamin D deficiency
C0042870|T047|PT|34713006|SNOMEDCT_CORE|Vitamin D deficiency|Vitamin D deficiency
C0042870|T047|FN|34713006|SNOMEDCT_CORE|Vitamin D deficiency|Vitamin D deficiency
C0042870|T047|IS|34713006|SNOMEDCT_CORE|Vitamin D deficiency, NOS|Vitamin D deficiency
C0042900|T047|PT|56727007|SNOMEDCT_CORE|Vitiligo|Vitiligo
C0042900|T047|FN|56727007|SNOMEDCT_CORE|Vitiligo|Vitiligo
C0042907|T047|PT|53772007|SNOMEDCT_CORE|Vitreous detachment|Vitreous detachment
C0042907|T047|FN|53772007|SNOMEDCT_CORE|Vitreous detachment|Vitreous detachment
C0042907|T047|SY|53772007|SNOMEDCT_CORE|Vitreous separation|Vitreous detachment
C0042909|T046|SYGB|31341008|SNOMEDCT_CORE|Intragel vitreous haemorrhage|Vitreous hemorrhage
C0042909|T046|SY|31341008|SNOMEDCT_CORE|Intragel vitreous hemorrhage|Vitreous hemorrhage
C0042909|T046|SYGB|31341008|SNOMEDCT_CORE|VH - Vitreous haemorrhage|Vitreous hemorrhage
C0042909|T046|SY|31341008|SNOMEDCT_CORE|VH - Vitreous hemorrhage|Vitreous hemorrhage
C0042909|T046|PTGB|31341008|SNOMEDCT_CORE|Vitreous haemorrhage|Vitreous hemorrhage
C0042909|T046|PT|31341008|SNOMEDCT_CORE|Vitreous hemorrhage|Vitreous hemorrhage
C0042909|T046|FN|31341008|SNOMEDCT_CORE|Vitreous hemorrhage|Vitreous hemorrhage
C0042928|T047|SY|302912005|SNOMEDCT_CORE|Paralysis of vocal cords|Vocal cord paralysis
C0042928|T047|SY|302912005|SNOMEDCT_CORE|VCP - Vocal cord palsy|Vocal cord paralysis
C0042928|T047|SY|302912005|SNOMEDCT_CORE|Vocal cord palsy|Vocal cord paralysis
C0042928|T047|FN|302912005|SNOMEDCT_CORE|Vocal cord palsy|Vocal cord paralysis
C0042928|T047|PT|302912005|SNOMEDCT_CORE|Vocal cord paralysis|Vocal cord paralysis
C0042928|T047|SY|302912005|SNOMEDCT_CORE|Vocal fold palsy|Vocal cord paralysis
C0042929|T191|PT|9078005|SNOMEDCT_CORE|Polyp of vocal cord|Polyp of vocal cord
C0042929|T191|FN|9078005|SNOMEDCT_CORE|Polyp of vocal cord|Polyp of vocal cord
C0042929|T191|SY|9078005|SNOMEDCT_CORE|Vocal fold polyp|Polyp of vocal cord
C0042940|T047|IS|47004009|SNOMEDCT_CORE|Disorder of voice|Voice impairment, NOS
C0042940|T047|IS|47004009|SNOMEDCT_CORE|Voice disorder|Voice impairment, NOS
C0042940|T047|IS|47004009|SNOMEDCT_CORE|Voice disorder, NOS|Voice impairment, NOS
C0042940|T047|IS|47004009|SNOMEDCT_CORE|Voice impairment|Voice impairment, NOS
C0042940|T047|IS|47004009|SNOMEDCT_CORE|Voice impairment, NOS|Voice impairment, NOS
C0042963|T184|SY|422400008|SNOMEDCT_CORE|Emesis|Vomiting
C0042963|T184|PT|422400008|SNOMEDCT_CORE|Vomiting|Vomiting
C0042963|T184|FN|422400008|SNOMEDCT_CORE|Vomiting|Vomiting
C0042974|T047|SYGB|128105004|SNOMEDCT_CORE|Angiohaemophilia|von Willebrand disorder
C0042974|T047|SY|128105004|SNOMEDCT_CORE|Angiohemophilia|von Willebrand disorder
C0042974|T047|SY|128105004|SNOMEDCT_CORE|Constitutional thrombopathy|von Willebrand disorder
C0042974|T047|SY|128105004|SNOMEDCT_CORE|Factor VIII deficiency with vascular defect|von Willebrand disorder
C0042974|T047|SYGB|128105004|SNOMEDCT_CORE|Pseudohaemophilia type B|von Willebrand disorder
C0042974|T047|SY|128105004|SNOMEDCT_CORE|Pseudohemophilia type B|von Willebrand disorder
C0042974|T047|SYGB|128105004|SNOMEDCT_CORE|Vascular haemophilia|von Willebrand disorder
C0042974|T047|SY|128105004|SNOMEDCT_CORE|Vascular hemophilia|von Willebrand disorder
C0042974|T047|SY|128105004|SNOMEDCT_CORE|von Willebrand disease|von Willebrand disorder
C0042974|T047|FN|128105004|SNOMEDCT_CORE|von Willebrand disorder|von Willebrand disorder
C0042974|T047|PT|128105004|SNOMEDCT_CORE|von Willebrand disorder|von Willebrand disorder
C0042974|T047|IS|128105004|SNOMEDCT_CORE|von Willebrand-J?rgens disease|von Willebrand disorder
C0042974|T047|SY|128105004|SNOMEDCT_CORE|von Willebrand-Jurgens disease|von Willebrand disorder
C0042974|T047|SY|128105004|SNOMEDCT_CORE|von Willebrand's disease|von Willebrand disorder
C0042974|T047|SY|128105004|SNOMEDCT_CORE|vWD - von Willebrand's disease|von Willebrand disorder
C0042996|T047|PT|63144007|SNOMEDCT_CORE|Vulvitis|Vulvitis
C0042996|T047|FN|63144007|SNOMEDCT_CORE|Vulvitis|Vulvitis
C0042996|T047|IS|63144007|SNOMEDCT_CORE|Vulvitis, NOS|Vulvitis
C0042998|T047|PT|53277000|SNOMEDCT_CORE|Vulvovaginitis|Vulvovaginitis
C0042998|T047|FN|53277000|SNOMEDCT_CORE|Vulvovaginitis|Vulvovaginitis
C0042998|T047|IS|53277000|SNOMEDCT_CORE|Vulvovaginitis, NOS|Vulvovaginitis
C0043037|T047|SY|57019003|SNOMEDCT_CORE|Common wart|Verruca vulgaris
C0043037|T047|SY|57019003|SNOMEDCT_CORE|Human papilloma virus infection of skin|Verruca vulgaris
C0043037|T047|SY|57019003|SNOMEDCT_CORE|Infectious warts|Verruca vulgaris
C0043037|T047|SY|57019003|SNOMEDCT_CORE|Verruca simplex|Verruca vulgaris
C0043037|T047|PT|57019003|SNOMEDCT_CORE|Verruca vulgaris|Verruca vulgaris
C0043037|T047|FN|57019003|SNOMEDCT_CORE|Verruca vulgaris|Verruca vulgaris
C0043037|T047|SY|57019003|SNOMEDCT_CORE|Viral wart|Verruca vulgaris
C0043037|T047|SY|57019003|SNOMEDCT_CORE|Viral warts|Verruca vulgaris
C0043037|T047|SY|57019003|SNOMEDCT_CORE|Viral warts due to papilloma virus|Verruca vulgaris
C0043066|T184|IS|16331000|SNOMEDCT_CORE|Waterbrash|Waterbrash
C0043094|T033|PT|262286000|SNOMEDCT_CORE|Weight increased|Weight increased
C0043094|T033|OF|262286000|SNOMEDCT_CORE|Weight increased|Weight increased
C0043094|T033|FN|262286000|SNOMEDCT_CORE|Weight increased|Weight increased
C0043144|T184|SY|56018004|SNOMEDCT_CORE|Wheeze|Wheezing
C0043144|T184|PT|56018004|SNOMEDCT_CORE|Wheezing|Wheezing
C0043144|T184|FN|56018004|SNOMEDCT_CORE|Wheezing|Wheezing
C0043144|T184|IS|56018004|SNOMEDCT_CORE|Wheezing, NOS|Wheezing
C0043144|T184|SY|56018004|SNOMEDCT_CORE|Wheezy|Wheezing
C0043145|T037|SY|39848009|SNOMEDCT_CORE|Acceleration-deceleration injury of neck|Whiplash injury to neck
C0043145|T037|SY|39848009|SNOMEDCT_CORE|Whiplash injury|Whiplash injury to neck
C0043145|T037|PT|39848009|SNOMEDCT_CORE|Whiplash injury to neck|Whiplash injury to neck
C0043145|T037|FN|39848009|SNOMEDCT_CORE|Whiplash injury to neck|Whiplash injury to neck
C0043167|T047|SY|27836007|SNOMEDCT_CORE|Infection due to Bordetella pertussis|Pertussis
C0043167|T047|PT|27836007|SNOMEDCT_CORE|Pertussis|Pertussis
C0043167|T047|FN|27836007|SNOMEDCT_CORE|Pertussis|Pertussis
C0043167|T047|SY|27836007|SNOMEDCT_CORE|WC - Whooping cough|Pertussis
C0043167|T047|SY|27836007|SNOMEDCT_CORE|Whooping cough|Pertussis
C0043167|T047|IS|27836007|SNOMEDCT_CORE|Whooping cough, NOS|Pertussis
C0043202|T047|SY|74390002|SNOMEDCT_CORE|Ventricular pre-excitation with arrhythmia|Wolff-Parkinson-White pattern
C0043202|T047|IS|74390002|SNOMEDCT_CORE|Ventricular pre-excitation with arrhythmia, NOS|Wolff-Parkinson-White pattern
C0043202|T047|SY|74390002|SNOMEDCT_CORE|Wolff Parkinson White syndrome|Wolff-Parkinson-White pattern
C0043202|T047|PT|74390002|SNOMEDCT_CORE|Wolff-Parkinson-White pattern|Wolff-Parkinson-White pattern
C0043202|T047|FN|74390002|SNOMEDCT_CORE|Wolff-Parkinson-White pattern|Wolff-Parkinson-White pattern
C0043202|T047|IS|74390002|SNOMEDCT_CORE|Wolff-Parkinson-White syndrome|Wolff-Parkinson-White pattern
C0043202|T047|SY|74390002|SNOMEDCT_CORE|WPW - Wolff-Parkinson-White pattern|Wolff-Parkinson-White pattern
C0043202|T047|SY|74390002|SNOMEDCT_CORE|WPW - Wolff-Parkinson-White syndrome|Wolff-Parkinson-White pattern
C0043241|T046|SY|76844004|SNOMEDCT_CORE|Infected wound|Local infection of wound
C0043241|T046|IS|76844004|SNOMEDCT_CORE|Infected wound, NOS|Local infection of wound
C0043241|T046|PT|76844004|SNOMEDCT_CORE|Local infection of wound|Local infection of wound
C0043241|T046|FN|76844004|SNOMEDCT_CORE|Local infection of wound|Local infection of wound
C0043241|T046|IS|76844004|SNOMEDCT_CORE|Local infection of wound, NOS|Local infection of wound
C0043241|T046|SY|76844004|SNOMEDCT_CORE|Septic wound|Local infection of wound
C0043241|T046|SY|76844004|SNOMEDCT_CORE|Wound infected|Local infection of wound
C0043241|T046|SY|76844004|SNOMEDCT_CORE|Wound infection|Local infection of wound
C0043246|T037|SY|312608009|SNOMEDCT_CORE|Laceration|Laceration - injury
C0043246|T037|PT|312608009|SNOMEDCT_CORE|Laceration - injury|Laceration - injury
C0043246|T037|FN|312608009|SNOMEDCT_CORE|Laceration - injury|Laceration - injury
C0043250|T037|PT|416462003|SNOMEDCT_CORE|Wound|Wound
C0043250|T037|FN|416462003|SNOMEDCT_CORE|Wound|Wound
C0043252|T037|IS|283545005|SNOMEDCT_CORE|GSW|Gunshot wound
C0043252|T037|SY|283545005|SNOMEDCT_CORE|GSW - Gun shot wound|Gunshot wound
C0043252|T037|SY|283545005|SNOMEDCT_CORE|Gun shot wound|Gunshot wound
C0043252|T037|OF|283545005|SNOMEDCT_CORE|Gun shot wound|Gunshot wound
C0043252|T037|PT|283545005|SNOMEDCT_CORE|Gunshot wound|Gunshot wound
C0043252|T037|FN|283545005|SNOMEDCT_CORE|Gunshot wound|Gunshot wound
C0043253|T037|PT|425359009|SNOMEDCT_CORE|Blunt injury|Blunt injury
C0043253|T037|FN|425359009|SNOMEDCT_CORE|Blunt injury|Blunt injury
C0043253|T037|SY|425359009|SNOMEDCT_CORE|Blunt trauma|Blunt injury
C0043255|T037|PT|425322008|SNOMEDCT_CORE|Stab wound|Stab wound
C0043255|T037|FN|425322008|SNOMEDCT_CORE|Stab wound|Stab wound
C0043264|T037|PT|125598003|SNOMEDCT_CORE|Injury of wrist|Injury of wrist
C0043264|T037|FN|125598003|SNOMEDCT_CORE|Injury of wrist|Injury of wrist
C0043264|T037|SY|125598003|SNOMEDCT_CORE|Wrist injury|Injury of wrist
C0043349|T047|PT|46152009|SNOMEDCT_CORE|Tear film insufficiency|Tear film insufficiency
C0043349|T047|FN|46152009|SNOMEDCT_CORE|Tear film insufficiency|Tear film insufficiency
C0043349|T047|IS|46152009|SNOMEDCT_CORE|Tear film insufficiency, NOS|Tear film insufficiency
C0043352|T033|SY|87715008|SNOMEDCT_CORE|Absent salivary secretion|Xerostomia
C0043352|T033|SY|87715008|SNOMEDCT_CORE|Aptyalia|Xerostomia
C0043352|T033|SY|87715008|SNOMEDCT_CORE|Aptyalism|Xerostomia
C0043352|T033|OF|87715008|SNOMEDCT_CORE|Aptyalism|Xerostomia
C0043352|T033|SY|87715008|SNOMEDCT_CORE|Asialia|Xerostomia
C0043352|T033|SY|87715008|SNOMEDCT_CORE|Clinical xerostomia|Xerostomia
C0043352|T033|SY|87715008|SNOMEDCT_CORE|Dry mouth|Xerostomia
C0043352|T033|PT|87715008|SNOMEDCT_CORE|Xerostomia|Xerostomia
C0043352|T033|FN|87715008|SNOMEDCT_CORE|Xerostomia|Xerostomia
C0078981|T047|PT|33595009|SNOMEDCT_CORE|Arachnoid cyst|Arachnoid cyst
C0078981|T047|FN|33595009|SNOMEDCT_CORE|Arachnoid cyst|Arachnoid cyst
C0079352|T019|SY|268240006|SNOMEDCT_CORE|Congenital sternomastoid torticollis|Congenital torticollis
C0079352|T019|PT|268240006|SNOMEDCT_CORE|Congenital torticollis|Congenital torticollis
C0079352|T019|FN|268240006|SNOMEDCT_CORE|Congenital torticollis|Congenital torticollis
C0079352|T019|SY|268240006|SNOMEDCT_CORE|Congenital wry neck|Congenital torticollis
C0079352|T019|SY|268240006|SNOMEDCT_CORE|Congenital wryneck|Congenital torticollis
C0079352|T019|SY|268240006|SNOMEDCT_CORE|Contracture of sternocleidomastoid muscle|Congenital torticollis
C0079745|T191|OAP|277641001|SNOMEDCT_CORE|Follicular malignant lymphoma - large cell|Malignant lymphoma - non-cleaved, follicular
C0079745|T191|OAF|277641001|SNOMEDCT_CORE|Follicular malignant lymphoma - large cell|Malignant lymphoma - non-cleaved, follicular
C0079745|T191|OAS|277641001|SNOMEDCT_CORE|Malignant lymphoma - histiocytic, nodular|Malignant lymphoma - non-cleaved, follicular
C0079745|T191|OAS|277641001|SNOMEDCT_CORE|Malignant lymphoma - non-cleaved, follicular|Malignant lymphoma - non-cleaved, follicular
C0079773|T191|SY|400122007|SNOMEDCT_CORE|CTCL - Cutaneous T-cell lymphoma|Primary cutaneous T-cell lymphoma
C0079773|T191|SY|400122007|SNOMEDCT_CORE|Cutaneous T-cell lymphoma|Primary cutaneous T-cell lymphoma
C0079773|T191|FN|400122007|SNOMEDCT_CORE|Primary cutaneous T-cell lymphoma|Primary cutaneous T-cell lymphoma
C0079773|T191|PT|400122007|SNOMEDCT_CORE|Primary cutaneous T-cell lymphoma|Primary cutaneous T-cell lymphoma
C0079924|T046|SY|59566000|SNOMEDCT_CORE|Deficient liquor|Oligohydramnios
C0079924|T046|PT|59566000|SNOMEDCT_CORE|Oligohydramnios|Oligohydramnios
C0079924|T046|FN|59566000|SNOMEDCT_CORE|Oligohydramnios|Oligohydramnios
C0079924|T046|IS|59566000|SNOMEDCT_CORE|Oligohydramnios, NOS|Oligohydramnios
C0079924|T046|SY|59566000|SNOMEDCT_CORE|Reduced liquor volume|Oligohydramnios
C0079924|T046|SY|59566000|SNOMEDCT_CORE|Scanty liquor|Oligohydramnios
C0080032|T047|SY|83270006|SNOMEDCT_CORE|Malignant effusion|Neoplastic pleural effusion
C0080032|T047|SY|83270006|SNOMEDCT_CORE|Malignant pleural effusion|Neoplastic pleural effusion
C0080032|T047|PT|83270006|SNOMEDCT_CORE|Neoplastic pleural effusion|Neoplastic pleural effusion
C0080032|T047|FN|83270006|SNOMEDCT_CORE|Neoplastic pleural effusion|Neoplastic pleural effusion
C0080032|T047|SY|83270006|SNOMEDCT_CORE|Pleural effusion due to malignancy|Neoplastic pleural effusion
C0080040|T047|PT|31097004|SNOMEDCT_CORE|Post poliomyelitis syndrome|Post poliomyelitis syndrome
C0080040|T047|FN|31097004|SNOMEDCT_CORE|Post poliomyelitis syndrome|Post poliomyelitis syndrome
C0080040|T047|SY|31097004|SNOMEDCT_CORE|Post-polio progressive muscular atrophy|Post poliomyelitis syndrome
C0080040|T047|SY|31097004|SNOMEDCT_CORE|Postpolio muscular atrophy|Post poliomyelitis syndrome
C0080040|T047|SY|31097004|SNOMEDCT_CORE|Postpolio syndrome|Post poliomyelitis syndrome
C0080040|T047|SY|31097004|SNOMEDCT_CORE|Progressive muscular atrophy following poliomyelitis|Post poliomyelitis syndrome
C0080178|T019|SY|67531005|SNOMEDCT_CORE|Posterior rachischisis|Spina bifida
C0080178|T019|SY|67531005|SNOMEDCT_CORE|SB - Spina bifida|Spina bifida
C0080178|T019|PT|67531005|SNOMEDCT_CORE|Spina bifida|Spina bifida
C0080178|T019|FN|67531005|SNOMEDCT_CORE|Spina bifida|Spina bifida
C0080178|T019|IS|67531005|SNOMEDCT_CORE|Spina bifida, NOS|Spina bifida
C0080178|T019|IS|67531005|SNOMEDCT_CORE|Spinal dysraphism|Spina bifida
C0080179|T037|SY|50448004|SNOMEDCT_CORE|Fracture of spinal vertebra|Fracture of vertebral column
C0080179|T037|SY|50448004|SNOMEDCT_CORE|Fracture of spine|Fracture of vertebral column
C0080179|T037|SY|50448004|SNOMEDCT_CORE|Fracture of vertebra|Fracture of vertebral column
C0080179|T037|PT|50448004|SNOMEDCT_CORE|Fracture of vertebral column|Fracture of vertebral column
C0080179|T037|FN|50448004|SNOMEDCT_CORE|Fracture of vertebral column|Fracture of vertebral column
C0080179|T037|IS|50448004|SNOMEDCT_CORE|Fracture of vertebral column, NOS|Fracture of vertebral column
C0080179|T037|SY|50448004|SNOMEDCT_CORE|Fractured spine|Fracture of vertebral column
C0080179|T037|SY|50448004|SNOMEDCT_CORE|Spinal fracture|Fracture of vertebral column
C0080194|T037|PT|48532005|SNOMEDCT_CORE|Muscle strain|Muscle strain
C0080194|T037|FN|48532005|SNOMEDCT_CORE|Muscle strain|Muscle strain
C0080194|T037|SY|48532005|SNOMEDCT_CORE|Pulled muscle|Muscle strain
C0080194|T037|SY|48532005|SNOMEDCT_CORE|Strain|Muscle strain
C0080194|T037|IS|48532005|SNOMEDCT_CORE|Strain, NOS|Muscle strain
C0080203|T033|PT|6285003|SNOMEDCT_CORE|Tachyarrhythmia|Tachyarrhythmia
C0080203|T033|FN|6285003|SNOMEDCT_CORE|Tachyarrhythmia|Tachyarrhythmia
C0080203|T033|IS|6285003|SNOMEDCT_CORE|Tachyarrhythmia, NOS|Tachyarrhythmia
C0080218|T047|SY|70534000|SNOMEDCT_CORE|Congenital tethering of spinal cord|Occult spinal dysraphism sequence
C0080218|T047|FN|70534000|SNOMEDCT_CORE|Occult spinal dysraphism sequence|Occult spinal dysraphism sequence
C0080218|T047|PT|70534000|SNOMEDCT_CORE|Occult spinal dysraphism sequence|Occult spinal dysraphism sequence
C0080218|T047|SY|70534000|SNOMEDCT_CORE|Tethered cord malformation sequence|Occult spinal dysraphism sequence
C0080218|T047|SY|70534000|SNOMEDCT_CORE|Tethered cord syndrome|Occult spinal dysraphism sequence
C0080233|T020|IS|37320007|SNOMEDCT_CORE|Absence of tooth - acquired|Acquired absence of teeth
C0080233|T020|PT|37320007|SNOMEDCT_CORE|Acquired absence of teeth|Acquired absence of teeth
C0080233|T020|FN|37320007|SNOMEDCT_CORE|Acquired absence of teeth|Acquired absence of teeth
C0080233|T020|IS|37320007|SNOMEDCT_CORE|Acquired absence of teeth, NOS|Acquired absence of teeth
C0080233|T020|SY|37320007|SNOMEDCT_CORE|Acquired edentia|Acquired absence of teeth
C0080233|T020|SY|37320007|SNOMEDCT_CORE|Loss of teeth|Acquired absence of teeth
C0080233|T020|SY|37320007|SNOMEDCT_CORE|Loss of teeth - acquired|Acquired absence of teeth
C0080233|T020|IS|37320007|SNOMEDCT_CORE|Loss of teeth, NOS|Acquired absence of teeth
C0080233|T020|IS|37320007|SNOMEDCT_CORE|Missing tooth - acquired|Acquired absence of teeth
C0080233|T020|SY|25540007|SNOMEDCT_CORE|Shedding of tooth|Acquired absence of teeth
C0080233|T020|SY|37320007|SNOMEDCT_CORE|Teeth missing|Acquired absence of teeth
C0080233|T020|PT|25540007|SNOMEDCT_CORE|Tooth loss|Acquired absence of teeth
C0080233|T020|FN|25540007|SNOMEDCT_CORE|Tooth loss|Acquired absence of teeth
C0080233|T020|IS|25540007|SNOMEDCT_CORE|Tooth loss, NOS|Acquired absence of teeth
C0080274|T033|SY|267064002|SNOMEDCT_CORE|Cannot pass urine - retention|Retention of urine
C0080274|T033|SY|267064002|SNOMEDCT_CORE|Not passing urine|Retention of urine
C0080274|T033|PT|267064002|SNOMEDCT_CORE|Retention of urine|Retention of urine
C0080274|T033|FN|267064002|SNOMEDCT_CORE|Retention of urine|Retention of urine
C0080274|T033|SY|267064002|SNOMEDCT_CORE|Unable to empty bladder|Retention of urine
C0080274|T033|SY|267064002|SNOMEDCT_CORE|Unable to pass urine|Retention of urine
C0080274|T033|SY|267064002|SNOMEDCT_CORE|Urinary retention|Retention of urine
C0085074|T047|SY|65508009|SNOMEDCT_CORE|GA - Granuloma annulare|Granuloma annulare
C0085074|T047|PT|65508009|SNOMEDCT_CORE|Granuloma annulare|Granuloma annulare
C0085074|T047|FN|65508009|SNOMEDCT_CORE|Granuloma annulare|Granuloma annulare
C0085083|T047|PT|129635004|SNOMEDCT_CORE|Ovarian hyperstimulation syndrome|Ovarian hyperstimulation syndrome
C0085083|T047|FN|129635004|SNOMEDCT_CORE|Ovarian hyperstimulation syndrome|Ovarian hyperstimulation syndrome
C0085083|T047|SY|129635004|SNOMEDCT_CORE|Secondary Meig's syndrome|Ovarian hyperstimulation syndrome
C0085084|T047|SY|37340000|SNOMEDCT_CORE|MND - Motor neurone disease|Motor neuron disease
C0085084|T047|PT|37340000|SNOMEDCT_CORE|Motor neuron disease|Motor neuron disease
C0085084|T047|FN|37340000|SNOMEDCT_CORE|Motor neuron disease|Motor neuron disease
C0085084|T047|IS|37340000|SNOMEDCT_CORE|Motor neuron disease, NOS|Motor neuron disease
C0085084|T047|SY|37340000|SNOMEDCT_CORE|Motor neurone disease|Motor neuron disease
C0085096|T047|SY|399957001|SNOMEDCT_CORE|Peripheral angiopathy|Peripheral vascular disease
C0085096|T047|PT|400047006|SNOMEDCT_CORE|Peripheral vascular disease|Peripheral vascular disease
C0085096|T047|FN|400047006|SNOMEDCT_CORE|Peripheral vascular disease|Peripheral vascular disease
C0085096|T047|SY|400047006|SNOMEDCT_CORE|PVD - peripheral vascular disease|Peripheral vascular disease
C0085096|T047|IS|399957001|SNOMEDCT_CORE|PVD - Peripheral vascular disease|Peripheral vascular disease
C0085096|T047|IS|400047006|SNOMEDCT_CORE|PVD-peripheral vascular disease|Peripheral vascular disease
C0085111|T037|SY|125603006|SNOMEDCT_CORE|Ankle injury|Injury of ankle
C0085111|T037|PT|125603006|SNOMEDCT_CORE|Injury of ankle|Injury of ankle
C0085111|T037|FN|125603006|SNOMEDCT_CORE|Injury of ankle|Injury of ankle
C0085119|T047|SY|95345008|SNOMEDCT_CORE|Foot ulcer|Ulcer of foot
C0085119|T047|PT|95345008|SNOMEDCT_CORE|Ulcer of foot|Ulcer of foot
C0085119|T047|FN|95345008|SNOMEDCT_CORE|Ulcer of foot|Ulcer of foot
C0085119|T047|IS|95345008|SNOMEDCT_CORE|Ulcer of foot, NOS|Ulcer of foot
C0085129|T047|SY|195967001|SNOMEDCT_CORE|BHR - Bronchial hyperreactivity|BHR - Bronchial hyperreactivity
C0085129|T047|SY|195967001|SNOMEDCT_CORE|Bronchial hyperreactivity|BHR - Bronchial hyperreactivity
C0085129|T047|SY|195967001|SNOMEDCT_CORE|Bronchial hyperresponsiveness|BHR - Bronchial hyperreactivity
C0085129|T047|SY|195967001|SNOMEDCT_CORE|Bronchial hypersensitivity|BHR - Bronchial hyperreactivity
C0085159|T048|SY|247803002|SNOMEDCT_CORE|SAD - Seasonal affective disorder|Seasonal affective disorder
C0085159|T048|PT|247803002|SNOMEDCT_CORE|Seasonal affective disorder|Seasonal affective disorder
C0085159|T048|FN|247803002|SNOMEDCT_CORE|Seasonal affective disorder|Seasonal affective disorder
C0085160|T047|PT|69741000|SNOMEDCT_CORE|Hidradenitis|Hidradenitis
C0085160|T047|FN|69741000|SNOMEDCT_CORE|Hidradenitis|Hidradenitis
C0085166|T047|IS|419760006|SNOMEDCT_CORE|AV - Anaerobic vaginosis|Bacterial vaginosis
C0085166|T047|SY|419760006|SNOMEDCT_CORE|Bacterial vaginitis|Bacterial vaginosis
C0085166|T047|PT|419760006|SNOMEDCT_CORE|Bacterial vaginosis|Bacterial vaginosis
C0085166|T047|FN|419760006|SNOMEDCT_CORE|Bacterial vaginosis|Bacterial vaginosis
C0085166|T047|SY|419760006|SNOMEDCT_CORE|BV - Bacterial vaginosis|Bacterial vaginosis
C0085166|T047|SY|419760006|SNOMEDCT_CORE|Nonspecific bacterial vaginosis|Bacterial vaginosis
C0085166|T047|IS|419760006|SNOMEDCT_CORE|Nonspecific vaginitis|Bacterial vaginosis
C0085166|T047|IS|419760006|SNOMEDCT_CORE|NSV - Nonspecific vaginitis|Bacterial vaginosis
C0085178|T037|OAS|283596007|SNOMEDCT_CORE|Needle prick injury|Needle prick injury
C0085178|T037|OAF|283596007|SNOMEDCT_CORE|Needle stick injury|Needle prick injury
C0085178|T037|OAP|283596007|SNOMEDCT_CORE|Needle stick injury|Needle prick injury
C0085207|T047|SY|11687002|SNOMEDCT_CORE|Diabetes mellitus arising in pregnancy|Gestational diabetes mellitus
C0085207|T047|SY|11687002|SNOMEDCT_CORE|GDM|Gestational diabetes mellitus
C0085207|T047|SY|11687002|SNOMEDCT_CORE|GDM - Gestational diabetes mellitus|Gestational diabetes mellitus
C0085207|T047|SY|11687002|SNOMEDCT_CORE|Gestational diabetes|Gestational diabetes mellitus
C0085207|T047|PT|11687002|SNOMEDCT_CORE|Gestational diabetes mellitus|Gestational diabetes mellitus
C0085207|T047|FN|11687002|SNOMEDCT_CORE|Gestational diabetes mellitus|Gestational diabetes mellitus
C0085207|T047|IS|11687002|SNOMEDCT_CORE|Gestational diabetes mellitus, NOS|Gestational diabetes mellitus
C0085207|T047|SY|11687002|SNOMEDCT_CORE|Maternal gestational diabetes mellitus|Gestational diabetes mellitus
C0085215|T047|SY|237788002|SNOMEDCT_CORE|POF - Premature ovarian failure|Premature ovarian failure
C0085215|T047|PT|237788002|SNOMEDCT_CORE|Premature ovarian failure|Premature ovarian failure
C0085215|T047|FN|237788002|SNOMEDCT_CORE|Premature ovarian failure|Premature ovarian failure
C0085222|T047|PT|266463007|SNOMEDCT_CORE|Iliopsoas abscess|Iliopsoas abscess
C0085222|T047|FN|266463007|SNOMEDCT_CORE|Iliopsoas abscess|Iliopsoas abscess
C0085222|T047|SY|266463007|SNOMEDCT_CORE|Psoas abscess|Iliopsoas abscess
C0085222|T047|SY|266463007|SNOMEDCT_CORE|Psoas muscle abscess|Iliopsoas abscess
C0085232|T047|SYGB|399291005|SNOMEDCT_CORE|Acquired pharyngo-oesophageal diverticulum|Zenker's diverticulum
C0085232|T047|SY|399291005|SNOMEDCT_CORE|Acquired pharyngoesophageal diverticulum|Zenker's diverticulum
C0085232|T047|SY|399291005|SNOMEDCT_CORE|Hypopharyngeal diverticulum|Zenker's diverticulum
C0085232|T047|SY|399291005|SNOMEDCT_CORE|Pharyngo-oesophageal diverticulum|Zenker's diverticulum
C0085232|T047|SY|399291005|SNOMEDCT_CORE|Pharyngoesophageal diverticulum|Zenker's diverticulum
C0085232|T047|FN|399291005|SNOMEDCT_CORE|Pharyngoesophageal diverticulum|Zenker's diverticulum
C0085232|T047|SY|399291005|SNOMEDCT_CORE|Zenker diverticulum|Zenker's diverticulum
C0085232|T047|PT|399291005|SNOMEDCT_CORE|Zenker's diverticulum|Zenker's diverticulum
C0085232|T047|OF|399291005|SNOMEDCT_CORE|Zenker's diverticulum|Zenker's diverticulum
C0085232|T047|SY|399291005|SNOMEDCT_CORE|Zenker's hypopharyngeal diverticulum|Zenker's diverticulum
C0085273|T047|SY|34730008|SNOMEDCT_CORE|Erythema contagiosum|Primate erythroparvovirus 1 infection
C0085273|T047|SY|34730008|SNOMEDCT_CORE|Erythema infectiosum|Primate erythroparvovirus 1 infection
C0085273|T047|OF|34730008|SNOMEDCT_CORE|Erythema infectiosum|Primate erythroparvovirus 1 infection
C0085273|T047|SY|34730008|SNOMEDCT_CORE|Fifth disease|Primate erythroparvovirus 1 infection
C0085273|T047|SY|34730008|SNOMEDCT_CORE|Parvovirus B19 infection|Primate erythroparvovirus 1 infection
C0085273|T047|PT|34730008|SNOMEDCT_CORE|Primate erythroparvovirus 1 infection|Primate erythroparvovirus 1 infection
C0085273|T047|FN|34730008|SNOMEDCT_CORE|Primate erythroparvovirus 1 infection|Primate erythroparvovirus 1 infection
C0085273|T047|SY|34730008|SNOMEDCT_CORE|Slapped cheek syndrome|Primate erythroparvovirus 1 infection
C0085278|T047|SY|26843008|SNOMEDCT_CORE|Anticardiolipin syndrome|Antiphospholipid syndrome
C0085278|T047|IS|19267009|SNOMEDCT_CORE|Antiphospholipid syndrome|Antiphospholipid syndrome
C0085278|T047|PT|26843008|SNOMEDCT_CORE|Antiphospholipid syndrome|Antiphospholipid syndrome
C0085278|T047|FN|26843008|SNOMEDCT_CORE|Antiphospholipid syndrome|Antiphospholipid syndrome
C0085278|T047|SY|26843008|SNOMEDCT_CORE|APL - Antiphospholipid syndrome|Antiphospholipid syndrome
C0085278|T047|SY|26843008|SNOMEDCT_CORE|APS - Antiphospholipid syndrome|Antiphospholipid syndrome
C0085292|T047|SY|5217008|SNOMEDCT_CORE|Gamma neuron overactivity syndrome|Stiff-man syndrome
C0085292|T047|SY|5217008|SNOMEDCT_CORE|Moersch-Woltman syndrome|Stiff-man syndrome
C0085292|T047|SY|5217008|SNOMEDCT_CORE|Moersch-Woltmann syndrome|Stiff-man syndrome
C0085292|T047|SY|5217008|SNOMEDCT_CORE|Stiff man syndrome|Stiff-man syndrome
C0085292|T047|PT|5217008|SNOMEDCT_CORE|Stiff-man syndrome|Stiff-man syndrome
C0085292|T047|FN|5217008|SNOMEDCT_CORE|Stiff-man syndrome|Stiff-man syndrome
C0085404|T047|SY|79268002|SNOMEDCT_CORE|POEMS - Polyneuropathy organomegaly endocrinopathy monoclonal and skin changes|POEMS syndrome
C0085404|T047|PT|79268002|SNOMEDCT_CORE|POEMS syndrome|POEMS syndrome
C0085404|T047|OF|79268002|SNOMEDCT_CORE|POEMS syndrome|POEMS syndrome
C0085404|T047|SY|79268002|SNOMEDCT_CORE|Polyneuropathy organomegaly endocrinopathy monoclonal gammopathy and skin changes|POEMS syndrome
C0085404|T047|IS|79268002|SNOMEDCT_CORE|Polyneuropathy organomegaly endocrinopathy monoclonal gammopathy and skin changes|POEMS syndrome
C0085404|T047|FN|79268002|SNOMEDCT_CORE|Polyneuropathy, organomegaly, endocrinopathy, monoclonal gammopathy, and skin changes syndrome|POEMS syndrome
C0085404|T047|SY|79268002|SNOMEDCT_CORE|Polyneuropathy, organomegaly, endocrinopathy, monoclonal gammopathy, and skin changes syndrome|POEMS syndrome
C0085404|T047|OF|79268002|SNOMEDCT_CORE|Polyneuropathy, organomegaly, endocrinopathy, monoclonal gammopathy, and skin changes syndrome|POEMS syndrome
C0085413|T047|SY|765330003|SNOMEDCT_CORE|ADPKD - autosomal dominant polycystic kidney disease|Autosomal dominant polycystic kidney disease
C0085413|T047|OAS|28728008|SNOMEDCT_CORE|ADPKD - Autosomal dominant polycystic kidney disease|Autosomal dominant polycystic kidney disease
C0085413|T047|OAS|28728008|SNOMEDCT_CORE|Autosomal dominant adult polycystic kidney disease|Autosomal dominant polycystic kidney disease
C0085413|T047|OAS|28728008|SNOMEDCT_CORE|Autosomal dominant polycystic kidney disease|Autosomal dominant polycystic kidney disease
C0085413|T047|PT|765330003|SNOMEDCT_CORE|Autosomal dominant polycystic kidney disease|Autosomal dominant polycystic kidney disease
C0085413|T047|FN|765330003|SNOMEDCT_CORE|Autosomal dominant polycystic kidney disease|Autosomal dominant polycystic kidney disease
C0085413|T047|OAP|28728008|SNOMEDCT_CORE|Polycystic kidney disease, adult type|Autosomal dominant polycystic kidney disease
C0085413|T047|OAF|28728008|SNOMEDCT_CORE|Polycystic kidney disease, adult type|Autosomal dominant polycystic kidney disease
C0085413|T047|OAS|28728008|SNOMEDCT_CORE|Polycystic kidneys - adult type|Autosomal dominant polycystic kidney disease
C0085417|T047|PT|361123003|SNOMEDCT_CORE|Psychomotor epilepsy|Psychomotor epilepsy
C0085417|T047|FN|361123003|SNOMEDCT_CORE|Psychomotor epilepsy|Psychomotor epilepsy
C0085435|T047|SY|239783001|SNOMEDCT_CORE|Arthritis occurring after infection|Post-infective arthritis
C0085435|T047|PT|239783001|SNOMEDCT_CORE|Post-infective arthritis|Post-infective arthritis
C0085435|T047|FN|239783001|SNOMEDCT_CORE|Post-infective arthritis|Post-infective arthritis
C0085435|T047|SY|239783001|SNOMEDCT_CORE|Post-infective arthropathy|Post-infective arthritis
C0085435|T047|IS|239783001|SNOMEDCT_CORE|Reactive arthritis|Post-infective arthritis
C0085576|T047|PTGB|234349007|SNOMEDCT_CORE|Microcytic anaemia|Microcytic anemia
C0085576|T047|PT|234349007|SNOMEDCT_CORE|Microcytic anemia|Microcytic anemia
C0085576|T047|FN|234349007|SNOMEDCT_CORE|Microcytic anemia|Microcytic anemia
C0085577|T047|PTGB|300980002|SNOMEDCT_CORE|Normocytic anaemia|Normocytic anemia
C0085577|T047|PT|300980002|SNOMEDCT_CORE|Normocytic anemia|Normocytic anemia
C0085577|T047|FN|300980002|SNOMEDCT_CORE|Normocytic anemia|Normocytic anemia
C0085578|T047|SYGB|19442009|SNOMEDCT_CORE|Thalassaemia minor|Thalassemia minor
C0085578|T047|SY|19442009|SNOMEDCT_CORE|Thalassemia minor|Thalassemia minor
C0085580|T047|PT|59621000|SNOMEDCT_CORE|Essential hypertension|Essential hypertension
C0085580|T047|FN|59621000|SNOMEDCT_CORE|Essential hypertension|Essential hypertension
C0085580|T047|IS|59621000|SNOMEDCT_CORE|Essential hypertension, NOS|Essential hypertension
C0085580|T047|SY|59621000|SNOMEDCT_CORE|Idiopathic hypertension|Essential hypertension
C0085580|T047|SY|59621000|SNOMEDCT_CORE|Primary hypertension|Essential hypertension
C0085580|T047|IS|59621000|SNOMEDCT_CORE|Primary hypertension, NOS|Essential hypertension
C0085580|T047|SY|59621000|SNOMEDCT_CORE|Systemic primary arterial hypertension|Essential hypertension
C0085581|T047|PT|36485005|SNOMEDCT_CORE|Restrictive lung disease|Restrictive lung disease
C0085581|T047|FN|36485005|SNOMEDCT_CORE|Restrictive lung disease|Restrictive lung disease
C0085581|T047|IS|36485005|SNOMEDCT_CORE|Restrictive lung disease, NOS|Restrictive lung disease
C0085584|T047|SY|81308009|SNOMEDCT_CORE|Encephalopathy|Encephalopathy
C0085593|T184|PT|43724002|SNOMEDCT_CORE|Chill|Chill
C0085593|T184|FN|43724002|SNOMEDCT_CORE|Chill|Chill
C0085593|T184|IS|43724002|SNOMEDCT_CORE|Chills|Chill
C0085598|T046|PT|199047001|SNOMEDCT_CORE|False labor|False labor
C0085598|T046|FN|199047001|SNOMEDCT_CORE|False labor|False labor
C0085598|T046|OF|199047001|SNOMEDCT_CORE|False labor|False labor
C0085598|T046|PTGB|199047001|SNOMEDCT_CORE|False labour|False labor
C0085598|T046|SY|199047001|SNOMEDCT_CORE|Spurious labor|False labor
C0085598|T046|SYGB|199047001|SNOMEDCT_CORE|Spurious labour|False labor
C0085602|T184|SY|17173007|SNOMEDCT_CORE|Always thirsty|Excessive thirst
C0085602|T184|SY|17173007|SNOMEDCT_CORE|Desperate to drink|Excessive thirst
C0085602|T184|PT|17173007|SNOMEDCT_CORE|Excessive thirst|Excessive thirst
C0085602|T184|FN|17173007|SNOMEDCT_CORE|Excessive thirst|Excessive thirst
C0085602|T184|SY|17173007|SNOMEDCT_CORE|Keen for fluids|Excessive thirst
C0085602|T184|IS|17173007|SNOMEDCT_CORE|Polydipsia|Excessive thirst
C0085605|T047|PT|59927004|SNOMEDCT_CORE|Hepatic failure|Hepatic failure
C0085605|T047|FN|59927004|SNOMEDCT_CORE|Hepatic failure|Hepatic failure
C0085605|T047|IS|59927004|SNOMEDCT_CORE|Hepatic failure, NOS|Hepatic failure
C0085605|T047|SY|59927004|SNOMEDCT_CORE|Liver decompensation|Hepatic failure
C0085605|T047|IS|59927004|SNOMEDCT_CORE|Liver decompensation, NOS|Hepatic failure
C0085605|T047|SY|59927004|SNOMEDCT_CORE|Liver failure|Hepatic failure
C0085605|T047|SY|59927004|SNOMEDCT_CORE|Liver function failure|Hepatic failure
C0085605|T047|IS|59927004|SNOMEDCT_CORE|Liver function failure, NOS|Hepatic failure
C0085606|T184|SY|75088002|SNOMEDCT_CORE|Must hurry to pass urine|Urgent desire to urinate
C0085606|T184|SY|75088002|SNOMEDCT_CORE|Precipitancy of micturition|Urgent desire to urinate
C0085606|T184|SY|75088002|SNOMEDCT_CORE|Precipitancy of urine|Urgent desire to urinate
C0085606|T184|SY|75088002|SNOMEDCT_CORE|Urgency - urination|Urgent desire to urinate
C0085606|T184|SY|75088002|SNOMEDCT_CORE|Urgency of micturition|Urgent desire to urinate
C0085606|T184|SY|75088002|SNOMEDCT_CORE|Urgency to micturate|Urgent desire to urinate
C0085606|T184|SY|75088002|SNOMEDCT_CORE|Urgency to pass urine|Urgent desire to urinate
C0085606|T184|PT|75088002|SNOMEDCT_CORE|Urgent desire to urinate|Urgent desire to urinate
C0085606|T184|FN|75088002|SNOMEDCT_CORE|Urgent desire to urinate|Urgent desire to urinate
C0085606|T184|SY|75088002|SNOMEDCT_CORE|Urging to urinate|Urgent desire to urinate
C0085606|T184|SY|75088002|SNOMEDCT_CORE|Urinary precipitancy|Urgent desire to urinate
C0085606|T184|IS|75088002|SNOMEDCT_CORE|Urinary urgency|Urgent desire to urinate
C0085610|T046|PT|49710005|SNOMEDCT_CORE|Sinus bradycardia|Sinus bradycardia
C0085610|T046|FN|49710005|SNOMEDCT_CORE|Sinus bradycardia|Sinus bradycardia
C0085611|T046|PT|17366009|SNOMEDCT_CORE|Atrial arrhythmia|Atrial arrhythmia
C0085611|T046|FN|17366009|SNOMEDCT_CORE|Atrial arrhythmia|Atrial arrhythmia
C0085611|T046|IS|17366009|SNOMEDCT_CORE|Atrial arrhythmia, NOS|Atrial arrhythmia
C0085612|T047|PT|44103008|SNOMEDCT_CORE|Ventricular arrhythmia|Ventricular arrhythmia
C0085612|T047|FN|44103008|SNOMEDCT_CORE|Ventricular arrhythmia|Ventricular arrhythmia
C0085612|T047|IS|44103008|SNOMEDCT_CORE|Ventricular arrhythmia, NOS|Ventricular arrhythmia
C0085614|T047|PT|270492004|SNOMEDCT_CORE|First degree atrioventricular block|First degree atrioventricular block
C0085614|T047|FN|270492004|SNOMEDCT_CORE|First degree atrioventricular block|First degree atrioventricular block
C0085614|T047|SY|270492004|SNOMEDCT_CORE|First degree heart block|First degree atrioventricular block
C0085614|T047|SY|270492004|SNOMEDCT_CORE|Incomplete atrioventricular block, first degree|First degree atrioventricular block
C0085615|T047|SY|59118001|SNOMEDCT_CORE|RBBB - Right bundle branch block|Right bundle branch block
C0085615|T047|PT|59118001|SNOMEDCT_CORE|Right bundle branch block|Right bundle branch block
C0085615|T047|FN|59118001|SNOMEDCT_CORE|Right bundle branch block|Right bundle branch block
C0085615|T047|SY|59118001|SNOMEDCT_CORE|Right fascicular block|Right bundle branch block
C0085616|T046|SY|71772004|SNOMEDCT_CORE|Angiospasm|Vasospasm
C0085616|T046|IS|71772004|SNOMEDCT_CORE|Angiospasm, NOS|Vasospasm
C0085616|T046|SY|71772004|SNOMEDCT_CORE|Blood vessel spasm|Vasospasm
C0085616|T046|SY|71772004|SNOMEDCT_CORE|Vascular spasm|Vasospasm
C0085616|T046|PT|71772004|SNOMEDCT_CORE|Vasospasm|Vasospasm
C0085616|T046|FN|71772004|SNOMEDCT_CORE|Vasospasm|Vasospasm
C0085616|T046|IS|71772004|SNOMEDCT_CORE|Vasospasm, NOS|Vasospasm
C0085619|T033|SY|62744007|SNOMEDCT_CORE|Breathlessness lying flat|Orthopnea
C0085619|T033|IS|62744007|SNOMEDCT_CORE|Must sit up to breath|Orthopnea
C0085619|T033|PT|62744007|SNOMEDCT_CORE|Orthopnea|Orthopnea
C0085619|T033|FN|62744007|SNOMEDCT_CORE|Orthopnea|Orthopnea
C0085619|T033|PTGB|62744007|SNOMEDCT_CORE|Orthopnoea|Orthopnea
C0085624|T184|PT|90673000|SNOMEDCT_CORE|Burning sensation|Burning sensation
C0085624|T184|FN|90673000|SNOMEDCT_CORE|Burning sensation|Burning sensation
C0085624|T184|IS|90673000|SNOMEDCT_CORE|Sensation of burning of skin|Burning sensation
C0085631|T184|SY|24199005|SNOMEDCT_CORE|Agitated|Feeling agitated
C0085631|T184|SY|24199005|SNOMEDCT_CORE|Agitated behavior|Feeling agitated
C0085631|T184|SYGB|24199005|SNOMEDCT_CORE|Agitated behaviour|Feeling agitated
C0085631|T184|SY|24199005|SNOMEDCT_CORE|Agitation|Feeling agitated
C0085631|T184|PT|24199005|SNOMEDCT_CORE|Feeling agitated|Feeling agitated
C0085631|T184|FN|24199005|SNOMEDCT_CORE|Feeling agitated|Feeling agitated
C0085631|T184|SY|24199005|SNOMEDCT_CORE|Unable to keep still|Feeling agitated
C0085633|T048|SY|18963009|SNOMEDCT_CORE|Changeable mood|Mood swings
C0085633|T048|SY|18963009|SNOMEDCT_CORE|Emotional instability|Mood swings
C0085633|T048|SY|18963009|SNOMEDCT_CORE|Emotional lability|Mood swings
C0085633|T048|SY|18963009|SNOMEDCT_CORE|Emotionally labile|Mood swings
C0085633|T048|SY|18963009|SNOMEDCT_CORE|Labile in mood|Mood swings
C0085633|T048|SY|18963009|SNOMEDCT_CORE|Labile mood|Mood swings
C0085633|T048|SY|18963009|SNOMEDCT_CORE|Mood swing|Mood swings
C0085633|T048|PT|18963009|SNOMEDCT_CORE|Mood swings|Mood swings
C0085633|T048|FN|18963009|SNOMEDCT_CORE|Mood swings|Mood swings
C0085633|T048|SY|18963009|SNOMEDCT_CORE|Unstable mood|Mood swings
C0085633|T048|SY|18963009|SNOMEDCT_CORE|Variable mood|Mood swings
C0085635|T047|SY|56170001|SNOMEDCT_CORE|Flashes|Photopsia
C0085635|T047|SY|56170001|SNOMEDCT_CORE|Light flashes|Photopsia
C0085635|T047|PT|56170001|SNOMEDCT_CORE|Photopsia|Photopsia
C0085635|T047|FN|56170001|SNOMEDCT_CORE|Photopsia|Photopsia
C0085639|T033|PT|1912002|SNOMEDCT_CORE|Fall|Falls
C0085639|T033|OF|1912002|SNOMEDCT_CORE|Fall|Falls
C0085639|T033|FN|1912002|SNOMEDCT_CORE|Fall|Falls
C0085639|T033|IS|1912002|SNOMEDCT_CORE|Fall, NOS|Falls
C0085639|T033|PT|161898004|SNOMEDCT_CORE|Falls|Falls
C0085639|T033|IS|1912002|SNOMEDCT_CORE|Falls|Falls
C0085639|T033|FN|161898004|SNOMEDCT_CORE|Falls|Falls
C0085642|T047|SY|238772004|SNOMEDCT_CORE|Livedo racemosa|Livedo reticularis
C0085642|T047|PT|238772004|SNOMEDCT_CORE|Livedo reticularis|Livedo reticularis
C0085642|T047|FN|238772004|SNOMEDCT_CORE|Livedo reticularis|Livedo reticularis
C0085648|T047|IS|71307009|SNOMEDCT_CORE|Synovial cyst|Synovial cyst
C0085648|T047|PT|240205003|SNOMEDCT_CORE|Synovial cyst|Synovial cyst
C0085648|T047|FN|240205003|SNOMEDCT_CORE|Synovial cyst|Synovial cyst
C0085648|T047|IS|71307009|SNOMEDCT_CORE|Synovial cyst, NOS|Synovial cyst
C0085649|T046|PT|271809000|SNOMEDCT_CORE|Peripheral edema|Peripheral edema
C0085649|T046|FN|271809000|SNOMEDCT_CORE|Peripheral edema|Peripheral edema
C0085649|T046|PTGB|271809000|SNOMEDCT_CORE|Peripheral oedema|Peripheral edema
C0085653|T191|SY|39629007|SNOMEDCT_CORE|PG - Pyogenic granuloma|Pyogenic granuloma
C0085653|T191|PT|200722003|SNOMEDCT_CORE|Pyogenic granuloma|Pyogenic granuloma
C0085653|T191|OF|200722003|SNOMEDCT_CORE|Pyogenic granuloma|Pyogenic granuloma
C0085653|T191|FN|200722003|SNOMEDCT_CORE|Pyogenic granuloma|Pyogenic granuloma
C0085655|T047|SY|31384009|SNOMEDCT_CORE|Neuromyositis|Polymyositis
C0085655|T047|SY|31384009|SNOMEDCT_CORE|PM - Polymyositis|Polymyositis
C0085655|T047|PT|31384009|SNOMEDCT_CORE|Polymyositis|Polymyositis
C0085655|T047|FN|31384009|SNOMEDCT_CORE|Polymyositis|Polymyositis
C0085656|T047|SY|81418003|SNOMEDCT_CORE|Discoid eczema|Nummular eczema
C0085656|T047|IS|81418003|SNOMEDCT_CORE|Exudative neurodermatitis|Nummular eczema
C0085656|T047|SY|81418003|SNOMEDCT_CORE|Nummular dermatitis|Nummular eczema
C0085656|T047|PT|81418003|SNOMEDCT_CORE|Nummular eczema|Nummular eczema
C0085656|T047|FN|81418003|SNOMEDCT_CORE|Nummular eczema|Nummular eczema
C0085656|T047|SY|81418003|SNOMEDCT_CORE|Nummular eczematous dermatitis|Nummular eczema
C0085656|T047|IS|81418003|SNOMEDCT_CORE|Nummular neurodermatitis|Nummular eczema
C0085657|T047|PT|402296004|SNOMEDCT_CORE|Pityriasis alba|Pityriasis alba
C0085657|T047|FN|402296004|SNOMEDCT_CORE|Pityriasis alba|Pityriasis alba
C0085658|T047|SY|414492009|SNOMEDCT_CORE|Dermatitis infectiosa eczematoides|Infectious eczematoid dermatitis
C0085658|T047|PT|414492009|SNOMEDCT_CORE|Infectious eczematoid dermatitis|Infectious eczematoid dermatitis
C0085658|T047|SY|414492009|SNOMEDCT_CORE|Infective eczematoid dermatitis|Infectious eczematoid dermatitis
C0085658|T047|FN|414492009|SNOMEDCT_CORE|Infective eczematoid dermatitis|Infectious eczematoid dermatitis
C0085661|T047|IS|75789001|SNOMEDCT_CORE|Detachment of nail|Onycholysis
C0085661|T047|SY|75789001|SNOMEDCT_CORE|Detachment of nail plate|Onycholysis
C0085661|T047|PT|75789001|SNOMEDCT_CORE|Onycholysis|Onycholysis
C0085661|T047|FN|75789001|SNOMEDCT_CORE|Onycholysis|Onycholysis
C0085661|T047|SY|75789001|SNOMEDCT_CORE|Separation of nail plate|Onycholysis
C0085666|T047|SY|195382003|SNOMEDCT_CORE|Arterial spider|Spider nevus
C0085666|T047|SY|195382003|SNOMEDCT_CORE|Arterial spider of skin|Spider nevus
C0085666|T047|SYGB|195382003|SNOMEDCT_CORE|Naevus araneus of skin|Spider nevus
C0085666|T047|SY|195382003|SNOMEDCT_CORE|Nevus araneus of skin|Spider nevus
C0085666|T047|SY|195382003|SNOMEDCT_CORE|Spider angioma|Spider nevus
C0085666|T047|SY|195382003|SNOMEDCT_CORE|Spider angioma of skin|Spider nevus
C0085666|T047|PTGB|195382003|SNOMEDCT_CORE|Spider naevus|Spider nevus
C0085666|T047|SYGB|195382003|SNOMEDCT_CORE|Spider naevus of skin|Spider nevus
C0085666|T047|PT|195382003|SNOMEDCT_CORE|Spider nevus|Spider nevus
C0085666|T047|FN|195382003|SNOMEDCT_CORE|Spider nevus|Spider nevus
C0085666|T047|SY|195382003|SNOMEDCT_CORE|Spider nevus of skin|Spider nevus
C0085666|T047|SY|195382003|SNOMEDCT_CORE|Spider telangiectasia|Spider nevus
C0085666|T047|SY|195382003|SNOMEDCT_CORE|Spider telangiectasis of skin|Spider nevus
C0085666|T047|SYGB|195382003|SNOMEDCT_CORE|Stellar naevus of skin|Spider nevus
C0085666|T047|SY|195382003|SNOMEDCT_CORE|Stellar nevus of skin|Spider nevus
C0085666|T047|SYGB|195382003|SNOMEDCT_CORE|Telangiectatic naevus|Spider nevus
C0085666|T047|SY|195382003|SNOMEDCT_CORE|Telangiectatic nevus|Spider nevus
C0085669|T191|PTGB|91855006|SNOMEDCT_CORE|Acute leukaemia|Acute leukemia
C0085669|T191|SYGB|91855006|SNOMEDCT_CORE|Acute leukaemia, disease|Acute leukemia
C0085669|T191|PT|91855006|SNOMEDCT_CORE|Acute leukemia|Acute leukemia
C0085669|T191|FN|91855006|SNOMEDCT_CORE|Acute leukemia, disease|Acute leukemia
C0085669|T191|SY|91855006|SNOMEDCT_CORE|Acute leukemia, disease|Acute leukemia
C0085677|T047|SY|7916009|SNOMEDCT_CORE|Alcohol-induced polyneuropathy|Alcoholic polyneuropathy
C0085677|T047|SY|7916009|SNOMEDCT_CORE|Alcoholic peripheral neuropathy|Alcoholic polyneuropathy
C0085677|T047|PT|7916009|SNOMEDCT_CORE|Alcoholic polyneuropathy|Alcoholic polyneuropathy
C0085677|T047|FN|7916009|SNOMEDCT_CORE|Alcoholic polyneuropathy|Alcoholic polyneuropathy
C0085681|T047|PTGB|20165001|SNOMEDCT_CORE|Hyperphosphataemia|Hyperphosphatemia
C0085681|T047|FN|20165001|SNOMEDCT_CORE|Hyperphosphatemia|Hyperphosphatemia
C0085681|T047|PT|20165001|SNOMEDCT_CORE|Hyperphosphatemia|Hyperphosphatemia
C0085682|T047|PTGB|4996001|SNOMEDCT_CORE|Hypophosphataemia|Hypophosphatemia
C0085682|T047|IS|4996001|SNOMEDCT_CORE|Hypophosphataemia, NOS|Hypophosphatemia
C0085682|T047|PT|4996001|SNOMEDCT_CORE|Hypophosphatemia|Hypophosphatemia
C0085682|T047|FN|4996001|SNOMEDCT_CORE|Hypophosphatemia|Hypophosphatemia
C0085682|T047|IS|4996001|SNOMEDCT_CORE|Hypophosphatemia, NOS|Hypophosphatemia
C0085684|T047|SY|6077001|SNOMEDCT_CORE|Dropfoot|Foot-drop
C0085684|T047|SY|6077001|SNOMEDCT_CORE|FD - Foot-drop|Foot-drop
C0085684|T047|PT|6077001|SNOMEDCT_CORE|Foot-drop|Foot-drop
C0085684|T047|FN|6077001|SNOMEDCT_CORE|Foot-drop|Foot-drop
C0085684|T047|SY|6077001|SNOMEDCT_CORE|Footdrop|Foot-drop
C0085690|T047|SY|414521009|SNOMEDCT_CORE|Hordeolum internum|Internal hordeolum
C0085690|T047|PT|414521009|SNOMEDCT_CORE|Internal hordeolum|Internal hordeolum
C0085690|T047|FN|414521009|SNOMEDCT_CORE|Internal hordeolum|Internal hordeolum
C0085692|T047|PTGB|87696004|SNOMEDCT_CORE|Haemorrhagic cystitis|Hemorrhagic cystitis
C0085692|T047|PT|87696004|SNOMEDCT_CORE|Hemorrhagic cystitis|Hemorrhagic cystitis
C0085692|T047|FN|87696004|SNOMEDCT_CORE|Hemorrhagic cystitis|Hemorrhagic cystitis
C0085693|T047|FN|85189001|SNOMEDCT_CORE|Acute appendicitis|Acute appendicitis
C0085693|T047|PT|85189001|SNOMEDCT_CORE|Acute appendicitis|Acute appendicitis
C0085693|T047|IS|85189001|SNOMEDCT_CORE|Acute appendicitis, NOS|Acute appendicitis
C0085694|T047|PT|20824003|SNOMEDCT_CORE|Chronic cholecystitis|Chronic cholecystitis
C0085694|T047|FN|20824003|SNOMEDCT_CORE|Chronic cholecystitis|Chronic cholecystitis
C0085694|T047|IS|20824003|SNOMEDCT_CORE|Chronic cholecystitis, NOS|Chronic cholecystitis
C0085695|T047|SY|8493009|SNOMEDCT_CORE|CG - Chronic gastritis|Chronic gastritis
C0085695|T047|PT|8493009|SNOMEDCT_CORE|Chronic gastritis|Chronic gastritis
C0085695|T047|FN|8493009|SNOMEDCT_CORE|Chronic gastritis|Chronic gastritis
C0085695|T047|IS|8493009|SNOMEDCT_CORE|Chronic gastritis, NOS|Chronic gastritis
C0085696|T047|PT|19905009|SNOMEDCT_CORE|Chronic prostatitis|Chronic prostatitis
C0085696|T047|FN|19905009|SNOMEDCT_CORE|Chronic prostatitis|Chronic prostatitis
C0085700|T047|PT|63198006|SNOMEDCT_CORE|Chondromalacia|Chondromalacia
C0085700|T047|FN|63198006|SNOMEDCT_CORE|Chondromalacia|Chondromalacia
C0085700|T047|IS|63198006|SNOMEDCT_CORE|Chondromalacia, NOS|Chondromalacia
C0085702|T047|PT|19636003|SNOMEDCT_CORE|Monocytosis|Monocytosis
C0085702|T047|FN|19636003|SNOMEDCT_CORE|Monocytosis|Monocytosis
C0085702|T047|IS|19636003|SNOMEDCT_CORE|Monocytosis, NOS|Monocytosis
C0085762|T048|SY|15167005|SNOMEDCT_CORE|AA - Alcohol abuse|Alcohol abuse
C0085762|T048|PT|15167005|SNOMEDCT_CORE|Alcohol abuse|Alcohol abuse
C0085762|T048|FN|15167005|SNOMEDCT_CORE|Alcohol abuse|Alcohol abuse
C0085762|T048|SY|15167005|SNOMEDCT_CORE|Ethanol abuse|Alcohol abuse
C0085786|T047|IS|45157009|SNOMEDCT_CORE|Diffuse idiopathic pulmonary fibrosis|Diffuse interstitial pulmonary fibrosis
C0085786|T047|IS|45157009|SNOMEDCT_CORE|Diffuse interstitial pulmonary fibrosis|Diffuse interstitial pulmonary fibrosis
C0085786|T047|PT|196125002|SNOMEDCT_CORE|Diffuse interstitial pulmonary fibrosis|Diffuse interstitial pulmonary fibrosis
C0085786|T047|FN|196125002|SNOMEDCT_CORE|Diffuse interstitial pulmonary fibrosis|Diffuse interstitial pulmonary fibrosis
C0085786|T047|SY|196125002|SNOMEDCT_CORE|DIPF - Diffuse interstitial pulmonary fibrosis|Diffuse interstitial pulmonary fibrosis
C0085786|T047|SY|196125002|SNOMEDCT_CORE|Fibrosing alveolitis|Diffuse interstitial pulmonary fibrosis
C0085786|T047|IS|45157009|SNOMEDCT_CORE|Hamman-Rich syndrome|Diffuse interstitial pulmonary fibrosis
C0085786|T047|OAS|45157009|SNOMEDCT_CORE|Idiopathic fibrosing alveolitis|Diffuse interstitial pulmonary fibrosis
C0085786|T047|OAF|45157009|SNOMEDCT_CORE|Idiopathic fibrosing alveolitis|Diffuse interstitial pulmonary fibrosis
C0085786|T047|SY|196125002|SNOMEDCT_CORE|UIP - Usual interstitial pneumonitis|Diffuse interstitial pulmonary fibrosis
C0085786|T047|SY|196125002|SNOMEDCT_CORE|Usual interstitial pneumonitis|Diffuse interstitial pulmonary fibrosis
C0085932|T047|SY|7231009|SNOMEDCT_CORE|Bullous dermatitis|Bullous dermatosis
C0085932|T047|IS|7231009|SNOMEDCT_CORE|Bullous dermatitis, NOS|Bullous dermatosis
C0085932|T047|SY|7231009|SNOMEDCT_CORE|Bullous dermatoses|Bullous dermatosis
C0085932|T047|PT|7231009|SNOMEDCT_CORE|Bullous dermatosis|Bullous dermatosis
C0085932|T047|FN|7231009|SNOMEDCT_CORE|Bullous dermatosis|Bullous dermatosis
C0085932|T047|IS|7231009|SNOMEDCT_CORE|Bullous dermatosis, NOS|Bullous dermatosis
C0085988|T033|PT|199397009|SNOMEDCT_CORE|Cephalopelvic disproportion|Cephalopelvic disproportion
C0085988|T033|FN|199397009|SNOMEDCT_CORE|Cephalopelvic disproportion|Cephalopelvic disproportion
C0085988|T033|SY|199397009|SNOMEDCT_CORE|CPD - Cephalopelvic disproportion|Cephalopelvic disproportion
C0085988|T033|SY|199397009|SNOMEDCT_CORE|Disproportion of mixed maternal AND fetal origin with normally formed fetus|Cephalopelvic disproportion
C0085988|T033|SY|199397009|SNOMEDCT_CORE|Disproportion of mixed maternal AND foetal origin with normally formed foetus|Cephalopelvic disproportion
C0086209|T048|PT|442347009|SNOMEDCT_CORE|Emotional stress|Emotional stress
C0086209|T048|FN|442347009|SNOMEDCT_CORE|Emotional stress|Emotional stress
C0086227|T047|PT|266162007|SNOMEDCT_CORE|Enterobiasis|Enterobiasis
C0086227|T047|FN|266162007|SNOMEDCT_CORE|Enterobiasis|Enterobiasis
C0086227|T047|SY|266162007|SNOMEDCT_CORE|Enterobiasis - threadworm|Enterobiasis
C0086227|T047|SY|266162007|SNOMEDCT_CORE|Enterobiosis|Enterobiasis
C0086227|T047|SY|266162007|SNOMEDCT_CORE|Pinworm disease|Enterobiasis
C0086227|T047|SY|266162007|SNOMEDCT_CORE|Pinworm infection|Enterobiasis
C0086227|T047|SY|266162007|SNOMEDCT_CORE|Threadworm infection|Enterobiasis
C0086438|T047|PTGB|119250001|SNOMEDCT_CORE|Hypogammaglobulinaemia|Hypogammaglobulinemia
C0086438|T047|IS|119250001|SNOMEDCT_CORE|Hypogammaglobulinemia|Hypogammaglobulinemia
C0086438|T047|PT|119250001|SNOMEDCT_CORE|Hypogammaglobulinemia|Hypogammaglobulinemia
C0086438|T047|FN|119250001|SNOMEDCT_CORE|Hypogammaglobulinemia|Hypogammaglobulinemia
C0086501|T020|SY|201040000|SNOMEDCT_CORE|Keratoma|Keratoma
C0086543|T020|IS|193570009|SNOMEDCT_CORE|Cat. - Cataract|Cataract
C0086543|T020|PT|193570009|SNOMEDCT_CORE|Cataract|Cataract
C0086543|T020|FN|193570009|SNOMEDCT_CORE|Cataract|Cataract
C0086565|T033|SY|75183008|SNOMEDCT_CORE|Abnormal hepatic function|Abnormal liver function
C0086565|T033|PT|75183008|SNOMEDCT_CORE|Abnormal liver function|Abnormal liver function
C0086565|T033|FN|75183008|SNOMEDCT_CORE|Abnormal liver function|Abnormal liver function
C0086666|T047|SY|4557003|SNOMEDCT_CORE|Pre-infarction syndrome|Preinfarction syndrome
C0086666|T047|SY|4557003|SNOMEDCT_CORE|Preinfarction angina|Preinfarction syndrome
C0086666|T047|PT|4557003|SNOMEDCT_CORE|Preinfarction syndrome|Preinfarction syndrome
C0086666|T047|FN|4557003|SNOMEDCT_CORE|Preinfarction syndrome|Preinfarction syndrome
C0086692|T191|PT|20376005|SNOMEDCT_CORE|Benign neoplastic disease|Benign neoplastic disease
C0086692|T191|FN|20376005|SNOMEDCT_CORE|Benign neoplastic disease|Benign neoplastic disease
C0086769|T048|PT|225624000|SNOMEDCT_CORE|Panic attack|Panic attack
C0086769|T048|FN|225624000|SNOMEDCT_CORE|Panic attack|Panic attack
C0086809|T190|SY|254677004|SNOMEDCT_CORE|Pilar cyst|Pilar cyst
C0086809|T190|IS|419603000|SNOMEDCT_CORE|Wen|Pilar cyst
C0086981|T047|SY|83901003|SNOMEDCT_CORE|Sicca syndrome|Sicca syndrome
C0087031|T047|SY|201796004|SNOMEDCT_CORE|Juvenile onset Still's disease|Still's disease
C0087031|T047|IS|201796004|SNOMEDCT_CORE|Still's disease|Still's disease
C0149507|T047|PT|194005002|SNOMEDCT_CORE|Orbital cellulitis|Orbital cellulitis
C0149507|T047|FN|194005002|SNOMEDCT_CORE|Orbital cellulitis|Orbital cellulitis
C0149507|T047|SY|194005002|SNOMEDCT_CORE|Postseptal orbital cellulitis|Orbital cellulitis
C0149512|T047|IS|15805002|SNOMEDCT_CORE|Acute infection of nasal sinus, NOS|Acute sinusitis
C0149512|T047|SY|15805002|SNOMEDCT_CORE|Acute infection of sinus|Acute sinusitis
C0149512|T047|SY|15805002|SNOMEDCT_CORE|Acute inflammation of nasal sinus|Acute sinusitis
C0149512|T047|IS|15805002|SNOMEDCT_CORE|Acute inflammation of nasal sinus, NOS|Acute sinusitis
C0149512|T047|SY|15805002|SNOMEDCT_CORE|Acute inflammation of sinus|Acute sinusitis
C0149512|T047|PT|15805002|SNOMEDCT_CORE|Acute sinusitis|Acute sinusitis
C0149512|T047|FN|15805002|SNOMEDCT_CORE|Acute sinusitis|Acute sinusitis
C0149512|T047|IS|15805002|SNOMEDCT_CORE|Acute sinusitis, NOS|Acute sinusitis
C0149514|T047|PT|10509002|SNOMEDCT_CORE|Acute bronchitis|Acute bronchitis
C0149514|T047|FN|10509002|SNOMEDCT_CORE|Acute bronchitis|Acute bronchitis
C0149514|T047|IS|10509002|SNOMEDCT_CORE|Acute bronchitis, NOS|Acute bronchitis
C0149516|T047|SY|40055000|SNOMEDCT_CORE|Chronic infection of sinus|Chronic sinusitis
C0149516|T047|IS|40055000|SNOMEDCT_CORE|Chronic infection of sinus, NOS|Chronic sinusitis
C0149516|T047|SY|40055000|SNOMEDCT_CORE|Chronic rhinosinusitis|Chronic sinusitis
C0149516|T047|PT|40055000|SNOMEDCT_CORE|Chronic sinusitis|Chronic sinusitis
C0149516|T047|FN|40055000|SNOMEDCT_CORE|Chronic sinusitis|Chronic sinusitis
C0149516|T047|IS|40055000|SNOMEDCT_CORE|Chronic sinusitis, NOS|Chronic sinusitis
C0149517|T047|PT|90979004|SNOMEDCT_CORE|Chronic tonsillitis|Chronic tonsillitis
C0149517|T047|FN|90979004|SNOMEDCT_CORE|Chronic tonsillitis|Chronic tonsillitis
C0149518|T047|PT|25458004|SNOMEDCT_CORE|Acute gastritis|Acute gastritis
C0149518|T047|FN|25458004|SNOMEDCT_CORE|Acute gastritis|Acute gastritis
C0149520|T047|PT|65275009|SNOMEDCT_CORE|Acute cholecystitis|Acute cholecystitis
C0149520|T047|FN|65275009|SNOMEDCT_CORE|Acute cholecystitis|Acute cholecystitis
C0149520|T047|IS|65275009|SNOMEDCT_CORE|Inflamed gallbladder|Acute cholecystitis
C0149521|T047|PT|235494005|SNOMEDCT_CORE|Chronic pancreatitis|Chronic pancreatitis
C0149521|T047|FN|235494005|SNOMEDCT_CORE|Chronic pancreatitis|Chronic pancreatitis
C0149521|T047|SY|235494005|SNOMEDCT_CORE|CP - Chronic pancreatitis|Chronic pancreatitis
C0149523|T047|PT|68226007|SNOMEDCT_CORE|Acute cystitis|Acute cystitis
C0149523|T047|FN|68226007|SNOMEDCT_CORE|Acute cystitis|Acute cystitis
C0149524|T047|PT|79411002|SNOMEDCT_CORE|Acute prostatitis|Acute prostatitis
C0149524|T047|FN|79411002|SNOMEDCT_CORE|Acute prostatitis|Acute prostatitis
C0149526|T047|PT|40178009|SNOMEDCT_CORE|Allergic urticaria|Allergic urticaria
C0149526|T047|FN|40178009|SNOMEDCT_CORE|Allergic urticaria|Allergic urticaria
C0149531|T037|PT|77493009|SNOMEDCT_CORE|Fracture of pelvis|Fracture of pelvis
C0149531|T037|FN|77493009|SNOMEDCT_CORE|Fracture of pelvis|Fracture of pelvis
C0149531|T037|IS|77493009|SNOMEDCT_CORE|Fracture of pelvis, NOS|Fracture of pelvis
C0149531|T037|SY|77493009|SNOMEDCT_CORE|Pelvic fracture|Fracture of pelvis
C0149532|T037|SY|47609003|SNOMEDCT_CORE|FB Esophagus|Foreign body in esophagus
C0149532|T037|SYGB|47609003|SNOMEDCT_CORE|FB Oesophagus|Foreign body in esophagus
C0149532|T037|PT|47609003|SNOMEDCT_CORE|Foreign body in esophagus|Foreign body in esophagus
C0149532|T037|FN|47609003|SNOMEDCT_CORE|Foreign body in esophagus|Foreign body in esophagus
C0149532|T037|PTGB|47609003|SNOMEDCT_CORE|Foreign body in oesophagus|Foreign body in esophagus
C0149612|T033|SY|165084003|SNOMEDCT_CORE|Exercise ECG abnormal|Exercise tolerance test abnormal
C0149612|T033|SY|165084003|SNOMEDCT_CORE|Exercise ECG positive|Exercise tolerance test abnormal
C0149612|T033|PT|165084003|SNOMEDCT_CORE|Exercise tolerance test abnormal|Exercise tolerance test abnormal
C0149612|T033|FN|165084003|SNOMEDCT_CORE|Exercise tolerance test abnormal|Exercise tolerance test abnormal
C0149612|T033|SY|165084003|SNOMEDCT_CORE|Positive exercise ECG test|Exercise tolerance test abnormal
C0149630|T019|PT|72352009|SNOMEDCT_CORE|Bicuspid aortic valve|Bicuspid aortic valve
C0149630|T019|FN|72352009|SNOMEDCT_CORE|Bicuspid aortic valve|Bicuspid aortic valve
C0149642|T047|SY|3502005|SNOMEDCT_CORE|Cervical adenitis|Cervical lymphadenitis
C0149642|T047|PT|3502005|SNOMEDCT_CORE|Cervical lymphadenitis|Cervical lymphadenitis
C0149642|T047|FN|3502005|SNOMEDCT_CORE|Cervical lymphadenitis|Cervical lymphadenitis
C0149645|T047|PT|202664003|SNOMEDCT_CORE|Cervical myelopathy|Cervical myelopathy
C0149645|T047|FN|202664003|SNOMEDCT_CORE|Cervical myelopathy|Cervical myelopathy
C0149653|T047|PT|398311004|SNOMEDCT_CORE|Diverticulosis of colon without diverticulitis|Diverticulosis of colon without diverticulitis
C0149653|T047|FN|398311004|SNOMEDCT_CORE|Diverticulosis of colon without diverticulitis|Diverticulosis of colon without diverticulitis
C0149653|T047|OF|398311004|SNOMEDCT_CORE|Diverticulosis of colon without diverticulitis|Diverticulosis of colon without diverticulitis
C0149671|T033|IS|58972000|SNOMEDCT_CORE|Dribbling|Dribbling of urine
C0149671|T033|PT|58972000|SNOMEDCT_CORE|Dribbling of urine|Dribbling of urine
C0149671|T033|FN|58972000|SNOMEDCT_CORE|Dribbling of urine|Dribbling of urine
C0149674|T037|SY|125596004|SNOMEDCT_CORE|Elbow injury|Injury of elbow
C0149674|T037|PT|125596004|SNOMEDCT_CORE|Injury of elbow|Injury of elbow
C0149674|T037|FN|125596004|SNOMEDCT_CORE|Injury of elbow|Injury of elbow
C0149678|T047|PT|240530001|SNOMEDCT_CORE|Epstein-Barr virus disease|Epstein-Barr virus disease
C0149678|T047|FN|240530001|SNOMEDCT_CORE|Epstein-Barr virus disease|Epstein-Barr virus disease
C0149678|T047|OAP|402121009|SNOMEDCT_CORE|Epstein-Barr virus infection|Epstein-Barr virus disease
C0149678|T047|OAF|402121009|SNOMEDCT_CORE|Epstein-Barr virus infection|Epstein-Barr virus disease
C0149696|T047|OF|235719002|SNOMEDCT_CORE|Food intolerance|Intolerance to food
C0149696|T047|SY|235719002|SNOMEDCT_CORE|Food intolerance|Intolerance to food
C0149696|T047|PT|235719002|SNOMEDCT_CORE|Intolerance to food|Intolerance to food
C0149696|T047|FN|235719002|SNOMEDCT_CORE|Intolerance to food|Intolerance to food
C0149696|T047|IS|235719002|SNOMEDCT_CORE|Malabsorption due to food intolerance|Intolerance to food
C0149697|T037|SY|125604000|SNOMEDCT_CORE|Foot injury|Injury of foot
C0149697|T037|PT|125604000|SNOMEDCT_CORE|Injury of foot|Injury of foot
C0149697|T037|FN|125604000|SNOMEDCT_CORE|Injury of foot|Injury of foot
C0149699|T037|PT|75591007|SNOMEDCT_CORE|Fracture of fibula|Fracture of fibula
C0149699|T037|FN|75591007|SNOMEDCT_CORE|Fracture of fibula|Fracture of fibula
C0149699|T037|IS|75591007|SNOMEDCT_CORE|Fracture of fibula, NOS|Fracture of fibula
C0149704|T047|PT|20607006|SNOMEDCT_CORE|Gingivostomatitis|Gingivostomatitis
C0149704|T047|FN|20607006|SNOMEDCT_CORE|Gingivostomatitis|Gingivostomatitis
C0149707|T033|SY|34615008|SNOMEDCT_CORE|Blood in semen|Hemospermia
C0149707|T033|PTGB|34615008|SNOMEDCT_CORE|Haemospermia|Hemospermia
C0149707|T033|IS|34615008|SNOMEDCT_CORE|Hematospermia|Hemospermia
C0149707|T033|PT|34615008|SNOMEDCT_CORE|Hemospermia|Hemospermia
C0149707|T033|FN|34615008|SNOMEDCT_CORE|Hemospermia|Hemospermia
C0149715|T048|SY|191956005|SNOMEDCT_CORE|HVS - Hyperventilation syndrome|Psychogenic hyperventilation
C0149715|T048|SY|191956005|SNOMEDCT_CORE|Hyperventilation syndrome|Psychogenic hyperventilation
C0149715|T048|IS|191956005|SNOMEDCT_CORE|Psychogenic hyperventilat|Psychogenic hyperventilation
C0149715|T048|PT|191956005|SNOMEDCT_CORE|Psychogenic hyperventilation|Psychogenic hyperventilation
C0149715|T048|FN|191956005|SNOMEDCT_CORE|Psychogenic hyperventilation|Psychogenic hyperventilation
C0149715|T048|SY|191956005|SNOMEDCT_CORE|Psychogenic overbreathing|Psychogenic hyperventilation
C0149721|T047|PT|55827005|SNOMEDCT_CORE|Left ventricular hypertrophy|Left ventricular hypertrophy
C0149721|T047|FN|55827005|SNOMEDCT_CORE|Left ventricular hypertrophy|Left ventricular hypertrophy
C0149721|T047|SY|55827005|SNOMEDCT_CORE|LV hypertrophy|Left ventricular hypertrophy
C0149721|T047|SY|55827005|SNOMEDCT_CORE|LV+ - Left ventricular hypertrophy|Left ventricular hypertrophy
C0149721|T047|SY|55827005|SNOMEDCT_CORE|LVH - Left ventricular hypertrophy|Left ventricular hypertrophy
C0149725|T047|SY|50417007|SNOMEDCT_CORE|Chest cold|Lower respiratory tract infection
C0149725|T047|IS|50417007|SNOMEDCT_CORE|Chest cold, NOS|Lower respiratory tract infection
C0149725|T047|SY|50417007|SNOMEDCT_CORE|Lower respiratory infection|Lower respiratory tract infection
C0149725|T047|IS|50417007|SNOMEDCT_CORE|Lower respiratory infection, NOS|Lower respiratory tract infection
C0149725|T047|PT|50417007|SNOMEDCT_CORE|Lower respiratory tract infection|Lower respiratory tract infection
C0149725|T047|FN|50417007|SNOMEDCT_CORE|Lower respiratory tract infection|Lower respiratory tract infection
C0149725|T047|IS|50417007|SNOMEDCT_CORE|Lower respiratory tract infection, NOS|Lower respiratory tract infection
C0149725|T047|SY|50417007|SNOMEDCT_CORE|LRTI - Lower respiratory tract infection|Lower respiratory tract infection
C0149726|T033|PT|309529002|SNOMEDCT_CORE|Lung mass|Lung mass
C0149726|T033|FN|309529002|SNOMEDCT_CORE|Lung mass|Lung mass
C0149732|T037|SY|262966007|SNOMEDCT_CORE|Muscle tear|Rupture of muscle
C0149732|T037|PT|262966007|SNOMEDCT_CORE|Rupture of muscle|Rupture of muscle
C0149732|T037|FN|262966007|SNOMEDCT_CORE|Rupture of muscle|Rupture of muscle
C0149732|T037|SY|262966007|SNOMEDCT_CORE|Torn muscle|Rupture of muscle
C0149736|T033|SY|299703001|SNOMEDCT_CORE|Lump on neck|Mass of neck
C0149736|T033|PT|299703001|SNOMEDCT_CORE|Mass of neck|Mass of neck
C0149736|T033|FN|299703001|SNOMEDCT_CORE|Mass of neck|Mass of neck
C0149741|T184|SY|54302000|SNOMEDCT_CORE|Breast discharge|Discharge from nipple
C0149741|T184|PT|54302000|SNOMEDCT_CORE|Discharge from nipple|Discharge from nipple
C0149741|T184|FN|54302000|SNOMEDCT_CORE|Discharge from nipple|Discharge from nipple
C0149741|T184|IS|54302000|SNOMEDCT_CORE|Nipple discharge|Discharge from nipple
C0149741|T184|SY|54302000|SNOMEDCT_CORE|Observation of nipple discharge|Discharge from nipple
C0149745|T047|SY|26284000|SNOMEDCT_CORE|Mouth ulcer|Ulcer of mouth
C0149745|T047|SY|26284000|SNOMEDCT_CORE|Mouth ulceration|Ulcer of mouth
C0149745|T047|SY|26284000|SNOMEDCT_CORE|Oral ulcer|Ulcer of mouth
C0149745|T047|PT|26284000|SNOMEDCT_CORE|Ulcer of mouth|Ulcer of mouth
C0149745|T047|FN|26284000|SNOMEDCT_CORE|Ulcer of mouth|Ulcer of mouth
C0149745|T047|SY|26284000|SNOMEDCT_CORE|Ulceration of oral mucosa|Ulcer of mouth
C0149751|T184|PT|300513000|SNOMEDCT_CORE|Lesion of penis|Lesion of penis
C0149751|T184|FN|300513000|SNOMEDCT_CORE|Lesion of penis|Lesion of penis
C0149751|T184|SY|300513000|SNOMEDCT_CORE|Lesion penis|Lesion of penis
C0149754|T047|PT|109245003|SNOMEDCT_CORE|Cellulitis of periorbital region|Cellulitis of periorbital region
C0149754|T047|FN|109245003|SNOMEDCT_CORE|Cellulitis of periorbital region|Cellulitis of periorbital region
C0149754|T047|SY|109245003|SNOMEDCT_CORE|Periorbital cellulitis|Cellulitis of periorbital region
C0149755|T037|PT|21351003|SNOMEDCT_CORE|Fracture of phalanx of foot|Fracture of phalanx of foot
C0149755|T037|FN|21351003|SNOMEDCT_CORE|Fracture of phalanx of foot|Fracture of phalanx of foot
C0149755|T037|IS|21351003|SNOMEDCT_CORE|Fracture of phalanx of foot, NOS|Fracture of phalanx of foot
C0149755|T037|SY|21351003|SNOMEDCT_CORE|Fracture of phalanx of toe|Fracture of phalanx of foot
C0149755|T037|SY|21351003|SNOMEDCT_CORE|Fracture of toe|Fracture of phalanx of foot
C0149755|T037|IS|21351003|SNOMEDCT_CORE|Fracture of toe, NOS|Fracture of phalanx of foot
C0149755|T037|SY|21351003|SNOMEDCT_CORE|Toe fracture|Fracture of phalanx of foot
C0149756|T047|PT|202882003|SNOMEDCT_CORE|Plantar fasciitis|Plantar fasciitis
C0149756|T047|FN|202882003|SNOMEDCT_CORE|Plantar fasciitis|Plantar fasciitis
C0149756|T047|SY|202882003|SNOMEDCT_CORE|Policeman's heel|Plantar fasciitis
C0149770|T046|PT|197166005|SNOMEDCT_CORE|Rectal abscess|Rectal abscess
C0149770|T046|FN|197166005|SNOMEDCT_CORE|Rectal abscess|Rectal abscess
C0149770|T046|SY|197166005|SNOMEDCT_CORE|Rectal boil|Rectal abscess
C0149771|T020|IS|62730001|SNOMEDCT_CORE|Proctocele|Rectocele
C0149771|T020|IS|62730001|SNOMEDCT_CORE|Proctocele, NOS|Rectocele
C0149771|T020|IS|62730001|SNOMEDCT_CORE|Rectocele|Rectocele
C0149771|T020|IS|62730001|SNOMEDCT_CORE|Rectocele, NOS|Rectocele
C0149771|T020|SY|62730001|SNOMEDCT_CORE|Rectovaginal hernia|Rectocele
C0149774|T033|SY|53929009|SNOMEDCT_CORE|Mass of scrotum|Scrotal mass
C0149774|T033|FN|53929009|SNOMEDCT_CORE|Mass of scrotum|Scrotal mass
C0149774|T033|PT|53929009|SNOMEDCT_CORE|Scrotal mass|Scrotal mass
C0149774|T033|OF|53929009|SNOMEDCT_CORE|Scrotal mass|Scrotal mass
C0149774|T033|IS|53929009|SNOMEDCT_CORE|Scrotal mass, NOS|Scrotal mass
C0149776|T037|PT|125594001|SNOMEDCT_CORE|Injury of shoulder region|Injury of shoulder region
C0149776|T037|FN|125594001|SNOMEDCT_CORE|Injury of shoulder region|Injury of shoulder region
C0149777|T046|IS|31928004|SNOMEDCT_CORE|Abscess of skin and subcutaneous tissue, NOS|Abscess of skin and/or subcutaneous tissue
C0149777|T046|OP|31928004|SNOMEDCT_CORE|Abscess of skin AND/OR subcutaneous tissue|Abscess of skin and/or subcutaneous tissue
C0149777|T046|PT|31928004|SNOMEDCT_CORE|Abscess of skin and/or subcutaneous tissue|Abscess of skin and/or subcutaneous tissue
C0149777|T046|FN|31928004|SNOMEDCT_CORE|Abscess of skin and/or subcutaneous tissue|Abscess of skin and/or subcutaneous tissue
C0149777|T046|OF|31928004|SNOMEDCT_CORE|Abscess of skin AND/OR subcutaneous tissue|Abscess of skin and/or subcutaneous tissue
C0149777|T046|SY|31928004|SNOMEDCT_CORE|Cutaneous abscess|Abscess of skin and/or subcutaneous tissue
C0149777|T046|SY|31928004|SNOMEDCT_CORE|Skin abscess|Abscess of skin and/or subcutaneous tissue
C0149778|T047|PT|95880003|SNOMEDCT_CORE|Soft tissue infection|Soft tissue infection
C0149778|T047|FN|95880003|SNOMEDCT_CORE|Soft tissue infection|Soft tissue infection
C0149778|T047|IS|95880003|SNOMEDCT_CORE|Soft tissue infection, NOS|Soft tissue infection
C0149781|T047|PT|80423007|SNOMEDCT_CORE|Spontaneous pneumothorax|Spontaneous pneumothorax
C0149781|T047|FN|80423007|SNOMEDCT_CORE|Spontaneous pneumothorax|Spontaneous pneumothorax
C0149782|T191|SY|254634000|SNOMEDCT_CORE|Epidermoid carcinoma of lung|Squamous cell carcinoma of lung
C0149782|T191|SY|254634000|SNOMEDCT_CORE|SCC - Squamous cell carcinoma of lung|Squamous cell carcinoma of lung
C0149782|T191|PT|254634000|SNOMEDCT_CORE|Squamous cell carcinoma of lung|Squamous cell carcinoma of lung
C0149782|T191|FN|254634000|SNOMEDCT_CORE|Squamous cell carcinoma of lung|Squamous cell carcinoma of lung
C0149793|T184|SY|88032003|SNOMEDCT_CORE|AF - Amaurosis fugax|Amaurosis fugax
C0149793|T184|SY|88032003|SNOMEDCT_CORE|AFx - Amaurosis fugax|Amaurosis fugax
C0149793|T184|PT|88032003|SNOMEDCT_CORE|Amaurosis fugax|Amaurosis fugax
C0149793|T184|FN|88032003|SNOMEDCT_CORE|Amaurosis fugax|Amaurosis fugax
C0149793|T184|SY|88032003|SNOMEDCT_CORE|Momentary blindness|Amaurosis fugax
C0149793|T184|SY|88032003|SNOMEDCT_CORE|Transient monocular blindness|Amaurosis fugax
C0149797|T047|PT|200724002|SNOMEDCT_CORE|Umbilical granuloma|Umbilical granuloma
C0149797|T047|FN|200724002|SNOMEDCT_CORE|Umbilical granuloma|Umbilical granuloma
C0149801|T047|OAP|371093006|SNOMEDCT_CORE|Sepsis due to urinary tract infection|Sepsis due to urinary tract infection
C0149801|T047|PT|721104000|SNOMEDCT_CORE|Sepsis due to urinary tract infection|Sepsis due to urinary tract infection
C0149801|T047|FN|721104000|SNOMEDCT_CORE|Sepsis due to urinary tract infection|Sepsis due to urinary tract infection
C0149801|T047|OAS|371093006|SNOMEDCT_CORE|Urinary sepsis|Sepsis due to urinary tract infection
C0149801|T047|OAS|371093006|SNOMEDCT_CORE|Urosepsis|Sepsis due to urinary tract infection
C0149801|T047|OAF|371093006|SNOMEDCT_CORE|Urosepsis|Sepsis due to urinary tract infection
C0149804|T037|PT|34124000|SNOMEDCT_CORE|Foreign body in vagina|Foreign body in vagina
C0149804|T037|FN|34124000|SNOMEDCT_CORE|Foreign body in vagina|Foreign body in vagina
C0149816|T047|PT|36046008|SNOMEDCT_CORE|Ischiorectal abscess|Ischiorectal abscess
C0149816|T047|FN|36046008|SNOMEDCT_CORE|Ischiorectal abscess|Ischiorectal abscess
C0149825|T047|SY|111591002|SNOMEDCT_CORE|Adenoidal enlargement|Hypertrophy of adenoids
C0149825|T047|SY|111591002|SNOMEDCT_CORE|Adenoidal hypertrophy|Hypertrophy of adenoids
C0149825|T047|SY|111591002|SNOMEDCT_CORE|Enlargement of adenoids|Hypertrophy of adenoids
C0149825|T047|PT|111591002|SNOMEDCT_CORE|Hypertrophy of adenoids|Hypertrophy of adenoids
C0149825|T047|FN|111591002|SNOMEDCT_CORE|Hypertrophy of adenoids|Hypertrophy of adenoids
C0149836|T047|PT|75993002|SNOMEDCT_CORE|Atrophic vulvovaginitis|Atrophic vulvovaginitis
C0149836|T047|FN|75993002|SNOMEDCT_CORE|Atrophic vulvovaginitis|Atrophic vulvovaginitis
C0149836|T047|SY|75993002|SNOMEDCT_CORE|Senile vulvovaginitis|Atrophic vulvovaginitis
C0149842|T047|SY|231797007|SNOMEDCT_CORE|Blepharitis in seborrheic eczema|Seborrheic blepharitis
C0149842|T047|SYGB|231797007|SNOMEDCT_CORE|Blepharitis in seborrhoeic eczema|Seborrheic blepharitis
C0149842|T047|PT|231797007|SNOMEDCT_CORE|Seborrheic blepharitis|Seborrheic blepharitis
C0149842|T047|FN|231797007|SNOMEDCT_CORE|Seborrheic blepharitis|Seborrheic blepharitis
C0149842|T047|PTGB|231797007|SNOMEDCT_CORE|Seborrhoeic blepharitis|Seborrheic blepharitis
C0149846|T047|PT|221695002|SNOMEDCT_CORE|Achilles bursitis|Achilles bursitis
C0149846|T047|OF|221695002|SNOMEDCT_CORE|Achilles bursitis|Achilles bursitis
C0149846|T047|SY|221695002|SNOMEDCT_CORE|Achillobursitis|Achilles bursitis
C0149846|T047|SY|221695002|SNOMEDCT_CORE|Albert's syndrome|Achilles bursitis
C0149846|T047|SY|221695002|SNOMEDCT_CORE|Bursitis of calcaneal tendon bursa|Achilles bursitis
C0149846|T047|FN|221695002|SNOMEDCT_CORE|Bursitis of calcaneal tendon bursa|Achilles bursitis
C0149846|T047|SY|221695002|SNOMEDCT_CORE|Capped hock|Achilles bursitis
C0149846|T047|IS|221695002|SNOMEDCT_CORE|Haglund's deformity|Achilles bursitis
C0149846|T047|IS|221695002|SNOMEDCT_CORE|Haglund's disease|Achilles bursitis
C0149846|T047|SY|221695002|SNOMEDCT_CORE|Swediaur's disease|Achilles bursitis
C0149848|T047|SY|399114005|SNOMEDCT_CORE|Duplay's periarthritis syndrome|Subdeltoid bursitis
C0149848|T047|PT|78715003|SNOMEDCT_CORE|Subdeltoid bursitis|Subdeltoid bursitis
C0149848|T047|IS|27741009|SNOMEDCT_CORE|Subdeltoid bursitis|Subdeltoid bursitis
C0149848|T047|FN|78715003|SNOMEDCT_CORE|Subdeltoid bursitis|Subdeltoid bursitis
C0149862|T191|PT|309084001|SNOMEDCT_CORE|Villous adenoma of colon|Villous adenoma of colon
C0149862|T191|FN|309084001|SNOMEDCT_CORE|Villous adenoma of colon|Villous adenoma of colon
C0149863|T046|PT|197060001|SNOMEDCT_CORE|Sigmoid volvulus|Sigmoid volvulus
C0149863|T046|FN|197060001|SNOMEDCT_CORE|Sigmoid volvulus|Sigmoid volvulus
C0149863|T046|SY|197060001|SNOMEDCT_CORE|Volvulus of sigmoid colon|Sigmoid volvulus
C0149870|T047|SY|21794005|SNOMEDCT_CORE|de Quervain's disease|Radial styloid tenosynovitis
C0149870|T047|PT|21794005|SNOMEDCT_CORE|Radial styloid tenosynovitis|Radial styloid tenosynovitis
C0149870|T047|FN|21794005|SNOMEDCT_CORE|Radial styloid tenosynovitis|Radial styloid tenosynovitis
C0149871|T047|SY|128053003|SNOMEDCT_CORE|Deep vein thrombosis|Deep venous thrombosis
C0149871|T047|PT|128053003|SNOMEDCT_CORE|Deep venous thrombosis|Deep venous thrombosis
C0149871|T047|FN|128053003|SNOMEDCT_CORE|Deep venous thrombosis|Deep venous thrombosis
C0149871|T047|IS|128053003|SNOMEDCT_CORE|DVT|Deep venous thrombosis
C0149871|T047|SY|128053003|SNOMEDCT_CORE|DVT - Deep vein thrombosis|Deep venous thrombosis
C0149880|T047|PT|43491000|SNOMEDCT_CORE|Acute epididymitis|Acute epididymitis
C0149880|T047|FN|43491000|SNOMEDCT_CORE|Acute epididymitis|Acute epididymitis
C0149881|T047|SY|197983000|SNOMEDCT_CORE|Epididymo-orchitis|Orchitis and epididymitis
C0149881|T047|SY|197983000|SNOMEDCT_CORE|Inflammation of testis and epididymis|Orchitis and epididymitis
C0149881|T047|PT|197983000|SNOMEDCT_CORE|Orchitis and epididymitis|Orchitis and epididymitis
C0149881|T047|FN|197983000|SNOMEDCT_CORE|Orchitis and epididymitis|Orchitis and epididymitis
C0149882|T047|PT|409656006|SNOMEDCT_CORE|Acute esophagitis|Acute esophagitis
C0149882|T047|FN|409656006|SNOMEDCT_CORE|Acute esophagitis|Acute esophagitis
C0149882|T047|PTGB|409656006|SNOMEDCT_CORE|Acute oesophagitis|Acute esophagitis
C0149889|T046|PT|72779005|SNOMEDCT_CORE|Anorectal fistula|Anorectal fistula
C0149889|T046|FN|72779005|SNOMEDCT_CORE|Anorectal fistula|Anorectal fistula
C0149893|T047|SY|95717004|SNOMEDCT_CORE|Glaucoma due to ocular disease|Secondary glaucoma
C0149893|T047|PT|95717004|SNOMEDCT_CORE|Secondary glaucoma|Secondary glaucoma
C0149893|T047|FN|95717004|SNOMEDCT_CORE|Secondary glaucoma|Secondary glaucoma
C0149893|T047|IS|95717004|SNOMEDCT_CORE|Secondary glaucoma, NOS|Secondary glaucoma
C0149896|T047|IS|24595009|SNOMEDCT_CORE|Acute gouty arthritis|Primary gout
C0149896|T047|IS|24595009|SNOMEDCT_CORE|Acute gouty arthropathy|Primary gout
C0149896|T047|SY|24595009|SNOMEDCT_CORE|Idiopathic gout|Primary gout
C0149896|T047|PT|24595009|SNOMEDCT_CORE|Primary gout|Primary gout
C0149896|T047|FN|24595009|SNOMEDCT_CORE|Primary gout|Primary gout
C0149908|T047|PT|301864002|SNOMEDCT_CORE|Transient synovitis of hip|Transient synovitis of hip
C0149908|T047|FN|301864002|SNOMEDCT_CORE|Transient synovitis of hip|Transient synovitis of hip
C0149922|T047|SY|53891004|SNOMEDCT_CORE|Circumscribed neurodermatitis|Lichen simplex chronicus
C0149922|T047|SY|53891004|SNOMEDCT_CORE|Lichen simplex|Lichen simplex chronicus
C0149922|T047|PT|53891004|SNOMEDCT_CORE|Lichen simplex chronicus|Lichen simplex chronicus
C0149922|T047|FN|53891004|SNOMEDCT_CORE|Lichen simplex chronicus|Lichen simplex chronicus
C0149922|T047|IS|53891004|SNOMEDCT_CORE|Lichenified eczema|Lichen simplex chronicus
C0149922|T047|SY|53891004|SNOMEDCT_CORE|Lichenoid dermatitis|Lichen simplex chronicus
C0149922|T047|SY|53891004|SNOMEDCT_CORE|Local neurodermatitis|Lichen simplex chronicus
C0149922|T047|SY|53891004|SNOMEDCT_CORE|LSC - Lichen simplex chronicus|Lichen simplex chronicus
C0149922|T047|SY|53891004|SNOMEDCT_CORE|Neurodermatitis circumscripta|Lichen simplex chronicus
C0149925|T191|SY|254632001|SNOMEDCT_CORE|SCLC - Small cell lung cancer|Small cell carcinoma of lung
C0149925|T191|PT|254632001|SNOMEDCT_CORE|Small cell carcinoma of lung|Small cell carcinoma of lung
C0149925|T191|FN|254632001|SNOMEDCT_CORE|Small cell carcinoma of lung|Small cell carcinoma of lung
C0149925|T191|SY|254632001|SNOMEDCT_CORE|Small cell lung cancer|Small cell carcinoma of lung
C0149931|T047|FN|37796009|SNOMEDCT_CORE|Migraine|Migraine
C0149931|T047|PT|37796009|SNOMEDCT_CORE|Migraine|Migraine
C0149931|T047|IS|37796009|SNOMEDCT_CORE|Migraine, NOS|Migraine
C0149940|T047|PT|52585001|SNOMEDCT_CORE|Sciatic neuropathy|Sciatic neuropathy
C0149940|T047|FN|52585001|SNOMEDCT_CORE|Sciatic neuropathy|Sciatic neuropathy
C0149944|T037|PT|207787008|SNOMEDCT_CORE|Fracture of orbital floor|Fracture of orbital floor
C0149944|T037|FN|207787008|SNOMEDCT_CORE|Fracture of orbital floor|Fracture of orbital floor
C0149944|T037|SY|207787008|SNOMEDCT_CORE|Orbital floor fracture|Fracture of orbital floor
C0149948|T047|PT|30250000|SNOMEDCT_CORE|Acute otitis externa|Acute otitis externa
C0149948|T047|FN|30250000|SNOMEDCT_CORE|Acute otitis externa|Acute otitis externa
C0149948|T047|IS|30250000|SNOMEDCT_CORE|Acute otitis externa, NOS|Acute otitis externa
C0149952|T190|SY|13595002|SNOMEDCT_CORE|Ovarian torsion|Torsion of ovary
C0149952|T190|PT|13595002|SNOMEDCT_CORE|Torsion of ovary|Torsion of ovary
C0149952|T190|FN|13595002|SNOMEDCT_CORE|Torsion of ovary|Torsion of ovary
C0149958|T047|SY|4103001|SNOMEDCT_CORE|Complex partial seizure|Psychomotor fit
C0149958|T047|SY|4103001|SNOMEDCT_CORE|Psychomotor fit|Psychomotor fit
C0149959|T047|PT|237037006|SNOMEDCT_CORE|Acute pelvic inflammatory disease|Acute pelvic inflammatory disease
C0149959|T047|FN|237037006|SNOMEDCT_CORE|Acute pelvic inflammatory disease|Acute pelvic inflammatory disease
C0149959|T047|IS|237037006|SNOMEDCT_CORE|Acute PID|Acute pelvic inflammatory disease
C0149959|T047|SY|237037006|SNOMEDCT_CORE|Acute PID - acute pelvic inflammatory disease|Acute pelvic inflammatory disease
C0149959|T047|SY|237037006|SNOMEDCT_CORE|PID - Acute pelvic inflammatory disease|Acute pelvic inflammatory disease
C0149960|T047|PT|237044002|SNOMEDCT_CORE|Chronic pelvic inflammatory disease|Chronic pelvic inflammatory disease
C0149960|T047|FN|237044002|SNOMEDCT_CORE|Chronic pelvic inflammatory disease|Chronic pelvic inflammatory disease
C0149960|T047|IS|237044002|SNOMEDCT_CORE|Chronic pelvic inflammatory disease of the female pelvic organs AND/OR tissues|Chronic pelvic inflammatory disease
C0149960|T047|IS|237044002|SNOMEDCT_CORE|Chronic PID|Chronic pelvic inflammatory disease
C0149960|T047|SY|237044002|SNOMEDCT_CORE|Chronic PID - Chronic pelvic inflammatory disease|Chronic pelvic inflammatory disease
C0149977|T037|OAS|95854004|SNOMEDCT_CORE|Goyrand's injury|Subluxation of radial head
C0149977|T037|SY|417109008|SNOMEDCT_CORE|Goyrand's injury|Subluxation of radial head
C0149977|T037|OAS|95854004|SNOMEDCT_CORE|Malgaigne's luxation|Subluxation of radial head
C0149977|T037|OAS|95854004|SNOMEDCT_CORE|Nursemaids' elbow|Subluxation of radial head
C0149977|T037|SY|417109008|SNOMEDCT_CORE|Nursemaids' elbow|Subluxation of radial head
C0149977|T037|OAP|95854004|SNOMEDCT_CORE|Pulled elbow|Subluxation of radial head
C0149977|T037|SY|417109008|SNOMEDCT_CORE|Pulled elbow|Subluxation of radial head
C0149977|T037|OAF|95854004|SNOMEDCT_CORE|Pulled elbow|Subluxation of radial head
C0149977|T037|PT|417109008|SNOMEDCT_CORE|Subluxation of radial head|Subluxation of radial head
C0149977|T037|FN|417109008|SNOMEDCT_CORE|Subluxation of radial head|Subluxation of radial head
C0149978|T191|PT|254582000|SNOMEDCT_CORE|Adenocarcinoma of rectum|Adenocarcinoma of rectum
C0149978|T191|FN|254582000|SNOMEDCT_CORE|Adenocarcinoma of rectum|Adenocarcinoma of rectum
C0149980|T047|PT|95239003|SNOMEDCT_CORE|Rhinitis medicamentosa|Rhinitis medicamentosa
C0149980|T047|FN|95239003|SNOMEDCT_CORE|Rhinitis medicamentosa|Rhinitis medicamentosa
C0149983|T047|PT|239880009|SNOMEDCT_CORE|Lumbar spondylosis|Lumbar spondylosis
C0149983|T047|FN|239880009|SNOMEDCT_CORE|Lumbar spondylosis|Lumbar spondylosis
C0149987|T047|PT|442048005|SNOMEDCT_CORE|Tenosynovitis of wrist|Tenosynovitis of wrist
C0149987|T047|FN|442048005|SNOMEDCT_CORE|Tenosynovitis of wrist|Tenosynovitis of wrist
C0150037|T033|PT|129823000|SNOMEDCT_CORE|Childhood growth AND/OR development alteration|Childhood growth AND/OR development alteration
C0150037|T033|FN|129823000|SNOMEDCT_CORE|Childhood growth AND/OR development alteration|Childhood growth AND/OR development alteration
C0150037|T033|IS|129823000|SNOMEDCT_CORE|Growth and development alteration|Childhood growth AND/OR development alteration
C0150037|T033|IS|129823000|SNOMEDCT_CORE|Growth and devlopment alteration|Childhood growth AND/OR development alteration
C0150044|T033|PT|129853007|SNOMEDCT_CORE|Total urinary incontinence|Total urinary incontinence
C0150044|T033|FN|129853007|SNOMEDCT_CORE|Total urinary incontinence|Total urinary incontinence
C0150044|T033|SY|129853007|SNOMEDCT_CORE|Urinary incontinence with continuous leakage|Total urinary incontinence
C0150045|T033|SY|87557004|SNOMEDCT_CORE|Lack of bladder control if desire resisted|Urge incontinence of urine
C0150045|T033|SY|87557004|SNOMEDCT_CORE|Lack of bladder control if desire urgent|Urge incontinence of urine
C0150045|T033|SY|87557004|SNOMEDCT_CORE|Must urinate at once with urge|Urge incontinence of urine
C0150045|T033|IS|87557004|SNOMEDCT_CORE|Urge incontinence|Urge incontinence of urine
C0150045|T033|PT|87557004|SNOMEDCT_CORE|Urge incontinence of urine|Urge incontinence of urine
C0150045|T033|FN|87557004|SNOMEDCT_CORE|Urge incontinence of urine|Urge incontinence of urine
C0150045|T033|SY|87557004|SNOMEDCT_CORE|Urge urinary incontinence|Urge incontinence of urine
C0150055|T184|PT|82423001|SNOMEDCT_CORE|Chronic pain|Chronic pain
C0150055|T184|FN|82423001|SNOMEDCT_CORE|Chronic pain|Chronic pain
C0150077|T033|PT|247442005|SNOMEDCT_CORE|Broken skin|Broken skin
C0150077|T033|FN|247442005|SNOMEDCT_CORE|Broken skin|Broken skin
C0150077|T033|SY|247442005|SNOMEDCT_CORE|Defect in skin surface|Broken skin
C0150077|T033|SY|247442005|SNOMEDCT_CORE|Skin breakdown|Broken skin
C0150618|T033|PT|63332003|SNOMEDCT_CORE|History AND physical examination|History AND physical examination
C0150618|T033|FN|63332003|SNOMEDCT_CORE|History AND physical examination|History AND physical examination
C0150618|T033|IS|63332003|SNOMEDCT_CORE|History and physical examination, NOS|History AND physical examination
C0151205|T046|SY|49563000|SNOMEDCT_CORE|Edema around eye|Periorbital edema
C0151205|T046|SYGB|49563000|SNOMEDCT_CORE|Oedema around eye|Periorbital edema
C0151205|T046|PT|49563000|SNOMEDCT_CORE|Periorbital edema|Periorbital edema
C0151205|T046|FN|49563000|SNOMEDCT_CORE|Periorbital edema|Periorbital edema
C0151205|T046|PTGB|49563000|SNOMEDCT_CORE|Periorbital oedema|Periorbital edema
C0151217|T047|PT|53295002|SNOMEDCT_CORE|Chronic otitis externa|Chronic otitis externa
C0151217|T047|FN|53295002|SNOMEDCT_CORE|Chronic otitis externa|Chronic otitis externa
C0151217|T047|IS|53295002|SNOMEDCT_CORE|Chronic otitis externa, NOS|Chronic otitis externa
C0151295|T047|PT|30292005|SNOMEDCT_CORE|Mononeuritis multiplex|Mononeuritis multiplex
C0151295|T047|FN|30292005|SNOMEDCT_CORE|Mononeuritis multiplex|Mononeuritis multiplex
C0151313|T047|PT|95662005|SNOMEDCT_CORE|Sensory neuropathy|Sensory neuropathy
C0151313|T047|FN|95662005|SNOMEDCT_CORE|Sensory neuropathy|Sensory neuropathy
C0151313|T047|IS|95662005|SNOMEDCT_CORE|Sensory peripheral neuropathy|Sensory neuropathy
C0151315|T184|SY|161882006|SNOMEDCT_CORE|Neck stiffness|Stiff neck
C0151315|T184|SY|161882006|SNOMEDCT_CORE|NS - Neck stiffness|Stiff neck
C0151315|T184|PT|161882006|SNOMEDCT_CORE|Stiff neck|Stiff neck
C0151315|T184|FN|161882006|SNOMEDCT_CORE|Stiff neck|Stiff neck
C0151332|T047|PT|427099000|SNOMEDCT_CORE|Active tuberculosis|Active tuberculosis
C0151332|T047|FN|427099000|SNOMEDCT_CORE|Active tuberculosis|Active tuberculosis
C0151434|T047|PT|202856007|SNOMEDCT_CORE|Biceps tendinitis|Biceps tendinitis
C0151434|T047|FN|202856007|SNOMEDCT_CORE|Biceps tendinitis|Biceps tendinitis
C0151434|T047|SY|202856007|SNOMEDCT_CORE|Bicipital tendinitis|Biceps tendinitis
C0151448|T047|PT|442520000|SNOMEDCT_CORE|Inflammation of rotator cuff tendon|Inflammation of rotator cuff tendon
C0151448|T047|FN|442520000|SNOMEDCT_CORE|Inflammation of rotator cuff tendon|Inflammation of rotator cuff tendon
C0151448|T047|IS|442520000|SNOMEDCT_CORE|Tendinitis of rotator cuff|Inflammation of rotator cuff tendon
C0151451|T047|SY|7674000|SNOMEDCT_CORE|GTPS - greater trochanteric pain syndrome|Trochanteric bursitis
C0151451|T047|PT|7674000|SNOMEDCT_CORE|Trochanteric bursitis|Trochanteric bursitis
C0151451|T047|FN|7674000|SNOMEDCT_CORE|Trochanteric bursitis|Trochanteric bursitis
C0151451|T047|IS|7674000|SNOMEDCT_CORE|Whirlbone lameness|Trochanteric bursitis
C0151463|T047|PT|28432003|SNOMEDCT_CORE|Abscess of breast|Abscess of breast
C0151463|T047|FN|28432003|SNOMEDCT_CORE|Abscess of breast|Abscess of breast
C0151463|T047|IS|28432003|SNOMEDCT_CORE|Abscess of breast, NOS|Abscess of breast
C0151467|T047|IS|24867002|SNOMEDCT_CORE|Acute adrenal insufficiency|Severe adrenal insufficiency
C0151467|T047|IS|24867002|SNOMEDCT_CORE|Addisonian crisis|Severe adrenal insufficiency
C0151467|T047|IS|24867002|SNOMEDCT_CORE|Adrenal crisis|Severe adrenal insufficiency
C0151467|T047|IS|24867002|SNOMEDCT_CORE|Adrenocortical crisis|Severe adrenal insufficiency
C0151467|T047|PT|24867002|SNOMEDCT_CORE|Severe adrenal insufficiency|Severe adrenal insufficiency
C0151467|T047|FN|24867002|SNOMEDCT_CORE|Severe adrenal insufficiency|Severe adrenal insufficiency
C0151468|T191|PT|255034006|SNOMEDCT_CORE|Thyroid follicular adenoma|Thyroid follicular adenoma
C0151468|T191|FN|255034006|SNOMEDCT_CORE|Thyroid follicular adenoma|Thyroid follicular adenoma
C0151482|T047|SYGB|85649008|SNOMEDCT_CORE|Folate deficiency anaemia|Megaloblastic anemia due to folate deficiency
C0151482|T047|SY|85649008|SNOMEDCT_CORE|Folate deficiency anemia|Megaloblastic anemia due to folate deficiency
C0151482|T047|SYGB|85649008|SNOMEDCT_CORE|Folic acid deficiency anaemia|Megaloblastic anemia due to folate deficiency
C0151482|T047|SY|85649008|SNOMEDCT_CORE|Folic acid deficiency anemia|Megaloblastic anemia due to folate deficiency
C0151482|T047|PTGB|85649008|SNOMEDCT_CORE|Megaloblastic anaemia due to folate deficiency|Megaloblastic anemia due to folate deficiency
C0151482|T047|PT|85649008|SNOMEDCT_CORE|Megaloblastic anemia due to folate deficiency|Megaloblastic anemia due to folate deficiency
C0151482|T047|FN|85649008|SNOMEDCT_CORE|Megaloblastic anemia due to folate deficiency|Megaloblastic anemia due to folate deficiency
C0151482|T047|IS|85649008|SNOMEDCT_CORE|Megaloblastic anemia due to folate deficiency, NOS|Megaloblastic anemia due to folate deficiency
C0151517|T047|SY|27885002|SNOMEDCT_CORE|CHB - Complete heart block|Complete atrioventricular block
C0151517|T047|FN|27885002|SNOMEDCT_CORE|Complete atrioventricular block|Complete atrioventricular block
C0151517|T047|PT|27885002|SNOMEDCT_CORE|Complete atrioventricular block|Complete atrioventricular block
C0151517|T047|SY|27885002|SNOMEDCT_CORE|Complete heart block|Complete atrioventricular block
C0151517|T047|SY|27885002|SNOMEDCT_CORE|High grade atrioventricular block|Complete atrioventricular block
C0151517|T047|SY|27885002|SNOMEDCT_CORE|Third degree atrioventricular block|Complete atrioventricular block
C0151517|T047|SY|27885002|SNOMEDCT_CORE|Third degree heart block|Complete atrioventricular block
C0151526|T046|PT|282020008|SNOMEDCT_CORE|Premature delivery|Premature delivery
C0151526|T046|FN|282020008|SNOMEDCT_CORE|Premature delivery|Premature delivery
C0151594|T047|SY|95545007|SNOMEDCT_CORE|Bloody diarrhea|Hemorrhagic diarrhea
C0151594|T047|SYGB|95545007|SNOMEDCT_CORE|Bloody diarrhoea|Hemorrhagic diarrhea
C0151594|T047|PTGB|95545007|SNOMEDCT_CORE|Haemorrhagic diarrhoea|Hemorrhagic diarrhea
C0151594|T047|PT|95545007|SNOMEDCT_CORE|Hemorrhagic diarrhea|Hemorrhagic diarrhea
C0151594|T047|FN|95545007|SNOMEDCT_CORE|Hemorrhagic diarrhea|Hemorrhagic diarrhea
C0151602|T033|FN|278528006|SNOMEDCT_CORE|Facial swelling|Facial swelling
C0151602|T033|PT|278528006|SNOMEDCT_CORE|Facial swelling|Facial swelling
C0151602|T033|SY|278528006|SNOMEDCT_CORE|Swollen face|Facial swelling
C0151611|T033|SY|274521009|SNOMEDCT_CORE|EEG abnormal|Electroencephalogram abnormal
C0151611|T033|PT|274521009|SNOMEDCT_CORE|Electroencephalogram abnormal|Electroencephalogram abnormal
C0151611|T033|FN|274521009|SNOMEDCT_CORE|Electroencephalogram abnormal|Electroencephalogram abnormal
C0151632|T033|OAP|416103000|SNOMEDCT_CORE|Elevated erythrocyte sedimentation rate|ESR raised
C0151632|T033|OAF|416103000|SNOMEDCT_CORE|Elevated erythrocyte sedimentation rate|ESR raised
C0151632|T033|SY|165468009|SNOMEDCT_CORE|Erythrocyte sedimentation rate raised|ESR raised
C0151632|T033|FN|165468009|SNOMEDCT_CORE|Erythrocyte sedimentation rate raised|ESR raised
C0151632|T033|OF|165468009|SNOMEDCT_CORE|Erythrocyte sedimentation rate raised|ESR raised
C0151632|T033|PT|165468009|SNOMEDCT_CORE|ESR raised|ESR raised
C0151632|T033|OF|165468009|SNOMEDCT_CORE|ESR raised|ESR raised
C0151636|T047|SY|251175005|SNOMEDCT_CORE|Premature ventricular complex|Ventricular premature complex
C0151636|T047|SY|251175005|SNOMEDCT_CORE|Ventricular ectopic complex|Ventricular premature complex
C0151636|T047|PT|251175005|SNOMEDCT_CORE|Ventricular premature complex|Ventricular premature complex
C0151636|T047|FN|251175005|SNOMEDCT_CORE|Ventricular premature complex|Ventricular premature complex
C0151636|T047|SYGB|251175005|SNOMEDCT_CORE|Ventricular premature depolarisation|Ventricular premature complex
C0151636|T047|SY|251175005|SNOMEDCT_CORE|Ventricular premature depolarization|Ventricular premature complex
C0151694|T046|SYGB|95540002|SNOMEDCT_CORE|Colonic haemorrhage|Hemorrhage of colon
C0151694|T046|SY|95540002|SNOMEDCT_CORE|Colonic hemorrhage|Hemorrhage of colon
C0151694|T046|PTGB|95540002|SNOMEDCT_CORE|Haemorrhage of colon|Hemorrhage of colon
C0151694|T046|PT|95540002|SNOMEDCT_CORE|Hemorrhage of colon|Hemorrhage of colon
C0151694|T046|FN|95540002|SNOMEDCT_CORE|Hemorrhage of colon|Hemorrhage of colon
C0151699|T046|PTGB|1386000|SNOMEDCT_CORE|Intracranial haemorrhage|Intracranial hemorrhage
C0151699|T046|PT|1386000|SNOMEDCT_CORE|Intracranial hemorrhage|Intracranial hemorrhage
C0151699|T046|FN|1386000|SNOMEDCT_CORE|Intracranial hemorrhage|Intracranial hemorrhage
C0151699|T046|IS|1386000|SNOMEDCT_CORE|Intracranial hemorrhage, NOS|Intracranial hemorrhage
C0151721|T047|SY|48723006|SNOMEDCT_CORE|Eunuchoidism|Male hypogonadism
C0151721|T047|SY|48723006|SNOMEDCT_CORE|Eunuchoidism hypogonadism|Male hypogonadism
C0151721|T047|SY|48723006|SNOMEDCT_CORE|Eunuchoidism, hypogonadism|Male hypogonadism
C0151721|T047|PT|48723006|SNOMEDCT_CORE|Male hypogonadism|Male hypogonadism
C0151721|T047|FN|48723006|SNOMEDCT_CORE|Male hypogonadism|Male hypogonadism
C0151721|T047|IS|48723006|SNOMEDCT_CORE|Male hypogonadism, NOS|Male hypogonadism
C0151721|T047|SY|48723006|SNOMEDCT_CORE|Testicular failure|Male hypogonadism
C0151721|T047|SY|48723006|SNOMEDCT_CORE|Testicular hypogonadism|Male hypogonadism
C0151723|T047|PTGB|190855004|SNOMEDCT_CORE|Hypomagnesaemia|Hypomagnesemia
C0151723|T047|PT|190855004|SNOMEDCT_CORE|Hypomagnesemia|Hypomagnesemia
C0151723|T047|FN|190855004|SNOMEDCT_CORE|Hypomagnesemia|Hypomagnesemia
C0151723|T047|IS|190855004|SNOMEDCT_CORE|Magnesium deficiency syndrome|Hypomagnesemia
C0151739|T046|PT|235741002|SNOMEDCT_CORE|Perforation of small intestine|Perforation of small intestine
C0151739|T046|FN|235741002|SNOMEDCT_CORE|Perforation of small intestine|Perforation of small intestine
C0151739|T046|SY|235741002|SNOMEDCT_CORE|Small bowel perforation|Perforation of small intestine
C0151744|T047|SY|414795007|SNOMEDCT_CORE|Cardiac ischemia|Myocardial ischemia
C0151744|T047|PTGB|414795007|SNOMEDCT_CORE|Myocardial ischaemia|Myocardial ischemia
C0151744|T047|PT|414795007|SNOMEDCT_CORE|Myocardial ischemia|Myocardial ischemia
C0151744|T047|FN|414795007|SNOMEDCT_CORE|Myocardial ischemia|Myocardial ischemia
C0151746|T046|PT|39539005|SNOMEDCT_CORE|Abnormal renal function|Abnormal renal function
C0151746|T046|FN|39539005|SNOMEDCT_CORE|Abnormal renal function|Abnormal renal function
C0151766|T033|SY|166603001|SNOMEDCT_CORE|Abnormal results of liver function studies|Liver function tests abnormal
C0151766|T033|FN|166603001|SNOMEDCT_CORE|Liver function tests abnormal|Liver function tests abnormal
C0151766|T033|PT|166603001|SNOMEDCT_CORE|Liver function tests abnormal|Liver function tests abnormal
C0151772|T048|SY|231494001|SNOMEDCT_CORE|Manic psychosis|Manic psychosis
C0151779|T191|SY|93655004|SNOMEDCT_CORE|Cutaneous malignant melanoma|Malignant melanoma of skin
C0151779|T191|PT|93655004|SNOMEDCT_CORE|Malignant melanoma of skin|Malignant melanoma of skin
C0151779|T191|FN|93655004|SNOMEDCT_CORE|Malignant melanoma of skin|Malignant melanoma of skin
C0151779|T191|IS|93655004|SNOMEDCT_CORE|Malignant melanoma of skin, NOS|Malignant melanoma of skin
C0151779|T191|SY|93655004|SNOMEDCT_CORE|Melanoma of skin|Malignant melanoma of skin
C0151779|T191|SY|93655004|SNOMEDCT_CORE|MM - Malignant melanoma of skin|Malignant melanoma of skin
C0151786|T184|SY|26544005|SNOMEDCT_CORE|Decreased muscle strength|Muscle weakness
C0151786|T184|SY|26544005|SNOMEDCT_CORE|Muscle strength reduced|Muscle weakness
C0151786|T184|PT|26544005|SNOMEDCT_CORE|Muscle weakness|Muscle weakness
C0151786|T184|FN|26544005|SNOMEDCT_CORE|Muscle weakness|Muscle weakness
C0151799|T046|SY|95347000|SNOMEDCT_CORE|Cutaneous necrosis|Skin necrosis
C0151799|T046|IS|95347000|SNOMEDCT_CORE|Necrosis of skin|Skin necrosis
C0151799|T046|PT|95347000|SNOMEDCT_CORE|Skin necrosis|Skin necrosis
C0151799|T046|FN|95347000|SNOMEDCT_CORE|Skin necrosis|Skin necrosis
C0151799|T046|SY|95347000|SNOMEDCT_CORE|Sloughing of skin|Skin necrosis
C0151811|T046|SY|95325000|SNOMEDCT_CORE|Nodule of subcutaneous tissue|Subcutaneous nodule
C0151811|T046|IS|95325000|SNOMEDCT_CORE|Nodule of subcutaneous tissue, NOS|Subcutaneous nodule
C0151811|T046|PT|95325000|SNOMEDCT_CORE|Subcutaneous nodule|Subcutaneous nodule
C0151811|T046|OF|95325000|SNOMEDCT_CORE|Subcutaneous nodule|Subcutaneous nodule
C0151811|T046|FN|95325000|SNOMEDCT_CORE|Subcutaneous nodule|Subcutaneous nodule
C0151811|T046|IS|95325000|SNOMEDCT_CORE|Subcutaneous nodule, NOS|Subcutaneous nodule
C0151824|T047|PT|37389005|SNOMEDCT_CORE|Biliary colic|Biliary colic
C0151824|T047|OF|37389005|SNOMEDCT_CORE|Biliary colic|Biliary colic
C0151824|T047|FN|37389005|SNOMEDCT_CORE|Biliary colic|Biliary colic
C0151824|T047|SY|37389005|SNOMEDCT_CORE|Biliary colic symptom|Biliary colic
C0151824|T047|SY|37389005|SNOMEDCT_CORE|Hepatic colic|Biliary colic
C0151825|T184|PT|12584003|SNOMEDCT_CORE|Bone pain|Bone pain
C0151825|T184|FN|12584003|SNOMEDCT_CORE|Bone pain|Bone pain
C0151825|T184|IS|12584003|SNOMEDCT_CORE|Ostealgia|Bone pain
C0151825|T184|SY|12584003|SNOMEDCT_CORE|Osteodynia|Bone pain
C0151826|T184|SY|4568003|SNOMEDCT_CORE|Retrosternal chest pain|Retrosternal pain
C0151826|T184|PT|4568003|SNOMEDCT_CORE|Retrosternal pain|Retrosternal pain
C0151826|T184|FN|4568003|SNOMEDCT_CORE|Retrosternal pain|Retrosternal pain
C0151826|T184|IS|4568003|SNOMEDCT_CORE|Substernal chest pain|Retrosternal pain
C0151827|T184|SY|41652007|SNOMEDCT_CORE|Eye pain|Pain in eye
C0151827|T184|SY|41652007|SNOMEDCT_CORE|Ocular pain|Pain in eye
C0151827|T184|PT|41652007|SNOMEDCT_CORE|Pain in eye|Pain in eye
C0151827|T184|FN|41652007|SNOMEDCT_CORE|Pain in eye|Pain in eye
C0151849|T033|PT|274770006|SNOMEDCT_CORE|Alkaline phosphatase raised|Alkaline phosphatase raised
C0151849|T033|FN|274770006|SNOMEDCT_CORE|Alkaline phosphatase raised|Alkaline phosphatase raised
C0151878|T033|IS|111975006|SNOMEDCT_CORE|Increased Q-T interval|Prolonged QT interval
C0151878|T033|SY|111975006|SNOMEDCT_CORE|Increased QT interval|Prolonged QT interval
C0151878|T033|PT|111975006|SNOMEDCT_CORE|Prolonged QT interval|Prolonged QT interval
C0151878|T033|FN|111975006|SNOMEDCT_CORE|Prolonged QT interval|Prolonged QT interval
C0151889|T033|SY|86854008|SNOMEDCT_CORE|Exaggeration of the deep reflexes|Hyperreflexia
C0151889|T033|PT|86854008|SNOMEDCT_CORE|Hyperreflexia|Hyperreflexia
C0151889|T033|FN|86854008|SNOMEDCT_CORE|Hyperreflexia|Hyperreflexia
C0151889|T033|SY|86854008|SNOMEDCT_CORE|Increased tendon reflexes|Hyperreflexia
C0151900|T033|PT|165624002|SNOMEDCT_CORE|Serum iron raised|Serum iron raised
C0151900|T033|FN|165624002|SNOMEDCT_CORE|Serum iron raised|Serum iron raised
C0151907|T033|PT|3253007|SNOMEDCT_CORE|Discoloration of skin|Discoloration of skin
C0151907|T033|FN|3253007|SNOMEDCT_CORE|Discoloration of skin|Discoloration of skin
C0151907|T033|PTGB|3253007|SNOMEDCT_CORE|Discolouration of skin|Discoloration of skin
C0151907|T033|SY|3253007|SNOMEDCT_CORE|Dyschromia|Discoloration of skin
C0151908|T184|SY|16386004|SNOMEDCT_CORE|Anhydrotic skin|Dry skin
C0151908|T184|PT|16386004|SNOMEDCT_CORE|Dry skin|Dry skin
C0151908|T184|FN|16386004|SNOMEDCT_CORE|Dry skin|Dry skin
C0151942|T046|PT|65198009|SNOMEDCT_CORE|Arterial thrombosis|Arterial thrombosis
C0151942|T046|FN|65198009|SNOMEDCT_CORE|Arterial thrombosis|Arterial thrombosis
C0151942|T046|IS|65198009|SNOMEDCT_CORE|Arterial thrombosis, NOS, of unspecified artery|Arterial thrombosis
C0151970|T047|SY|30811009|SNOMEDCT_CORE|Esophageal ulcer|Ulcer of esophagus
C0151970|T047|SYGB|30811009|SNOMEDCT_CORE|Oesophageal ulcer|Ulcer of esophagus
C0151970|T047|SY|30811009|SNOMEDCT_CORE|OU - Esophageal ulcer|Ulcer of esophagus
C0151970|T047|SYGB|30811009|SNOMEDCT_CORE|OU - Oesophageal ulcer|Ulcer of esophagus
C0151970|T047|SY|30811009|SNOMEDCT_CORE|Peptic ulcer of esophagus|Ulcer of esophagus
C0151970|T047|SYGB|30811009|SNOMEDCT_CORE|Peptic ulcer of oesophagus|Ulcer of esophagus
C0151970|T047|SY|30811009|SNOMEDCT_CORE|Peptic ulceration of esophagus|Ulcer of esophagus
C0151970|T047|SYGB|30811009|SNOMEDCT_CORE|Peptic ulceration of oesophagus|Ulcer of esophagus
C0151970|T047|PT|30811009|SNOMEDCT_CORE|Ulcer of esophagus|Ulcer of esophagus
C0151970|T047|FN|30811009|SNOMEDCT_CORE|Ulcer of esophagus|Ulcer of esophagus
C0151970|T047|IS|30811009|SNOMEDCT_CORE|Ulcer of esophagus, NOS|Ulcer of esophagus
C0151970|T047|PTGB|30811009|SNOMEDCT_CORE|Ulcer of oesophagus|Ulcer of esophagus
C0151971|T047|IS|85942002|SNOMEDCT_CORE|Primary ulcer of intestine|Ulceration of intestine
C0151971|T047|IS|85942002|SNOMEDCT_CORE|Primary ulcer of intestine, NOS|Ulceration of intestine
C0151971|T047|PT|85942002|SNOMEDCT_CORE|Ulceration of intestine|Ulceration of intestine
C0151971|T047|FN|85942002|SNOMEDCT_CORE|Ulceration of intestine|Ulceration of intestine
C0151971|T047|IS|85942002|SNOMEDCT_CORE|Ulceration of intestine, NOS|Ulceration of intestine
C0151994|T033|PT|198319004|SNOMEDCT_CORE|Enlarged uterus|Enlarged uterus
C0151994|T033|FN|198319004|SNOMEDCT_CORE|Enlarged uterus|Enlarged uterus
C0151994|T033|SY|198319004|SNOMEDCT_CORE|Large uterus|Enlarged uterus
C0151994|T033|SY|198319004|SNOMEDCT_CORE|Uterine enlargement|Enlarged uterus
C0152013|T191|FN|254626006|SNOMEDCT_CORE|Adenocarcinoma of lung|Adenocarcinoma of lung
C0152013|T191|PT|254626006|SNOMEDCT_CORE|Adenocarcinoma of lung|Adenocarcinoma of lung
C0152018|T191|PT|372138000|SNOMEDCT_CORE|Carcinoma of esophagus|Carcinoma of esophagus
C0152018|T191|FN|372138000|SNOMEDCT_CORE|Carcinoma of esophagus|Carcinoma of esophagus
C0152018|T191|PTGB|372138000|SNOMEDCT_CORE|Carcinoma of oesophagus|Carcinoma of esophagus
C0152020|T047|SY|235675006|SNOMEDCT_CORE|Gastric atony|Gastroparesis syndrome
C0152020|T047|SY|235675006|SNOMEDCT_CORE|Gastric stasis|Gastroparesis syndrome
C0152020|T047|SY|235675006|SNOMEDCT_CORE|Gastroparesis|Gastroparesis syndrome
C0152020|T047|FN|235675006|SNOMEDCT_CORE|Gastroparesis|Gastroparesis syndrome
C0152020|T047|PT|235675006|SNOMEDCT_CORE|Gastroparesis syndrome|Gastroparesis syndrome
C0152021|T019|SY|13213009|SNOMEDCT_CORE|CHD - Congenital heart disease|Congenital heart disease
C0152021|T019|PT|13213009|SNOMEDCT_CORE|Congenital heart disease|Congenital heart disease
C0152021|T019|FN|13213009|SNOMEDCT_CORE|Congenital heart disease|Congenital heart disease
C0152021|T019|IS|13213009|SNOMEDCT_CORE|Congenital heart disease, NOS|Congenital heart disease
C0152025|T047|PT|42345000|SNOMEDCT_CORE|Polyneuropathy|Polyneuropathy
C0152025|T047|SY|42345000|SNOMEDCT_CORE|Polyneuropathy|Polyneuropathy
C0152025|T047|FN|42345000|SNOMEDCT_CORE|Polyneuropathy|Polyneuropathy
C0152025|T047|IS|42345000|SNOMEDCT_CORE|Polyneuropathy, NOS|Polyneuropathy
C0152029|T184|PT|82297005|SNOMEDCT_CORE|Congestion of nasal sinus|Congestion of nasal sinus
C0152029|T184|FN|82297005|SNOMEDCT_CORE|Congestion of nasal sinus|Congestion of nasal sinus
C0152029|T184|IS|82297005|SNOMEDCT_CORE|Congestion of nasal sinus, NOS|Congestion of nasal sinus
C0152029|T184|SY|82297005|SNOMEDCT_CORE|Sinus congestion|Congestion of nasal sinus
C0152029|T184|IS|82297005|SNOMEDCT_CORE|Sinus congestion, NOS|Congestion of nasal sinus
C0152030|T033|PT|367466007|SNOMEDCT_CORE|Skin irritation|Skin irritation
C0152030|T033|FN|367466007|SNOMEDCT_CORE|Skin irritation|Skin irritation
C0152031|T033|PT|271771009|SNOMEDCT_CORE|Joint swelling|Joint swelling
C0152031|T033|FN|271771009|SNOMEDCT_CORE|Joint swelling|Joint swelling
C0152031|T033|SY|271771009|SNOMEDCT_CORE|Observation of joint swelling|Joint swelling
C0152031|T033|SY|271771009|SNOMEDCT_CORE|Swollen joint|Joint swelling
C0152032|T184|PT|5972002|SNOMEDCT_CORE|Delay when starting to pass urine|Delay when starting to pass urine
C0152032|T184|FN|5972002|SNOMEDCT_CORE|Delay when starting to pass urine|Delay when starting to pass urine
C0152032|T184|SY|5972002|SNOMEDCT_CORE|Hesitancy|Delay when starting to pass urine
C0152032|T184|SY|5972002|SNOMEDCT_CORE|Hesitancy of micturition|Delay when starting to pass urine
C0152032|T184|SY|5972002|SNOMEDCT_CORE|Urinary hesitancy|Delay when starting to pass urine
C0152032|T184|SY|5972002|SNOMEDCT_CORE|Urinary hesitation|Delay when starting to pass urine
C0152086|T037|SY|58188004|SNOMEDCT_CORE|Posttraumatic arthropathy|Traumatic arthropathy
C0152086|T037|SY|58188004|SNOMEDCT_CORE|Traumatic arthritis|Traumatic arthropathy
C0152086|T037|PT|58188004|SNOMEDCT_CORE|Traumatic arthropathy|Traumatic arthropathy
C0152086|T037|FN|58188004|SNOMEDCT_CORE|Traumatic arthropathy|Traumatic arthropathy
C0152089|T047|SY|27151001|SNOMEDCT_CORE|Failed back syndrome|Post-laminectomy syndrome
C0152089|T047|PT|27151001|SNOMEDCT_CORE|Post-laminectomy syndrome|Post-laminectomy syndrome
C0152089|T047|FN|27151001|SNOMEDCT_CORE|Post-laminectomy syndrome|Post-laminectomy syndrome
C0152089|T047|IS|27151001|SNOMEDCT_CORE|Postlaminectomy syndrome|Post-laminectomy syndrome
C0152089|T047|IS|27151001|SNOMEDCT_CORE|Postlaminectomy syndrome, NOS|Post-laminectomy syndrome
C0152097|T047|SY|48475001|SNOMEDCT_CORE|Diaphragmatic disease|Disorder of diaphragm
C0152097|T047|SY|48475001|SNOMEDCT_CORE|Diaphragmatic disorder|Disorder of diaphragm
C0152097|T047|IS|48475001|SNOMEDCT_CORE|Disease of diaphragm|Disorder of diaphragm
C0152097|T047|OF|48475001|SNOMEDCT_CORE|Disease of diaphragm|Disorder of diaphragm
C0152097|T047|IS|48475001|SNOMEDCT_CORE|Disease of diaphragm, NOS|Disorder of diaphragm
C0152097|T047|PT|48475001|SNOMEDCT_CORE|Disorder of diaphragm|Disorder of diaphragm
C0152097|T047|FN|48475001|SNOMEDCT_CORE|Disorder of diaphragm|Disorder of diaphragm
C0152105|T047|SY|64715009|SNOMEDCT_CORE|HHD - Hypertensive heart disease|Hypertensive heart disease
C0152105|T047|SY|64715009|SNOMEDCT_CORE|Hypertensive cardiopathy|Hypertensive heart disease
C0152105|T047|SY|64715009|SNOMEDCT_CORE|Hypertensive cardiovascular disease|Hypertensive heart disease
C0152105|T047|FN|64715009|SNOMEDCT_CORE|Hypertensive heart disease|Hypertensive heart disease
C0152105|T047|PT|64715009|SNOMEDCT_CORE|Hypertensive heart disease|Hypertensive heart disease
C0152105|T047|IS|64715009|SNOMEDCT_CORE|Hypertensive heart disease, NOS|Hypertensive heart disease
C0152110|T047|SY|85007004|SNOMEDCT_CORE|Bernhardt-Rot syndrome|Meralgia paresthetica
C0152110|T047|SYGB|85007004|SNOMEDCT_CORE|Bernhardt's paraesthesia|Meralgia paresthetica
C0152110|T047|SY|85007004|SNOMEDCT_CORE|Bernhardt's paresthesia|Meralgia paresthetica
C0152110|T047|SY|85007004|SNOMEDCT_CORE|Compression of lateral cutaneous femoral nerve of thigh|Meralgia paresthetica
C0152110|T047|SY|85007004|SNOMEDCT_CORE|Entrapment of lateral cutaneous nerve of thigh|Meralgia paresthetica
C0152110|T047|SY|85007004|SNOMEDCT_CORE|Lateral cutaneous femoral nerve of thigh syndrome|Meralgia paresthetica
C0152110|T047|PTGB|85007004|SNOMEDCT_CORE|Meralgia paraesthetica|Meralgia paresthetica
C0152110|T047|PT|85007004|SNOMEDCT_CORE|Meralgia paresthetica|Meralgia paresthetica
C0152110|T047|FN|85007004|SNOMEDCT_CORE|Meralgia paresthetica|Meralgia paresthetica
C0152116|T184|SY|74333002|SNOMEDCT_CORE|Cervical dystonia|Spasmodic torticollis
C0152116|T184|PT|74333002|SNOMEDCT_CORE|Spasmodic torticollis|Spasmodic torticollis
C0152116|T184|FN|74333002|SNOMEDCT_CORE|Spasmodic torticollis|Spasmodic torticollis
C0152121|T047|OAP|19033007|SNOMEDCT_CORE|Pseudoclaudication syndrome|Pseudoclaudication syndrome
C0152121|T047|OAF|19033007|SNOMEDCT_CORE|Pseudoclaudication syndrome|Pseudoclaudication syndrome
C0152132|T047|PT|6962006|SNOMEDCT_CORE|Hypertensive retinopathy|Hypertensive retinopathy
C0152132|T047|FN|6962006|SNOMEDCT_CORE|Hypertensive retinopathy|Hypertensive retinopathy
C0152136|T047|PT|50485007|SNOMEDCT_CORE|Low tension glaucoma|Low tension glaucoma
C0152136|T047|FN|50485007|SNOMEDCT_CORE|Low tension glaucoma|Low tension glaucoma
C0152136|T047|SY|50485007|SNOMEDCT_CORE|LTG - Low tension glaucoma|Low tension glaucoma
C0152136|T047|SY|50485007|SNOMEDCT_CORE|Normal pressure glaucoma|Low tension glaucoma
C0152136|T047|SY|50485007|SNOMEDCT_CORE|Normal tension glaucoma|Low tension glaucoma
C0152150|T033|PT|65147003|SNOMEDCT_CORE|Twin pregnancy|Twin pregnancy
C0152150|T033|FN|65147003|SNOMEDCT_CORE|Twin pregnancy|Twin pregnancy
C0152162|T033|SY|402410006|SNOMEDCT_CORE|Factitious urticaria|Factitious urticaria
C0152164|T047|SY|18773000|SNOMEDCT_CORE|Cyclical vomiting|Cyclical vomiting syndrome
C0152164|T047|FN|18773000|SNOMEDCT_CORE|Cyclical vomiting syndrome|Cyclical vomiting syndrome
C0152164|T047|PT|18773000|SNOMEDCT_CORE|Cyclical vomiting syndrome|Cyclical vomiting syndrome
C0152164|T047|SY|18773000|SNOMEDCT_CORE|Periodic vomiting|Cyclical vomiting syndrome
C0152165|T184|SY|196746003|SNOMEDCT_CORE|Emesis - persistent|Persistent vomiting
C0152165|T184|PT|196746003|SNOMEDCT_CORE|Persistent vomiting|Persistent vomiting
C0152165|T184|FN|196746003|SNOMEDCT_CORE|Persistent vomiting|Persistent vomiting
C0152169|T184|PT|7093002|SNOMEDCT_CORE|Renal colic|Ureteric colic
C0152169|T184|FN|7093002|SNOMEDCT_CORE|Renal colic|Ureteric colic
C0152169|T184|IS|17329003|SNOMEDCT_CORE|Ureteral colic|Ureteric colic
C0152169|T184|PT|17329003|SNOMEDCT_CORE|Ureteric colic|Ureteric colic
C0152169|T184|FN|17329003|SNOMEDCT_CORE|Ureteric colic|Ureteric colic
C0152171|T047|OAS|26174007|SNOMEDCT_CORE|Essential pulmonary hypertension|Primary pulmonary hypertension
C0152171|T047|IS|26174007|SNOMEDCT_CORE|Idiopathic pulmonary hypertension|Primary pulmonary hypertension
C0152171|T047|OAS|26174007|SNOMEDCT_CORE|PPHT - Primary pulmonary hypertension|Primary pulmonary hypertension
C0152171|T047|OAP|26174007|SNOMEDCT_CORE|Primary pulmonary hypertension|Primary pulmonary hypertension
C0152171|T047|OAF|26174007|SNOMEDCT_CORE|Primary pulmonary hypertension|Primary pulmonary hypertension
C0152172|T047|SY|59021001|SNOMEDCT_CORE|Angina at rest|Angina decubitus
C0152172|T047|PT|59021001|SNOMEDCT_CORE|Angina decubitus|Angina decubitus
C0152172|T047|FN|59021001|SNOMEDCT_CORE|Angina decubitus|Angina decubitus
C0152172|T047|SY|59021001|SNOMEDCT_CORE|Anginal chest pain at rest|Angina decubitus
C0152174|T048|SY|8971008|SNOMEDCT_CORE|Algopsychalia|Psychalgia
C0152174|T048|PT|8971008|SNOMEDCT_CORE|Psychalgia|Psychalgia
C0152174|T048|FN|8971008|SNOMEDCT_CORE|Psychalgia|Psychalgia
C0152174|T048|SY|8971008|SNOMEDCT_CORE|Psychogenic pain|Psychalgia
C0152177|T047|SY|64309007|SNOMEDCT_CORE|Disorder of the fifth cranial nerve|Trigeminal nerve disorder
C0152177|T047|IS|64309007|SNOMEDCT_CORE|Disorder of the fifth cranial nerve, NOS|Trigeminal nerve disorder
C0152177|T047|SY|64309007|SNOMEDCT_CORE|Disorders of the fifth nerve|Trigeminal nerve disorder
C0152177|T047|SY|64309007|SNOMEDCT_CORE|Disorders of the Vth cranial nerve|Trigeminal nerve disorder
C0152177|T047|PT|64309007|SNOMEDCT_CORE|Trigeminal nerve disorder|Trigeminal nerve disorder
C0152177|T047|FN|64309007|SNOMEDCT_CORE|Trigeminal nerve disorder|Trigeminal nerve disorder
C0152177|T047|IS|64309007|SNOMEDCT_CORE|Trigeminal nerve disorder, NOS|Trigeminal nerve disorder
C0152187|T020|SY|193638002|SNOMEDCT_CORE|Amblyopia ex anopsia|Amblyopia ex anopsia
C0152189|T047|SY|193638002|SNOMEDCT_CORE|Deprivation amblyopia|Stimulus deprivation amblyopia
C0152189|T047|SY|193638002|SNOMEDCT_CORE|Disuse amblyopia|Stimulus deprivation amblyopia
C0152189|T047|IS|193638002|SNOMEDCT_CORE|Disuse ambylopia|Stimulus deprivation amblyopia
C0152189|T047|PT|193638002|SNOMEDCT_CORE|Stimulus deprivation amblyopia|Stimulus deprivation amblyopia
C0152189|T047|FN|193638002|SNOMEDCT_CORE|Stimulus deprivation amblyopia|Stimulus deprivation amblyopia
C0152190|T047|SY|90927000|SNOMEDCT_CORE|Ametropic amblyopia|Refractive amblyopia
C0152190|T047|SY|90927000|SNOMEDCT_CORE|Meridional amblyopia|Refractive amblyopia
C0152190|T047|PT|90927000|SNOMEDCT_CORE|Refractive amblyopia|Refractive amblyopia
C0152190|T047|FN|90927000|SNOMEDCT_CORE|Refractive amblyopia|Refractive amblyopia
C0152193|T047|PT|68905002|SNOMEDCT_CORE|Regular astigmatism|Regular astigmatism
C0152193|T047|FN|68905002|SNOMEDCT_CORE|Regular astigmatism|Regular astigmatism
C0152194|T047|PT|47099006|SNOMEDCT_CORE|Irregular astigmatism|Irregular astigmatism
C0152194|T047|FN|47099006|SNOMEDCT_CORE|Irregular astigmatism|Irregular astigmatism
C0152205|T047|PT|39837002|SNOMEDCT_CORE|Alternating esotropia|Alternating esotropia
C0152205|T047|FN|39837002|SNOMEDCT_CORE|Alternating esotropia|Alternating esotropia
C0152205|T047|IS|39837002|SNOMEDCT_CORE|Alternating esotropia, NOS|Alternating esotropia
C0152207|T047|PT|37214009|SNOMEDCT_CORE|Alternating exotropia|Alternating exotropia
C0152207|T047|FN|37214009|SNOMEDCT_CORE|Alternating exotropia|Alternating exotropia
C0152207|T047|IS|37214009|SNOMEDCT_CORE|Alternating exotropia, NOS|Alternating exotropia
C0152218|T047|PT|20636006|SNOMEDCT_CORE|Vertical heterophoria|Vertical heterophoria
C0152218|T047|FN|20636006|SNOMEDCT_CORE|Vertical heterophoria|Vertical heterophoria
C0152218|T047|IS|20636006|SNOMEDCT_CORE|Vertical heterophoria, NOS|Vertical heterophoria
C0152226|T047|SY|60735000|SNOMEDCT_CORE|Defective lid closure|Lagophthalmos
C0152226|T047|PT|60735000|SNOMEDCT_CORE|Lagophthalmos|Lagophthalmos
C0152226|T047|OF|60735000|SNOMEDCT_CORE|Lagophthalmos|Lagophthalmos
C0152226|T047|FN|60735000|SNOMEDCT_CORE|Lagophthalmos|Lagophthalmos
C0152226|T047|IS|60735000|SNOMEDCT_CORE|Lagophthalmos, NOS|Lagophthalmos
C0152226|T047|SY|60735000|SNOMEDCT_CORE|Poor closure eyelids|Lagophthalmos
C0152227|T047|OF|193982009|SNOMEDCT_CORE|Epiphora|Epiphora
C0152227|T047|PT|193982009|SNOMEDCT_CORE|Epiphora|Epiphora
C0152227|T047|FN|193982009|SNOMEDCT_CORE|Epiphora|Epiphora
C0152227|T047|SY|193982009|SNOMEDCT_CORE|Tearing|Epiphora
C0152244|T047|SY|203468000|SNOMEDCT_CORE|ABC - Aneurysmal bone cyst|Aneurysmal bone cyst
C0152244|T047|PT|203468000|SNOMEDCT_CORE|Aneurysmal bone cyst|Aneurysmal bone cyst
C0152244|T047|FN|203468000|SNOMEDCT_CORE|Aneurysmal bone cyst|Aneurysmal bone cyst
C0152247|T020|PT|6929003|SNOMEDCT_CORE|Urethral caruncle|Urethral caruncle
C0152247|T020|FN|6929003|SNOMEDCT_CORE|Urethral caruncle|Urethral caruncle
C0152255|T047|PT|87614000|SNOMEDCT_CORE|Pinguecula|Pinguecula
C0152255|T047|FN|87614000|SNOMEDCT_CORE|Pinguecula|Pinguecula
C0152255|T047|SY|87614000|SNOMEDCT_CORE|Pinguicula|Pinguecula
C0152257|T020|PT|193590000|SNOMEDCT_CORE|Total, mature senile cataract|Total, mature senile cataract
C0152257|T020|FN|193590000|SNOMEDCT_CORE|Total, mature senile cataract|Total, mature senile cataract
C0152259|T047|PT|193600001|SNOMEDCT_CORE|Cataract secondary to ocular disease|Cataract secondary to ocular disease
C0152259|T047|FN|193600001|SNOMEDCT_CORE|Cataract secondary to ocular disease|Cataract secondary to ocular disease
C0152259|T047|SY|193600001|SNOMEDCT_CORE|Cataracta complicata|Cataract secondary to ocular disease
C0152259|T047|SY|193600001|SNOMEDCT_CORE|Complicated cataract|Cataract secondary to ocular disease
C0152268|T191|SY|118608000|SNOMEDCT_CORE|Hodgkin disease, nodular sclerosis|Hodgkin's disease, nodular sclerosis
C0152268|T191|SY|118608000|SNOMEDCT_CORE|Hodgkin's disease, nodular sclerosis|Hodgkin's disease, nodular sclerosis
C0152268|T191|PT|118608000|SNOMEDCT_CORE|Hodgkin's disease, nodular sclerosis|Hodgkin's disease, nodular sclerosis
C0152268|T191|FN|118608000|SNOMEDCT_CORE|Hodgkin's disease, nodular sclerosis|Hodgkin's disease, nodular sclerosis
C0152413|T047|FN|195881003|SNOMEDCT_CORE|Pneumonia caused by respiratory syncytial virus|Pneumonia due to respiratory syncytial virus
C0152413|T047|SY|195881003|SNOMEDCT_CORE|Pneumonia caused by respiratory syncytial virus|Pneumonia due to respiratory syncytial virus
C0152413|T047|PT|195881003|SNOMEDCT_CORE|Pneumonia due to respiratory syncytial virus|Pneumonia due to respiratory syncytial virus
C0152413|T047|OF|195881003|SNOMEDCT_CORE|Pneumonia due to respiratory syncytial virus|Pneumonia due to respiratory syncytial virus
C0152415|T019|SY|67787004|SNOMEDCT_CORE|Ankyloglossia|Tongue tie
C0152415|T019|PT|67787004|SNOMEDCT_CORE|Tongue tie|Tongue tie
C0152415|T019|FN|67787004|SNOMEDCT_CORE|Tongue tie|Tongue tie
C0152415|T019|SY|67787004|SNOMEDCT_CORE|Tongue-tie|Tongue tie
C0152417|T019|PT|18546004|SNOMEDCT_CORE|Congenital stenosis of aortic valve|Congenital stenosis of aortic valve
C0152417|T019|FN|18546004|SNOMEDCT_CORE|Congenital stenosis of aortic valve|Congenital stenosis of aortic valve
C0152424|T019|IS|30288003|SNOMEDCT_CORE|Absence of interventricular septum|Common ventricle
C0152424|T019|SY|45503006|SNOMEDCT_CORE|Absence of interventricular septum|Common ventricle
C0152424|T019|PT|45503006|SNOMEDCT_CORE|Common ventricle|Common ventricle
C0152424|T019|FN|45503006|SNOMEDCT_CORE|Common ventricle|Common ventricle
C0152424|T019|SY|45503006|SNOMEDCT_CORE|Cor triloculare biatriatum|Common ventricle
C0152424|T019|SY|45503006|SNOMEDCT_CORE|Single ventricle|Common ventricle
C0152432|T019|SY|79168008|SNOMEDCT_CORE|Congenital bow leg|Congenital genu varum
C0152432|T019|SY|79168008|SNOMEDCT_CORE|Congenital bowed limb|Congenital genu varum
C0152432|T019|SY|79168008|SNOMEDCT_CORE|Congenital bowleg|Congenital genu varum
C0152432|T019|PT|79168008|SNOMEDCT_CORE|Congenital genu varum|Congenital genu varum
C0152432|T019|FN|79168008|SNOMEDCT_CORE|Congenital genu varum|Congenital genu varum
C0152432|T019|SY|79168008|SNOMEDCT_CORE|Congenital varus deformity of knee|Congenital genu varum
C0152439|T047|PT|44268007|SNOMEDCT_CORE|Retinoschisis|Retinoschisis
C0152439|T047|FN|44268007|SNOMEDCT_CORE|Retinoschisis|Retinoschisis
C0152439|T047|IS|44268007|SNOMEDCT_CORE|Retinoschisis, NOS|Retinoschisis
C0152439|T047|SY|44268007|SNOMEDCT_CORE|RS - Retinoschisis|Retinoschisis
C0152439|T047|SY|44268007|SNOMEDCT_CORE|Schisis of retina|Retinoschisis
C0152447|T184|SY|9957009|SNOMEDCT_CORE|Observation of urethral discharge|Urethral discharge
C0152447|T184|SY|9957009|SNOMEDCT_CORE|UD - Urethral discharge|Urethral discharge
C0152447|T184|PT|9957009|SNOMEDCT_CORE|Urethral discharge|Urethral discharge
C0152447|T184|FN|9957009|SNOMEDCT_CORE|Urethral discharge|Urethral discharge
C0152447|T184|SY|9957009|SNOMEDCT_CORE|Urethrorrhea|Urethral discharge
C0152447|T184|SYGB|9957009|SNOMEDCT_CORE|Urethrorrhoea|Urethral discharge
C0152451|T047|SY|20917003|SNOMEDCT_CORE|CGN - Chronic glomerulonephritis|Chronic glomerulonephritis
C0152451|T047|PT|20917003|SNOMEDCT_CORE|Chronic glomerulonephritis|Chronic glomerulonephritis
C0152451|T047|FN|20917003|SNOMEDCT_CORE|Chronic glomerulonephritis|Chronic glomerulonephritis
C0152451|T047|IS|20917003|SNOMEDCT_CORE|Chronic glomerulonephritis, NOS|Chronic glomerulonephritis
C0152459|T020|PT|201067006|SNOMEDCT_CORE|Physiological striae|Physiological striae
C0152459|T020|FN|201067006|SNOMEDCT_CORE|Physiological striae|Physiological striae
C0152459|T020|SY|201067006|SNOMEDCT_CORE|Stretch marks|Physiological striae
C0152459|T020|SY|201067006|SNOMEDCT_CORE|Striae distensae|Physiological striae
C0152516|T047|PT|75375008|SNOMEDCT_CORE|Bacterial enteritis|Bacterial enteritis
C0152516|T047|FN|75375008|SNOMEDCT_CORE|Bacterial enteritis|Bacterial enteritis
C0152516|T047|IS|75375008|SNOMEDCT_CORE|Bacterial enteritis, NOS|Bacterial enteritis
C0152516|T047|SY|75375008|SNOMEDCT_CORE|Intestinal infection due to bacteria|Bacterial enteritis
C0152516|T047|SY|75375008|SNOMEDCT_CORE|Septic enteritis|Bacterial enteritis
C0152517|T047|SY|111843007|SNOMEDCT_CORE|Viral diarrhea|Viral gastroenteritis
C0152517|T047|SYGB|111843007|SNOMEDCT_CORE|Viral diarrhoea|Viral gastroenteritis
C0152517|T047|PT|111843007|SNOMEDCT_CORE|Viral gastroenteritis|Viral gastroenteritis
C0152517|T047|FN|111843007|SNOMEDCT_CORE|Viral gastroenteritis|Viral gastroenteritis
C0152517|T047|SY|111843007|SNOMEDCT_CORE|Viral vomiting|Viral gastroenteritis
C0152522|T047|PT|43240000|SNOMEDCT_CORE|Diarrhea of presumed infectious origin|Diarrhea of presumed infectious origin
C0152522|T047|FN|43240000|SNOMEDCT_CORE|Diarrhea of presumed infectious origin|Diarrhea of presumed infectious origin
C0152522|T047|PTGB|43240000|SNOMEDCT_CORE|Diarrhoea of presumed infectious origin|Diarrhea of presumed infectious origin
C0152964|T047|OAP|29577008|SNOMEDCT_CORE|Streptococcal septicaemia|Streptococcal septicemia
C0152964|T047|OAP|29577008|SNOMEDCT_CORE|Streptococcal septicemia|Streptococcal septicemia
C0152964|T047|OAF|29577008|SNOMEDCT_CORE|Streptococcal septicemia|Streptococcal septicemia
C0152965|T047|OAP|111821004|SNOMEDCT_CORE|Staphylococcal septicaemia|Staphylococcal septicemia
C0152965|T047|OAP|111821004|SNOMEDCT_CORE|Staphylococcal septicemia|Staphylococcal septicemia
C0152965|T047|OAF|111821004|SNOMEDCT_CORE|Staphylococcal septicemia|Staphylococcal septicemia
C0153027|T047|IS|42448002|SNOMEDCT_CORE|Herpes zoster keratitis|Herpes zoster keratoconjunctivitis
C0153027|T047|PT|42448002|SNOMEDCT_CORE|Herpes zoster keratoconjunctivitis|Herpes zoster keratoconjunctivitis
C0153027|T047|FN|42448002|SNOMEDCT_CORE|Herpes zoster keratoconjunctivitis|Herpes zoster keratoconjunctivitis
C0153027|T047|SY|42448002|SNOMEDCT_CORE|Herpes zoster with keratoconjunctivitis|Herpes zoster keratoconjunctivitis
C0153033|T047|SY|59819007|SNOMEDCT_CORE|Herpes simplex vulvitis|Herpetic ulceration of vulva
C0153033|T047|PT|59819007|SNOMEDCT_CORE|Herpetic ulceration of vulva|Herpetic ulceration of vulva
C0153033|T047|FN|59819007|SNOMEDCT_CORE|Herpetic ulceration of vulva|Herpetic ulceration of vulva
C0153038|T047|PT|59523007|SNOMEDCT_CORE|Herpes simplex disciform keratitis|Herpes simplex disciform keratitis
C0153038|T047|FN|59523007|SNOMEDCT_CORE|Herpes simplex disciform keratitis|Herpes simplex disciform keratitis
C0153038|T047|SY|59523007|SNOMEDCT_CORE|HSV disciform keratitis|Herpes simplex disciform keratitis
C0153062|T047|IS|186504007|SNOMEDCT_CORE|Nonspecific viral rash|Viral exanthem
C0153062|T047|OAP|186504007|SNOMEDCT_CORE|Viral disease characterised by exanthem|Viral exanthem
C0153062|T047|OAP|186504007|SNOMEDCT_CORE|Viral disease characterized by exanthem|Viral exanthem
C0153062|T047|OAF|186504007|SNOMEDCT_CORE|Viral disease characterized by exanthem|Viral exanthem
C0153062|T047|PT|49882001|SNOMEDCT_CORE|Viral exanthem|Viral exanthem
C0153062|T047|FN|49882001|SNOMEDCT_CORE|Viral exanthem|Viral exanthem
C0153062|T047|SY|49882001|SNOMEDCT_CORE|Viral exanthemata|Viral exanthem
C0153062|T047|SY|49882001|SNOMEDCT_CORE|Viral rash|Viral exanthem
C0153113|T047|SY|186738001|SNOMEDCT_CORE|Acute peripheral vestibulopathy|Acute peripheral vestibulopathy
C0153278|T047|PT|187058000|SNOMEDCT_CORE|Histoplasmosis with retinitis|Histoplasmosis with retinitis
C0153278|T047|FN|187058000|SNOMEDCT_CORE|Histoplasmosis with retinitis|Histoplasmosis with retinitis
C0153349|T191|SY|363375006|SNOMEDCT_CORE|CA - Cancer of tongue|Malignant tumor of tongue
C0153349|T191|SY|363375006|SNOMEDCT_CORE|Cancer of tongue|Malignant tumor of tongue
C0153349|T191|PT|363375006|SNOMEDCT_CORE|Malignant tumor of tongue|Malignant tumor of tongue
C0153349|T191|FN|363375006|SNOMEDCT_CORE|Malignant tumor of tongue|Malignant tumor of tongue
C0153349|T191|PTGB|363375006|SNOMEDCT_CORE|Malignant tumour of tongue|Malignant tumor of tongue
C0153354|T191|PT|363360003|SNOMEDCT_CORE|Malignant tumor of anterior two-thirds of tongue|Malignant tumor of anterior two-thirds of tongue
C0153354|T191|FN|363360003|SNOMEDCT_CORE|Malignant tumor of anterior two-thirds of tongue|Malignant tumor of anterior two-thirds of tongue
C0153354|T191|PTGB|363360003|SNOMEDCT_CORE|Malignant tumour of anterior two-thirds of tongue|Malignant tumor of anterior two-thirds of tongue
C0153368|T191|SY|363385007|SNOMEDCT_CORE|CA - Cancer of floor of mouth|Malignant tumor of floor of mouth
C0153368|T191|SY|363385007|SNOMEDCT_CORE|Cancer of floor of mouth|Malignant tumor of floor of mouth
C0153368|T191|SY|363385007|SNOMEDCT_CORE|FOM - Cancer of floor of mouth|Malignant tumor of floor of mouth
C0153368|T191|SY|363385007|SNOMEDCT_CORE|FOM - Malignant tumor of floor of mouth|Malignant tumor of floor of mouth
C0153368|T191|SYGB|363385007|SNOMEDCT_CORE|FOM - Malignant tumour of floor of mouth|Malignant tumor of floor of mouth
C0153368|T191|SY|363385007|SNOMEDCT_CORE|Malignant neoplasm of floor of mouth|Malignant tumor of floor of mouth
C0153368|T191|PT|363385007|SNOMEDCT_CORE|Malignant tumor of floor of mouth|Malignant tumor of floor of mouth
C0153368|T191|FN|363385007|SNOMEDCT_CORE|Malignant tumor of floor of mouth|Malignant tumor of floor of mouth
C0153368|T191|PTGB|363385007|SNOMEDCT_CORE|Malignant tumour of floor of mouth|Malignant tumor of floor of mouth
C0153378|T191|SY|363390005|SNOMEDCT_CORE|CA - Cancer of palate|Malignant tumor of palate
C0153378|T191|SY|363390005|SNOMEDCT_CORE|Cancer of palate|Malignant tumor of palate
C0153378|T191|SY|363390005|SNOMEDCT_CORE|Malignant neoplasm of roof of mouth|Malignant tumor of palate
C0153378|T191|PT|363390005|SNOMEDCT_CORE|Malignant tumor of palate|Malignant tumor of palate
C0153378|T191|FN|363390005|SNOMEDCT_CORE|Malignant tumor of palate|Malignant tumor of palate
C0153378|T191|SY|363390005|SNOMEDCT_CORE|Malignant tumor of roof of mouth|Malignant tumor of palate
C0153378|T191|PTGB|363390005|SNOMEDCT_CORE|Malignant tumour of palate|Malignant tumor of palate
C0153378|T191|SYGB|363390005|SNOMEDCT_CORE|Malignant tumour of roof of mouth|Malignant tumor of palate
C0153381|T191|SY|363505006|SNOMEDCT_CORE|CA - Mouth cancer|Malignant tumor of oral cavity
C0153381|T191|SY|363505006|SNOMEDCT_CORE|Cancer of oral cavity|Malignant tumor of oral cavity
C0153381|T191|SY|363505006|SNOMEDCT_CORE|Malignant neoplasm of mouth|Malignant tumor of oral cavity
C0153381|T191|SY|363505006|SNOMEDCT_CORE|Malignant tumor of mouth|Malignant tumor of oral cavity
C0153381|T191|PT|363505006|SNOMEDCT_CORE|Malignant tumor of oral cavity|Malignant tumor of oral cavity
C0153381|T191|FN|363505006|SNOMEDCT_CORE|Malignant tumor of oral cavity|Malignant tumor of oral cavity
C0153381|T191|SYGB|363505006|SNOMEDCT_CORE|Malignant tumour of mouth|Malignant tumor of oral cavity
C0153381|T191|PTGB|363505006|SNOMEDCT_CORE|Malignant tumour of oral cavity|Malignant tumor of oral cavity
C0153381|T191|SY|363505006|SNOMEDCT_CORE|Mouth cancer|Malignant tumor of oral cavity
C0153382|T191|SY|363392002|SNOMEDCT_CORE|CA - Cancer of oropharynx|Malignant tumor of oropharynx
C0153382|T191|SY|363392002|SNOMEDCT_CORE|Cancer of oropharynx|Malignant tumor of oropharynx
C0153382|T191|SY|363392002|SNOMEDCT_CORE|Malignant tumor of mesopharynx|Malignant tumor of oropharynx
C0153382|T191|PT|363392002|SNOMEDCT_CORE|Malignant tumor of oropharynx|Malignant tumor of oropharynx
C0153382|T191|FN|363392002|SNOMEDCT_CORE|Malignant tumor of oropharynx|Malignant tumor of oropharynx
C0153382|T191|SYGB|363392002|SNOMEDCT_CORE|Malignant tumour of mesopharynx|Malignant tumor of oropharynx
C0153382|T191|PTGB|363392002|SNOMEDCT_CORE|Malignant tumour of oropharynx|Malignant tumor of oropharynx
C0153392|T191|SY|187692001|SNOMEDCT_CORE|Malignant neoplasm of nasopharynx|Malignant tumor of nasopharynx
C0153392|T191|SY|187692001|SNOMEDCT_CORE|Malignant tumor of epipharynx|Malignant tumor of nasopharynx
C0153392|T191|PT|187692001|SNOMEDCT_CORE|Malignant tumor of nasopharynx|Malignant tumor of nasopharynx
C0153392|T191|FN|187692001|SNOMEDCT_CORE|Malignant tumor of nasopharynx|Malignant tumor of nasopharynx
C0153392|T191|SY|187692001|SNOMEDCT_CORE|Malignant tumor of postnasal space|Malignant tumor of nasopharynx
C0153392|T191|SYGB|187692001|SNOMEDCT_CORE|Malignant tumour of epipharynx|Malignant tumor of nasopharynx
C0153392|T191|PTGB|187692001|SNOMEDCT_CORE|Malignant tumour of nasopharynx|Malignant tumor of nasopharynx
C0153392|T191|SYGB|187692001|SNOMEDCT_CORE|Malignant tumour of postnasal space|Malignant tumor of nasopharynx
C0153398|T191|SY|363399006|SNOMEDCT_CORE|Malignant neoplasm of laryngopharynx|Malignant tumor of hypopharynx
C0153398|T191|PT|363399006|SNOMEDCT_CORE|Malignant tumor of hypopharynx|Malignant tumor of hypopharynx
C0153398|T191|FN|363399006|SNOMEDCT_CORE|Malignant tumor of hypopharynx|Malignant tumor of hypopharynx
C0153398|T191|SY|363399006|SNOMEDCT_CORE|Malignant tumor of laryngopharynx|Malignant tumor of hypopharynx
C0153398|T191|PTGB|363399006|SNOMEDCT_CORE|Malignant tumour of hypopharynx|Malignant tumor of hypopharynx
C0153398|T191|SYGB|363399006|SNOMEDCT_CORE|Malignant tumour of laryngopharynx|Malignant tumor of hypopharynx
C0153411|T191|SY|187723009|SNOMEDCT_CORE|Malignant neoplasm of thoracic esophagus|Malignant tumor of thoracic part of esophagus
C0153411|T191|SYGB|187723009|SNOMEDCT_CORE|Malignant neoplasm of thoracic oesophagus|Malignant tumor of thoracic part of esophagus
C0153411|T191|PT|187723009|SNOMEDCT_CORE|Malignant tumor of thoracic part of esophagus|Malignant tumor of thoracic part of esophagus
C0153411|T191|FN|187723009|SNOMEDCT_CORE|Malignant tumor of thoracic part of esophagus|Malignant tumor of thoracic part of esophagus
C0153411|T191|PTGB|187723009|SNOMEDCT_CORE|Malignant tumour of thoracic part of oesophagus|Malignant tumor of thoracic part of esophagus
C0153414|T191|SY|187726001|SNOMEDCT_CORE|Ca middle third esophagus|Malignant tumor of middle third of esophagus
C0153414|T191|SYGB|187726001|SNOMEDCT_CORE|Ca middle third oesophagus|Malignant tumor of middle third of esophagus
C0153414|T191|SY|187726001|SNOMEDCT_CORE|Malignant neoplasm of middle third of esophagus|Malignant tumor of middle third of esophagus
C0153414|T191|SYGB|187726001|SNOMEDCT_CORE|Malignant neoplasm of middle third of oesophagus|Malignant tumor of middle third of esophagus
C0153414|T191|PT|187726001|SNOMEDCT_CORE|Malignant tumor of middle third of esophagus|Malignant tumor of middle third of esophagus
C0153414|T191|FN|187726001|SNOMEDCT_CORE|Malignant tumor of middle third of esophagus|Malignant tumor of middle third of esophagus
C0153414|T191|PTGB|187726001|SNOMEDCT_CORE|Malignant tumour of middle third of oesophagus|Malignant tumor of middle third of esophagus
C0153415|T191|SY|187727005|SNOMEDCT_CORE|Ca lower third esophagus|Malignant tumor of lower third of esophagus
C0153415|T191|SYGB|187727005|SNOMEDCT_CORE|Ca lower third oesophagus|Malignant tumor of lower third of esophagus
C0153415|T191|SY|187727005|SNOMEDCT_CORE|Malignant neoplasm of lower third of esophagus|Malignant tumor of lower third of esophagus
C0153415|T191|SYGB|187727005|SNOMEDCT_CORE|Malignant neoplasm of lower third of oesophagus|Malignant tumor of lower third of esophagus
C0153415|T191|PT|187727005|SNOMEDCT_CORE|Malignant tumor of lower third of esophagus|Malignant tumor of lower third of esophagus
C0153415|T191|FN|187727005|SNOMEDCT_CORE|Malignant tumor of lower third of esophagus|Malignant tumor of lower third of esophagus
C0153415|T191|PTGB|187727005|SNOMEDCT_CORE|Malignant tumour of lower third of oesophagus|Malignant tumor of lower third of esophagus
C0153417|T191|SY|187732006|SNOMEDCT_CORE|Ca cardia - stomach|Malignant tumor of cardia
C0153417|T191|SY|187732006|SNOMEDCT_CORE|Malignant neoplasm of cardia of stomach|Malignant tumor of cardia
C0153417|T191|PT|187732006|SNOMEDCT_CORE|Malignant tumor of cardia|Malignant tumor of cardia
C0153417|T191|FN|187732006|SNOMEDCT_CORE|Malignant tumor of cardia|Malignant tumor of cardia
C0153417|T191|PTGB|187732006|SNOMEDCT_CORE|Malignant tumour of cardia|Malignant tumor of cardia
C0153422|T191|SY|269459004|SNOMEDCT_CORE|Ca lesser curvature - stomach|Malignant tumor of lesser curve of stomach
C0153422|T191|PT|269459004|SNOMEDCT_CORE|Malignant tumor of lesser curve of stomach|Malignant tumor of lesser curve of stomach
C0153422|T191|FN|269459004|SNOMEDCT_CORE|Malignant tumor of lesser curve of stomach|Malignant tumor of lesser curve of stomach
C0153422|T191|PTGB|269459004|SNOMEDCT_CORE|Malignant tumour of lesser curve of stomach|Malignant tumor of lesser curve of stomach
C0153423|T191|SY|269460009|SNOMEDCT_CORE|Ca greater curvature - stomach|Malignant tumor of greater curve of stomach
C0153423|T191|PT|269460009|SNOMEDCT_CORE|Malignant tumor of greater curve of stomach|Malignant tumor of greater curve of stomach
C0153423|T191|FN|269460009|SNOMEDCT_CORE|Malignant tumor of greater curve of stomach|Malignant tumor of greater curve of stomach
C0153423|T191|PTGB|269460009|SNOMEDCT_CORE|Malignant tumour of greater curve of stomach|Malignant tumor of greater curve of stomach
C0153433|T191|SY|363407001|SNOMEDCT_CORE|Ca hepatic flexure - colon|Malignant tumor of hepatic flexure
C0153433|T191|SY|363407001|SNOMEDCT_CORE|Hepatic flexure colon cancer|Malignant tumor of hepatic flexure
C0153433|T191|PT|363407001|SNOMEDCT_CORE|Malignant tumor of hepatic flexure|Malignant tumor of hepatic flexure
C0153433|T191|FN|363407001|SNOMEDCT_CORE|Malignant tumor of hepatic flexure|Malignant tumor of hepatic flexure
C0153433|T191|PTGB|363407001|SNOMEDCT_CORE|Malignant tumour of hepatic flexure|Malignant tumor of hepatic flexure
C0153434|T191|SY|363408006|SNOMEDCT_CORE|Ca transverse colon|Malignant tumor of transverse colon
C0153434|T191|PT|363408006|SNOMEDCT_CORE|Malignant tumor of transverse colon|Malignant tumor of transverse colon
C0153434|T191|FN|363408006|SNOMEDCT_CORE|Malignant tumor of transverse colon|Malignant tumor of transverse colon
C0153434|T191|PTGB|363408006|SNOMEDCT_CORE|Malignant tumour of transverse colon|Malignant tumor of transverse colon
C0153434|T191|SY|363408006|SNOMEDCT_CORE|Transverse colon cancer|Malignant tumor of transverse colon
C0153435|T191|IS|363409003|SNOMEDCT_CORE|Ca descending colon|Malignant tumor of descending colon
C0153435|T191|SY|363409003|SNOMEDCT_CORE|Descending colon cancer|Malignant tumor of descending colon
C0153435|T191|PT|363409003|SNOMEDCT_CORE|Malignant tumor of descending colon|Malignant tumor of descending colon
C0153435|T191|FN|363409003|SNOMEDCT_CORE|Malignant tumor of descending colon|Malignant tumor of descending colon
C0153435|T191|PTGB|363409003|SNOMEDCT_CORE|Malignant tumour of descending colon|Malignant tumor of descending colon
C0153436|T191|IS|363410008|SNOMEDCT_CORE|Ca sigmoid colon|Malignant tumor of sigmoid colon
C0153436|T191|PT|363410008|SNOMEDCT_CORE|Malignant tumor of sigmoid colon|Malignant tumor of sigmoid colon
C0153436|T191|FN|363410008|SNOMEDCT_CORE|Malignant tumor of sigmoid colon|Malignant tumor of sigmoid colon
C0153436|T191|PTGB|363410008|SNOMEDCT_CORE|Malignant tumour of sigmoid colon|Malignant tumor of sigmoid colon
C0153436|T191|SY|363410008|SNOMEDCT_CORE|Sigmoid colon cancer|Malignant tumor of sigmoid colon
C0153437|T191|SYGB|363350007|SNOMEDCT_CORE|CA - Cancer of caecum|Malignant tumor of cecum
C0153437|T191|SY|363350007|SNOMEDCT_CORE|CA - Cancer of cecum|Malignant tumor of cecum
C0153437|T191|SYGB|363350007|SNOMEDCT_CORE|Cancer of caecum|Malignant tumor of cecum
C0153437|T191|SY|363350007|SNOMEDCT_CORE|Cancer of cecum|Malignant tumor of cecum
C0153437|T191|SY|363350007|SNOMEDCT_CORE|Cecal cancer|Malignant tumor of cecum
C0153437|T191|SYGB|363350007|SNOMEDCT_CORE|Malignant neoplasm of caecum|Malignant tumor of cecum
C0153437|T191|SY|363350007|SNOMEDCT_CORE|Malignant neoplasm of cecum|Malignant tumor of cecum
C0153437|T191|PT|363350007|SNOMEDCT_CORE|Malignant tumor of cecum|Malignant tumor of cecum
C0153437|T191|FN|363350007|SNOMEDCT_CORE|Malignant tumor of cecum|Malignant tumor of cecum
C0153437|T191|PTGB|363350007|SNOMEDCT_CORE|Malignant tumour of caecum|Malignant tumor of cecum
C0153439|T191|SY|363412000|SNOMEDCT_CORE|Ascending colon cancer|Malignant tumor of ascending colon
C0153439|T191|IS|363412000|SNOMEDCT_CORE|Ca ascending colon|Malignant tumor of ascending colon
C0153439|T191|PT|363412000|SNOMEDCT_CORE|Malignant tumor of ascending colon|Malignant tumor of ascending colon
C0153439|T191|FN|363412000|SNOMEDCT_CORE|Malignant tumor of ascending colon|Malignant tumor of ascending colon
C0153439|T191|PTGB|363412000|SNOMEDCT_CORE|Malignant tumour of ascending colon|Malignant tumor of ascending colon
C0153440|T191|SY|363413005|SNOMEDCT_CORE|Ca splenic flexure - colon|Malignant tumor of splenic flexure
C0153440|T191|PT|363413005|SNOMEDCT_CORE|Malignant tumor of splenic flexure|Malignant tumor of splenic flexure
C0153440|T191|FN|363413005|SNOMEDCT_CORE|Malignant tumor of splenic flexure|Malignant tumor of splenic flexure
C0153440|T191|PTGB|363413005|SNOMEDCT_CORE|Malignant tumour of splenic flexure|Malignant tumor of splenic flexure
C0153440|T191|SY|363413005|SNOMEDCT_CORE|Splenic flexure colon cancer|Malignant tumor of splenic flexure
C0153443|T191|IS|363414004|SNOMEDCT_CORE|Ca rectosigmoid junction|Malignant tumor of rectosigmoid junction
C0153443|T191|IS|93980002|SNOMEDCT_CORE|Malignant neoplasm of rectosigmoid junction|Malignant tumor of rectosigmoid junction
C0153443|T191|PT|363414004|SNOMEDCT_CORE|Malignant tumor of rectosigmoid junction|Malignant tumor of rectosigmoid junction
C0153443|T191|FN|363414004|SNOMEDCT_CORE|Malignant tumor of rectosigmoid junction|Malignant tumor of rectosigmoid junction
C0153443|T191|PTGB|363414004|SNOMEDCT_CORE|Malignant tumour of rectosigmoid junction|Malignant tumor of rectosigmoid junction
C0153443|T191|SY|363414004|SNOMEDCT_CORE|Rectosigmoid colon cancer|Malignant tumor of rectosigmoid junction
C0153445|T191|SY|363352004|SNOMEDCT_CORE|Cancer of anal canal|Malignant tumor of anal canal
C0153445|T191|PT|363352004|SNOMEDCT_CORE|Malignant tumor of anal canal|Malignant tumor of anal canal
C0153445|T191|FN|363352004|SNOMEDCT_CORE|Malignant tumor of anal canal|Malignant tumor of anal canal
C0153445|T191|PTGB|363352004|SNOMEDCT_CORE|Malignant tumour of anal canal|Malignant tumor of anal canal
C0153452|T191|SY|363353009|SNOMEDCT_CORE|Gallbladder Ca|Malignant tumor of gallbladder
C0153452|T191|PT|363353009|SNOMEDCT_CORE|Malignant tumor of gallbladder|Malignant tumor of gallbladder
C0153452|T191|FN|363353009|SNOMEDCT_CORE|Malignant tumor of gallbladder|Malignant tumor of gallbladder
C0153452|T191|PTGB|363353009|SNOMEDCT_CORE|Malignant tumour of gallbladder|Malignant tumor of gallbladder
C0153458|T191|SY|363419009|SNOMEDCT_CORE|Ca head of pancreas|Malignant tumor of head of pancreas
C0153458|T191|PT|363419009|SNOMEDCT_CORE|Malignant tumor of head of pancreas|Malignant tumor of head of pancreas
C0153458|T191|FN|363419009|SNOMEDCT_CORE|Malignant tumor of head of pancreas|Malignant tumor of head of pancreas
C0153458|T191|PTGB|363419009|SNOMEDCT_CORE|Malignant tumour of head of pancreas|Malignant tumor of head of pancreas
C0153459|T191|SY|187791002|SNOMEDCT_CORE|Ca body of pancreas|Malignant tumor of body of pancreas
C0153459|T191|SY|187791002|SNOMEDCT_CORE|Malignant neoplasm of body of pancreas|Malignant tumor of body of pancreas
C0153459|T191|PT|187791002|SNOMEDCT_CORE|Malignant tumor of body of pancreas|Malignant tumor of body of pancreas
C0153459|T191|FN|187791002|SNOMEDCT_CORE|Malignant tumor of body of pancreas|Malignant tumor of body of pancreas
C0153459|T191|PTGB|187791002|SNOMEDCT_CORE|Malignant tumour of body of pancreas|Malignant tumor of body of pancreas
C0153460|T191|SY|187792009|SNOMEDCT_CORE|Ca tail of pancreas|Malignant tumor of tail of pancreas
C0153460|T191|SY|187792009|SNOMEDCT_CORE|Malignant neoplasm of tail of pancreas|Malignant tumor of tail of pancreas
C0153460|T191|PT|187792009|SNOMEDCT_CORE|Malignant tumor of tail of pancreas|Malignant tumor of tail of pancreas
C0153460|T191|FN|187792009|SNOMEDCT_CORE|Malignant tumor of tail of pancreas|Malignant tumor of tail of pancreas
C0153460|T191|PTGB|187792009|SNOMEDCT_CORE|Malignant tumour of tail of pancreas|Malignant tumor of tail of pancreas
C0153461|T191|SY|187793004|SNOMEDCT_CORE|Malignant neoplasm of pancreatic duct|Malignant tumor of pancreatic duct
C0153461|T191|PT|187793004|SNOMEDCT_CORE|Malignant tumor of pancreatic duct|Malignant tumor of pancreatic duct
C0153461|T191|FN|187793004|SNOMEDCT_CORE|Malignant tumor of pancreatic duct|Malignant tumor of pancreatic duct
C0153461|T191|PTGB|187793004|SNOMEDCT_CORE|Malignant tumour of pancreatic duct|Malignant tumor of pancreatic duct
C0153467|T191|SY|363492001|SNOMEDCT_CORE|CA - Cancer of peritoneum|Malignant tumor of peritoneum
C0153467|T191|SY|363492001|SNOMEDCT_CORE|Cancer of peritoneum|Malignant tumor of peritoneum
C0153467|T191|PT|363492001|SNOMEDCT_CORE|Malignant tumor of peritoneum|Malignant tumor of peritoneum
C0153467|T191|FN|363492001|SNOMEDCT_CORE|Malignant tumor of peritoneum|Malignant tumor of peritoneum
C0153467|T191|PTGB|363492001|SNOMEDCT_CORE|Malignant tumour of peritoneum|Malignant tumor of peritoneum
C0153467|T191|SY|363492001|SNOMEDCT_CORE|Peritoneal cancer|Malignant tumor of peritoneum
C0153476|T191|SY|363425008|SNOMEDCT_CORE|Malignant tumor of maxillary antrum|Malignant tumor of maxillary sinus
C0153476|T191|PT|363425008|SNOMEDCT_CORE|Malignant tumor of maxillary sinus|Malignant tumor of maxillary sinus
C0153476|T191|FN|363425008|SNOMEDCT_CORE|Malignant tumor of maxillary sinus|Malignant tumor of maxillary sinus
C0153476|T191|SYGB|363425008|SNOMEDCT_CORE|Malignant tumour of maxillary antrum|Malignant tumor of maxillary sinus
C0153476|T191|PTGB|363425008|SNOMEDCT_CORE|Malignant tumour of maxillary sinus|Malignant tumor of maxillary sinus
C0153483|T191|SY|187841006|SNOMEDCT_CORE|Ca larynx - glottis|Malignant tumor of glottis
C0153483|T191|IS|187841006|SNOMEDCT_CORE|Ca larynx - glottis|Malignant tumor of glottis
C0153483|T191|SY|187841006|SNOMEDCT_CORE|Malignant neoplasm of glottis|Malignant tumor of glottis
C0153483|T191|PT|187841006|SNOMEDCT_CORE|Malignant tumor of glottis|Malignant tumor of glottis
C0153483|T191|FN|187841006|SNOMEDCT_CORE|Malignant tumor of glottis|Malignant tumor of glottis
C0153483|T191|PTGB|187841006|SNOMEDCT_CORE|Malignant tumour of glottis|Malignant tumor of glottis
C0153484|T191|SY|187842004|SNOMEDCT_CORE|Ca larynx - supraglottis|Malignant tumor of supraglottis
C0153484|T191|SY|187842004|SNOMEDCT_CORE|Malignant neoplasm of supraglottis|Malignant tumor of supraglottis
C0153484|T191|PT|187842004|SNOMEDCT_CORE|Malignant tumor of supraglottis|Malignant tumor of supraglottis
C0153484|T191|FN|187842004|SNOMEDCT_CORE|Malignant tumor of supraglottis|Malignant tumor of supraglottis
C0153484|T191|PTGB|187842004|SNOMEDCT_CORE|Malignant tumour of supraglottis|Malignant tumor of supraglottis
C0153504|T191|SY|363494000|SNOMEDCT_CORE|Malignant mediastinal tumor|Malignant tumor of mediastinum
C0153504|T191|SYGB|363494000|SNOMEDCT_CORE|Malignant mediastinal tumour|Malignant tumor of mediastinum
C0153504|T191|SY|363494000|SNOMEDCT_CORE|Malignant neoplasm of mediastinum|Malignant tumor of mediastinum
C0153504|T191|PT|363494000|SNOMEDCT_CORE|Malignant tumor of mediastinum|Malignant tumor of mediastinum
C0153504|T191|FN|363494000|SNOMEDCT_CORE|Malignant tumor of mediastinum|Malignant tumor of mediastinum
C0153504|T191|PTGB|363494000|SNOMEDCT_CORE|Malignant tumour of mediastinum|Malignant tumor of mediastinum
C0153549|T191|PT|188151006|SNOMEDCT_CORE|Malignant neoplasm of central part of female breast|Malignant neoplasm of central part of female breast
C0153549|T191|FN|188151006|SNOMEDCT_CORE|Malignant neoplasm of central part of female breast|Malignant neoplasm of central part of female breast
C0153550|T191|PT|188152004|SNOMEDCT_CORE|Malignant neoplasm of upper-inner quadrant of female breast|Malignant neoplasm of upper-inner quadrant of female breast
C0153550|T191|FN|188152004|SNOMEDCT_CORE|Malignant neoplasm of upper-inner quadrant of female breast|Malignant neoplasm of upper-inner quadrant of female breast
C0153551|T191|PT|188153009|SNOMEDCT_CORE|Malignant neoplasm of lower-inner quadrant of female breast|Malignant neoplasm of lower-inner quadrant of female breast
C0153551|T191|FN|188153009|SNOMEDCT_CORE|Malignant neoplasm of lower-inner quadrant of female breast|Malignant neoplasm of lower-inner quadrant of female breast
C0153552|T191|PT|188154003|SNOMEDCT_CORE|Malignant neoplasm of upper-outer quadrant of female breast|Malignant neoplasm of upper-outer quadrant of female breast
C0153552|T191|FN|188154003|SNOMEDCT_CORE|Malignant neoplasm of upper-outer quadrant of female breast|Malignant neoplasm of upper-outer quadrant of female breast
C0153553|T191|PT|188155002|SNOMEDCT_CORE|Malignant neoplasm of lower-outer quadrant of female breast|Malignant neoplasm of lower-outer quadrant of female breast
C0153553|T191|FN|188155002|SNOMEDCT_CORE|Malignant neoplasm of lower-outer quadrant of female breast|Malignant neoplasm of lower-outer quadrant of female breast
C0153567|T191|SY|371973000|SNOMEDCT_CORE|CA - Cancer of uterus|Malignant neoplasm of uterus
C0153567|T191|SY|371973000|SNOMEDCT_CORE|Cancer of uterus|Malignant neoplasm of uterus
C0153567|T191|PT|371973000|SNOMEDCT_CORE|Malignant neoplasm of uterus|Malignant neoplasm of uterus
C0153567|T191|FN|371973000|SNOMEDCT_CORE|Malignant neoplasm of uterus|Malignant neoplasm of uterus
C0153567|T191|SY|371973000|SNOMEDCT_CORE|Malignant tumor of uterus|Malignant neoplasm of uterus
C0153567|T191|SYGB|371973000|SNOMEDCT_CORE|Malignant tumour of uterus|Malignant neoplasm of uterus
C0153567|T191|SY|371973000|SNOMEDCT_CORE|Uterine cancer|Malignant neoplasm of uterus
C0153594|T191|PT|363449006|SNOMEDCT_CORE|Malignant tumor of testis|Malignant tumor of testis
C0153594|T191|FN|363449006|SNOMEDCT_CORE|Malignant tumor of testis|Malignant tumor of testis
C0153594|T191|PTGB|363449006|SNOMEDCT_CORE|Malignant tumour of testis|Malignant tumor of testis
C0153601|T191|SY|363516004|SNOMEDCT_CORE|CA - Cancer of penis|Malignant tumor of penis
C0153601|T191|SY|363516004|SNOMEDCT_CORE|Ca penis|Malignant tumor of penis
C0153601|T191|SY|363516004|SNOMEDCT_CORE|Cancer of penis|Malignant tumor of penis
C0153601|T191|PT|363516004|SNOMEDCT_CORE|Malignant tumor of penis|Malignant tumor of penis
C0153601|T191|FN|363516004|SNOMEDCT_CORE|Malignant tumor of penis|Malignant tumor of penis
C0153601|T191|PTGB|363516004|SNOMEDCT_CORE|Malignant tumour of penis|Malignant tumor of penis
C0153601|T191|SY|363516004|SNOMEDCT_CORE|Penile Ca|Malignant tumor of penis
C0153612|T191|PT|188243001|SNOMEDCT_CORE|Malignant neoplasm of posterior wall of urinary bladder|Malignant neoplasm of posterior wall of urinary bladder
C0153612|T191|FN|188243001|SNOMEDCT_CORE|Malignant neoplasm of posterior wall of urinary bladder|Malignant neoplasm of posterior wall of urinary bladder
C0153618|T191|PT|363457009|SNOMEDCT_CORE|Malignant tumor of renal pelvis|Malignant tumor of renal pelvis
C0153618|T191|FN|363457009|SNOMEDCT_CORE|Malignant tumor of renal pelvis|Malignant tumor of renal pelvis
C0153618|T191|PTGB|363457009|SNOMEDCT_CORE|Malignant tumour of renal pelvis|Malignant tumor of renal pelvis
C0153619|T191|SY|363458004|SNOMEDCT_CORE|Cancer of ureter|Malignant tumor of ureter
C0153619|T191|PT|363458004|SNOMEDCT_CORE|Malignant tumor of ureter|Malignant tumor of ureter
C0153619|T191|FN|363458004|SNOMEDCT_CORE|Malignant tumor of ureter|Malignant tumor of ureter
C0153619|T191|PTGB|363458004|SNOMEDCT_CORE|Malignant tumour of ureter|Malignant tumor of ureter
C0153619|T191|SY|363458004|SNOMEDCT_CORE|Ureter Ca|Malignant tumor of ureter
C0153620|T191|PT|363459007|SNOMEDCT_CORE|Malignant tumor of urethra|Malignant tumor of urethra
C0153620|T191|FN|363459007|SNOMEDCT_CORE|Malignant tumor of urethra|Malignant tumor of urethra
C0153620|T191|PTGB|363459007|SNOMEDCT_CORE|Malignant tumour of urethra|Malignant tumor of urethra
C0153620|T191|SY|363459007|SNOMEDCT_CORE|Malignant urethral tumor|Malignant tumor of urethra
C0153620|T191|SYGB|363459007|SNOMEDCT_CORE|Malignant urethral tumour|Malignant tumor of urethra
C0153633|T191|PT|428061005|SNOMEDCT_CORE|Malignant neoplasm of brain|Malignant neoplasm of brain
C0153633|T191|FN|428061005|SNOMEDCT_CORE|Malignant neoplasm of brain|Malignant neoplasm of brain
C0153646|T191|PT|363475005|SNOMEDCT_CORE|Malignant tumor of spinal cord|Malignant tumor of spinal cord
C0153646|T191|FN|363475005|SNOMEDCT_CORE|Malignant tumor of spinal cord|Malignant tumor of spinal cord
C0153646|T191|PTGB|363475005|SNOMEDCT_CORE|Malignant tumour of spinal cord|Malignant tumor of spinal cord
C0153660|T191|OAP|188353002|SNOMEDCT_CORE|Malignant neoplasm of head, neck and face|Malignant neoplasm of head, neck and face
C0153660|T191|OAF|188353002|SNOMEDCT_CORE|Malignant neoplasm of head, neck and face|Malignant neoplasm of head, neck and face
C0153676|T191|SY|94391008|SNOMEDCT_CORE|Cancer metastatic to lung|Secondary malignant neoplasm of lung
C0153676|T191|SY|94391008|SNOMEDCT_CORE|Metastatic malignant neoplasm to lung|Secondary malignant neoplasm of lung
C0153676|T191|IS|94391008|SNOMEDCT_CORE|Metastatic malignant neoplasm to lung, NOS|Secondary malignant neoplasm of lung
C0153676|T191|SY|94391008|SNOMEDCT_CORE|Pulmonary metastasis|Secondary malignant neoplasm of lung
C0153676|T191|SY|94391008|SNOMEDCT_CORE|Secondary cancer of lung|Secondary malignant neoplasm of lung
C0153676|T191|PT|94391008|SNOMEDCT_CORE|Secondary malignant neoplasm of lung|Secondary malignant neoplasm of lung
C0153676|T191|FN|94391008|SNOMEDCT_CORE|Secondary malignant neoplasm of lung|Secondary malignant neoplasm of lung
C0153676|T191|IS|94391008|SNOMEDCT_CORE|Secondary malignant neoplasm of lung, NOS|Secondary malignant neoplasm of lung
C0153676|T191|SY|94391008|SNOMEDCT_CORE|Secondary malignant tumor of lung|Secondary malignant neoplasm of lung
C0153676|T191|SYGB|94391008|SNOMEDCT_CORE|Secondary malignant tumour of lung|Secondary malignant neoplasm of lung
C0153677|T191|SY|94409002|SNOMEDCT_CORE|Cancer metastatic to mediastinum|Secondary malignant neoplasm of mediastinum
C0153677|T191|SY|94409002|SNOMEDCT_CORE|Mediastinal metastasis|Secondary malignant neoplasm of mediastinum
C0153677|T191|SY|94409002|SNOMEDCT_CORE|Metastasis to mediastinum|Secondary malignant neoplasm of mediastinum
C0153677|T191|SY|94409002|SNOMEDCT_CORE|Metastatic malignant neoplasm to mediastinum|Secondary malignant neoplasm of mediastinum
C0153677|T191|IS|94409002|SNOMEDCT_CORE|Metastatic malignant neoplasm to mediastinum, NOS|Secondary malignant neoplasm of mediastinum
C0153677|T191|PT|94409002|SNOMEDCT_CORE|Secondary malignant neoplasm of mediastinum|Secondary malignant neoplasm of mediastinum
C0153677|T191|FN|94409002|SNOMEDCT_CORE|Secondary malignant neoplasm of mediastinum|Secondary malignant neoplasm of mediastinum
C0153677|T191|IS|94409002|SNOMEDCT_CORE|Secondary malignant neoplasm of mediastinum, NOS|Secondary malignant neoplasm of mediastinum
C0153677|T191|SY|94409002|SNOMEDCT_CORE|Secondary malignant tumor of mediastinum|Secondary malignant neoplasm of mediastinum
C0153677|T191|SYGB|94409002|SNOMEDCT_CORE|Secondary malignant tumour of mediastinum|Secondary malignant neoplasm of mediastinum
C0153678|T191|SY|94493005|SNOMEDCT_CORE|Cancer metastatic to pleura|Secondary malignant neoplasm of pleura
C0153678|T191|SY|94493005|SNOMEDCT_CORE|Metastasis to pleura|Secondary malignant neoplasm of pleura
C0153678|T191|SY|94493005|SNOMEDCT_CORE|Metastatic malignant neoplasm to pleura|Secondary malignant neoplasm of pleura
C0153678|T191|IS|94493005|SNOMEDCT_CORE|Metastatic malignant neoplasm to pleura, NOS|Secondary malignant neoplasm of pleura
C0153678|T191|SY|94493005|SNOMEDCT_CORE|Pleural seedling|Secondary malignant neoplasm of pleura
C0153678|T191|PT|94493005|SNOMEDCT_CORE|Secondary malignant neoplasm of pleura|Secondary malignant neoplasm of pleura
C0153678|T191|FN|94493005|SNOMEDCT_CORE|Secondary malignant neoplasm of pleura|Secondary malignant neoplasm of pleura
C0153678|T191|IS|94493005|SNOMEDCT_CORE|Secondary malignant neoplasm of pleura, NOS|Secondary malignant neoplasm of pleura
C0153678|T191|SY|94493005|SNOMEDCT_CORE|Secondary malignant tumor of pleura|Secondary malignant neoplasm of pleura
C0153678|T191|SYGB|94493005|SNOMEDCT_CORE|Secondary malignant tumour of pleura|Secondary malignant neoplasm of pleura
C0153685|T191|SY|94360002|SNOMEDCT_CORE|Cancer metastatic to kidney|Secondary malignant neoplasm of kidney
C0153685|T191|SY|94360002|SNOMEDCT_CORE|Metastasis to renal parenchyma|Secondary malignant neoplasm of kidney
C0153685|T191|SY|94360002|SNOMEDCT_CORE|Metastatic malignant neoplasm to kidney|Secondary malignant neoplasm of kidney
C0153685|T191|IS|94360002|SNOMEDCT_CORE|Metastatic malignant neoplasm to kidney, NOS|Secondary malignant neoplasm of kidney
C0153685|T191|SY|94360002|SNOMEDCT_CORE|Metastatic tumor in kidney|Secondary malignant neoplasm of kidney
C0153685|T191|SYGB|94360002|SNOMEDCT_CORE|Metastatic tumour in kidney|Secondary malignant neoplasm of kidney
C0153685|T191|SY|94360002|SNOMEDCT_CORE|Renal metastasis|Secondary malignant neoplasm of kidney
C0153685|T191|SY|94360002|SNOMEDCT_CORE|Secondary cancer of kidney|Secondary malignant neoplasm of kidney
C0153685|T191|PT|94360002|SNOMEDCT_CORE|Secondary malignant neoplasm of kidney|Secondary malignant neoplasm of kidney
C0153685|T191|FN|94360002|SNOMEDCT_CORE|Secondary malignant neoplasm of kidney|Secondary malignant neoplasm of kidney
C0153685|T191|IS|94360002|SNOMEDCT_CORE|Secondary malignant neoplasm of kidney, NOS|Secondary malignant neoplasm of kidney
C0153685|T191|SY|94360002|SNOMEDCT_CORE|Secondary renal cancer|Secondary malignant neoplasm of kidney
C0153687|T191|SY|94579000|SNOMEDCT_CORE|Cancer metastatic to skin|Secondary malignant neoplasm of skin
C0153687|T191|SY|94579000|SNOMEDCT_CORE|Cutaneous metastasis|Secondary malignant neoplasm of skin
C0153687|T191|SY|94579000|SNOMEDCT_CORE|Dermal metastasis|Secondary malignant neoplasm of skin
C0153687|T191|SY|94579000|SNOMEDCT_CORE|Malignant infiltration of skin|Secondary malignant neoplasm of skin
C0153687|T191|SY|94579000|SNOMEDCT_CORE|Metastasis to skin|Secondary malignant neoplasm of skin
C0153687|T191|SY|94579000|SNOMEDCT_CORE|Metastatic malignant neoplasm to skin|Secondary malignant neoplasm of skin
C0153687|T191|IS|94579000|SNOMEDCT_CORE|Metastatic malignant neoplasm to skin, NOS|Secondary malignant neoplasm of skin
C0153687|T191|SY|94579000|SNOMEDCT_CORE|Secondary cancer of skin|Secondary malignant neoplasm of skin
C0153687|T191|PT|94579000|SNOMEDCT_CORE|Secondary malignant neoplasm of skin|Secondary malignant neoplasm of skin
C0153687|T191|FN|94579000|SNOMEDCT_CORE|Secondary malignant neoplasm of skin|Secondary malignant neoplasm of skin
C0153687|T191|IS|94579000|SNOMEDCT_CORE|Secondary malignant neoplasm of skin, NOS|Secondary malignant neoplasm of skin
C0153687|T191|SY|94579000|SNOMEDCT_CORE|Skin secondaries|Secondary malignant neoplasm of skin
C0153688|T191|PT|188462001|SNOMEDCT_CORE|Secondary malignant neoplasm of brain and spinal cord|Secondary malignant neoplasm of brain and spinal cord
C0153688|T191|FN|188462001|SNOMEDCT_CORE|Secondary malignant neoplasm of brain and spinal cord|Secondary malignant neoplasm of brain and spinal cord
C0153690|T191|SY|94222008|SNOMEDCT_CORE|Bony metastasis|Secondary malignant neoplasm of bone
C0153690|T191|SY|94222008|SNOMEDCT_CORE|Cancer metastatic to bone|Secondary malignant neoplasm of bone
C0153690|T191|SY|94222008|SNOMEDCT_CORE|Metastatic malignant neoplasm to bone|Secondary malignant neoplasm of bone
C0153690|T191|IS|94222008|SNOMEDCT_CORE|Metastatic malignant neoplasm to bone, NOS|Secondary malignant neoplasm of bone
C0153690|T191|SY|94222008|SNOMEDCT_CORE|Metastatic tumor of bone|Secondary malignant neoplasm of bone
C0153690|T191|SYGB|94222008|SNOMEDCT_CORE|Metastatic tumour of bone|Secondary malignant neoplasm of bone
C0153690|T191|SY|94222008|SNOMEDCT_CORE|Osseous metastasis|Secondary malignant neoplasm of bone
C0153690|T191|SY|94222008|SNOMEDCT_CORE|Secondary cancer of bone|Secondary malignant neoplasm of bone
C0153690|T191|PT|94222008|SNOMEDCT_CORE|Secondary malignant neoplasm of bone|Secondary malignant neoplasm of bone
C0153690|T191|FN|94222008|SNOMEDCT_CORE|Secondary malignant neoplasm of bone|Secondary malignant neoplasm of bone
C0153690|T191|SY|94222008|SNOMEDCT_CORE|Secondary malignant neoplasm of bone and bone marrow|Secondary malignant neoplasm of bone
C0153690|T191|IS|94222008|SNOMEDCT_CORE|Secondary malignant neoplasm of bone, NOS|Secondary malignant neoplasm of bone
C0153690|T191|SY|94222008|SNOMEDCT_CORE|Tumor metastatic to bone|Secondary malignant neoplasm of bone
C0153690|T191|SYGB|94222008|SNOMEDCT_CORE|Tumour metastatic to bone|Secondary malignant neoplasm of bone
C0153691|T191|SY|94161006|SNOMEDCT_CORE|Cancer metastatic to adrenal gland|Secondary malignant neoplasm of adrenal gland
C0153691|T191|SY|94161006|SNOMEDCT_CORE|Metastasis to adrenal gland|Secondary malignant neoplasm of adrenal gland
C0153691|T191|SY|94161006|SNOMEDCT_CORE|Metastatic malignant neoplasm to adrenal gland|Secondary malignant neoplasm of adrenal gland
C0153691|T191|PT|94161006|SNOMEDCT_CORE|Secondary malignant neoplasm of adrenal gland|Secondary malignant neoplasm of adrenal gland
C0153691|T191|FN|94161006|SNOMEDCT_CORE|Secondary malignant neoplasm of adrenal gland|Secondary malignant neoplasm of adrenal gland
C0153691|T191|SY|94161006|SNOMEDCT_CORE|Suprarenal metastasis|Secondary malignant neoplasm of adrenal gland
C0153711|T191|PT|188507008|SNOMEDCT_CORE|Lymphosarcoma of lymph nodes of multiple sites|Lymphosarcoma of lymph nodes of multiple sites
C0153711|T191|FN|188507008|SNOMEDCT_CORE|Lymphosarcoma of lymph nodes of multiple sites|Lymphosarcoma of lymph nodes of multiple sites
C0153801|T191|PT|95192000|SNOMEDCT_CORE|Nodular lymphoma of lymph nodes of multiple sites|Nodular lymphoma of lymph nodes of multiple sites
C0153801|T191|FN|95192000|SNOMEDCT_CORE|Nodular lymphoma of lymph nodes of multiple sites|Nodular lymphoma of lymph nodes of multiple sites
C0153817|T191|SY|188637007|SNOMEDCT_CORE|Sézary disease of lymph nodes of multiple sites|Sézary's disease of lymph nodes of multiple sites
C0153817|T191|PT|188637007|SNOMEDCT_CORE|Sézary's disease of lymph nodes of multiple sites|Sézary's disease of lymph nodes of multiple sites
C0153817|T191|SY|188637007|SNOMEDCT_CORE|Sezary's disease of lymph nodes of multiple sites|Sézary's disease of lymph nodes of multiple sites
C0153817|T191|FN|188637007|SNOMEDCT_CORE|Sézary's disease of lymph nodes of multiple sites|Sézary's disease of lymph nodes of multiple sites
C0153817|T191|OF|188637007|SNOMEDCT_CORE|Sezary's disease of lymph nodes of multiple sites|Sézary's disease of lymph nodes of multiple sites
C0153869|T191|PT|94704006|SNOMEDCT_CORE|Multiple myeloma in remission|Multiple myeloma in remission
C0153869|T191|FN|94704006|SNOMEDCT_CORE|Multiple myeloma in remission|Multiple myeloma in remission
C0153875|T191|IS|91857003|SNOMEDCT_CORE|Acute lymphoid leukemia without mention of remission|Acute lymphoid leukemia without mention of remission
C0153876|T191|PTGB|91856007|SNOMEDCT_CORE|Acute lymphoid leukaemia in remission|Acute lymphoid leukemia in remission
C0153876|T191|PT|91856007|SNOMEDCT_CORE|Acute lymphoid leukemia in remission|Acute lymphoid leukemia in remission
C0153876|T191|FN|91856007|SNOMEDCT_CORE|Acute lymphoid leukemia in remission|Acute lymphoid leukemia in remission
C0153877|T191|IS|92814006|SNOMEDCT_CORE|Chronic lymphoid leukemia without mention of remission|Chronic lymphoid leukemia without mention of remission
C0153878|T191|PTGB|92813000|SNOMEDCT_CORE|Chronic lymphoid leukaemia in remission|Chronic lymphoid leukemia in remission
C0153878|T191|PT|92813000|SNOMEDCT_CORE|Chronic lymphoid leukemia in remission|Chronic lymphoid leukemia in remission
C0153878|T191|FN|92813000|SNOMEDCT_CORE|Chronic lymphoid leukemia in remission|Chronic lymphoid leukemia in remission
C0153885|T191|IS|91861009|SNOMEDCT_CORE|Acute myeloid leukemia without mention of remission|Acute myeloid leukemia without mention of remission
C0153886|T191|PTGB|91860005|SNOMEDCT_CORE|Acute myeloid leukaemia in remission|Acute myeloid leukemia in remission
C0153886|T191|PT|91860005|SNOMEDCT_CORE|Acute myeloid leukemia in remission|Acute myeloid leukemia in remission
C0153886|T191|FN|91860005|SNOMEDCT_CORE|Acute myeloid leukemia in remission|Acute myeloid leukemia in remission
C0153887|T191|IS|92818009|SNOMEDCT_CORE|Chronic myeloid leukemia without mention of remission|Chronic myeloid leukemia without mention of remission
C0153972|T191|PT|93162007|SNOMEDCT_CORE|Lipoma of spermatic cord|Lipoma of spermatic cord
C0153972|T191|FN|93162007|SNOMEDCT_CORE|Lipoma of spermatic cord|Lipoma of spermatic cord
C0153982|T191|PT|92369000|SNOMEDCT_CORE|Benign neoplasm of skin of lip|Benign neoplasm of skin of lip
C0153982|T191|FN|92369000|SNOMEDCT_CORE|Benign neoplasm of skin of lip|Benign neoplasm of skin of lip
C0153983|T191|OAP|189053003|SNOMEDCT_CORE|Benign neoplasm of eyelid including canthus|Benign neoplasm of eyelid including canthus
C0153983|T191|OAF|189053003|SNOMEDCT_CORE|Benign neoplasm of eyelid including canthus|Benign neoplasm of eyelid including canthus
C0153988|T191|IS|189078004|SNOMEDCT_CORE|Benign neoplasm of skin of arm|Benign neoplasm of skin of upper limb
C0153988|T191|PT|92382008|SNOMEDCT_CORE|Benign neoplasm of skin of upper limb|Benign neoplasm of skin of upper limb
C0153988|T191|FN|92382008|SNOMEDCT_CORE|Benign neoplasm of skin of upper limb|Benign neoplasm of skin of upper limb
C0153988|T191|OAP|189078004|SNOMEDCT_CORE|Benign neoplasm of skin of upper limb and shoulder|Benign neoplasm of skin of upper limb
C0153988|T191|OAF|189078004|SNOMEDCT_CORE|Benign neoplasm of skin of upper limb and shoulder|Benign neoplasm of skin of upper limb
C0153988|T191|IS|92382008|SNOMEDCT_CORE|Benign neoplasm of skin of upper limb, NOS|Benign neoplasm of skin of upper limb
C0153989|T191|SY|92370004|SNOMEDCT_CORE|Benign neoplasm of skin of hip and lower limb|Benign neoplasm of skin of hip and lower limb
C0153993|T191|PT|95279007|SNOMEDCT_CORE|Submucous leiomyoma of uterus|Submucous leiomyoma of uterus
C0153993|T191|FN|95279007|SNOMEDCT_CORE|Submucous leiomyoma of uterus|Submucous leiomyoma of uterus
C0153993|T191|SY|95279007|SNOMEDCT_CORE|Submucous uterine fibroid|Submucous leiomyoma of uterus
C0153993|T191|SY|95279007|SNOMEDCT_CORE|Submucous uterine leiomyoma|Submucous leiomyoma of uterus
C0153994|T191|SY|93616000|SNOMEDCT_CORE|Interstitial uterine fibroid|Intramural leiomyoma of uterus
C0153994|T191|PT|93616000|SNOMEDCT_CORE|Intramural leiomyoma of uterus|Intramural leiomyoma of uterus
C0153994|T191|FN|93616000|SNOMEDCT_CORE|Intramural leiomyoma of uterus|Intramural leiomyoma of uterus
C0153994|T191|SY|93616000|SNOMEDCT_CORE|Intramural uterine fibroid|Intramural leiomyoma of uterus
C0153994|T191|SY|93616000|SNOMEDCT_CORE|Intramural uterine leiomyoma|Intramural leiomyoma of uterus
C0153995|T191|PT|95280005|SNOMEDCT_CORE|Subserous leiomyoma of uterus|Subserous leiomyoma of uterus
C0153995|T191|FN|95280005|SNOMEDCT_CORE|Subserous leiomyoma of uterus|Subserous leiomyoma of uterus
C0153995|T191|SY|95280005|SNOMEDCT_CORE|Subserous uterine fibroid|Subserous leiomyoma of uterus
C0153995|T191|SY|95280005|SNOMEDCT_CORE|Subserous uterine leiomyoma|Subserous leiomyoma of uterus
C0154009|T191|PT|92308005|SNOMEDCT_CORE|Benign neoplasm of prostate|Benign neoplasm of prostate
C0154009|T191|FN|92308005|SNOMEDCT_CORE|Benign neoplasm of prostate|Benign neoplasm of prostate
C0154009|T191|SY|92308005|SNOMEDCT_CORE|Benign prostatic tumor|Benign neoplasm of prostate
C0154009|T191|SYGB|92308005|SNOMEDCT_CORE|Benign prostatic tumour|Benign neoplasm of prostate
C0154009|T191|SY|92308005|SNOMEDCT_CORE|Benign tumor of prostate|Benign neoplasm of prostate
C0154009|T191|SYGB|92308005|SNOMEDCT_CORE|Benign tumour of prostate|Benign neoplasm of prostate
C0154023|T191|PT|92258000|SNOMEDCT_CORE|Benign neoplasm of orbit|Benign neoplasm of orbit
C0154023|T191|FN|92258000|SNOMEDCT_CORE|Benign neoplasm of orbit|Benign neoplasm of orbit
C0154023|T191|SY|92258000|SNOMEDCT_CORE|Benign orbital tumor|Benign neoplasm of orbit
C0154023|T191|SYGB|92258000|SNOMEDCT_CORE|Benign orbital tumour|Benign neoplasm of orbit
C0154023|T191|SY|92258000|SNOMEDCT_CORE|Benign tumor of orbit|Benign neoplasm of orbit
C0154023|T191|SYGB|92258000|SNOMEDCT_CORE|Benign tumour of orbit|Benign neoplasm of orbit
C0154028|T191|PT|92059004|SNOMEDCT_CORE|Benign neoplasm of choroid|Benign neoplasm of choroid
C0154028|T191|FN|92059004|SNOMEDCT_CORE|Benign neoplasm of choroid|Benign neoplasm of choroid
C0154028|T191|SY|92059004|SNOMEDCT_CORE|Benign tumor of choroid|Benign neoplasm of choroid
C0154028|T191|SYGB|92059004|SNOMEDCT_CORE|Benign tumour of choroid|Benign neoplasm of choroid
C0154033|T191|PT|92051001|SNOMEDCT_CORE|Benign neoplasm of cerebral meninges|Benign neoplasm of cerebral meninges
C0154033|T191|FN|92051001|SNOMEDCT_CORE|Benign neoplasm of cerebral meninges|Benign neoplasm of cerebral meninges
C0154038|T191|PT|92439006|SNOMEDCT_CORE|Benign neoplasm of thyroid gland|Benign neoplasm of thyroid gland
C0154038|T191|FN|92439006|SNOMEDCT_CORE|Benign neoplasm of thyroid gland|Benign neoplasm of thyroid gland
C0154038|T191|SY|92439006|SNOMEDCT_CORE|Benign tumor of thyroid gland|Benign neoplasm of thyroid gland
C0154038|T191|SYGB|92439006|SNOMEDCT_CORE|Benign tumour of thyroid gland|Benign neoplasm of thyroid gland
C0154040|T191|PT|91967007|SNOMEDCT_CORE|Benign neoplasm of adrenal gland|Benign neoplasm of adrenal gland
C0154040|T191|FN|91967007|SNOMEDCT_CORE|Benign neoplasm of adrenal gland|Benign neoplasm of adrenal gland
C0154040|T191|SY|91967007|SNOMEDCT_CORE|Benign tumor of adrenal gland|Benign neoplasm of adrenal gland
C0154040|T191|SYGB|91967007|SNOMEDCT_CORE|Benign tumour of adrenal gland|Benign neoplasm of adrenal gland
C0154049|T191|PTGB|271481007|SNOMEDCT_CORE|Haemangioma of skin and subcutaneous tissue|Hemangioma of skin and subcutaneous tissue
C0154049|T191|PT|271481007|SNOMEDCT_CORE|Hemangioma of skin and subcutaneous tissue|Hemangioma of skin and subcutaneous tissue
C0154049|T191|FN|271481007|SNOMEDCT_CORE|Hemangioma of skin and subcutaneous tissue|Hemangioma of skin and subcutaneous tissue
C0154052|T191|PTGB|189197001|SNOMEDCT_CORE|Haemangioma of intra-abdominal structure|Hemangioma of intra-abdominal structure
C0154052|T191|SYGB|189197001|SNOMEDCT_CORE|Haemangioma of intra-abdominal structures|Hemangioma of intra-abdominal structure
C0154052|T191|PT|189197001|SNOMEDCT_CORE|Hemangioma of intra-abdominal structure|Hemangioma of intra-abdominal structure
C0154052|T191|FN|189197001|SNOMEDCT_CORE|Hemangioma of intra-abdominal structure|Hemangioma of intra-abdominal structure
C0154052|T191|SY|189197001|SNOMEDCT_CORE|Hemangioma of intra-abdominal structures|Hemangioma of intra-abdominal structure
C0154052|T191|OF|189197001|SNOMEDCT_CORE|Hemangioma of intra-abdominal structures|Hemangioma of intra-abdominal structure
C0154084|T191|IS|189336000|SNOMEDCT_CORE|Breast Ca in situ|Carcinoma in situ of breast
C0154084|T191|PT|189336000|SNOMEDCT_CORE|Carcinoma in situ of breast|Carcinoma in situ of breast
C0154084|T191|FN|189336000|SNOMEDCT_CORE|Carcinoma in situ of breast|Carcinoma in situ of breast
C0154084|T191|SY|189336000|SNOMEDCT_CORE|Non-invasive carcinoma of breast|Carcinoma in situ of breast
C0154091|T191|PT|92546004|SNOMEDCT_CORE|Cancer in situ of urinary bladder|Cancer in situ of urinary bladder
C0154091|T191|SY|92546004|SNOMEDCT_CORE|Carcinoma in situ of bladder|Cancer in situ of urinary bladder
C0154091|T191|FN|92546004|SNOMEDCT_CORE|Carcinoma in situ of bladder|Cancer in situ of urinary bladder
C0154091|T191|IS|92546004|SNOMEDCT_CORE|Carcinoma in situ of bladder, NOS|Cancer in situ of urinary bladder
C0154091|T191|IS|92546004|SNOMEDCT_CORE|CIS - Carcinoma in situ of bladder|Cancer in situ of urinary bladder
C0154119|T191|PT|189484008|SNOMEDCT_CORE|Neoplasm of uncertain behavior of brain and spinal cord|Neoplasm of uncertain behavior of brain and spinal cord
C0154119|T191|OF|189484008|SNOMEDCT_CORE|Neoplasm of uncertain behavior of brain and spinal cord|Neoplasm of uncertain behavior of brain and spinal cord
C0154119|T191|SY|189484008|SNOMEDCT_CORE|Neoplasm of uncertain behavior of brain and/or spinal cord|Neoplasm of uncertain behavior of brain and spinal cord
C0154119|T191|FN|189484008|SNOMEDCT_CORE|Neoplasm of uncertain behavior of brain and/or spinal cord|Neoplasm of uncertain behavior of brain and spinal cord
C0154119|T191|PTGB|189484008|SNOMEDCT_CORE|Neoplasm of uncertain behaviour of brain and spinal cord|Neoplasm of uncertain behavior of brain and spinal cord
C0154120|T191|PT|109914007|SNOMEDCT_CORE|Neoplasm of uncertain behavior of meninges|Neoplasm of uncertain behavior of meninges
C0154120|T191|FN|109914007|SNOMEDCT_CORE|Neoplasm of uncertain behavior of meninges|Neoplasm of uncertain behavior of meninges
C0154120|T191|PTGB|109914007|SNOMEDCT_CORE|Neoplasm of uncertain behaviour of meninges|Neoplasm of uncertain behavior of meninges
C0154125|T191|SY|94805002|SNOMEDCT_CORE|Neoplasm of uncertain behavior of connective and other soft tissues|Neoplasm of uncertain behavior of soft tissues
C0154125|T191|IS|94805002|SNOMEDCT_CORE|Neoplasm of uncertain behavior of connective and other soft tissues, NOS|Neoplasm of uncertain behavior of soft tissues
C0154125|T191|PT|94805002|SNOMEDCT_CORE|Neoplasm of uncertain behavior of soft tissues|Neoplasm of uncertain behavior of soft tissues
C0154125|T191|FN|94805002|SNOMEDCT_CORE|Neoplasm of uncertain behavior of soft tissues|Neoplasm of uncertain behavior of soft tissues
C0154125|T191|SYGB|94805002|SNOMEDCT_CORE|Neoplasm of uncertain behaviour of connective and other soft tissues|Neoplasm of uncertain behavior of soft tissues
C0154125|T191|PTGB|94805002|SNOMEDCT_CORE|Neoplasm of uncertain behaviour of soft tissues|Neoplasm of uncertain behavior of soft tissues
C0154143|T047|SY|26389007|SNOMEDCT_CORE|Secondary thyroid hyperplasia|Toxic multinodular goiter
C0154143|T047|SY|26389007|SNOMEDCT_CORE|Thyrotoxicosis due to multinodular goiter|Toxic multinodular goiter
C0154143|T047|SYGB|26389007|SNOMEDCT_CORE|Thyrotoxicosis due to multinodular goitre|Toxic multinodular goiter
C0154143|T047|SY|26389007|SNOMEDCT_CORE|Thyrotoxicosis with toxic multinodular goiter|Toxic multinodular goiter
C0154143|T047|SYGB|26389007|SNOMEDCT_CORE|Thyrotoxicosis with toxic multinodular goitre|Toxic multinodular goiter
C0154143|T047|PT|26389007|SNOMEDCT_CORE|Toxic multinodular goiter|Toxic multinodular goiter
C0154143|T047|FN|26389007|SNOMEDCT_CORE|Toxic multinodular goiter|Toxic multinodular goiter
C0154143|T047|PTGB|26389007|SNOMEDCT_CORE|Toxic multinodular goitre|Toxic multinodular goiter
C0154143|T047|SY|26389007|SNOMEDCT_CORE|Toxic multinodular thyroid goiter|Toxic multinodular goiter
C0154143|T047|SYGB|26389007|SNOMEDCT_CORE|Toxic multinodular thyroid goitre|Toxic multinodular goiter
C0154157|T047|SY|27059002|SNOMEDCT_CORE|Hypothyroidism after surgery|Postoperative hypothyroidism
C0154157|T047|OF|27059002|SNOMEDCT_CORE|Post-operative hypothyroidism|Postoperative hypothyroidism
C0154157|T047|IS|27059002|SNOMEDCT_CORE|Post-operative hypothyroidism|Postoperative hypothyroidism
C0154157|T047|IS|27059002|SNOMEDCT_CORE|Post-surgical hypothyroidism|Postoperative hypothyroidism
C0154157|T047|PT|27059002|SNOMEDCT_CORE|Postoperative hypothyroidism|Postoperative hypothyroidism
C0154157|T047|FN|27059002|SNOMEDCT_CORE|Postoperative hypothyroidism|Postoperative hypothyroidism
C0154157|T047|SY|27059002|SNOMEDCT_CORE|Postsurgical hypothyroidism|Postoperative hypothyroidism
C0154159|T047|PT|190279008|SNOMEDCT_CORE|Iodine hypothyroidism|Iodine hypothyroidism
C0154159|T047|FN|190279008|SNOMEDCT_CORE|Iodine hypothyroidism|Iodine hypothyroidism
C0154208|T047|PT|37102008|SNOMEDCT_CORE|Disorder of endocrine ovary|Disorder of endocrine ovary
C0154208|T047|FN|37102008|SNOMEDCT_CORE|Disorder of endocrine ovary|Disorder of endocrine ovary
C0154208|T047|IS|37102008|SNOMEDCT_CORE|Disorder of endocrine ovary, NOS|Disorder of endocrine ovary
C0154208|T047|SY|37102008|SNOMEDCT_CORE|Ovarian dysfunction|Disorder of endocrine ovary
C0154208|T047|IS|37102008|SNOMEDCT_CORE|Ovarian dysfunction, NOS|Disorder of endocrine ovary
C0154251|T047|PT|267431006|SNOMEDCT_CORE|Disorder of lipid metabolism|Disorder of lipid metabolism
C0154251|T047|FN|267431006|SNOMEDCT_CORE|Disorder of lipid metabolism|Disorder of lipid metabolism
C0154251|T047|IS|267431006|SNOMEDCT_CORE|Disorders of lipoid metabolism|Disorder of lipid metabolism
C0154251|T047|SY|267431006|SNOMEDCT_CORE|Lipid metabolism disorder|Disorder of lipid metabolism
C0154286|T047|PTGB|413533008|SNOMEDCT_CORE|Anaemia due to chronic blood loss|Anemia due to chronic blood loss
C0154286|T047|PT|413533008|SNOMEDCT_CORE|Anemia due to chronic blood loss|Anemia due to chronic blood loss
C0154286|T047|FN|413533008|SNOMEDCT_CORE|Anemia due to chronic blood loss|Anemia due to chronic blood loss
C0154286|T047|SYGB|413533008|SNOMEDCT_CORE|Chronic blood loss anaemia|Anemia due to chronic blood loss
C0154286|T047|SY|413533008|SNOMEDCT_CORE|Chronic blood loss anemia|Anemia due to chronic blood loss
C0154286|T047|SY|413533008|SNOMEDCT_CORE|Chronic hemorrhagic anemia|Anemia due to chronic blood loss
C0154286|T047|SY|413533008|SNOMEDCT_CORE|Iron deficiency anemia due to chronic blood loss|Anemia due to chronic blood loss
C0154287|T047|PTGB|371315009|SNOMEDCT_CORE|Iron deficiency anaemia secondary to inadequate dietary iron intake|Iron deficiency anemia secondary to inadequate dietary iron intake
C0154287|T047|PT|371315009|SNOMEDCT_CORE|Iron deficiency anemia secondary to inadequate dietary iron intake|Iron deficiency anemia secondary to inadequate dietary iron intake
C0154287|T047|FN|371315009|SNOMEDCT_CORE|Iron deficiency anemia secondary to inadequate dietary iron intake|Iron deficiency anemia secondary to inadequate dietary iron intake
C0154301|T047|PT|74576004|SNOMEDCT_CORE|Acquired thrombocytopenia|Acquired thrombocytopenia
C0154301|T047|FN|74576004|SNOMEDCT_CORE|Acquired thrombocytopenia|Acquired thrombocytopenia
C0154301|T047|IS|74576004|SNOMEDCT_CORE|Secondary thrombocytopenia|Acquired thrombocytopenia
C0154315|T048|SY|191461002|SNOMEDCT_CORE|Senile delirium|Senile dementia with delirium
C0154315|T048|PT|191461002|SNOMEDCT_CORE|Senile dementia with delirium|Senile dementia with delirium
C0154315|T048|FN|191461002|SNOMEDCT_CORE|Senile dementia with delirium|Senile dementia with delirium
C0154378|T048|PT|191572009|SNOMEDCT_CORE|Acute exacerbation of chronic schizoaffective schizophrenia|Acute exacerbation of chronic schizoaffective schizophrenia
C0154378|T048|FN|191572009|SNOMEDCT_CORE|Acute exacerbation of chronic schizoaffective schizophrenia|Acute exacerbation of chronic schizoaffective schizophrenia
C0154403|T048|PT|79298009|SNOMEDCT_CORE|Mild major depression, single episode|Mild major depression, single episode
C0154403|T048|FN|79298009|SNOMEDCT_CORE|Mild major depression, single episode|Mild major depression, single episode
C0154404|T048|PT|15639000|SNOMEDCT_CORE|Moderate major depression, single episode|Moderate major depression, single episode
C0154404|T048|FN|15639000|SNOMEDCT_CORE|Moderate major depression, single episode|Moderate major depression, single episode
C0154405|T048|PT|76441001|SNOMEDCT_CORE|Severe major depression, single episode, without psychotic features|Severe major depression, single episode, without psychotic features
C0154405|T048|FN|76441001|SNOMEDCT_CORE|Severe major depression, single episode, without psychotic features|Severe major depression, single episode, without psychotic features
C0154406|T048|SY|430852001|SNOMEDCT_CORE|Major depressive disorder, single episode, severe with psychotic features|Severe major depression, single episode, with psychotic features
C0154406|T048|PT|430852001|SNOMEDCT_CORE|Severe major depression, single episode, with psychotic features|Severe major depression, single episode, with psychotic features
C0154406|T048|FN|430852001|SNOMEDCT_CORE|Severe major depression, single episode, with psychotic features|Severe major depression, single episode, with psychotic features
C0154408|T048|OAF|191606003|SNOMEDCT_CORE|Single major depressive episode, in full remission|Single major depressive episode, in full remission
C0154408|T048|OAP|191606003|SNOMEDCT_CORE|Single major depressive episode, in full remission|Single major depressive episode, in full remission
C0154409|T048|PT|66344007|SNOMEDCT_CORE|Recurrent major depression|Recurrent major depressive episodes
C0154409|T048|FN|66344007|SNOMEDCT_CORE|Recurrent major depression|Recurrent major depressive episodes
C0154409|T048|IS|66344007|SNOMEDCT_CORE|Recurrent major depression, NOS|Recurrent major depressive episodes
C0154409|T048|SY|66344007|SNOMEDCT_CORE|Recurrent major depressive disorder|Recurrent major depressive episodes
C0154409|T048|IS|66344007|SNOMEDCT_CORE|Recurrent major depressive disorder, NOS|Recurrent major depressive episodes
C0154409|T048|PT|268621008|SNOMEDCT_CORE|Recurrent major depressive episodes|Recurrent major depressive episodes
C0154409|T048|FN|268621008|SNOMEDCT_CORE|Recurrent major depressive episodes|Recurrent major depressive episodes
C0154410|T048|PT|40379007|SNOMEDCT_CORE|Mild recurrent major depression|Mild recurrent major depression
C0154410|T048|FN|40379007|SNOMEDCT_CORE|Mild recurrent major depression|Mild recurrent major depression
C0154411|T048|PT|18818009|SNOMEDCT_CORE|Moderate recurrent major depression|Moderate recurrent major depression
C0154411|T048|FN|18818009|SNOMEDCT_CORE|Moderate recurrent major depression|Moderate recurrent major depression
C0154412|T048|PT|36474008|SNOMEDCT_CORE|Severe recurrent major depression without psychotic features|Severe recurrent major depression without psychotic features
C0154412|T048|FN|36474008|SNOMEDCT_CORE|Severe recurrent major depression without psychotic features|Severe recurrent major depression without psychotic features
C0154413|T048|PT|28475009|SNOMEDCT_CORE|Severe recurrent major depression with psychotic features|Severe recurrent major depression with psychotic features
C0154413|T048|FN|28475009|SNOMEDCT_CORE|Severe recurrent major depression with psychotic features|Severe recurrent major depression with psychotic features
C0154437|T048|PT|191659001|SNOMEDCT_CORE|Atypical depressive disorder|Atypical depressive disorder
C0154437|T048|FN|191659001|SNOMEDCT_CORE|Atypical depressive disorder|Atypical depressive disorder
C0154487|T048|PT|191833002|SNOMEDCT_CORE|Cocaine dependence in remission|Cocaine dependence in remission
C0154487|T048|FN|191833002|SNOMEDCT_CORE|Cocaine dependence in remission|Cocaine dependence in remission
C0154490|T047|PT|191839003|SNOMEDCT_CORE|Cannabis dependence in remission|Cannabis dependence in remission
C0154490|T047|FN|191839003|SNOMEDCT_CORE|Cannabis dependence in remission|Cannabis dependence in remission
C0154575|T048|PT|37941009|SNOMEDCT_CORE|Rumination disorder|Rumination disorder
C0154575|T048|FN|37941009|SNOMEDCT_CORE|Rumination disorder|Rumination disorder
C0154575|T048|IS|37941009|SNOMEDCT_CORE|Rumination disorder, NOS|Rumination disorder
C0154583|T048|PT|192049004|SNOMEDCT_CORE|Prolonged depressive adjustment reaction|Prolonged depressive adjustment reaction
C0154583|T048|FN|192049004|SNOMEDCT_CORE|Prolonged depressive adjustment reaction|Prolonged depressive adjustment reaction
C0154587|T048|SY|47372000|SNOMEDCT_CORE|Adjustment disorder with anxiety|Adjustment disorder with anxious mood
C0154587|T048|PT|47372000|SNOMEDCT_CORE|Adjustment disorder with anxious mood|Adjustment disorder with anxious mood
C0154587|T048|FN|47372000|SNOMEDCT_CORE|Adjustment disorder with anxious mood|Adjustment disorder with anxious mood
C0154587|T048|SY|47372000|SNOMEDCT_CORE|Adjustment reaction with anxious mood|Adjustment disorder with anxious mood
C0154653|T047|PT|21664006|SNOMEDCT_CORE|Chronic meningitis|Chronic meningitis
C0154653|T047|FN|21664006|SNOMEDCT_CORE|Chronic meningitis|Chronic meningitis
C0154653|T047|IS|21664006|SNOMEDCT_CORE|Chronic meningitis, NOS|Chronic meningitis
C0154663|T047|PT|192775006|SNOMEDCT_CORE|Late effects of intracranial abscess or pyogenic infection|Late effects of intracranial abscess or pyogenic infection
C0154663|T047|FN|192775006|SNOMEDCT_CORE|Late effects of intracranial abscess or pyogenic infection|Late effects of intracranial abscess or pyogenic infection
C0154681|T047|PT|85672005|SNOMEDCT_CORE|Anterior horn cell disease|Anterior horn cell disease
C0154681|T047|FN|85672005|SNOMEDCT_CORE|Anterior horn cell disease|Anterior horn cell disease
C0154681|T047|IS|85672005|SNOMEDCT_CORE|Anterior horn cell disease, NOS|Anterior horn cell disease
C0154690|T047|PT|86489003|SNOMEDCT_CORE|Idiopathic peripheral autonomic neuropathy|Idiopathic peripheral autonomic neuropathy
C0154690|T047|FN|86489003|SNOMEDCT_CORE|Idiopathic peripheral autonomic neuropathy|Idiopathic peripheral autonomic neuropathy
C0154695|T047|OAP|275469001|SNOMEDCT_CORE|Congenital diplegia|Congenital diplegia
C0154697|T019|PT|275468009|SNOMEDCT_CORE|Congenital quadriplegia|Congenital quadriplegia
C0154697|T047|PT|275468009|SNOMEDCT_CORE|Congenital quadriplegia|Congenital quadriplegia
C0154697|T019|FN|275468009|SNOMEDCT_CORE|Congenital quadriplegia|Congenital quadriplegia
C0154697|T047|FN|275468009|SNOMEDCT_CORE|Congenital quadriplegia|Congenital quadriplegia
C0154697|T019|SY|275468009|SNOMEDCT_CORE|Congenital tetraplegia|Congenital quadriplegia
C0154697|T047|SY|275468009|SNOMEDCT_CORE|Congenital tetraplegia|Congenital quadriplegia
C0154723|T047|PT|4473006|SNOMEDCT_CORE|Migraine with aura|Migraine with aura
C0154723|T047|FN|4473006|SNOMEDCT_CORE|Migraine with aura|Migraine with aura
C0154729|T184|IS|71303008|SNOMEDCT_CORE|Atypical face pain|Atypical facial pain
C0154729|T184|PT|71303008|SNOMEDCT_CORE|Atypical facial pain|Atypical facial pain
C0154729|T184|FN|71303008|SNOMEDCT_CORE|Atypical facial pain|Atypical facial pain
C0154733|T047|PT|78152008|SNOMEDCT_CORE|Multiple cranial nerve palsy|Multiple cranial nerve palsy
C0154733|T047|FN|78152008|SNOMEDCT_CORE|Multiple cranial nerve palsy|Multiple cranial nerve palsy
C0154733|T047|IS|78152008|SNOMEDCT_CORE|Multiple cranial nerve palsy, NOS|Multiple cranial nerve palsy
C0154737|T047|PT|42452002|SNOMEDCT_CORE|Thoracic radiculopathy|Thoracic radiculopathy
C0154737|T047|FN|42452002|SNOMEDCT_CORE|Thoracic radiculopathy|Thoracic radiculopathy
C0154737|T047|SY|42452002|SNOMEDCT_CORE|Thoracic root lesion|Thoracic radiculopathy
C0154737|T047|IS|42452002|SNOMEDCT_CORE|Thoracic root lesion, NOS|Thoracic radiculopathy
C0154738|T047|PT|2415007|SNOMEDCT_CORE|Lumbosacral radiculopathy|Lumbosacral radiculopathy
C0154738|T047|FN|2415007|SNOMEDCT_CORE|Lumbosacral radiculopathy|Lumbosacral radiculopathy
C0154738|T047|IS|2415007|SNOMEDCT_CORE|Lumbosacral radiculopathy, NOS|Lumbosacral radiculopathy
C0154738|T047|SY|2415007|SNOMEDCT_CORE|Lumbosacral root lesion|Lumbosacral radiculopathy
C0154738|T047|IS|2415007|SNOMEDCT_CORE|Lumbosacral root lesion, NOS|Lumbosacral radiculopathy
C0154743|T047|PT|359837005|SNOMEDCT_CORE|Ulnar neuropathy|Ulnar neuropathy
C0154743|T047|FN|359837005|SNOMEDCT_CORE|Ulnar neuropathy|Ulnar neuropathy
C0154744|T047|IS|16644004|SNOMEDCT_CORE|Lesion of radial nerve|Lesion of radial nerve
C0154744|T047|PT|193137006|SNOMEDCT_CORE|Lesion of radial nerve|Lesion of radial nerve
C0154744|T047|FN|193137006|SNOMEDCT_CORE|Lesion of radial nerve|Lesion of radial nerve
C0154744|T047|IS|16644004|SNOMEDCT_CORE|Lesion of radial nerve, NOS|Lesion of radial nerve
C0154744|T047|IS|16644004|SNOMEDCT_CORE|Radial nerve lesion|Lesion of radial nerve
C0154744|T047|SY|193137006|SNOMEDCT_CORE|Radial nerve lesion|Lesion of radial nerve
C0154744|T047|IS|193137006|SNOMEDCT_CORE|Radial nerve lesions|Lesion of radial nerve
C0154744|T047|OF|193137006|SNOMEDCT_CORE|Radial nerve lesions|Lesion of radial nerve
C0154748|T047|IS|52585001|SNOMEDCT_CORE|Lesion of sciatic nerve|Lesion of sciatic nerve
C0154748|T047|IS|52585001|SNOMEDCT_CORE|Lesion of sciatic nerve, NOS|Lesion of sciatic nerve, NOS
C0154756|T047|PT|33209009|SNOMEDCT_CORE|Idiopathic progressive polyneuropathy|Idiopathic progressive polyneuropathy
C0154756|T047|FN|33209009|SNOMEDCT_CORE|Idiopathic progressive polyneuropathy|Idiopathic progressive polyneuropathy
C0154762|T047|SY|7339009|SNOMEDCT_CORE|Drug-related polyneuropathy|Polyneuropathy due to drug
C0154762|T047|FN|7339009|SNOMEDCT_CORE|Polyneuropathy caused by drug|Polyneuropathy due to drug
C0154762|T047|SY|7339009|SNOMEDCT_CORE|Polyneuropathy caused by drug|Polyneuropathy due to drug
C0154762|T047|PT|7339009|SNOMEDCT_CORE|Polyneuropathy due to drug|Polyneuropathy due to drug
C0154762|T047|OF|7339009|SNOMEDCT_CORE|Polyneuropathy due to drug|Polyneuropathy due to drug
C0154762|T047|IS|7339009|SNOMEDCT_CORE|Polyneuropathy due to drug, NOS|Polyneuropathy due to drug
C0154778|T047|SY|32022003|SNOMEDCT_CORE|Degenerative myopia|Degenerative progressive high myopia
C0154778|T047|PT|32022003|SNOMEDCT_CORE|Degenerative progressive high myopia|Degenerative progressive high myopia
C0154778|T047|FN|32022003|SNOMEDCT_CORE|Degenerative progressive high myopia|Degenerative progressive high myopia
C0154778|T047|IS|32022003|SNOMEDCT_CORE|Malignant myopia|Degenerative progressive high myopia
C0154808|T047|PT|56202001|SNOMEDCT_CORE|Retinal detachment with retinal defect|Retinal detachment with retinal defect
C0154808|T047|FN|56202001|SNOMEDCT_CORE|Retinal detachment with retinal defect|Retinal detachment with retinal defect
C0154808|T047|IS|56202001|SNOMEDCT_CORE|Retinal detachment with retinal defect, NOS|Retinal detachment with retinal defect
C0154823|T190|PT|40024006|SNOMEDCT_CORE|Retinal defect|Retinal defect
C0154823|T190|FN|40024006|SNOMEDCT_CORE|Retinal defect|Retinal defect
C0154823|T190|IS|40024006|SNOMEDCT_CORE|Retinal defect, NOS|Retinal defect
C0154825|T047|OAP|193340000|SNOMEDCT_CORE|Retinal round hole without detachment|Round hole of retina without detachment
C0154825|T047|OAF|193340000|SNOMEDCT_CORE|Retinal round hole without detachment|Round hole of retina without detachment
C0154825|T047|PT|51226000|SNOMEDCT_CORE|Round hole of retina without detachment|Round hole of retina without detachment
C0154825|T047|FN|51226000|SNOMEDCT_CORE|Round hole of retina without detachment|Round hole of retina without detachment
C0154826|T047|FN|193341001|SNOMEDCT_CORE|Horseshoe retinal tear without detachment|Horseshoe retinal tear without detachment
C0154826|T047|PT|193341001|SNOMEDCT_CORE|Horseshoe retinal tear without detachment|Horseshoe retinal tear without detachment
C0154828|T046|PT|34711008|SNOMEDCT_CORE|Traction detachment of retina|Traction detachment of retina
C0154828|T046|FN|34711008|SNOMEDCT_CORE|Traction detachment of retina|Traction detachment of retina
C0154828|T046|SY|34711008|SNOMEDCT_CORE|Traction retinal detachment|Traction detachment of retina
C0154828|T046|SY|34711008|SNOMEDCT_CORE|TRD - Traction retinal detachment|Traction detachment of retina
C0154830|T047|IS|59276001|SNOMEDCT_CORE|PDR|Proliferative retinopathy due to diabetes mellitus
C0154830|T047|SY|59276001|SNOMEDCT_CORE|PDR - proliferative diabetic retinopathy|Proliferative retinopathy due to diabetes mellitus
C0154830|T047|IS|59276001|SNOMEDCT_CORE|PDR - Proliferative diabetic retinopathy|Proliferative retinopathy due to diabetes mellitus
C0154830|T047|SY|59276001|SNOMEDCT_CORE|Proliferative diabetic retinopathy|Proliferative retinopathy due to diabetes mellitus
C0154830|T047|OF|59276001|SNOMEDCT_CORE|Proliferative diabetic retinopathy|Proliferative retinopathy due to diabetes mellitus
C0154830|T047|OF|59276001|SNOMEDCT_CORE|Proliferative retinopathy co-occurrent and due to diabetes mellitus|Proliferative retinopathy due to diabetes mellitus
C0154830|T047|IS|59276001|SNOMEDCT_CORE|Proliferative retinopathy co-occurrent and due to diabetes mellitus|Proliferative retinopathy due to diabetes mellitus
C0154830|T047|FN|59276001|SNOMEDCT_CORE|Proliferative retinopathy due to diabetes mellitus|Proliferative retinopathy due to diabetes mellitus
C0154830|T047|PT|59276001|SNOMEDCT_CORE|Proliferative retinopathy due to diabetes mellitus|Proliferative retinopathy due to diabetes mellitus
C0154830|T047|SY|59276001|SNOMEDCT_CORE|Proliferative retinopathy with diabetes mellitus|Proliferative retinopathy due to diabetes mellitus
C0154833|T047|PT|57534004|SNOMEDCT_CORE|Retinal vascular disorder|Retinal vascular disorder
C0154833|T047|FN|57534004|SNOMEDCT_CORE|Retinal vascular disorder|Retinal vascular disorder
C0154841|T047|PT|68478007|SNOMEDCT_CORE|Central retinal vein occlusion|Central retinal vein occlusion
C0154841|T047|FN|68478007|SNOMEDCT_CORE|Central retinal vein occlusion|Central retinal vein occlusion
C0154841|T047|SY|68478007|SNOMEDCT_CORE|Central retinal vein thrombosis|Central retinal vein occlusion
C0154841|T047|SY|68478007|SNOMEDCT_CORE|CRVO - Central retinal vein occlusion|Central retinal vein occlusion
C0154841|T047|SY|68478007|SNOMEDCT_CORE|CRVT - Central retinal vein thrombosis|Central retinal vein occlusion
C0154844|T020|SY|42059000|SNOMEDCT_CORE|Separation of retinal layers|Separation of retinal layers
C0154845|T047|SY|52002008|SNOMEDCT_CORE|Retinal pigment epithelium serous detachment|Serous detachment of retinal pigment epithelium
C0154845|T047|PT|52002008|SNOMEDCT_CORE|Serous detachment of retinal pigment epithelium|Serous detachment of retinal pigment epithelium
C0154845|T047|FN|52002008|SNOMEDCT_CORE|Serous detachment of retinal pigment epithelium|Serous detachment of retinal pigment epithelium
C0154856|T047|SY|3577000|SNOMEDCT_CORE|Lattice degeneration|Retinal lattice degeneration
C0154856|T047|SY|3577000|SNOMEDCT_CORE|Lattice retinal degeneration|Retinal lattice degeneration
C0154856|T047|SY|3577000|SNOMEDCT_CORE|LD - Lattice degeneration|Retinal lattice degeneration
C0154856|T047|SY|3577000|SNOMEDCT_CORE|Palisade degeneration of retina|Retinal lattice degeneration
C0154856|T047|PT|3577000|SNOMEDCT_CORE|Retinal lattice degeneration|Retinal lattice degeneration
C0154856|T047|FN|3577000|SNOMEDCT_CORE|Retinal lattice degeneration|Retinal lattice degeneration
C0154916|T047|SYGB|51995000|SNOMEDCT_CORE|Iris neovascularisation|Rubeosis iridis
C0154916|T047|SY|51995000|SNOMEDCT_CORE|Iris neovascularization|Rubeosis iridis
C0154916|T047|SY|51995000|SNOMEDCT_CORE|New vessels in iris|Rubeosis iridis
C0154916|T047|SY|51995000|SNOMEDCT_CORE|NVI - New vessels iris|Rubeosis iridis
C0154916|T047|PT|51995000|SNOMEDCT_CORE|Rubeosis iridis|Rubeosis iridis
C0154916|T047|FN|51995000|SNOMEDCT_CORE|Rubeosis iridis|Rubeosis iridis
C0154916|T047|SY|51995000|SNOMEDCT_CORE|Rubeotic iris|Rubeosis iridis
C0154946|T047|SY|30041005|SNOMEDCT_CORE|AACG - Acute angle closure glaucoma|Acute angle-closure glaucoma
C0154946|T047|PT|30041005|SNOMEDCT_CORE|Acute angle-closure glaucoma|Acute angle-closure glaucoma
C0154946|T047|FN|30041005|SNOMEDCT_CORE|Acute angle-closure glaucoma|Acute angle-closure glaucoma
C0154946|T047|SY|30041005|SNOMEDCT_CORE|Acute closed-angle glaucoma|Acute angle-closure glaucoma
C0154947|T047|SY|33647009|SNOMEDCT_CORE|Anatomical narrow angle glaucoma|Chronic angle-closure glaucoma
C0154947|T047|FN|33647009|SNOMEDCT_CORE|Anatomical narrow angle glaucoma|Chronic angle-closure glaucoma
C0154947|T047|PT|33647009|SNOMEDCT_CORE|Chronic angle-closure glaucoma|Chronic angle-closure glaucoma
C0154947|T047|SY|33647009|SNOMEDCT_CORE|Chronic closed-angle glaucoma|Chronic angle-closure glaucoma
C0154947|T047|SY|33647009|SNOMEDCT_CORE|Chronic narrow angle glaucoma|Chronic angle-closure glaucoma
C0154947|T047|SY|33647009|SNOMEDCT_CORE|CNAG - Chronic narrow angle glaucoma|Chronic angle-closure glaucoma
C0154964|T047|PT|19309007|SNOMEDCT_CORE|Glaucoma associated with vascular disorder|Glaucoma associated with vascular disorder
C0154964|T047|FN|19309007|SNOMEDCT_CORE|Glaucoma associated with vascular disorder|Glaucoma associated with vascular disorder
C0154964|T047|IS|19309007|SNOMEDCT_CORE|Glaucoma associated with vascular disorders|Glaucoma associated with vascular disorder
C0154979|T047|PT|5318001|SNOMEDCT_CORE|Posterior subcapsular polar senile cataract|Posterior subcapsular polar senile cataract
C0154979|T047|FN|5318001|SNOMEDCT_CORE|Posterior subcapsular polar senile cataract|Posterior subcapsular polar senile cataract
C0154980|T047|PT|78875003|SNOMEDCT_CORE|Cortical senile cataract|Cortical senile cataract
C0154980|T047|FN|78875003|SNOMEDCT_CORE|Cortical senile cataract|Cortical senile cataract
C0154983|T037|PT|34361001|SNOMEDCT_CORE|Traumatic cataract|Traumatic cataract
C0154983|T037|FN|34361001|SNOMEDCT_CORE|Traumatic cataract|Traumatic cataract
C0154983|T037|IS|34361001|SNOMEDCT_CORE|Traumatic cataract, NOS|Traumatic cataract
C0154998|T020|SY|193615000|SNOMEDCT_CORE|After-cataract with vision obscured|After-cataract with vision obscured following extraction of cataract
C0154998|T020|OF|193615000|SNOMEDCT_CORE|After-cataract with vision obscured|After-cataract with vision obscured following extraction of cataract
C0154998|T020|PT|193615000|SNOMEDCT_CORE|After-cataract with vision obscured following extraction of cataract|After-cataract with vision obscured following extraction of cataract
C0154998|T020|FN|193615000|SNOMEDCT_CORE|After-cataract with vision obscured following extraction of cataract|After-cataract with vision obscured following extraction of cataract
C0155003|T046|PT|83785004|SNOMEDCT_CORE|Transient blindness|Transient blindness
C0155003|T046|FN|83785004|SNOMEDCT_CORE|Transient blindness|Transient blindness
C0155003|T046|IS|83785004|SNOMEDCT_CORE|Transient blindness, NOS|Transient blindness
C0155069|T047|PT|7426009|SNOMEDCT_CORE|Central corneal ulcer|Central corneal ulcer
C0155069|T047|FN|7426009|SNOMEDCT_CORE|Central corneal ulcer|Central corneal ulcer
C0155084|T047|PT|77080005|SNOMEDCT_CORE|Neurotrophic keratoconjunctivitis|Neurotrophic keratoconjunctivitis
C0155084|T047|FN|77080005|SNOMEDCT_CORE|Neurotrophic keratoconjunctivitis|Neurotrophic keratoconjunctivitis
C0155111|T047|SY|57207003|SNOMEDCT_CORE|BK - Bullous keratopathy|Bullous keratopathy
C0155111|T047|PT|57207003|SNOMEDCT_CORE|Bullous keratopathy|Bullous keratopathy
C0155111|T047|FN|57207003|SNOMEDCT_CORE|Bullous keratopathy|Bullous keratopathy
C0155119|T047|SY|2055003|SNOMEDCT_CORE|Recurrent corneal erosion|Recurrent erosion of cornea
C0155119|T047|PT|2055003|SNOMEDCT_CORE|Recurrent erosion of cornea|Recurrent erosion of cornea
C0155119|T047|FN|2055003|SNOMEDCT_CORE|Recurrent erosion of cornea|Recurrent erosion of cornea
C0155119|T047|SY|2055003|SNOMEDCT_CORE|Recurrent erosion syndrome|Recurrent erosion of cornea
C0155120|T047|SY|35055000|SNOMEDCT_CORE|Band keratopathy|Band-shaped keratopathy
C0155120|T047|SY|35055000|SNOMEDCT_CORE|Band shaped keratopathy|Band-shaped keratopathy
C0155120|T047|PT|35055000|SNOMEDCT_CORE|Band-shaped keratopathy|Band-shaped keratopathy
C0155120|T047|FN|35055000|SNOMEDCT_CORE|Band-shaped keratopathy|Band-shaped keratopathy
C0155120|T047|SY|35055000|SNOMEDCT_CORE|BK - Band keratopathy|Band-shaped keratopathy
C0155122|T047|PT|72620002|SNOMEDCT_CORE|Nodular degeneration of cornea|Nodular degeneration of cornea
C0155122|T047|FN|72620002|SNOMEDCT_CORE|Nodular degeneration of cornea|Nodular degeneration of cornea
C0155141|T047|PT|53726008|SNOMEDCT_CORE|Acute conjunctivitis|Acute conjunctivitis
C0155141|T047|FN|53726008|SNOMEDCT_CORE|Acute conjunctivitis|Acute conjunctivitis
C0155141|T047|IS|53726008|SNOMEDCT_CORE|Acute conjunctivitis, NOS|Acute conjunctivitis
C0155143|T047|PT|41308008|SNOMEDCT_CORE|Acute follicular conjunctivitis|Acute follicular conjunctivitis
C0155143|T047|FN|41308008|SNOMEDCT_CORE|Acute follicular conjunctivitis|Acute follicular conjunctivitis
C0155143|T047|IS|41308008|SNOMEDCT_CORE|Acute follicular conjunctivitis, NOS|Acute follicular conjunctivitis
C0155143|T047|SY|41308008|SNOMEDCT_CORE|Conjunctival folliculosis|Acute follicular conjunctivitis
C0155143|T047|IS|41308008|SNOMEDCT_CORE|Conjunctival folliculosis, NOS|Acute follicular conjunctivitis
C0155158|T047|PT|73181007|SNOMEDCT_CORE|Recurrent pterygium|Recurrent pterygium
C0155158|T047|FN|73181007|SNOMEDCT_CORE|Recurrent pterygium|Recurrent pterygium
C0155169|T047|SY|781682005|SNOMEDCT_CORE|Bloodshot eye|Hyperemia of eye
C0155169|T047|PTGB|781682005|SNOMEDCT_CORE|Hyperaemia of eye|Hyperemia of eye
C0155169|T047|PT|781682005|SNOMEDCT_CORE|Hyperemia of eye|Hyperemia of eye
C0155169|T047|FN|781682005|SNOMEDCT_CORE|Hyperemia of eye|Hyperemia of eye
C0155188|T047|SY|55408009|SNOMEDCT_CORE|Age-related entropion|Senile entropion
C0155188|T047|SY|55408009|SNOMEDCT_CORE|Involutional entropion|Senile entropion
C0155188|T047|PT|55408009|SNOMEDCT_CORE|Senile entropion|Senile entropion
C0155188|T047|FN|55408009|SNOMEDCT_CORE|Senile entropion|Senile entropion
C0155197|T047|PT|59890007|SNOMEDCT_CORE|Paralytic lagophthalmos|Paralytic lagophthalmos
C0155197|T047|OF|59890007|SNOMEDCT_CORE|Paralytic lagophthalmos|Paralytic lagophthalmos
C0155197|T047|FN|59890007|SNOMEDCT_CORE|Paralytic lagophthalmos|Paralytic lagophthalmos
C0155198|T047|PT|21783006|SNOMEDCT_CORE|Mechanical lagophthalmos|Mechanical lagophthalmos
C0155198|T047|FN|21783006|SNOMEDCT_CORE|Mechanical lagophthalmos|Mechanical lagophthalmos
C0155202|T020|PT|76201007|SNOMEDCT_CORE|Mechanical ptosis|Mechanical ptosis
C0155202|T020|FN|76201007|SNOMEDCT_CORE|Mechanical ptosis|Mechanical ptosis
C0155218|T047|PT|46210008|SNOMEDCT_CORE|Cyst of eyelid|Cyst of eyelid
C0155218|T047|FN|46210008|SNOMEDCT_CORE|Cyst of eyelid|Cyst of eyelid
C0155218|T047|IS|46210008|SNOMEDCT_CORE|Cyst of eyelid, NOS|Cyst of eyelid
C0155234|T047|PT|85042000|SNOMEDCT_CORE|Epiphora due to insufficient drainage|Epiphora due to insufficient drainage
C0155234|T047|FN|85042000|SNOMEDCT_CORE|Epiphora due to insufficient drainage|Epiphora due to insufficient drainage
C0155244|T047|SY|74783009|SNOMEDCT_CORE|Punctal stenosis|Stenosis of lacrimal punctum
C0155244|T047|PT|74783009|SNOMEDCT_CORE|Stenosis of lacrimal punctum|Stenosis of lacrimal punctum
C0155244|T047|FN|74783009|SNOMEDCT_CORE|Stenosis of lacrimal punctum|Stenosis of lacrimal punctum
C0155245|T190|PT|81345003|SNOMEDCT_CORE|Stenosis of lacrimal canaliculi|Stenosis of lacrimal canaliculi
C0155245|T190|FN|81345003|SNOMEDCT_CORE|Stenosis of lacrimal canaliculi|Stenosis of lacrimal canaliculi
C0155245|T190|SY|81345003|SNOMEDCT_CORE|Stenosis of lacrimal canaliculus|Stenosis of lacrimal canaliculi
C0155245|T190|SY|81345003|SNOMEDCT_CORE|Stenosis of lacrimal passage|Stenosis of lacrimal canaliculi
C0155247|T047|SY|193994000|SNOMEDCT_CORE|CNDO - Congenital nasolacrimal duct obstruction|Congenital nasolacrimal duct obstruction
C0155247|T047|SY|193994000|SNOMEDCT_CORE|CNLDO - Congenital nasolacrimal duct obstruction|Congenital nasolacrimal duct obstruction
C0155247|T047|PT|193994000|SNOMEDCT_CORE|Congenital nasolacrimal duct obstruction|Congenital nasolacrimal duct obstruction
C0155247|T047|FN|193994000|SNOMEDCT_CORE|Congenital nasolacrimal duct obstruction|Congenital nasolacrimal duct obstruction
C0155247|T047|SY|193994000|SNOMEDCT_CORE|Neonatal nasolacrimal duct obstruction|Congenital nasolacrimal duct obstruction
C0155248|T020|SY|193995004|SNOMEDCT_CORE|Acquired dacryostenosis|Acquired stenosis of nasolacrimal duct
C0155248|T020|SY|193995004|SNOMEDCT_CORE|Acquired nasolacrimal duct stenosis|Acquired stenosis of nasolacrimal duct
C0155248|T020|FN|193995004|SNOMEDCT_CORE|Acquired nasolacrimal duct stenosis|Acquired stenosis of nasolacrimal duct
C0155248|T020|PT|193995004|SNOMEDCT_CORE|Acquired stenosis of nasolacrimal duct|Acquired stenosis of nasolacrimal duct
C0155248|T020|SY|193995004|SNOMEDCT_CORE|Acquired tear duct stenosis|Acquired stenosis of nasolacrimal duct
C0155264|T047|SY|276177000|SNOMEDCT_CORE|Endocrine exophthalmos|Endocrine exophthalmos
C0155305|T047|IS|14357004|SNOMEDCT_CORE|AION - Acute ischaemic optic neuropathy|Ischemic optic neuropathy
C0155305|T047|IS|14357004|SNOMEDCT_CORE|AION - Acute ischemic optic neuropathy|Ischemic optic neuropathy
C0155305|T047|SYGB|14357004|SNOMEDCT_CORE|ION - Ischaemic optic neuropathy|Ischemic optic neuropathy
C0155305|T047|SY|14357004|SNOMEDCT_CORE|ION - Ischemic optic neuropathy|Ischemic optic neuropathy
C0155305|T047|PTGB|14357004|SNOMEDCT_CORE|Ischaemic optic neuropathy|Ischemic optic neuropathy
C0155305|T047|PT|14357004|SNOMEDCT_CORE|Ischemic optic neuropathy|Ischemic optic neuropathy
C0155305|T047|FN|14357004|SNOMEDCT_CORE|Ischemic optic neuropathy|Ischemic optic neuropathy
C0155332|T047|PT|57805002|SNOMEDCT_CORE|Alternating exotropia with V pattern|Alternating exotropia with V pattern
C0155332|T047|FN|57805002|SNOMEDCT_CORE|Alternating exotropia with V pattern|Alternating exotropia with V pattern
C0155336|T047|PT|194112008|SNOMEDCT_CORE|Esotropia with accommodative compensation|Esotropia with accommodative compensation
C0155336|T047|FN|194112008|SNOMEDCT_CORE|Esotropia with accommodative compensation|Esotropia with accommodative compensation
C0155366|T047|PT|60189009|SNOMEDCT_CORE|Vitreous degeneration|Vitreous degeneration
C0155366|T047|FN|60189009|SNOMEDCT_CORE|Vitreous degeneration|Vitreous degeneration
C0155366|T047|IS|60189009|SNOMEDCT_CORE|Vitreous degeneration, NOS|Vitreous degeneration
C0155388|T047|PT|49130001|SNOMEDCT_CORE|Disorder of external ear|Disorder of external ear
C0155388|T047|FN|49130001|SNOMEDCT_CORE|Disorder of external ear|Disorder of external ear
C0155388|T047|IS|49130001|SNOMEDCT_CORE|Disorder of external ear, NOS|Disorder of external ear
C0155393|T047|IS|30250000|SNOMEDCT_CORE|Acute swimmer's ear|Acute swimmer's ear
C0155402|T047|PT|41663005|SNOMEDCT_CORE|Disorder of pinna|Disorder of pinna
C0155402|T047|FN|41663005|SNOMEDCT_CORE|Disorder of pinna|Disorder of pinna
C0155402|T047|IS|41663005|SNOMEDCT_CORE|Disorder of pinna, NOS|Disorder of pinna
C0155415|T047|PT|194240006|SNOMEDCT_CORE|Acute non-suppurative otitis media - serous|Acute non-suppurative otitis media - serous
C0155415|T047|FN|194240006|SNOMEDCT_CORE|Acute non-suppurative otitis media - serous|Acute non-suppurative otitis media - serous
C0155415|T047|OP|194240006|SNOMEDCT_CORE|Acute serous otitis media|Acute non-suppurative otitis media - serous
C0155421|T047|SY|81564005|SNOMEDCT_CORE|Chronic non-suppurative otitis media with effusion - serous|Chronic serous otitis media
C0155421|T047|SY|81564005|SNOMEDCT_CORE|Chronic secretory otitis media, serous|Chronic serous otitis media
C0155421|T047|PT|81564005|SNOMEDCT_CORE|Chronic serous otitis media|Chronic serous otitis media
C0155421|T047|FN|81564005|SNOMEDCT_CORE|Chronic serous otitis media|Chronic serous otitis media
C0155421|T047|IS|81564005|SNOMEDCT_CORE|Chronic serous otitis media, NOS|Chronic serous otitis media
C0155421|T047|SY|81564005|SNOMEDCT_CORE|Glue ear - serous|Chronic serous otitis media
C0155421|T047|SY|81564005|SNOMEDCT_CORE|Otitis media with effusion - serous|Chronic serous otitis media
C0155421|T047|SY|81564005|SNOMEDCT_CORE|Simple chronic serous otitis media|Chronic serous otitis media
C0155421|T047|IS|81564005|SNOMEDCT_CORE|Simple chronic serous otitis media, NOS|Chronic serous otitis media
C0155440|T047|SY|87665008|SNOMEDCT_CORE|Chronic suppurative otitis media - tubotympanic|Chronic tubotympanic suppurative otitis media
C0155440|T047|PT|87665008|SNOMEDCT_CORE|Chronic tubotympanic suppurative otitis media|Chronic tubotympanic suppurative otitis media
C0155440|T047|FN|87665008|SNOMEDCT_CORE|Chronic tubotympanic suppurative otitis media|Chronic tubotympanic suppurative otitis media
C0155447|T047|PT|80645004|SNOMEDCT_CORE|Chronic mastoiditis|Chronic mastoiditis
C0155447|T047|FN|80645004|SNOMEDCT_CORE|Chronic mastoiditis|Chronic mastoiditis
C0155461|T047|PT|33528003|SNOMEDCT_CORE|Bullous myringitis|Bullous myringitis
C0155461|T047|FN|33528003|SNOMEDCT_CORE|Bullous myringitis|Bullous myringitis
C0155461|T047|SY|33528003|SNOMEDCT_CORE|Myringitis bullosa|Bullous myringitis
C0155461|T047|SYGB|33528003|SNOMEDCT_CORE|Myringitis bullosa haemorrhagica|Bullous myringitis
C0155461|T047|SY|33528003|SNOMEDCT_CORE|Myringitis bullosa hemorrhagica|Bullous myringitis
C0155478|T047|PT|7699004|SNOMEDCT_CORE|Adhesive middle ear disease|Adhesive middle ear disease
C0155478|T047|FN|7699004|SNOMEDCT_CORE|Adhesive middle ear disease|Adhesive middle ear disease
C0155478|T047|IS|7699004|SNOMEDCT_CORE|Adhesive middle ear disease, NOS|Adhesive middle ear disease
C0155478|T047|SY|7699004|SNOMEDCT_CORE|Adhesive otitis media|Adhesive middle ear disease
C0155478|T047|IS|7699004|SNOMEDCT_CORE|Adhesive otitis media, NOS|Adhesive middle ear disease
C0155478|T047|SY|7699004|SNOMEDCT_CORE|Chronic adhesive otitis media|Adhesive middle ear disease
C0155478|T047|SY|7699004|SNOMEDCT_CORE|Fibrotic adhesive otitis media|Adhesive middle ear disease
C0155489|T047|PT|38708003|SNOMEDCT_CORE|Cholesteatoma of attic|Cholesteatoma of attic
C0155489|T047|FN|38708003|SNOMEDCT_CORE|Cholesteatoma of attic|Cholesteatoma of attic
C0155490|T047|PT|87688009|SNOMEDCT_CORE|Cholesteatoma of middle ear|Cholesteatoma of middle ear
C0155490|T047|FN|87688009|SNOMEDCT_CORE|Cholesteatoma of middle ear|Cholesteatoma of middle ear
C0155490|T047|SY|87688009|SNOMEDCT_CORE|Epidermosis of middle ear|Cholesteatoma of middle ear
C0155501|T047|PT|50438001|SNOMEDCT_CORE|Peripheral vertigo|Peripheral vertigo
C0155501|T047|FN|50438001|SNOMEDCT_CORE|Peripheral vertigo|Peripheral vertigo
C0155501|T047|IS|50438001|SNOMEDCT_CORE|Peripheral vertigo, NOS|Peripheral vertigo
C0155501|T047|SY|50438001|SNOMEDCT_CORE|Peripheral vestibular vertigo|Peripheral vertigo
C0155501|T047|SY|50438001|SNOMEDCT_CORE|Vestibular vertigo|Peripheral vertigo
C0155502|T047|SY|111541001|SNOMEDCT_CORE|Benign paroxysmal positional nystagmus|Benign paroxysmal positional vertigo
C0155502|T047|PT|111541001|SNOMEDCT_CORE|Benign paroxysmal positional vertigo|Benign paroxysmal positional vertigo
C0155502|T047|FN|111541001|SNOMEDCT_CORE|Benign paroxysmal positional vertigo|Benign paroxysmal positional vertigo
C0155502|T047|SY|111541001|SNOMEDCT_CORE|BPPV - Benign paroxysmal positional vertigo|Benign paroxysmal positional vertigo
C0155503|T047|SY|20425006|SNOMEDCT_CORE|Central vestibular vertigo|Vertigo of central origin
C0155503|T047|IS|20425006|SNOMEDCT_CORE|Vertigo of central origin|Vertigo of central origin
C0155508|T047|PT|409711008|SNOMEDCT_CORE|Viral labyrinthitis|Viral labyrinthitis
C0155508|T047|FN|409711008|SNOMEDCT_CORE|Viral labyrinthitis|Viral labyrinthitis
C0155508|T047|SY|409711008|SNOMEDCT_CORE|Viral otitis interna|Viral labyrinthitis
C0155524|T047|SY|62856000|SNOMEDCT_CORE|Non-obliterative otosclerosis|Nonobliterative otosclerosis involving oval window
C0155524|T047|PT|62856000|SNOMEDCT_CORE|Nonobliterative otosclerosis involving oval window|Nonobliterative otosclerosis involving oval window
C0155524|T047|FN|62856000|SNOMEDCT_CORE|Nonobliterative otosclerosis involving oval window|Nonobliterative otosclerosis involving oval window
C0155524|T047|SY|62856000|SNOMEDCT_CORE|Otosclerosis involving oval window - non-obliterative|Nonobliterative otosclerosis involving oval window
C0155533|T184|PT|62452009|SNOMEDCT_CORE|Subjective tinnitus|Subjective tinnitus
C0155533|T184|FN|62452009|SNOMEDCT_CORE|Subjective tinnitus|Subjective tinnitus
C0155533|T184|SY|62452009|SNOMEDCT_CORE|Tinnitus aurium|Subjective tinnitus
C0155534|T184|PT|28715001|SNOMEDCT_CORE|Objective tinnitus|Objective tinnitus
C0155534|T184|FN|28715001|SNOMEDCT_CORE|Objective tinnitus|Objective tinnitus
C0155540|T033|SY|65668001|SNOMEDCT_CORE|Discharge of ear|Otorrhea
C0155540|T033|IS|65668001|SNOMEDCT_CORE|Discharge of ear, NOS|Otorrhea
C0155540|T033|SY|65668001|SNOMEDCT_CORE|Drainage from external ear canal|Otorrhea
C0155540|T033|IS|65668001|SNOMEDCT_CORE|Drainage from external ear canal, NOS|Otorrhea
C0155540|T033|PT|65668001|SNOMEDCT_CORE|Otorrhea|Otorrhea
C0155540|T033|FN|65668001|SNOMEDCT_CORE|Otorrhea|Otorrhea
C0155540|T033|IS|65668001|SNOMEDCT_CORE|Otorrhea, NOS|Otorrhea
C0155540|T033|PTGB|65668001|SNOMEDCT_CORE|Otorrhoea|Otorrhea
C0155552|T047|SY|77507001|SNOMEDCT_CORE|MHL - Mixed hearing loss|Mixed conductive AND sensorineural hearing loss
C0155552|T047|SY|77507001|SNOMEDCT_CORE|Mixed conductive and sensorineural deafness|Mixed conductive AND sensorineural hearing loss
C0155552|T047|PT|77507001|SNOMEDCT_CORE|Mixed conductive AND sensorineural hearing loss|Mixed conductive AND sensorineural hearing loss
C0155552|T047|IS|77507001|SNOMEDCT_CORE|Mixed conductive and sensorineural hearing loss|Mixed conductive AND sensorineural hearing loss
C0155552|T047|OF|77507001|SNOMEDCT_CORE|Mixed conductive AND sensorineural hearing loss|Mixed conductive AND sensorineural hearing loss
C0155552|T047|FN|77507001|SNOMEDCT_CORE|Mixed conductive AND sensorineural hearing loss|Mixed conductive AND sensorineural hearing loss
C0155552|T047|SY|77507001|SNOMEDCT_CORE|Mixed deafness|Mixed conductive AND sensorineural hearing loss
C0155552|T047|SY|77507001|SNOMEDCT_CORE|Mixed hearing loss|Mixed conductive AND sensorineural hearing loss
C0155552|T047|SY|77507001|SNOMEDCT_CORE|Mixed type deafness|Mixed conductive AND sensorineural hearing loss
C0155563|T047|SY|31085000|SNOMEDCT_CORE|Mitral incompetence - rheumatic|Rheumatic mitral regurgitation
C0155563|T047|SY|31085000|SNOMEDCT_CORE|Rheumatic mitral incompetence|Rheumatic mitral regurgitation
C0155563|T047|SY|31085000|SNOMEDCT_CORE|Rheumatic mitral insufficiency|Rheumatic mitral regurgitation
C0155563|T047|PT|31085000|SNOMEDCT_CORE|Rheumatic mitral regurgitation|Rheumatic mitral regurgitation
C0155563|T047|FN|31085000|SNOMEDCT_CORE|Rheumatic mitral regurgitation|Rheumatic mitral regurgitation
C0155567|T047|PT|72011007|SNOMEDCT_CORE|Rheumatic aortic stenosis|Rheumatic aortic stenosis
C0155567|T047|FN|72011007|SNOMEDCT_CORE|Rheumatic aortic stenosis|Rheumatic aortic stenosis
C0155567|T047|SY|72011007|SNOMEDCT_CORE|Rheumatic aortic valve obstruction|Rheumatic aortic stenosis
C0155568|T047|SY|78031003|SNOMEDCT_CORE|Aortic incompetence - rheumatic|Rheumatic aortic regurgitation
C0155568|T047|SY|78031003|SNOMEDCT_CORE|Rheumatic aortic incompetence|Rheumatic aortic regurgitation
C0155568|T047|SY|78031003|SNOMEDCT_CORE|Rheumatic aortic insufficiency|Rheumatic aortic regurgitation
C0155568|T047|PT|78031003|SNOMEDCT_CORE|Rheumatic aortic regurgitation|Rheumatic aortic regurgitation
C0155568|T047|FN|78031003|SNOMEDCT_CORE|Rheumatic aortic regurgitation|Rheumatic aortic regurgitation
C0155569|T047|SY|17759006|SNOMEDCT_CORE|Rheumatic aortic stenosis with incompetence|Rheumatic aortic stenosis with regurgitation
C0155569|T047|SY|17759006|SNOMEDCT_CORE|Rheumatic aortic stenosis with insufficiency|Rheumatic aortic stenosis with regurgitation
C0155569|T047|PT|17759006|SNOMEDCT_CORE|Rheumatic aortic stenosis with regurgitation|Rheumatic aortic stenosis with regurgitation
C0155569|T047|FN|17759006|SNOMEDCT_CORE|Rheumatic aortic stenosis with regurgitation|Rheumatic aortic stenosis with regurgitation
C0155582|T047|PT|82523003|SNOMEDCT_CORE|Congestive rheumatic heart failure|Congestive rheumatic heart failure
C0155582|T047|FN|82523003|SNOMEDCT_CORE|Congestive rheumatic heart failure|Congestive rheumatic heart failure
C0155583|T047|FN|1201005|SNOMEDCT_CORE|Benign essential hypertension|Benign essential hypertension
C0155583|T047|PT|1201005|SNOMEDCT_CORE|Benign essential hypertension|Benign essential hypertension
C0155591|T047|PT|60899001|SNOMEDCT_CORE|Hypertensive heart disease without congestive heart failure|Hypertensive heart disease without congestive heart failure
C0155591|T047|FN|60899001|SNOMEDCT_CORE|Hypertensive heart disease without congestive heart failure|Hypertensive heart disease without congestive heart failure
C0155601|T047|SY|86234004|SNOMEDCT_CORE|Cardiorenal disease|Hypertensive heart AND renal disease
C0155601|T047|IS|86234004|SNOMEDCT_CORE|Cardiorenal disease, NOS|Hypertensive heart AND renal disease
C0155601|T047|PT|86234004|SNOMEDCT_CORE|Hypertensive heart AND renal disease|Hypertensive heart AND renal disease
C0155601|T047|FN|86234004|SNOMEDCT_CORE|Hypertensive heart AND renal disease|Hypertensive heart AND renal disease
C0155601|T047|IS|86234004|SNOMEDCT_CORE|Hypertensive heart and renal disease, NOS|Hypertensive heart AND renal disease
C0155616|T047|PT|31992008|SNOMEDCT_CORE|Secondary hypertension|Secondary hypertension
C0155616|T047|FN|31992008|SNOMEDCT_CORE|Secondary hypertension|Secondary hypertension
C0155616|T047|IS|31992008|SNOMEDCT_CORE|Secondary hypertension, NOS|Secondary hypertension
C0155620|T047|PT|194785008|SNOMEDCT_CORE|Benign secondary hypertension|Benign secondary hypertension
C0155620|T047|SY|194785008|SNOMEDCT_CORE|Secondary benign hypertension|Benign secondary hypertension
C0155620|T047|FN|194785008|SNOMEDCT_CORE|Secondary benign hypertension|Benign secondary hypertension
C0155626|T047|PT|57054005|SNOMEDCT_CORE|Acute myocardial infarction|Acute myocardial infarction
C0155626|T047|FN|57054005|SNOMEDCT_CORE|Acute myocardial infarction|Acute myocardial infarction
C0155626|T047|IS|57054005|SNOMEDCT_CORE|Acute myocardial infarction, NOS|Acute myocardial infarction
C0155626|T047|SY|57054005|SNOMEDCT_CORE|AMI - Acute myocardial infarction|Acute myocardial infarction
C0155668|T047|SY|1755008|SNOMEDCT_CORE|Healed coronary|Old myocardial infarction
C0155668|T047|SY|1755008|SNOMEDCT_CORE|Healed myocardial infarction|Old myocardial infarction
C0155668|T047|PT|1755008|SNOMEDCT_CORE|Old myocardial infarction|Old myocardial infarction
C0155668|T047|FN|1755008|SNOMEDCT_CORE|Old myocardial infarction|Old myocardial infarction
C0155672|T047|PT|49584005|SNOMEDCT_CORE|Acute cor pulmonale|Acute cor pulmonale
C0155672|T047|FN|49584005|SNOMEDCT_CORE|Acute cor pulmonale|Acute cor pulmonale
C0155679|T047|PT|15555002|SNOMEDCT_CORE|Acute pericarditis|Acute pericarditis
C0155679|T047|FN|15555002|SNOMEDCT_CORE|Acute pericarditis|Acute pericarditis
C0155679|T047|IS|15555002|SNOMEDCT_CORE|Acute pericarditis, NOS|Acute pericarditis
C0155700|T047|SY|28189009|SNOMEDCT_CORE|Mobitz type 2 second degree atrioventricular block|Mobitz type II atrioventricular block
C0155700|T047|PT|28189009|SNOMEDCT_CORE|Mobitz type II atrioventricular block|Mobitz type II atrioventricular block
C0155700|T047|FN|28189009|SNOMEDCT_CORE|Mobitz type II atrioventricular block|Mobitz type II atrioventricular block
C0155700|T047|SY|28189009|SNOMEDCT_CORE|Mobitz type II incomplete atrioventricular block|Mobitz type II atrioventricular block
C0155700|T047|SY|28189009|SNOMEDCT_CORE|Second degree Mobitz type II incomplete atrioventricular block|Mobitz type II atrioventricular block
C0155709|T046|PT|195080001|SNOMEDCT_CORE|Atrial fibrillation and flutter|Atrial fibrillation and flutter
C0155709|T046|FN|195080001|SNOMEDCT_CORE|Atrial fibrillation and flutter|Atrial fibrillation and flutter
C0155730|T190|OAS|42994005|SNOMEDCT_CORE|Cerebral aneurysm, nonruptured|Cerebral aneurysm, nonruptured
C0155730|T190|OAP|42994005|SNOMEDCT_CORE|Nonruptured cerebral aneurysm|Cerebral aneurysm, nonruptured
C0155730|T190|OAF|42994005|SNOMEDCT_CORE|Nonruptured cerebral aneurysm|Cerebral aneurysm, nonruptured
C0155730|T190|OAS|42994005|SNOMEDCT_CORE|Unruptured cerebral aneurysm|Cerebral aneurysm, nonruptured
C0155732|T046|PT|195239002|SNOMEDCT_CORE|Late effects of cerebrovascular disease|Late effects of cerebrovascular disease
C0155732|T046|FN|195239002|SNOMEDCT_CORE|Late effects of cerebrovascular disease|Late effects of cerebrovascular disease
C0155732|T046|SY|195239002|SNOMEDCT_CORE|Sequelae of cerebrovascular disease|Late effects of cerebrovascular disease
C0155733|T047|SY|81817003|SNOMEDCT_CORE|Atherosclerosis aorta|Atherosclerosis of aorta
C0155733|T047|PT|81817003|SNOMEDCT_CORE|Atherosclerosis of aorta|Atherosclerosis of aorta
C0155733|T047|FN|81817003|SNOMEDCT_CORE|Atherosclerosis of aorta|Atherosclerosis of aorta
C0155734|T047|PT|45281005|SNOMEDCT_CORE|Atherosclerosis of renal artery|Atherosclerosis of renal artery
C0155734|T047|FN|45281005|SNOMEDCT_CORE|Atherosclerosis of renal artery|Atherosclerosis of renal artery
C0155734|T047|SY|45281005|SNOMEDCT_CORE|Atherosclerosis renal artery|Atherosclerosis of renal artery
C0155734|T047|SY|45281005|SNOMEDCT_CORE|Renal artery atheroma|Atherosclerosis of renal artery
C0155734|T047|SY|45281005|SNOMEDCT_CORE|Renal artery atherosclerosis|Atherosclerosis of renal artery
C0155735|T047|PT|51274000|SNOMEDCT_CORE|Atherosclerosis of arteries of the extremities|Atherosclerosis of arteries of the extremities
C0155735|T047|FN|51274000|SNOMEDCT_CORE|Atherosclerosis of arteries of the extremities|Atherosclerosis of arteries of the extremities
C0155742|T190|PT|36184004|SNOMEDCT_CORE|Aneurysm of renal artery|Aneurysm of renal artery
C0155742|T190|FN|36184004|SNOMEDCT_CORE|Aneurysm of renal artery|Aneurysm of renal artery
C0155773|T047|SY|17920008|SNOMEDCT_CORE|Deep vein thrombosis of portal vein|Portal vein thrombosis
C0155773|T047|PT|17920008|SNOMEDCT_CORE|Portal vein thrombosis|Portal vein thrombosis
C0155773|T047|FN|17920008|SNOMEDCT_CORE|Portal vein thrombosis|Portal vein thrombosis
C0155773|T047|SY|17920008|SNOMEDCT_CORE|PVT - Portal vein thrombosis|Portal vein thrombosis
C0155778|T047|SY|72866009|SNOMEDCT_CORE|Phlebectasia of lower extremity|Varicose veins of lower extremity
C0155778|T047|IS|72866009|SNOMEDCT_CORE|Phlebectasia of lower extremity, NOS|Varicose veins of lower extremity
C0155778|T047|PT|72866009|SNOMEDCT_CORE|Varicose veins of lower extremity|Varicose veins of lower extremity
C0155778|T047|FN|72866009|SNOMEDCT_CORE|Varicose veins of lower extremity|Varicose veins of lower extremity
C0155778|T047|IS|72866009|SNOMEDCT_CORE|Varicose veins of lower extremity, NOS|Varicose veins of lower extremity
C0155778|T047|SY|72866009|SNOMEDCT_CORE|Varicose veins of lower limb|Varicose veins of lower extremity
C0155778|T047|SY|72866009|SNOMEDCT_CORE|Varix of lower extremity|Varicose veins of lower extremity
C0155778|T047|IS|72866009|SNOMEDCT_CORE|Varix of lower extremity, NOS|Varicose veins of lower extremity
C0155778|T047|SY|72866009|SNOMEDCT_CORE|VV - Varicose veins of leg|Varicose veins of lower extremity
C0155779|T047|PT|69352009|SNOMEDCT_CORE|Varicose veins of lower extremity with ulcer AND inflammation|Varicose veins of lower extremity with ulcer AND inflammation
C0155779|T047|IS|69352009|SNOMEDCT_CORE|Varicose veins of lower extremity with ulcer and inflammation|Varicose veins of lower extremity with ulcer AND inflammation
C0155779|T047|FN|69352009|SNOMEDCT_CORE|Varicose veins of lower extremity with ulcer AND inflammation|Varicose veins of lower extremity with ulcer AND inflammation
C0155781|T047|PTGB|52931009|SNOMEDCT_CORE|Thrombosed internal haemorrhoids|Thrombosed internal hemorrhoids
C0155781|T047|PT|52931009|SNOMEDCT_CORE|Thrombosed internal hemorrhoids|Thrombosed internal hemorrhoids
C0155781|T047|FN|52931009|SNOMEDCT_CORE|Thrombosed internal hemorrhoids|Thrombosed internal hemorrhoids
C0155784|T020|SYGB|26373009|SNOMEDCT_CORE|External thrombosed haemorrhoids|Thrombosed external hemorrhoids
C0155784|T020|SY|26373009|SNOMEDCT_CORE|External thrombosed hemorrhoids|Thrombosed external hemorrhoids
C0155784|T020|IS|26373009|SNOMEDCT_CORE|Perianal haematoma|Thrombosed external hemorrhoids
C0155784|T020|IS|26373009|SNOMEDCT_CORE|Perianal hematoma|Thrombosed external hemorrhoids
C0155784|T020|SYGB|26373009|SNOMEDCT_CORE|Thrombosed external haemorrhoid|Thrombosed external hemorrhoids
C0155784|T020|PTGB|26373009|SNOMEDCT_CORE|Thrombosed external haemorrhoids|Thrombosed external hemorrhoids
C0155784|T020|SY|26373009|SNOMEDCT_CORE|Thrombosed external hemorrhoid|Thrombosed external hemorrhoids
C0155784|T020|PT|26373009|SNOMEDCT_CORE|Thrombosed external hemorrhoids|Thrombosed external hemorrhoids
C0155784|T020|FN|26373009|SNOMEDCT_CORE|Thrombosed external hemorrhoids|Thrombosed external hemorrhoids
C0155784|T020|SY|26373009|SNOMEDCT_CORE|Thrombosed external pile|Thrombosed external hemorrhoids
C0155789|T047|PT|17709002|SNOMEDCT_CORE|Bleeding esophageal varices|Bleeding esophageal varices
C0155789|T047|FN|17709002|SNOMEDCT_CORE|Bleeding esophageal varices|Bleeding esophageal varices
C0155789|T047|PTGB|17709002|SNOMEDCT_CORE|Bleeding oesophageal varices|Bleeding esophageal varices
C0155789|T047|SY|17709002|SNOMEDCT_CORE|BOV - Bleeding esophageal varices|Bleeding esophageal varices
C0155789|T047|SYGB|17709002|SNOMEDCT_CORE|BOV - Bleeding oesophageal varices|Bleeding esophageal varices
C0155789|T047|SY|17709002|SNOMEDCT_CORE|Esophageal varices with bleeding|Bleeding esophageal varices
C0155789|T047|SY|17709002|SNOMEDCT_CORE|Esophageal varices with hemorrhage|Bleeding esophageal varices
C0155789|T047|SYGB|17709002|SNOMEDCT_CORE|Oesophageal varices with bleeding|Bleeding esophageal varices
C0155789|T047|SYGB|17709002|SNOMEDCT_CORE|Oesophageal varices with haemorrhage|Bleeding esophageal varices
C0155791|T047|IS|195474004|SNOMEDCT_CORE|Esophageal varices in diseases EC|Oesophageal varices in diseases EC
C0155791|T047|OF|195474004|SNOMEDCT_CORE|Esophageal varices in diseases EC|Oesophageal varices in diseases EC
C0155791|T047|IS|195474004|SNOMEDCT_CORE|Oesophageal varices in diseases EC|Oesophageal varices in diseases EC
C0155804|T047|SY|68272006|SNOMEDCT_CORE|Acute antritis|Acute maxillary sinusitis
C0155804|T047|PT|68272006|SNOMEDCT_CORE|Acute maxillary sinusitis|Acute maxillary sinusitis
C0155804|T047|FN|68272006|SNOMEDCT_CORE|Acute maxillary sinusitis|Acute maxillary sinusitis
C0155805|T047|PT|91038008|SNOMEDCT_CORE|Acute frontal sinusitis|Acute frontal sinusitis
C0155805|T047|FN|91038008|SNOMEDCT_CORE|Acute frontal sinusitis|Acute frontal sinusitis
C0155814|T047|PT|29608009|SNOMEDCT_CORE|Acute epiglottitis|Acute epiglottitis
C0155814|T047|FN|29608009|SNOMEDCT_CORE|Acute epiglottitis|Acute epiglottitis
C0155814|T047|SY|29608009|SNOMEDCT_CORE|Acute epiglottitis and supraglottitis|Acute epiglottitis
C0155825|T047|FN|140004|SNOMEDCT_CORE|Chronic pharyngitis|Chronic pharyngitis
C0155825|T047|SY|140004|SNOMEDCT_CORE|Chronic sore throat|Chronic sore throat
C0155826|T047|PT|47841006|SNOMEDCT_CORE|Chronic nasopharyngitis|Chronic nasopharyngitis
C0155826|T047|FN|47841006|SNOMEDCT_CORE|Chronic nasopharyngitis|Chronic nasopharyngitis
C0155827|T047|PT|88850006|SNOMEDCT_CORE|Chronic pansinusitis|Chronic pansinusitis
C0155827|T047|FN|88850006|SNOMEDCT_CORE|Chronic pansinusitis|Chronic pansinusitis
C0155828|T047|IS|16358007|SNOMEDCT_CORE|Chronic disease of tonsils and adenoids, NOS|Chronic disease of tonsils AND/OR adenoids
C0155828|T047|PT|16358007|SNOMEDCT_CORE|Chronic disease of tonsils AND/OR adenoids|Chronic disease of tonsils AND/OR adenoids
C0155828|T047|FN|16358007|SNOMEDCT_CORE|Chronic disease of tonsils AND/OR adenoids|Chronic disease of tonsils AND/OR adenoids
C0155829|T047|PT|232419008|SNOMEDCT_CORE|Enlargement of tonsil or adenoid|Enlargement of tonsil or adenoid
C0155829|T047|FN|232419008|SNOMEDCT_CORE|Enlargement of tonsil or adenoid|Enlargement of tonsil or adenoid
C0155836|T047|PT|29951006|SNOMEDCT_CORE|Chronic laryngitis|Chronic laryngitis
C0155836|T047|FN|29951006|SNOMEDCT_CORE|Chronic laryngitis|Chronic laryngitis
C0155836|T047|IS|29951006|SNOMEDCT_CORE|Chronic laryngitis, NOS|Chronic laryngitis
C0155840|T047|PT|17467004|SNOMEDCT_CORE|Hypertrophy of nasal turbinates|Hypertrophy of nasal turbinates
C0155840|T047|FN|17467004|SNOMEDCT_CORE|Hypertrophy of nasal turbinates|Hypertrophy of nasal turbinates
C0155842|T047|SY|84889008|SNOMEDCT_CORE|Abscess of lateral pharyngeal space|Parapharyngeal abscess
C0155842|T047|SY|84889008|SNOMEDCT_CORE|Abscess of parapharyngeal space|Parapharyngeal abscess
C0155842|T047|PT|84889008|SNOMEDCT_CORE|Parapharyngeal abscess|Parapharyngeal abscess
C0155842|T047|FN|84889008|SNOMEDCT_CORE|Parapharyngeal abscess|Parapharyngeal abscess
C0155842|T047|SY|84889008|SNOMEDCT_CORE|Peripharyngeal abscess|Parapharyngeal abscess
C0155847|T047|SY|195842003|SNOMEDCT_CORE|Partial paralysis of one vocal cord|Unilateral partial vocal cord paralysis
C0155847|T047|SY|195842003|SNOMEDCT_CORE|Partial unilateral paralysis of vocal cords|Unilateral partial vocal cord paralysis
C0155847|T047|PT|195842003|SNOMEDCT_CORE|Unilateral partial vocal cord paralysis|Unilateral partial vocal cord paralysis
C0155847|T047|OF|195842003|SNOMEDCT_CORE|Unilateral partial vocal cord paralysis|Unilateral partial vocal cord paralysis
C0155847|T047|FN|195842003|SNOMEDCT_CORE|Unilateral partial vocal cord paralysis|Unilateral partial vocal cord paralysis
C0155848|T047|OAP|195843008|SNOMEDCT_CORE|Unilateral total vocal cord paralysis|Unilateral total vocal cord paralysis
C0155848|T047|OF|195843008|SNOMEDCT_CORE|Unilateral total vocal cord paralysis|Unilateral total vocal cord paralysis
C0155848|T047|OAF|195843008|SNOMEDCT_CORE|Unilateral total vocal cord paralysis|Unilateral total vocal cord paralysis
C0155850|T047|OAP|195845001|SNOMEDCT_CORE|Bilateral total vocal cord paralysis|Complete bilateral paralysis of vocal cords
C0155850|T047|SY|42655007|SNOMEDCT_CORE|Bilateral total vocal cord paralysis|Complete bilateral paralysis of vocal cords
C0155850|T047|OAF|195845001|SNOMEDCT_CORE|Bilateral total vocal cord paralysis|Complete bilateral paralysis of vocal cords
C0155850|T047|SY|42655007|SNOMEDCT_CORE|BVCP - bilateral vocal cord paralysis|Complete bilateral paralysis of vocal cords
C0155850|T047|SY|42655007|SNOMEDCT_CORE|BVFP- bilateral vocal fold paralysis|Complete bilateral paralysis of vocal cords
C0155850|T047|PT|42655007|SNOMEDCT_CORE|Complete bilateral paralysis of vocal cords|Complete bilateral paralysis of vocal cords
C0155850|T047|FN|42655007|SNOMEDCT_CORE|Complete bilateral paralysis of vocal cords|Complete bilateral paralysis of vocal cords
C0155850|T047|SY|42655007|SNOMEDCT_CORE|Complete paralysis of both vocal cords|Complete bilateral paralysis of vocal cords
C0155851|T047|PT|195847009|SNOMEDCT_CORE|Polyp of vocal cord or larynx|Polyp of vocal cord or larynx
C0155851|T047|FN|195847009|SNOMEDCT_CORE|Polyp of vocal cord or larynx|Polyp of vocal cord or larynx
C0155860|T047|FN|41381004|SNOMEDCT_CORE|Pneumonia caused by Pseudomonas|Pneumonia due to Pseudomonas
C0155860|T047|SY|41381004|SNOMEDCT_CORE|Pneumonia caused by Pseudomonas|Pneumonia due to Pseudomonas
C0155860|T047|PT|41381004|SNOMEDCT_CORE|Pneumonia due to Pseudomonas|Pneumonia due to Pseudomonas
C0155860|T047|OF|41381004|SNOMEDCT_CORE|Pneumonia due to Pseudomonas|Pneumonia due to Pseudomonas
C0155860|T047|SY|41381004|SNOMEDCT_CORE|Pseudomonal pneumonia|Pneumonia due to Pseudomonas
C0155862|T047|SY|34020007|SNOMEDCT_CORE|Pneumonia caused by Streptococcus|Pneumonia due to Streptococcus
C0155862|T047|FN|34020007|SNOMEDCT_CORE|Pneumonia caused by Streptococcus|Pneumonia due to Streptococcus
C0155862|T047|PT|34020007|SNOMEDCT_CORE|Pneumonia due to Streptococcus|Pneumonia due to Streptococcus
C0155862|T047|OF|34020007|SNOMEDCT_CORE|Pneumonia due to Streptococcus|Pneumonia due to Streptococcus
C0155862|T047|SY|34020007|SNOMEDCT_CORE|Streptococcal pneumonia|Pneumonia due to Streptococcus
C0155870|T047|PT|195878008|SNOMEDCT_CORE|Pneumonia and influenza|Pneumonia and influenza
C0155870|T047|FN|195878008|SNOMEDCT_CORE|Pneumonia and influenza|Pneumonia and influenza
C0155871|T047|PT|61700007|SNOMEDCT_CORE|Influenza with non-respiratory manifestation|Influenza with non-respiratory manifestation
C0155871|T047|FN|61700007|SNOMEDCT_CORE|Influenza with non-respiratory manifestation|Influenza with non-respiratory manifestation
C0155871|T047|IS|61700007|SNOMEDCT_CORE|Influenza with other manifestations|Influenza with non-respiratory manifestation
C0155872|T047|IS|61937009|SNOMEDCT_CORE|Chronic catarrhal bronchitis|Simple chronic bronchitis
C0155872|T047|IS|74417001|SNOMEDCT_CORE|Chronic catarrhal bronchitis|Simple chronic bronchitis
C0155872|T047|FN|61937009|SNOMEDCT_CORE|Simple chronic bronchitis|Simple chronic bronchitis
C0155872|T047|PT|61937009|SNOMEDCT_CORE|Simple chronic bronchitis|Simple chronic bronchitis
C0155873|T047|PT|74417001|SNOMEDCT_CORE|Mucopurulent chronic bronchitis|Mucopurulent chronic bronchitis
C0155873|T047|FN|74417001|SNOMEDCT_CORE|Mucopurulent chronic bronchitis|Mucopurulent chronic bronchitis
C0155874|T047|SY|185086009|SNOMEDCT_CORE|Bronchitis with airway obstruction|Emphysematous bronchitis
C0155874|T047|SY|185086009|SNOMEDCT_CORE|Chronic bronchitis with emphysema|Emphysematous bronchitis
C0155874|T047|SY|185086009|SNOMEDCT_CORE|Chronic obstructive bronchitis|Emphysematous bronchitis
C0155874|T047|FN|185086009|SNOMEDCT_CORE|Chronic obstructive bronchitis|Emphysematous bronchitis
C0155874|T047|SY|185086009|SNOMEDCT_CORE|COB - Chronic obstructive bronchitis|Emphysematous bronchitis
C0155874|T047|PT|185086009|SNOMEDCT_CORE|Emphysematous bronchitis|Emphysematous bronchitis
C0155874|T047|SY|185086009|SNOMEDCT_CORE|Obstructive chronic bronchitis|Emphysematous bronchitis
C0155877|T047|PT|389145006|SNOMEDCT_CORE|Allergic asthma|Allergic asthma
C0155877|T047|FN|389145006|SNOMEDCT_CORE|Allergic asthma|Allergic asthma
C0155877|T047|IS|389145006|SNOMEDCT_CORE|Allergic atopic asthma|Allergic asthma
C0155877|T047|IS|389145006|SNOMEDCT_CORE|Atopic asthma|Allergic asthma
C0155880|T047|SY|266361008|SNOMEDCT_CORE|Asthma due to internal immunological process|Intrinsic asthma
C0155880|T047|PT|266361008|SNOMEDCT_CORE|Intrinsic asthma|Intrinsic asthma
C0155880|T047|SY|266361008|SNOMEDCT_CORE|Non-allergic asthma|Intrinsic asthma
C0155880|T047|FN|266361008|SNOMEDCT_CORE|Non-allergic asthma|Intrinsic asthma
C0155907|T047|PT|196102003|SNOMEDCT_CORE|Spontaneous tension pneumothorax|Spontaneous tension pneumothorax
C0155907|T047|FN|196102003|SNOMEDCT_CORE|Spontaneous tension pneumothorax|Spontaneous tension pneumothorax
C0155918|T047|PT|33325001|SNOMEDCT_CORE|Compensatory emphysema|Compensatory emphysema
C0155918|T047|FN|33325001|SNOMEDCT_CORE|Compensatory emphysema|Compensatory emphysema
C0155919|T047|SY|40541001|SNOMEDCT_CORE|Acute edema of lung|Acute pulmonary edema
C0155919|T047|IS|40541001|SNOMEDCT_CORE|Acute edema of lung, NOS|Acute pulmonary edema
C0155919|T047|SYGB|40541001|SNOMEDCT_CORE|Acute oedema of lung|Acute pulmonary edema
C0155919|T047|PT|40541001|SNOMEDCT_CORE|Acute pulmonary edema|Acute pulmonary edema
C0155919|T047|FN|40541001|SNOMEDCT_CORE|Acute pulmonary edema|Acute pulmonary edema
C0155919|T047|IS|40541001|SNOMEDCT_CORE|Acute pulmonary edema, NOS|Acute pulmonary edema
C0155919|T047|PTGB|40541001|SNOMEDCT_CORE|Acute pulmonary oedema|Acute pulmonary edema
C0155919|T047|SY|40541001|SNOMEDCT_CORE|Pulmonary edema - acute|Acute pulmonary edema
C0155919|T047|SYGB|40541001|SNOMEDCT_CORE|Pulmonary oedema - acute|Acute pulmonary edema
C0155921|T046|SY|68033004|SNOMEDCT_CORE|Disorder of tracheostomy|Tracheostomy complication
C0155921|T046|PT|68033004|SNOMEDCT_CORE|Tracheostomy complication|Tracheostomy complication
C0155921|T046|FN|68033004|SNOMEDCT_CORE|Tracheostomy complication|Tracheostomy complication
C0155921|T046|IS|68033004|SNOMEDCT_CORE|Tracheostomy complication, NOS|Tracheostomy complication
C0155922|T047|OAS|266413002|SNOMEDCT_CORE|Disorder of tooth development AND/OR eruption|Disorder of tooth development AND/OR eruption
C0155922|T047|OAS|266413002|SNOMEDCT_CORE|Teeth development and eruption disorder|Disorder of tooth development AND/OR eruption
C0155922|T047|IS|266413002|SNOMEDCT_CORE|Teeth development and eruption disorders|Disorder of tooth development AND/OR eruption
C0155922|T047|OAP|266413002|SNOMEDCT_CORE|Tooth development and eruption disorder|Disorder of tooth development AND/OR eruption
C0155922|T047|OAF|266413002|SNOMEDCT_CORE|Tooth development and eruption disorder|Disorder of tooth development AND/OR eruption
C0155922|T047|IS|266413002|SNOMEDCT_CORE|Tooth development and eruption disorders|Disorder of tooth development AND/OR eruption
C0155922|T047|OF|266413002|SNOMEDCT_CORE|Tooth development and eruption disorders|Disorder of tooth development AND/OR eruption
C0155937|T047|SY|31642005|SNOMEDCT_CORE|Acute gingival inflammation|Acute gingivitis
C0155937|T047|PT|31642005|SNOMEDCT_CORE|Acute gingivitis|Acute gingivitis
C0155937|T047|FN|31642005|SNOMEDCT_CORE|Acute gingivitis|Acute gingivitis
C0155940|T190|PT|81256000|SNOMEDCT_CORE|Anomaly of tooth position|Anomaly of tooth position
C0155940|T190|FN|81256000|SNOMEDCT_CORE|Anomaly of tooth position|Anomaly of tooth position
C0155940|T190|SY|81256000|SNOMEDCT_CORE|Malpositioned tooth|Anomaly of tooth position
C0155943|T047|PT|91943004|SNOMEDCT_CORE|Arthralgia of temporomandibular joint|Arthralgia of temporomandibular joint
C0155943|T047|FN|91943004|SNOMEDCT_CORE|Arthralgia of temporomandibular joint|Arthralgia of temporomandibular joint
C0155951|T047|PT|91950000|SNOMEDCT_CORE|Atrophy of edentulous alveolar ridge|Atrophy of edentulous alveolar ridge
C0155951|T047|FN|91950000|SNOMEDCT_CORE|Atrophy of edentulous alveolar ridge|Atrophy of edentulous alveolar ridge
C0155951|T047|SY|91950000|SNOMEDCT_CORE|Edentulous alveolar ridge atrophy|Atrophy of edentulous alveolar ridge
C0155952|T047|PT|66569006|SNOMEDCT_CORE|Retained dental root|Retained dental root
C0155952|T047|FN|66569006|SNOMEDCT_CORE|Retained dental root|Retained dental root
C0155955|T047|PT|111347003|SNOMEDCT_CORE|Exostosis of jaw|Exostosis of jaw
C0155955|T047|FN|111347003|SNOMEDCT_CORE|Exostosis of jaw|Exostosis of jaw
C0155955|T047|IS|111347003|SNOMEDCT_CORE|Exostosis of jaw, NOS|Exostosis of jaw
C0155967|T047|SY|89748001|SNOMEDCT_CORE|Acute gastric ulcer with bleeding|Acute gastric ulcer with hemorrhage
C0155967|T047|PTGB|89748001|SNOMEDCT_CORE|Acute gastric ulcer with haemorrhage|Acute gastric ulcer with hemorrhage
C0155967|T047|PT|89748001|SNOMEDCT_CORE|Acute gastric ulcer with hemorrhage|Acute gastric ulcer with hemorrhage
C0155967|T047|FN|89748001|SNOMEDCT_CORE|Acute gastric ulcer with hemorrhage|Acute gastric ulcer with hemorrhage
C0155967|T047|SY|89748001|SNOMEDCT_CORE|Bleeding acute gastric ulcer|Acute gastric ulcer with hemorrhage
C0155970|T047|PT|19850005|SNOMEDCT_CORE|Acute gastric ulcer with perforation|Acute gastric ulcer with perforation
C0155970|T047|FN|19850005|SNOMEDCT_CORE|Acute gastric ulcer with perforation|Acute gastric ulcer with perforation
C0155992|T047|PTGB|12847006|SNOMEDCT_CORE|Acute duodenal ulcer with haemorrhage|Acute duodenal ulcer with hemorrhage
C0155992|T047|PT|12847006|SNOMEDCT_CORE|Acute duodenal ulcer with hemorrhage|Acute duodenal ulcer with hemorrhage
C0155992|T047|FN|12847006|SNOMEDCT_CORE|Acute duodenal ulcer with hemorrhage|Acute duodenal ulcer with hemorrhage
C0155995|T047|PT|61347001|SNOMEDCT_CORE|Acute duodenal ulcer with perforation|Acute duodenal ulcer with perforation
C0155995|T047|FN|61347001|SNOMEDCT_CORE|Acute duodenal ulcer with perforation|Acute duodenal ulcer with perforation
C0156076|T047|PT|2043009|SNOMEDCT_CORE|Alcoholic gastritis|Alcoholic gastritis
C0156076|T047|FN|2043009|SNOMEDCT_CORE|Alcoholic gastritis|Alcoholic gastritis
C0156084|T047|PT|386211005|SNOMEDCT_CORE|Disorder of function of stomach|Disorder of function of stomach
C0156084|T047|FN|386211005|SNOMEDCT_CORE|Disorder of function of stomach|Disorder of function of stomach
C0156084|T047|SY|386211005|SNOMEDCT_CORE|Disorder of gastric function|Disorder of function of stomach
C0156084|T047|SY|386211005|SNOMEDCT_CORE|Disorder of stomach function|Disorder of function of stomach
C0156084|T047|SY|386211005|SNOMEDCT_CORE|Functional gastric disorder|Disorder of function of stomach
C0156084|T047|SY|386211005|SNOMEDCT_CORE|Functional gastric disturbance|Disorder of function of stomach
C0156092|T047|PTGB|28845006|SNOMEDCT_CORE|Acute appendicitis with generalised peritonitis|Acute appendicitis with generalized peritonitis
C0156092|T047|PT|28845006|SNOMEDCT_CORE|Acute appendicitis with generalized peritonitis|Acute appendicitis with generalized peritonitis
C0156092|T047|FN|28845006|SNOMEDCT_CORE|Acute appendicitis with generalized peritonitis|Acute appendicitis with generalized peritonitis
C0156093|T047|FN|51036000|SNOMEDCT_CORE|Acute appendicitis with peritoneal abscess|Acute appendicitis with peritoneal abscess
C0156093|T047|PT|51036000|SNOMEDCT_CORE|Acute appendicitis with peritoneal abscess|Acute appendicitis with peritoneal abscess
C0156146|T047|SY|56689002|SNOMEDCT_CORE|Crohn disease of small intestine|Crohn's disease of small intestine
C0156146|T047|PT|56689002|SNOMEDCT_CORE|Crohn's disease of small intestine|Crohn's disease of small intestine
C0156146|T047|FN|56689002|SNOMEDCT_CORE|Crohn's disease of small intestine|Crohn's disease of small intestine
C0156146|T047|SY|56689002|SNOMEDCT_CORE|Crohns disease, small intestine|Crohn's disease of small intestine
C0156146|T047|SY|56689002|SNOMEDCT_CORE|Regional enteritis of small intestine|Crohn's disease of small intestine
C0156146|T047|SY|56689002|SNOMEDCT_CORE|Regional ileitis of small intestine|Crohn's disease of small intestine
C0156146|T047|SY|56689002|SNOMEDCT_CORE|Segmental ileitis of small intestine|Crohn's disease of small intestine
C0156146|T047|IS|56689002|SNOMEDCT_CORE|Terminal ileitis of small intestine|Crohn's disease of small intestine
C0156147|T047|SY|7620006|SNOMEDCT_CORE|Crohn disease of large bowel|Crohn's disease of large bowel
C0156147|T047|PT|7620006|SNOMEDCT_CORE|Crohn's disease of large bowel|Crohn's disease of large bowel
C0156147|T047|FN|7620006|SNOMEDCT_CORE|Crohn's disease of large bowel|Crohn's disease of large bowel
C0156147|T047|SY|7620006|SNOMEDCT_CORE|Crohns disease, large intestine|Crohn's disease of large bowel
C0156147|T047|SY|7620006|SNOMEDCT_CORE|Regional enteritis of the large bowel|Crohn's disease of large bowel
C0156181|T020|SY|70190001|SNOMEDCT_CORE|Adhesive peritoneal band|Peritoneal adhesion
C0156181|T020|IS|70190001|SNOMEDCT_CORE|Adhesive peritoneal band, NOS|Peritoneal adhesion
C0156181|T020|PT|70190001|SNOMEDCT_CORE|Peritoneal adhesion|Peritoneal adhesion
C0156181|T020|FN|70190001|SNOMEDCT_CORE|Peritoneal adhesion|Peritoneal adhesion
C0156181|T020|IS|70190001|SNOMEDCT_CORE|Peritoneal adhesion, NOS|Peritoneal adhesion
C0156181|T020|SY|70190001|SNOMEDCT_CORE|Peritoneal band|Peritoneal adhesion
C0156189|T047|PT|197279005|SNOMEDCT_CORE|Cirrhosis and chronic liver disease|Cirrhosis and chronic liver disease
C0156189|T047|FN|197279005|SNOMEDCT_CORE|Cirrhosis and chronic liver disease|Cirrhosis and chronic liver disease
C0156257|T047|PT|266556005|SNOMEDCT_CORE|Calculus of kidney and ureter|Calculus of kidney and ureter
C0156257|T047|FN|266556005|SNOMEDCT_CORE|Calculus of kidney and ureter|Calculus of kidney and ureter
C0156257|T047|SY|266556005|SNOMEDCT_CORE|Calculus of kidney with calculus of ureter|Calculus of kidney and ureter
C0156270|T047|PT|11251000|SNOMEDCT_CORE|Irradiation cystitis|Irradiation cystitis
C0156270|T047|FN|11251000|SNOMEDCT_CORE|Irradiation cystitis|Irradiation cystitis
C0156270|T047|SY|11251000|SNOMEDCT_CORE|Radiation cystitis|Irradiation cystitis
C0156273|T020|SY|197866008|SNOMEDCT_CORE|Bladder diverticulum|Diverticulum of bladder
C0156273|T020|PT|197866008|SNOMEDCT_CORE|Diverticulum of bladder|Diverticulum of bladder
C0156273|T020|FN|197866008|SNOMEDCT_CORE|Diverticulum of bladder|Diverticulum of bladder
C0156284|T020|PT|111411000|SNOMEDCT_CORE|Postoperative urethral stricture|Postoperative urethral stricture
C0156284|T020|FN|111411000|SNOMEDCT_CORE|Postoperative urethral stricture|Postoperative urethral stricture
C0156309|T046|PT|198036002|SNOMEDCT_CORE|Impotence of organic origin|Impotence of organic origin
C0156309|T046|FN|198036002|SNOMEDCT_CORE|Impotence of organic origin|Impotence of organic origin
C0156309|T046|SY|198036002|SNOMEDCT_CORE|Organic erectile dysfunction|Impotence of organic origin
C0156331|T047|PT|62394006|SNOMEDCT_CORE|Female pelvic peritoneal adhesions|Female pelvic peritoneal adhesions
C0156331|T047|FN|62394006|SNOMEDCT_CORE|Female pelvic peritoneal adhesions|Female pelvic peritoneal adhesions
C0156344|T047|PT|266589005|SNOMEDCT_CORE|Endometriosis of ovary|Endometriosis of ovary
C0156344|T047|FN|266589005|SNOMEDCT_CORE|Endometriosis of ovary|Endometriosis of ovary
C0156345|T047|PT|198251001|SNOMEDCT_CORE|Endometriosis of pelvic peritoneum|Endometriosis of pelvic peritoneum
C0156345|T047|FN|198251001|SNOMEDCT_CORE|Endometriosis of pelvic peritoneum|Endometriosis of pelvic peritoneum
C0156349|T047|SY|73998008|SNOMEDCT_CORE|Female pelvic organ prolapse|Prolapse of female genital organs
C0156349|T047|SY|73998008|SNOMEDCT_CORE|Genital prolapse|Prolapse of female genital organs
C0156349|T047|IS|73998008|SNOMEDCT_CORE|Genital prolapse, NOS|Prolapse of female genital organs
C0156349|T047|PT|73998008|SNOMEDCT_CORE|Prolapse of female genital organs|Prolapse of female genital organs
C0156349|T047|FN|73998008|SNOMEDCT_CORE|Prolapse of female genital organs|Prolapse of female genital organs
C0156349|T047|IS|73998008|SNOMEDCT_CORE|Prolapse of female genital organs, NOS|Prolapse of female genital organs
C0156353|T020|PT|18973006|SNOMEDCT_CORE|Uterovaginal prolapse|Uterovaginal prolapse
C0156353|T020|FN|18973006|SNOMEDCT_CORE|Uterovaginal prolapse|Uterovaginal prolapse
C0156353|T020|IS|18973006|SNOMEDCT_CORE|Uterovaginal prolapse, NOS|Uterovaginal prolapse
C0156353|T020|SY|18973006|SNOMEDCT_CORE|Vaginal AND cervical prolapse|Uterovaginal prolapse
C0156353|T020|IS|18973006|SNOMEDCT_CORE|Vaginal and cervical prolapse|Uterovaginal prolapse
C0156354|T020|SY|42116007|SNOMEDCT_CORE|Post-hysterectomy vaginal vault prolapse|Prolapse of vaginal vault after hysterectomy
C0156354|T020|PT|42116007|SNOMEDCT_CORE|Prolapse of vaginal vault after hysterectomy|Prolapse of vaginal vault after hysterectomy
C0156354|T020|FN|42116007|SNOMEDCT_CORE|Prolapse of vaginal vault after hysterectomy|Prolapse of vaginal vault after hysterectomy
C0156367|T047|OAP|266591002|SNOMEDCT_CORE|Noninflammatory disorders of the ovary, fallopian tube and broad ligament|Noninflammatory disorders of the ovary, fallopian tube and broad ligament
C0156367|T047|OAF|266591002|SNOMEDCT_CORE|Noninflammatory disorders of the ovary, fallopian tube and broad ligament|Noninflammatory disorders of the ovary, fallopian tube and broad ligament
C0156369|T191|SY|11314008|SNOMEDCT_CORE|Intrauterine polyp|Polyp of corpus uteri
C0156369|T191|PT|11314008|SNOMEDCT_CORE|Polyp of corpus uteri|Polyp of corpus uteri
C0156369|T191|FN|11314008|SNOMEDCT_CORE|Polyp of corpus uteri|Polyp of corpus uteri
C0156369|T191|SY|11314008|SNOMEDCT_CORE|Uterine polyp|Polyp of corpus uteri
C0156377|T047|SY|198336007|SNOMEDCT_CORE|Non inflammatory disorder of cervix|Noninflammatory cervical disorder
C0156377|T047|PT|198336007|SNOMEDCT_CORE|Noninflammatory cervical disorder|Noninflammatory cervical disorder
C0156377|T047|FN|198336007|SNOMEDCT_CORE|Noninflammatory cervical disorder|Noninflammatory cervical disorder
C0156384|T046|PT|3754002|SNOMEDCT_CORE|Dysplasia of vagina|Dysplasia of vagina
C0156384|T046|FN|3754002|SNOMEDCT_CORE|Dysplasia of vagina|Dysplasia of vagina
C0156393|T047|PT|248861000|SNOMEDCT_CORE|Atrophic vulva|Atrophic vulva
C0156393|T047|FN|248861000|SNOMEDCT_CORE|Atrophic vulva|Atrophic vulva
C0156393|T047|SY|248861000|SNOMEDCT_CORE|Atrophic vulvitis|Atrophic vulva
C0156393|T047|SY|248861000|SNOMEDCT_CORE|Atrophy of vulva|Atrophic vulva
C0156404|T033|SY|80182007|SNOMEDCT_CORE|Irregular menstrual bleeding|Irregular periods
C0156404|T033|SY|80182007|SNOMEDCT_CORE|Irregular menstrual cycle|Irregular periods
C0156404|T033|SY|80182007|SNOMEDCT_CORE|Irregular menstruation|Irregular periods
C0156404|T033|PT|80182007|SNOMEDCT_CORE|Irregular periods|Irregular periods
C0156404|T033|FN|80182007|SNOMEDCT_CORE|Irregular periods|Irregular periods
C0156404|T033|SY|80182007|SNOMEDCT_CORE|Irregular uterine bleeding|Irregular periods
C0156404|T033|SY|80182007|SNOMEDCT_CORE|Menstrual periods irregular|Irregular periods
C0156404|T033|SY|80182007|SNOMEDCT_CORE|Variable menstrual cycle|Irregular periods
C0156406|T046|SY|48880000|SNOMEDCT_CORE|Bleeding after intercourse|Postcoital bleeding
C0156406|T046|SY|48880000|SNOMEDCT_CORE|PCB - Postcoital bleeding|Postcoital bleeding
C0156406|T046|PT|48880000|SNOMEDCT_CORE|Postcoital bleeding|Postcoital bleeding
C0156406|T046|FN|48880000|SNOMEDCT_CORE|Postcoital bleeding|Postcoital bleeding
C0156407|T047|PT|266677000|SNOMEDCT_CORE|Menopausal and postmenopausal disorders|Menopausal and postmenopausal disorders
C0156407|T047|FN|266677000|SNOMEDCT_CORE|Menopausal and postmenopausal disorders|Menopausal and postmenopausal disorders
C0156408|T046|OAS|88424000|SNOMEDCT_CORE|Climacteric menorrhagia|Premenopausal menorrhagia
C0156408|T046|OAS|88424000|SNOMEDCT_CORE|Excessive bleeding at onset of menopause|Premenopausal menorrhagia
C0156408|T046|OAS|88424000|SNOMEDCT_CORE|Menopausal menorrhagia|Premenopausal menorrhagia
C0156408|T046|OAS|88424000|SNOMEDCT_CORE|Preclimacteric menorrhagia|Premenopausal menorrhagia
C0156408|T046|OAP|88424000|SNOMEDCT_CORE|Premenopausal menorrhagia|Premenopausal menorrhagia
C0156408|T046|OAF|88424000|SNOMEDCT_CORE|Premenopausal menorrhagia|Premenopausal menorrhagia
C0156409|T047|SY|52441000|SNOMEDCT_CORE|Postmenopausal atrophic vaginitis|Postmenopausal atrophic vaginitis
C0156409|T047|SY|52441000|SNOMEDCT_CORE|Senile atrophic vaginitis|Postmenopausal atrophic vaginitis
C0156409|T047|SY|52441000|SNOMEDCT_CORE|Senile vaginitis|Postmenopausal atrophic vaginitis
C0156415|T047|PT|39446004|SNOMEDCT_CORE|Female infertility of tubal origin|Female infertility of tubal origin
C0156415|T047|FN|39446004|SNOMEDCT_CORE|Female infertility of tubal origin|Female infertility of tubal origin
C0156415|T047|IS|39446004|SNOMEDCT_CORE|Female infertility of tubal origin, NOS|Female infertility of tubal origin
C0156415|T047|SY|39446004|SNOMEDCT_CORE|Infertility of tubal origin|Female infertility of tubal origin
C0156604|T046|OAS|25825004|SNOMEDCT_CORE|Bleeding in early pregnancy|Hemorrhage in early pregnancy
C0156604|T046|OAS|25825004|SNOMEDCT_CORE|Haemorrhage before 22 weeks gestation|Hemorrhage in early pregnancy
C0156604|T046|IS|25825004|SNOMEDCT_CORE|Haemorrhage before 22 weeks gestation, NOS|Hemorrhage in early pregnancy
C0156604|T046|OAP|25825004|SNOMEDCT_CORE|Haemorrhage in early pregnancy|Hemorrhage in early pregnancy
C0156604|T046|IS|25825004|SNOMEDCT_CORE|Haemorrhage in early pregnancy, NOS|Hemorrhage in early pregnancy
C0156604|T046|OAS|25825004|SNOMEDCT_CORE|Hemorrhage before 22 weeks gestation|Hemorrhage in early pregnancy
C0156604|T046|IS|25825004|SNOMEDCT_CORE|Hemorrhage before 22 weeks gestation, NOS|Hemorrhage in early pregnancy
C0156604|T046|OAP|25825004|SNOMEDCT_CORE|Hemorrhage in early pregnancy|Hemorrhage in early pregnancy
C0156604|T046|OAF|25825004|SNOMEDCT_CORE|Hemorrhage in early pregnancy|Hemorrhage in early pregnancy
C0156604|T046|IS|25825004|SNOMEDCT_CORE|Hemorrhage in early pregnancy, NOS|Hemorrhage in early pregnancy
C0156617|T046|SYGB|7792000|SNOMEDCT_CORE|Low implantation of placenta without haemorrhage|Placenta previa without hemorrhage
C0156617|T046|SY|7792000|SNOMEDCT_CORE|Low implantation of placenta without hemorrhage|Placenta previa without hemorrhage
C0156617|T046|SYGB|7792000|SNOMEDCT_CORE|Placenta praevia found during pregnancy without haemorrhage|Placenta previa without hemorrhage
C0156617|T046|PTGB|7792000|SNOMEDCT_CORE|Placenta praevia without haemorrhage|Placenta previa without hemorrhage
C0156617|T046|SY|7792000|SNOMEDCT_CORE|Placenta previa found during pregnancy without hemorrhage|Placenta previa without hemorrhage
C0156617|T046|PT|7792000|SNOMEDCT_CORE|Placenta previa without hemorrhage|Placenta previa without hemorrhage
C0156617|T046|FN|7792000|SNOMEDCT_CORE|Placenta previa without hemorrhage|Placenta previa without hemorrhage
C0156621|T046|SYGB|198903000|SNOMEDCT_CORE|Haemorrhage from placenta praevia|Placenta previa with hemorrhage
C0156621|T046|IS|198903000|SNOMEDCT_CORE|Haemorrhage from placenta previa|Placenta previa with hemorrhage
C0156621|T046|SY|198903000|SNOMEDCT_CORE|Hemorrhage from placenta previa|Placenta previa with hemorrhage
C0156621|T046|PTGB|198903000|SNOMEDCT_CORE|Placenta praevia with haemorrhage|Placenta previa with hemorrhage
C0156621|T046|PT|198903000|SNOMEDCT_CORE|Placenta previa with hemorrhage|Placenta previa with hemorrhage
C0156621|T046|FN|198903000|SNOMEDCT_CORE|Placenta previa with hemorrhage|Placenta previa with hemorrhage
C0156924|T033|PT|270498000|SNOMEDCT_CORE|Malposition and malpresentation of fetus|Malposition and malpresentation of fetus
C0156924|T033|FN|270498000|SNOMEDCT_CORE|Malposition and malpresentation of fetus|Malposition and malpresentation of fetus
C0156924|T033|SY|270498000|SNOMEDCT_CORE|Malposition and malpresentation of foetus|Malposition and malpresentation of fetus
C0157063|T046|OAP|66064007|SNOMEDCT_CORE|Known OR suspected fetal abnormality affecting management of mother|Known OR suspected fetal abnormality affecting management of mother
C0157063|T046|OAF|66064007|SNOMEDCT_CORE|Known OR suspected fetal abnormality affecting management of mother|Known OR suspected fetal abnormality affecting management of mother
C0157063|T046|IS|66064007|SNOMEDCT_CORE|Known or suspected fetal abnormality affecting management of mother, NOS|Known or suspected fetal abnormality affecting management of mother, NOS
C0157063|T046|OAS|66064007|SNOMEDCT_CORE|Known OR suspected foetal abnormality affecting management of mother|Known OR suspected foetal abnormality affecting management of mother
C0157123|T046|PT|22173004|SNOMEDCT_CORE|Excessive fetal growth affecting management of mother|Excessive fetal growth affecting management of mother
C0157123|T046|FN|22173004|SNOMEDCT_CORE|Excessive fetal growth affecting management of mother|Excessive fetal growth affecting management of mother
C0157123|T046|PTGB|22173004|SNOMEDCT_CORE|Excessive foetal growth affecting management of mother|Excessive fetal growth affecting management of mother
C0157123|T046|SY|22173004|SNOMEDCT_CORE|Large for dates affecting management of mother|Excessive fetal growth affecting management of mother
C0157187|T033|PT|29399001|SNOMEDCT_CORE|Elderly primigravida|Elderly primigravida
C0157187|T033|FN|29399001|SNOMEDCT_CORE|Elderly primigravida|Elderly primigravida
C0157187|T033|SY|29399001|SNOMEDCT_CORE|Elderly primip|Elderly primigravida
C0157266|T046|PT|77259008|SNOMEDCT_CORE|Prolonged second stage of labor|Prolonged second stage of labor
C0157266|T046|FN|77259008|SNOMEDCT_CORE|Prolonged second stage of labor|Prolonged second stage of labor
C0157266|T046|PTGB|77259008|SNOMEDCT_CORE|Prolonged second stage of labour|Prolonged second stage of labor
C0157691|T047|PT|200630006|SNOMEDCT_CORE|Cellulitis and abscess of finger|Cellulitis and abscess of finger
C0157691|T047|FN|200630006|SNOMEDCT_CORE|Cellulitis and abscess of finger|Cellulitis and abscess of finger
C0157693|T047|PT|200638004|SNOMEDCT_CORE|Cellulitis and abscess of toe|Cellulitis and abscess of toe
C0157693|T047|FN|200638004|SNOMEDCT_CORE|Cellulitis and abscess of toe|Cellulitis and abscess of toe
C0157696|T047|PT|200645004|SNOMEDCT_CORE|Cellulitis and abscess of face|Cellulitis and abscess of face
C0157696|T047|FN|200645004|SNOMEDCT_CORE|Cellulitis and abscess of face|Cellulitis and abscess of face
C0157697|T047|PT|267779003|SNOMEDCT_CORE|Cellulitis and abscess of neck|Cellulitis and abscess of neck
C0157697|T047|FN|267779003|SNOMEDCT_CORE|Cellulitis and abscess of neck|Cellulitis and abscess of neck
C0157698|T047|PT|200655000|SNOMEDCT_CORE|Cellulitis and abscess of trunk|Cellulitis and abscess of trunk
C0157698|T047|FN|200655000|SNOMEDCT_CORE|Cellulitis and abscess of trunk|Cellulitis and abscess of trunk
C0157701|T047|PT|200676005|SNOMEDCT_CORE|Cellulitis and abscess of buttock|Cellulitis and abscess of buttock
C0157701|T047|FN|200676005|SNOMEDCT_CORE|Cellulitis and abscess of buttock|Cellulitis and abscess of buttock
C0157706|T047|IS|85224001|SNOMEDCT_CORE|Infected pilonidal cyst|Infected pilonidal sinus
C0157706|T047|IS|85224001|SNOMEDCT_CORE|Infected pilonidal sinus|Infected pilonidal sinus
C0157721|T047|SY|34250006|SNOMEDCT_CORE|Ocular pemphigoid|Ocular pemphigoid
C0157726|T020|OAS|201037000|SNOMEDCT_CORE|Corns and callosities|Corns and callosities
C0157726|T020|OAP|201037000|SNOMEDCT_CORE|Corns and callus|Corns and callosities
C0157726|T020|OAF|201037000|SNOMEDCT_CORE|Corns and callus|Corns and callosities
C0157738|T047|SY|19429009|SNOMEDCT_CORE|Chronic skin ulcer|Chronic ulcer of skin
C0157738|T047|PT|19429009|SNOMEDCT_CORE|Chronic ulcer of skin|Chronic ulcer of skin
C0157738|T047|FN|19429009|SNOMEDCT_CORE|Chronic ulcer of skin|Chronic ulcer of skin
C0157738|T047|IS|19429009|SNOMEDCT_CORE|Chronic ulcer of skin, NOS|Chronic ulcer of skin
C0157741|T047|SYGB|42265009|SNOMEDCT_CORE|Idiopathic angio-oedema-urticaria|Idiopathic urticaria
C0157741|T047|SY|42265009|SNOMEDCT_CORE|Idiopathic angioedema-urticaria|Idiopathic urticaria
C0157741|T047|PT|42265009|SNOMEDCT_CORE|Idiopathic urticaria|Idiopathic urticaria
C0157741|T047|FN|42265009|SNOMEDCT_CORE|Idiopathic urticaria|Idiopathic urticaria
C0157917|T047|SY|74391003|SNOMEDCT_CORE|JCA - Pauciarticular onset juvenile chronic arthritis|Pauciarticular juvenile rheumatoid arthritis
C0157917|T047|PT|74391003|SNOMEDCT_CORE|Pauciarticular juvenile rheumatoid arthritis|Pauciarticular juvenile rheumatoid arthritis
C0157917|T047|FN|74391003|SNOMEDCT_CORE|Pauciarticular juvenile rheumatoid arthritis|Pauciarticular juvenile rheumatoid arthritis
C0157917|T047|SY|74391003|SNOMEDCT_CORE|Pauciarticular onset juvenile arthritis|Pauciarticular juvenile rheumatoid arthritis
C0157917|T047|SY|74391003|SNOMEDCT_CORE|Pauciarticular onset juvenile chronic arthritis|Pauciarticular juvenile rheumatoid arthritis
C0158026|T047|OAS|220000|SNOMEDCT_CORE|Monoarthritis|Monoarthritis
C0158026|T047|PT|699462004|SNOMEDCT_CORE|Monoarthritis|Monoarthritis
C0158026|T047|FN|699462004|SNOMEDCT_CORE|Monoarthritis|Monoarthritis
C0158026|T047|IS|220000|SNOMEDCT_CORE|Monoarthritis, NOS|Monoarthritis
C0158026|T047|OAP|220000|SNOMEDCT_CORE|Unspecified monoarthritis|Monoarthritis
C0158026|T047|OAF|220000|SNOMEDCT_CORE|Unspecified monoarthritis|Monoarthritis
C0158053|T047|PT|63643000|SNOMEDCT_CORE|Derangement of knee|Derangement of knee
C0158053|T047|FN|63643000|SNOMEDCT_CORE|Derangement of knee|Derangement of knee
C0158053|T047|IS|63643000|SNOMEDCT_CORE|Derangement of knee, NOS|Derangement of knee
C0158053|T047|SY|63643000|SNOMEDCT_CORE|IDK - Internal derangement of knee joint|Derangement of knee
C0158053|T047|SY|63643000|SNOMEDCT_CORE|Internal derangement of knee|Derangement of knee
C0158053|T047|SY|63643000|SNOMEDCT_CORE|Internal derangement of knee joint|Derangement of knee
C0158053|T047|IS|63643000|SNOMEDCT_CORE|Internal derangement of knee, NOS|Derangement of knee
C0158054|T033|PT|86378006|SNOMEDCT_CORE|Old bucket handle tear of medial meniscus|Old bucket handle tear of medial meniscus
C0158054|T033|FN|86378006|SNOMEDCT_CORE|Old bucket handle tear of medial meniscus|Old bucket handle tear of medial meniscus
C0158056|T037|PT|5313005|SNOMEDCT_CORE|Derangement of posterior horn of medial meniscus|Derangement of posterior horn of medial meniscus
C0158056|T037|FN|5313005|SNOMEDCT_CORE|Derangement of posterior horn of medial meniscus|Derangement of posterior horn of medial meniscus
C0158056|T037|SY|5313005|SNOMEDCT_CORE|Medial meniscus, posterior horn derangement|Derangement of posterior horn of medial meniscus
C0158058|T037|PT|21333004|SNOMEDCT_CORE|Derangement of lateral meniscus|Derangement of lateral meniscus
C0158058|T037|FN|21333004|SNOMEDCT_CORE|Derangement of lateral meniscus|Derangement of lateral meniscus
C0158058|T037|SY|21333004|SNOMEDCT_CORE|Derangement of lateral meniscus of knee|Derangement of lateral meniscus
C0158058|T037|IS|21333004|SNOMEDCT_CORE|Derangement of lateral meniscus, NOS|Derangement of lateral meniscus
C0158058|T037|SY|21333004|SNOMEDCT_CORE|Lateral meniscus derangement|Derangement of lateral meniscus
C0158061|T037|PT|77860008|SNOMEDCT_CORE|Derangement of posterior horn of lateral meniscus|Derangement of posterior horn of lateral meniscus
C0158061|T037|FN|77860008|SNOMEDCT_CORE|Derangement of posterior horn of lateral meniscus|Derangement of posterior horn of lateral meniscus
C0158061|T037|SY|77860008|SNOMEDCT_CORE|Lateral meniscus, posterior horn derangement|Derangement of posterior horn of lateral meniscus
C0158067|T037|SY|202109007|SNOMEDCT_CORE|Old disruption of medial collateral ligament|Old medial collateral ligament disruption
C0158067|T037|PT|202109007|SNOMEDCT_CORE|Old medial collateral ligament disruption|Old medial collateral ligament disruption
C0158067|T037|FN|202109007|SNOMEDCT_CORE|Old medial collateral ligament disruption|Old medial collateral ligament disruption
C0158068|T037|PT|202110002|SNOMEDCT_CORE|Old anterior cruciate ligament disruption|Old anterior cruciate ligament disruption
C0158068|T037|FN|202110002|SNOMEDCT_CORE|Old anterior cruciate ligament disruption|Old anterior cruciate ligament disruption
C0158068|T037|SY|202110002|SNOMEDCT_CORE|Old disruption of anterior cruciate ligament|Old anterior cruciate ligament disruption
C0158073|T047|SY|53417006|SNOMEDCT_CORE|Articular cartilage disease|Articular cartilage disorder
C0158073|T047|IS|53417006|SNOMEDCT_CORE|Articular cartilage disease, NOS|Articular cartilage disorder
C0158073|T047|PT|53417006|SNOMEDCT_CORE|Articular cartilage disorder|Articular cartilage disorder
C0158073|T047|FN|53417006|SNOMEDCT_CORE|Articular cartilage disorder|Articular cartilage disorder
C0158073|T047|IS|53417006|SNOMEDCT_CORE|Articular cartilage disorder, NOS|Articular cartilage disorder
C0158073|T047|SY|53417006|SNOMEDCT_CORE|Disorder of articular cartilage|Articular cartilage disorder
C0158110|T020|PT|90116003|SNOMEDCT_CORE|Contracture of joint of shoulder region|Contracture of joint of shoulder region
C0158110|T020|FN|90116003|SNOMEDCT_CORE|Contracture of joint of shoulder region|Contracture of joint of shoulder region
C0158110|T020|SY|90116003|SNOMEDCT_CORE|Contracture of shoulder joint|Contracture of joint of shoulder region
C0158110|T020|SY|90116003|SNOMEDCT_CORE|Joint contracture of shoulder|Contracture of joint of shoulder region
C0158113|T190|SY|86414002|SNOMEDCT_CORE|Contracture of hand joint|Contracture of joint of hand
C0158113|T190|PT|86414002|SNOMEDCT_CORE|Contracture of joint of hand|Contracture of joint of hand
C0158113|T190|FN|86414002|SNOMEDCT_CORE|Contracture of joint of hand|Contracture of joint of hand
C0158113|T190|SY|86414002|SNOMEDCT_CORE|Joint contracture of hand|Contracture of joint of hand
C0158118|T020|PT|202264009|SNOMEDCT_CORE|Contracture of multiple joints|Contracture of multiple joints
C0158118|T020|FN|202264009|SNOMEDCT_CORE|Contracture of multiple joints|Contracture of multiple joints
C0158241|T047|PT|267970006|SNOMEDCT_CORE|Cervical spondylosis without myelopathy|Cervical spondylosis without myelopathy
C0158241|T047|FN|267970006|SNOMEDCT_CORE|Cervical spondylosis without myelopathy|Cervical spondylosis without myelopathy
C0158242|T047|SY|65260001|SNOMEDCT_CORE|Cervical spinal cord compression|Cervical spondylosis with myelopathy
C0158242|T047|SY|65260001|SNOMEDCT_CORE|Cervical spondylitic cord compression|Cervical spondylosis with myelopathy
C0158242|T047|PT|65260001|SNOMEDCT_CORE|Cervical spondylosis with myelopathy|Cervical spondylosis with myelopathy
C0158242|T047|FN|65260001|SNOMEDCT_CORE|Cervical spondylosis with myelopathy|Cervical spondylosis with myelopathy
C0158242|T047|SY|65260001|SNOMEDCT_CORE|Spondylogenic compression of cervical spinal cord|Cervical spondylosis with myelopathy
C0158243|T047|SY|267971005|SNOMEDCT_CORE|Dorsal spondylosis without myelopathy|Thoracic spondylosis without myelopathy
C0158243|T047|PT|267971005|SNOMEDCT_CORE|Thoracic spondylosis without myelopathy|Thoracic spondylosis without myelopathy
C0158243|T047|FN|267971005|SNOMEDCT_CORE|Thoracic spondylosis without myelopathy|Thoracic spondylosis without myelopathy
C0158244|T047|PT|48210000|SNOMEDCT_CORE|Lumbosacral spondylosis without myelopathy|Lumbosacral spondylosis without myelopathy
C0158244|T047|FN|48210000|SNOMEDCT_CORE|Lumbosacral spondylosis without myelopathy|Lumbosacral spondylosis without myelopathy
C0158247|T047|PT|67437007|SNOMEDCT_CORE|Lumbar spondylosis with myelopathy|Lumbar spondylosis with myelopathy
C0158247|T047|FN|67437007|SNOMEDCT_CORE|Lumbar spondylosis with myelopathy|Lumbar spondylosis with myelopathy
C0158247|T047|SY|67437007|SNOMEDCT_CORE|Spondylogenic compression of lumbar spinal cord|Lumbar spondylosis with myelopathy
C0158252|T047|SY|36427004|SNOMEDCT_CORE|Disorder of intervertebral disc|Intervertebral disc disorder
C0158252|T047|PT|36427004|SNOMEDCT_CORE|Intervertebral disc disorder|Intervertebral disc disorder
C0158252|T047|FN|36427004|SNOMEDCT_CORE|Intervertebral disc disorder|Intervertebral disc disorder
C0158252|T047|IS|36427004|SNOMEDCT_CORE|Intervertebral disc disorder, NOS|Intervertebral disc disorder
C0158253|T047|PT|85216006|SNOMEDCT_CORE|Displacement of cervical intervertebral disc without myelopathy|Displacement of cervical intervertebral disc without myelopathy
C0158253|T047|FN|85216006|SNOMEDCT_CORE|Displacement of cervical intervertebral disc without myelopathy|Displacement of cervical intervertebral disc without myelopathy
C0158255|T047|PT|20021007|SNOMEDCT_CORE|Displacement of lumbar intervertebral disc without myelopathy|Displacement of lumbar intervertebral disc without myelopathy
C0158255|T047|FN|20021007|SNOMEDCT_CORE|Displacement of lumbar intervertebral disc without myelopathy|Displacement of lumbar intervertebral disc without myelopathy
C0158262|T047|PT|69195002|SNOMEDCT_CORE|Degeneration of cervical intervertebral disc|Degeneration of cervical intervertebral disc
C0158262|T047|FN|69195002|SNOMEDCT_CORE|Degeneration of cervical intervertebral disc|Degeneration of cervical intervertebral disc
C0158266|T047|PT|77547008|SNOMEDCT_CORE|Degeneration of intervertebral disc|Degeneration of intervertebral disc
C0158266|T047|FN|77547008|SNOMEDCT_CORE|Degeneration of intervertebral disc|Degeneration of intervertebral disc
C0158266|T047|IS|77547008|SNOMEDCT_CORE|Degeneration of intervertebral disc, NOS|Degeneration of intervertebral disc
C0158266|T047|SY|77547008|SNOMEDCT_CORE|Degenerative disc disease|Degeneration of intervertebral disc
C0158266|T047|IS|77547008|SNOMEDCT_CORE|Degenerative disc disease, NOS|Degeneration of intervertebral disc
C0158266|T047|SY|77547008|SNOMEDCT_CORE|Intervertebral disc degeneration|Degeneration of intervertebral disc
C0158268|T047|PT|75467001|SNOMEDCT_CORE|Intervertebral disc disorder of cervical region with myelopathy|Intervertebral disc disorder of cervical region with myelopathy
C0158268|T047|FN|75467001|SNOMEDCT_CORE|Intervertebral disc disorder of cervical region with myelopathy|Intervertebral disc disorder of cervical region with myelopathy
C0158270|T047|SY|34139004|SNOMEDCT_CORE|Disorder of lumbar intervertebral disc with myelopathy|Intervertebral disc disorder of lumbar region with myelopathy
C0158270|T047|PT|34139004|SNOMEDCT_CORE|Intervertebral disc disorder of lumbar region with myelopathy|Intervertebral disc disorder of lumbar region with myelopathy
C0158270|T047|FN|34139004|SNOMEDCT_CORE|Intervertebral disc disorder of lumbar region with myelopathy|Intervertebral disc disorder of lumbar region with myelopathy
C0158272|T047|PT|202723000|SNOMEDCT_CORE|Cervical post-laminectomy syndrome|Cervical post-laminectomy syndrome
C0158272|T047|FN|202723000|SNOMEDCT_CORE|Cervical post-laminectomy syndrome|Cervical post-laminectomy syndrome
C0158274|T047|PT|202725007|SNOMEDCT_CORE|Lumbar post-laminectomy syndrome|Lumbar post-laminectomy syndrome
C0158274|T047|FN|202725007|SNOMEDCT_CORE|Lumbar post-laminectomy syndrome|Lumbar post-laminectomy syndrome
C0158280|T047|SY|83561009|SNOMEDCT_CORE|Cervical spinal stenosis|Spinal stenosis in cervical region
C0158280|T047|PT|83561009|SNOMEDCT_CORE|Spinal stenosis in cervical region|Spinal stenosis in cervical region
C0158280|T047|FN|83561009|SNOMEDCT_CORE|Spinal stenosis in cervical region|Spinal stenosis in cervical region
C0158288|T047|SY|18347007|SNOMEDCT_CORE|Lumbar spinal stenosis|Spinal stenosis of lumbar region
C0158288|T047|PT|18347007|SNOMEDCT_CORE|Spinal stenosis of lumbar region|Spinal stenosis of lumbar region
C0158288|T047|FN|18347007|SNOMEDCT_CORE|Spinal stenosis of lumbar region|Spinal stenosis of lumbar region
C0158292|T047|PT|12820001|SNOMEDCT_CORE|Disorder of sacrum|Disorder of sacrum
C0158292|T047|FN|12820001|SNOMEDCT_CORE|Disorder of sacrum|Disorder of sacrum
C0158292|T047|IS|12820001|SNOMEDCT_CORE|Disorder of sacrum, NOS|Disorder of sacrum
C0158301|T047|OAP|202838007|SNOMEDCT_CORE|Rotator cuff shoulder syndrome and allied disorders|Rotator cuff shoulder syndrome and allied disorders
C0158301|T047|OAF|202838007|SNOMEDCT_CORE|Rotator cuff shoulder syndrome and allied disorders|Rotator cuff shoulder syndrome and allied disorders
C0158303|T047|PT|27741009|SNOMEDCT_CORE|Calcific tendinitis of shoulder|Calcific tendinitis of shoulder
C0158303|T047|FN|27741009|SNOMEDCT_CORE|Calcific tendinitis of shoulder|Calcific tendinitis of shoulder
C0158303|T047|SY|27741009|SNOMEDCT_CORE|Calcific tendonitis of shoulder|Calcific tendinitis of shoulder
C0158303|T047|SY|27741009|SNOMEDCT_CORE|Calcifying tendinitis of shoulder|Calcific tendinitis of shoulder
C0158303|T047|SY|27741009|SNOMEDCT_CORE|Calcifying tendinitis of the shoulder|Calcific tendinitis of shoulder
C0158303|T047|IS|27741009|SNOMEDCT_CORE|Milwaukee shoulder|Calcific tendinitis of shoulder
C0158309|T020|IS|53286005|SNOMEDCT_CORE|Golfer's elbow|Medial epicondylitis
C0158309|T020|PT|53286005|SNOMEDCT_CORE|Medial epicondylitis|Medial epicondylitis
C0158309|T020|SY|53286005|SNOMEDCT_CORE|Medial epicondylitis of elbow|Medial epicondylitis
C0158309|T020|FN|53286005|SNOMEDCT_CORE|Medial epicondylitis of elbow joint|Medial epicondylitis
C0158309|T020|SY|53286005|SNOMEDCT_CORE|Medial epicondylitis of elbow joint|Medial epicondylitis
C0158311|T047|IS|33439002|SNOMEDCT_CORE|Enthesopathy of wrist and carpus, NOS|Enthesopathy of wrist AND/OR carpus
C0158311|T047|PT|33439002|SNOMEDCT_CORE|Enthesopathy of wrist AND/OR carpus|Enthesopathy of wrist AND/OR carpus
C0158311|T047|FN|33439002|SNOMEDCT_CORE|Enthesopathy of wrist AND/OR carpus|Enthesopathy of wrist AND/OR carpus
C0158317|T047|PT|37785001|SNOMEDCT_CORE|Patellar tendonitis|Patellar tendonitis
C0158317|T047|FN|37785001|SNOMEDCT_CORE|Patellar tendonitis|Patellar tendonitis
C0158319|T047|IS|21409006|SNOMEDCT_CORE|Enthesopathy of ankle and tarsus, NOS|Enthesopathy of ankle AND/OR tarsus
C0158319|T047|PT|21409006|SNOMEDCT_CORE|Enthesopathy of ankle AND/OR tarsus|Enthesopathy of ankle AND/OR tarsus
C0158319|T047|FN|21409006|SNOMEDCT_CORE|Enthesopathy of ankle AND/OR tarsus|Enthesopathy of ankle AND/OR tarsus
C0158321|T047|PT|50127006|SNOMEDCT_CORE|Tibialis tendinitis|Tibialis tendinitis
C0158321|T047|FN|50127006|SNOMEDCT_CORE|Tibialis tendinitis|Tibialis tendinitis
C0158321|T047|IS|50127006|SNOMEDCT_CORE|Tibialis tendinitis, NOS|Tibialis tendinitis
C0158321|T047|SY|50127006|SNOMEDCT_CORE|Tibialis tendonitis|Tibialis tendinitis
C0158322|T047|PT|55260003|SNOMEDCT_CORE|Calcaneal spur|Calcaneal spur
C0158322|T047|FN|55260003|SNOMEDCT_CORE|Calcaneal spur|Calcaneal spur
C0158322|T047|OF|55260003|SNOMEDCT_CORE|Calcaneal spur|Calcaneal spur
C0158334|T047|SY|78435003|SNOMEDCT_CORE|Ganglion cyst of joint|Ganglion of joint
C0158334|T047|PT|78435003|SNOMEDCT_CORE|Ganglion of joint|Ganglion of joint
C0158334|T047|FN|78435003|SNOMEDCT_CORE|Ganglion of joint|Ganglion of joint
C0158334|T047|IS|78435003|SNOMEDCT_CORE|Ganglion of joint, NOS|Ganglion of joint
C0158335|T020|PT|19354008|SNOMEDCT_CORE|Ganglion cyst of tendon sheath|Ganglion cyst of tendon sheath
C0158335|T020|FN|19354008|SNOMEDCT_CORE|Ganglion cyst of tendon sheath|Ganglion cyst of tendon sheath
C0158335|T020|SY|19354008|SNOMEDCT_CORE|Ganglion of tendon sheath|Ganglion cyst of tendon sheath
C0158335|T020|OF|19354008|SNOMEDCT_CORE|Ganglion of tendon sheath|Ganglion cyst of tendon sheath
C0158335|T020|IS|19354008|SNOMEDCT_CORE|Ganglion of tendon sheath, NOS|Ganglion cyst of tendon sheath
C0158347|T037|PT|202964000|SNOMEDCT_CORE|Non-traumatic rupture of Achilles tendon|Non-traumatic rupture of Achilles tendon
C0158347|T037|FN|202964000|SNOMEDCT_CORE|Non-traumatic rupture of Achilles tendon|Non-traumatic rupture of Achilles tendon
C0158350|T046|PT|274141009|SNOMEDCT_CORE|Tendon contracture|Tendon contracture
C0158350|T046|FN|274141009|SNOMEDCT_CORE|Tendon contracture|Tendon contracture
C0158360|T047|SY|13370002|SNOMEDCT_CORE|Dupuytren disease of foot|Plantar fascial fibromatosis
C0158360|T047|IS|13370002|SNOMEDCT_CORE|Dupuytren's contracture of foot|Plantar fascial fibromatosis
C0158360|T047|SY|13370002|SNOMEDCT_CORE|Ledderhose's disease|Plantar fascial fibromatosis
C0158360|T047|PT|13370002|SNOMEDCT_CORE|Plantar fascial fibromatosis|Plantar fascial fibromatosis
C0158360|T047|FN|13370002|SNOMEDCT_CORE|Plantar fascial fibromatosis|Plantar fascial fibromatosis
C0158360|T047|IS|202882003|SNOMEDCT_CORE|Plantar fascial fibromatosis|Plantar fascial fibromatosis
C0158360|T047|SY|13370002|SNOMEDCT_CORE|Plantar fibromatosis|Plantar fascial fibromatosis
C0158364|T190|PT|111248006|SNOMEDCT_CORE|Diastasis of muscle|Diastasis of muscle
C0158364|T190|FN|111248006|SNOMEDCT_CORE|Diastasis of muscle|Diastasis of muscle
C0158364|T190|IS|111248006|SNOMEDCT_CORE|Diastasis of muscle, NOS|Diastasis of muscle
C0158368|T020|PT|6058003|SNOMEDCT_CORE|Residual foreign body in soft tissue|Residual foreign body in soft tissue
C0158368|T020|FN|6058003|SNOMEDCT_CORE|Residual foreign body in soft tissue|Residual foreign body in soft tissue
C0158369|T184|PT|80068009|SNOMEDCT_CORE|Swelling of limb|Swelling of limb
C0158369|T184|FN|80068009|SNOMEDCT_CORE|Swelling of limb|Swelling of limb
C0158369|T184|IS|80068009|SNOMEDCT_CORE|Swelling of limb, NOS|Swelling of limb
C0158371|T047|PT|409780002|SNOMEDCT_CORE|Acute osteomyelitis|Acute osteomyelitis
C0158371|T047|FN|409780002|SNOMEDCT_CORE|Acute osteomyelitis|Acute osteomyelitis
C0158441|T037|SY|26460006|SNOMEDCT_CORE|Non-traumatic slipped upper femoral epiphysis|Slipped upper femoral epiphysis
C0158441|T037|SY|26460006|SNOMEDCT_CORE|Nontraumatic slipped upper femoral epiphysis|Slipped upper femoral epiphysis
C0158441|T037|IS|26460006|SNOMEDCT_CORE|Nontraumatic slipped upper femoral epiphysis, NOS|Slipped upper femoral epiphysis
C0158441|T037|SY|26460006|SNOMEDCT_CORE|Slipped femoral epiphysis|Slipped upper femoral epiphysis
C0158441|T037|IS|26460006|SNOMEDCT_CORE|Slipped femoral epiphysis, NOS|Slipped upper femoral epiphysis
C0158441|T037|PT|26460006|SNOMEDCT_CORE|Slipped upper femoral epiphysis|Slipped upper femoral epiphysis
C0158441|T037|FN|26460006|SNOMEDCT_CORE|Slipped upper femoral epiphysis|Slipped upper femoral epiphysis
C0158441|T037|IS|26460006|SNOMEDCT_CORE|Slipped upper femoral epiphysis, NOS|Slipped upper femoral epiphysis
C0158441|T037|SY|26460006|SNOMEDCT_CORE|SUFE - Slipped upper femoral epiphysis|Slipped upper femoral epiphysis
C0158447|T047|PT|3345002|SNOMEDCT_CORE|Idiopathic osteoporosis|Idiopathic osteoporosis
C0158447|T047|FN|3345002|SNOMEDCT_CORE|Idiopathic osteoporosis|Idiopathic osteoporosis
C0158454|T046|PT|425852005|SNOMEDCT_CORE|Fracture malunion|Fracture malunion
C0158454|T046|FN|425852005|SNOMEDCT_CORE|Fracture malunion|Fracture malunion
C0158454|T046|SY|425852005|SNOMEDCT_CORE|Malunion of fracture|Fracture malunion
C0158458|T020|PT|65358001|SNOMEDCT_CORE|Acquired hallux valgus|Acquired hallux valgus
C0158458|T020|FN|65358001|SNOMEDCT_CORE|Acquired hallux valgus|Acquired hallux valgus
C0158473|T020|FN|64298006|SNOMEDCT_CORE|Acquired deformity of distal interphalangeal joint of finger due to trauma|Mallet finger
C0158473|T020|SY|64298006|SNOMEDCT_CORE|Acquired deformity of distal interphalangeal joint of finger due to trauma|Mallet finger
C0158473|T020|SY|64298006|SNOMEDCT_CORE|Acquired deformity of finger due to trauma|Mallet finger
C0158473|T020|OF|64298006|SNOMEDCT_CORE|Acquired deformity of finger due to trauma|Mallet finger
C0158473|T020|SY|64298006|SNOMEDCT_CORE|Baseball finger|Mallet finger
C0158473|T020|PT|64298006|SNOMEDCT_CORE|Mallet finger|Mallet finger
C0158473|T020|OF|64298006|SNOMEDCT_CORE|Mallet finger|Mallet finger
C0158478|T020|PT|67321002|SNOMEDCT_CORE|Acquired deformity of hip|Acquired deformity of hip
C0158478|T020|FN|67321002|SNOMEDCT_CORE|Acquired deformity of hip|Acquired deformity of hip
C0158478|T020|IS|67321002|SNOMEDCT_CORE|Acquired deformity of hip, NOS|Acquired deformity of hip
C0158484|T020|PT|52012001|SNOMEDCT_CORE|Acquired genu valgum|Acquired genu valgum
C0158484|T020|FN|52012001|SNOMEDCT_CORE|Acquired genu valgum|Acquired genu valgum
C0158484|T020|SY|52012001|SNOMEDCT_CORE|Acquired knock knee|Acquired genu valgum
C0158484|T020|SY|52012001|SNOMEDCT_CORE|Acquired knock-knee|Acquired genu valgum
C0158484|T020|SY|52012001|SNOMEDCT_CORE|Acquired valgus deformity of knee|Acquired genu valgum
C0158484|T020|IS|52012001|SNOMEDCT_CORE|Knock-knees - acquired|Acquired genu valgum
C0158493|T020|PT|65362007|SNOMEDCT_CORE|Acquired cavovarus deformity of foot|Acquired cavovarus deformity of foot
C0158493|T020|FN|65362007|SNOMEDCT_CORE|Acquired cavovarus deformity of foot|Acquired cavovarus deformity of foot
C0158493|T020|SY|65362007|SNOMEDCT_CORE|Acquired cavovarus foot deformity|Acquired cavovarus deformity of foot
C0158513|T020|PT|245867000|SNOMEDCT_CORE|Acquired spondylolysis|Acquired spondylolysis
C0158513|T020|FN|245867000|SNOMEDCT_CORE|Acquired spondylolysis|Acquired spondylolysis
C0158598|T047|OAP|204270004|SNOMEDCT_CORE|Preauricular sinus and fistula|Preauricular sinus and fistula
C0158598|T047|OAF|204270004|SNOMEDCT_CORE|Preauricular sinus and fistula|Preauricular sinus and fistula
C0158621|T019|PT|73660006|SNOMEDCT_CORE|Congenital subaortic stenosis|Congenital subaortic stenosis
C0158621|T019|FN|73660006|SNOMEDCT_CORE|Congenital subaortic stenosis|Congenital subaortic stenosis
C0158621|T019|SY|73660006|SNOMEDCT_CORE|Congenital subvalvular aortic stenosis|Congenital subaortic stenosis
C0158638|T019|SY|65587001|SNOMEDCT_CORE|Congenital anomaly of cerebral vessels|Congenital anomaly of cerebrovascular system
C0158638|T019|IS|65587001|SNOMEDCT_CORE|Congenital anomaly of cerebral vessels, NOS|Congenital anomaly of cerebrovascular system
C0158638|T019|PT|65587001|SNOMEDCT_CORE|Congenital anomaly of cerebrovascular system|Congenital anomaly of cerebrovascular system
C0158638|T019|FN|65587001|SNOMEDCT_CORE|Congenital anomaly of cerebrovascular system|Congenital anomaly of cerebrovascular system
C0158638|T019|IS|65587001|SNOMEDCT_CORE|Congenital anomaly of cerebrovascular system, NOS|Congenital anomaly of cerebrovascular system
C0158646|T019|SY|66948001|SNOMEDCT_CORE|Cleft palate and lip|Cleft palate with cleft lip
C0158646|T019|PT|66948001|SNOMEDCT_CORE|Cleft palate with cleft lip|Cleft palate with cleft lip
C0158646|T019|FN|66948001|SNOMEDCT_CORE|Cleft palate with cleft lip|Cleft palate with cleft lip
C0158646|T019|IS|66948001|SNOMEDCT_CORE|Cleft palate with cleft lip, NOS|Cleft palate with cleft lip
C0158655|T019|OAP|204612005|SNOMEDCT_CORE|Unilateral complete cleft palate with cleft lip|Unilateral complete cleft palate with cleft lip
C0158655|T019|OF|204612005|SNOMEDCT_CORE|Unilateral complete cleft palate with cleft lip|Unilateral complete cleft palate with cleft lip
C0158655|T019|OAF|204612005|SNOMEDCT_CORE|Unilateral complete cleft palate with cleft lip|Unilateral complete cleft palate with cleft lip
C0158683|T047|PT|72925005|SNOMEDCT_CORE|Congenital cystic disease of liver|Congenital cystic disease of liver
C0158683|T047|FN|72925005|SNOMEDCT_CORE|Congenital cystic disease of liver|Congenital cystic disease of liver
C0158683|T047|SY|72925005|SNOMEDCT_CORE|Congenital cystic liver|Congenital cystic disease of liver
C0158683|T047|SY|72925005|SNOMEDCT_CORE|Congenital hepatic cyst|Congenital cystic disease of liver
C0158683|T047|SY|72925005|SNOMEDCT_CORE|Congenital polycystic disease of liver|Congenital cystic disease of liver
C0158683|T047|SY|72925005|SNOMEDCT_CORE|Congenital polycystic liver disease|Congenital cystic disease of liver
C0158683|T047|SY|72925005|SNOMEDCT_CORE|Cystic disease of liver|Congenital cystic disease of liver
C0158683|T047|SY|72925005|SNOMEDCT_CORE|Fibrocystic disease of liver|Congenital cystic disease of liver
C0158683|T047|SY|72925005|SNOMEDCT_CORE|Fibrocystic liver disease|Congenital cystic disease of liver
C0158683|T047|SY|72925005|SNOMEDCT_CORE|PLD - Polycystic liver disease|Congenital cystic disease of liver
C0158683|T047|SY|72925005|SNOMEDCT_CORE|Polycystic liver disease|Congenital cystic disease of liver
C0158687|T019|SY|204821009|SNOMEDCT_CORE|Congenital anomaly of genital organ|Congenital malformation of genital organs
C0158687|T019|SY|204821009|SNOMEDCT_CORE|Congenital deformity of genital organ|Congenital malformation of genital organs
C0158687|T019|SY|204821009|SNOMEDCT_CORE|Congenital genital organ anomalies|Congenital malformation of genital organs
C0158687|T019|PT|204821009|SNOMEDCT_CORE|Congenital malformation of genital organs|Congenital malformation of genital organs
C0158687|T019|FN|204821009|SNOMEDCT_CORE|Congenital malformation of genital organs|Congenital malformation of genital organs
C0158775|T019|PT|74877002|SNOMEDCT_CORE|Congenital anomaly of spine|Congenital anomaly of spine
C0158775|T019|FN|74877002|SNOMEDCT_CORE|Congenital anomaly of spine|Congenital anomaly of spine
C0158775|T019|IS|74877002|SNOMEDCT_CORE|Congenital anomaly of spine, NOS|Congenital anomaly of spine
C0158775|T019|SY|74877002|SNOMEDCT_CORE|Congenital anomaly of vertebral column|Congenital anomaly of spine
C0158775|T019|IS|74877002|SNOMEDCT_CORE|Congenital anomaly of vertebral column, NOS|Congenital anomaly of spine
C0158775|T019|SY|74877002|SNOMEDCT_CORE|Congenital malformation of spine|Congenital anomaly of spine
C0158775|T019|SY|74877002|SNOMEDCT_CORE|Congenital spine malformation|Congenital anomaly of spine
C0158775|T019|IS|74877002|SNOMEDCT_CORE|Congenital spine malformation, NOS|Congenital anomaly of spine
C0158816|T046|IS|68983007|SNOMEDCT_CORE|Complication of pregnancy affecting fetus OR newborn|Fetal or neonatal effect of maternal complication of pregnancy
C0158816|T046|PT|206035009|SNOMEDCT_CORE|Fetal or neonatal effect of maternal complication of pregnancy|Fetal or neonatal effect of maternal complication of pregnancy
C0158816|T046|FN|206035009|SNOMEDCT_CORE|Fetal or neonatal effect of maternal complication of pregnancy|Fetal or neonatal effect of maternal complication of pregnancy
C0158816|T046|OAP|68983007|SNOMEDCT_CORE|Fetal or neonatal effects of maternal complication of pregnancy|Fetal or neonatal effect of maternal complication of pregnancy
C0158816|T046|OAF|68983007|SNOMEDCT_CORE|Fetal or neonatal effects of maternal complication of pregnancy|Fetal or neonatal effect of maternal complication of pregnancy
C0158816|T046|OP|206035009|SNOMEDCT_CORE|Fetus or neonate affected by maternal complication of pregnancy|Fetal or neonatal effect of maternal complication of pregnancy
C0158816|T046|OF|206035009|SNOMEDCT_CORE|Fetus or neonate affected by maternal complication of pregnancy|Fetal or neonatal effect of maternal complication of pregnancy
C0158816|T046|OP|68983007|SNOMEDCT_CORE|Fetus OR newborn affected by maternal complication of pregnancy|Fetal or neonatal effect of maternal complication of pregnancy
C0158816|T046|OF|68983007|SNOMEDCT_CORE|Fetus OR newborn affected by maternal complication of pregnancy|Fetal or neonatal effect of maternal complication of pregnancy
C0158816|T046|IS|68983007|SNOMEDCT_CORE|Fetus or newborn affected by maternal complication of pregnancy, NOS|Fetal or neonatal effect of maternal complication of pregnancy
C0158816|T046|SY|206035009|SNOMEDCT_CORE|Foetal or neonatal effect of maternal complication of pregnancy|Fetal or neonatal effect of maternal complication of pregnancy
C0158816|T046|OAP|68983007|SNOMEDCT_CORE|Foetal or neonatal effects of maternal complication of pregnancy|Fetal or neonatal effect of maternal complication of pregnancy
C0158816|T046|IS|68983007|SNOMEDCT_CORE|Foetus or newborn affected by maternal complication of pregnancy, NOS|Fetal or neonatal effect of maternal complication of pregnancy
C0158816|T046|IS|68983007|SNOMEDCT_CORE|Maternal complication affecting fetus OR newborn|Fetal or neonatal effect of maternal complication of pregnancy
C0158816|T046|IS|68983007|SNOMEDCT_CORE|Unspecified complication of pregnancy affecting fetus or newborn|Fetal or neonatal effect of maternal complication of pregnancy
C0158819|T046|IS|65599008|SNOMEDCT_CORE|Fetus or newborn affected by oligohydramnios|Fetus or newborn affected by oligohydramnios
C0158819|T046|OP|65599008|SNOMEDCT_CORE|Fetus OR newborn affected by oligohydramnios|Fetus OR newborn affected by oligohydramnios
C0158819|T046|OF|65599008|SNOMEDCT_CORE|Fetus OR newborn affected by oligohydramnios|Fetus OR newborn affected by oligohydramnios
C0158820|T046|OAS|66215008|SNOMEDCT_CORE|Fetal or neonatal effect of hydramnios|Fetal or neonatal effect of polyhydramnios
C0158820|T046|OAP|66215008|SNOMEDCT_CORE|Fetal or neonatal effect of polyhydramnios|Fetal or neonatal effect of polyhydramnios
C0158820|T046|OAF|66215008|SNOMEDCT_CORE|Fetal or neonatal effect of polyhydramnios|Fetal or neonatal effect of polyhydramnios
C0158820|T046|IS|66215008|SNOMEDCT_CORE|Fetus or newborn affected by hydramnios|Fetal or neonatal effect of polyhydramnios
C0158820|T046|IS|66215008|SNOMEDCT_CORE|Fetus or newborn affected by polyhydramnios|Fetal or neonatal effect of polyhydramnios
C0158820|T046|OP|66215008|SNOMEDCT_CORE|Fetus OR newborn affected by polyhydramnios|Fetal or neonatal effect of polyhydramnios
C0158820|T046|OF|66215008|SNOMEDCT_CORE|Fetus OR newborn affected by polyhydramnios|Fetal or neonatal effect of polyhydramnios
C0158832|T046|PT|206087008|SNOMEDCT_CORE|Fetal or neonatal effect of prolapsed cord|Fetal or neonatal effect of prolapsed cord
C0158832|T046|FN|206087008|SNOMEDCT_CORE|Fetal or neonatal effect of prolapsed cord|Fetal or neonatal effect of prolapsed cord
C0158832|T046|OP|206087008|SNOMEDCT_CORE|Fetus or neonate affected by prolapsed cord|Fetal or neonatal effect of prolapsed cord
C0158832|T046|OF|206087008|SNOMEDCT_CORE|Fetus or neonate affected by prolapsed cord|Fetal or neonatal effect of prolapsed cord
C0158832|T046|IS|206087008|SNOMEDCT_CORE|Fetus OR newborn affected by prolapsed cord|Fetal or neonatal effect of prolapsed cord
C0158832|T046|SY|206087008|SNOMEDCT_CORE|Foetal or neonatal effect of prolapsed cord|Fetal or neonatal effect of prolapsed cord
C0158839|T047|IS|268808004|SNOMEDCT_CORE|Fetus affected by breech delivery|Fetus or neonate affected by breech delivery and extraction
C0158839|T047|OP|268808004|SNOMEDCT_CORE|Fetus or neonate affected by breech delivery and extraction|Fetus or neonate affected by breech delivery and extraction
C0158839|T047|OF|268808004|SNOMEDCT_CORE|Fetus or neonate affected by breech delivery and extraction|Fetus or neonate affected by breech delivery and extraction
C0158839|T047|IS|268808004|SNOMEDCT_CORE|Fetus or newborn affected by breech delivery|Fetus or neonate affected by breech delivery and extraction
C0158839|T047|IS|4787007|SNOMEDCT_CORE|Fetus or newborn affected by breech delivery and extraction|Fetus or neonate affected by breech delivery and extraction
C0158839|T047|OP|4787007|SNOMEDCT_CORE|Fetus OR newborn affected by breech delivery AND extraction|Fetus or neonate affected by breech delivery and extraction
C0158839|T047|OF|4787007|SNOMEDCT_CORE|Fetus OR newborn affected by breech delivery AND extraction|Fetus or neonate affected by breech delivery and extraction
C0158842|T033|OP|206122002|SNOMEDCT_CORE|Fetus or neonate affected by vacuum extraction delivery|Fetus or neonate affected by vacuum extraction delivery
C0158842|T033|OF|206122002|SNOMEDCT_CORE|Fetus or neonate affected by vacuum extraction delivery|Fetus or neonate affected by vacuum extraction delivery
C0158842|T033|IS|73890002|SNOMEDCT_CORE|Fetus or newborn affected by delivery by vacuum extractor|Fetus or neonate affected by vacuum extraction delivery
C0158842|T033|OP|73890002|SNOMEDCT_CORE|Fetus OR newborn affected by delivery by vacuum extractor|Fetus or neonate affected by vacuum extraction delivery
C0158842|T033|OF|73890002|SNOMEDCT_CORE|Fetus OR newborn affected by delivery by vacuum extractor|Fetus or neonate affected by vacuum extraction delivery
C0158935|T047|PT|78895009|SNOMEDCT_CORE|Congenital pneumonia|Congenital pneumonia
C0158935|T047|FN|78895009|SNOMEDCT_CORE|Congenital pneumonia|Congenital pneumonia
C0158935|T047|IS|78895009|SNOMEDCT_CORE|Congenital pneumonia, NOS|Congenital pneumonia
C0158940|T047|SY|7550008|SNOMEDCT_CORE|Idiopathic tachypnea of newborn|Transitory tachypnea of newborn
C0158940|T047|SYGB|7550008|SNOMEDCT_CORE|Idiopathic tachypnoea of newborn|Transitory tachypnea of newborn
C0158940|T047|SY|7550008|SNOMEDCT_CORE|Newborn transitory tachypnea|Transitory tachypnea of newborn
C0158940|T047|SYGB|7550008|SNOMEDCT_CORE|Newborn transitory tachypnoea|Transitory tachypnea of newborn
C0158940|T047|SY|7550008|SNOMEDCT_CORE|Tachypnea resolving about 6 hours postnatally|Transitory tachypnea of newborn
C0158940|T047|SYGB|7550008|SNOMEDCT_CORE|Tachypnoea resolving about 6 hours postnatally|Transitory tachypnea of newborn
C0158940|T047|SY|7550008|SNOMEDCT_CORE|Transient tachypnea of newborn|Transitory tachypnea of newborn
C0158940|T047|SYGB|7550008|SNOMEDCT_CORE|Transient tachypnoea of newborn|Transitory tachypnea of newborn
C0158940|T047|PT|7550008|SNOMEDCT_CORE|Transitory tachypnea of newborn|Transitory tachypnea of newborn
C0158940|T047|FN|7550008|SNOMEDCT_CORE|Transitory tachypnea of newborn|Transitory tachypnea of newborn
C0158940|T047|PTGB|7550008|SNOMEDCT_CORE|Transitory tachypnoea of newborn|Transitory tachypnea of newborn
C0158940|T047|SY|7550008|SNOMEDCT_CORE|TTN - Transient tachypnea of newborn|Transitory tachypnea of newborn
C0158940|T047|SYGB|7550008|SNOMEDCT_CORE|TTN - Transient tachypnoea of newborn|Transitory tachypnea of newborn
C0158940|T047|SY|7550008|SNOMEDCT_CORE|Wet lung syndrome in newborn|Transitory tachypnea of newborn
C0158944|T047|PT|206331005|SNOMEDCT_CORE|Infections specific to perinatal period|Infections specific to perinatal period
C0158944|T047|FN|206331005|SNOMEDCT_CORE|Infections specific to perinatal period|Infections specific to perinatal period
C0158969|T047|PTGB|56921004|SNOMEDCT_CORE|Perinatal jaundice due to hereditary haemolytic anaemia|Perinatal jaundice due to hereditary hemolytic anemia
C0158969|T047|PT|56921004|SNOMEDCT_CORE|Perinatal jaundice due to hereditary hemolytic anemia|Perinatal jaundice due to hereditary hemolytic anemia
C0158969|T047|FN|56921004|SNOMEDCT_CORE|Perinatal jaundice due to hereditary hemolytic anemia|Perinatal jaundice due to hereditary hemolytic anemia
C0158969|T047|OP|56921004|SNOMEDCT_CORE|Perinatal jaundice from hereditary haemolytic anaemia|Perinatal jaundice due to hereditary hemolytic anemia
C0158969|T047|IS|56921004|SNOMEDCT_CORE|Perinatal jaundice from hereditary haemolytic anaemias|Perinatal jaundice due to hereditary hemolytic anemia
C0158969|T047|OP|56921004|SNOMEDCT_CORE|Perinatal jaundice from hereditary hemolytic anemia|Perinatal jaundice due to hereditary hemolytic anemia
C0158969|T047|OF|56921004|SNOMEDCT_CORE|Perinatal jaundice from hereditary hemolytic anemia|Perinatal jaundice due to hereditary hemolytic anemia
C0158969|T047|IS|56921004|SNOMEDCT_CORE|Perinatal jaundice from hereditary hemolytic anemias|Perinatal jaundice due to hereditary hemolytic anemia
C0158971|T046|SYGB|73749009|SNOMEDCT_CORE|Hyperbilirubinaemia of prematurity|Neonatal jaundice associated with preterm delivery
C0158971|T046|SY|73749009|SNOMEDCT_CORE|Hyperbilirubinemia of prematurity|Neonatal jaundice associated with preterm delivery
C0158971|T046|SY|73749009|SNOMEDCT_CORE|Jaundice due to delayed conjugation associated with preterm delivery|Neonatal jaundice associated with preterm delivery
C0158971|T046|SY|73749009|SNOMEDCT_CORE|Neonatal jaundice after preterm delivery|Neonatal jaundice associated with preterm delivery
C0158971|T046|PT|73749009|SNOMEDCT_CORE|Neonatal jaundice associated with preterm delivery|Neonatal jaundice associated with preterm delivery
C0158971|T046|FN|73749009|SNOMEDCT_CORE|Neonatal jaundice associated with preterm delivery|Neonatal jaundice associated with preterm delivery
C0158971|T046|SY|73749009|SNOMEDCT_CORE|Preterm delivery-associated jaundice|Neonatal jaundice associated with preterm delivery
C0158986|T047|PTGB|52767006|SNOMEDCT_CORE|Neonatal hypoglycaemia|Neonatal hypoglycemia
C0158986|T047|PT|52767006|SNOMEDCT_CORE|Neonatal hypoglycemia|Neonatal hypoglycemia
C0158986|T047|FN|52767006|SNOMEDCT_CORE|Neonatal hypoglycemia|Neonatal hypoglycemia
C0158996|T047|PTGB|47100003|SNOMEDCT_CORE|Anaemia of prematurity|Anemia of prematurity
C0158996|T047|PT|47100003|SNOMEDCT_CORE|Anemia of prematurity|Anemia of prematurity
C0158996|T047|FN|47100003|SNOMEDCT_CORE|Anemia of prematurity|Anemia of prematurity
C0159015|T019|PT|82062003|SNOMEDCT_CORE|Congenital hydrocele|Congenital hydrocele
C0159015|T019|FN|82062003|SNOMEDCT_CORE|Congenital hydrocele|Congenital hydrocele
C0159015|T019|SY|82062003|SNOMEDCT_CORE|Congenital hydrocele of tunica vaginalis|Congenital hydrocele
C0159015|T019|IS|82062003|SNOMEDCT_CORE|Congenital hydrocele, NOS|Congenital hydrocele
C0159015|T019|PTGB|82062003|SNOMEDCT_CORE|Congenital hydrocoele|Congenital hydrocele
C0159015|T019|SYGB|82062003|SNOMEDCT_CORE|Congenital hydrocoele of tunica vaginalis|Congenital hydrocele
C0159020|T047|PT|87476004|SNOMEDCT_CORE|Convulsions in the newborn|Convulsions in the newborn
C0159020|T047|FN|87476004|SNOMEDCT_CORE|Convulsions in the newborn|Convulsions in the newborn
C0159020|T047|SY|87476004|SNOMEDCT_CORE|Fits in newborn|Convulsions in the newborn
C0159020|T047|SY|87476004|SNOMEDCT_CORE|Fits in the newborn|Convulsions in the newborn
C0159020|T047|SY|87476004|SNOMEDCT_CORE|Neonatal convulsions|Convulsions in the newborn
C0159020|T047|SY|87476004|SNOMEDCT_CORE|Neonatal seizures|Convulsions in the newborn
C0159020|T047|SY|87476004|SNOMEDCT_CORE|Seizures in newborn|Convulsions in the newborn
C0159020|T047|SY|87476004|SNOMEDCT_CORE|Seizures in the newborn|Convulsions in the newborn
C0159023|T033|SY|72552008|SNOMEDCT_CORE|Feeding difficulties in newborn|Feeding problems in newborn
C0159023|T033|IS|72552008|SNOMEDCT_CORE|Feeding problem in newborn|Feeding problems in newborn
C0159023|T033|IS|72552008|SNOMEDCT_CORE|Feeding problem in newborn, NOS|Feeding problems in newborn
C0159023|T033|PT|72552008|SNOMEDCT_CORE|Feeding problems in newborn|Feeding problems in newborn
C0159023|T033|FN|72552008|SNOMEDCT_CORE|Feeding problems in newborn|Feeding problems in newborn
C0159028|T184|PT|267022002|SNOMEDCT_CORE|General symptom|General symptom
C0159028|T184|FN|267022002|SNOMEDCT_CORE|General symptom|General symptom
C0159028|T184|IS|267022002|SNOMEDCT_CORE|General symptoms|General symptom
C0159028|T184|OF|267022002|SNOMEDCT_CORE|General symptoms|General symptom
C0159030|T184|PT|41975002|SNOMEDCT_CORE|Insomnia with sleep apnea|Insomnia with sleep apnea
C0159030|T184|FN|41975002|SNOMEDCT_CORE|Insomnia with sleep apnea|Insomnia with sleep apnea
C0159030|T184|PTGB|41975002|SNOMEDCT_CORE|Insomnia with sleep apnoea|Insomnia with sleep apnea
C0159047|T048|PT|271721006|SNOMEDCT_CORE|Symbolic dysfunction|Symbolic dysfunction
C0159047|T048|FN|271721006|SNOMEDCT_CORE|Symbolic dysfunction|Symbolic dysfunction
C0159054|T033|PT|274708000|SNOMEDCT_CORE|Abnormal sputum|Abnormal sputum
C0159054|T033|FN|274708000|SNOMEDCT_CORE|Abnormal sputum|Abnormal sputum
C0159127|T033|PT|441846005|SNOMEDCT_CORE|Nonspecific tuberculin test reaction|Nonspecific tuberculin test reaction
C0159127|T033|FN|441846005|SNOMEDCT_CORE|Nonspecific tuberculin test reaction|Nonspecific tuberculin test reaction
C0159158|T037|IS|57998008|SNOMEDCT_CORE|Closed fracture of vault of skull with subarachnoid, subdural and extradural hemorrhage|Closed fracture of vault of skull with subarachnoid, subdural and extradural hemorrhage
C0159158|T037|OAP|57998008|SNOMEDCT_CORE|Closed fracture of vault of skull with subarachnoid, subdural AND/OR extradural haemorrhage|Closed fracture of vault of skull with subarachnoid, subdural AND/OR extradural haemorrhage
C0159158|T037|OAP|57998008|SNOMEDCT_CORE|Closed fracture of vault of skull with subarachnoid, subdural AND/OR extradural hemorrhage|Closed fracture of vault of skull with subarachnoid, subdural AND/OR extradural hemorrhage
C0159158|T037|OAF|57998008|SNOMEDCT_CORE|Closed fracture of vault of skull with subarachnoid, subdural AND/OR extradural hemorrhage|Closed fracture of vault of skull with subarachnoid, subdural AND/OR extradural hemorrhage
C0159321|T037|PT|27477003|SNOMEDCT_CORE|Fracture of face bones|Fracture of face bones
C0159321|T037|FN|27477003|SNOMEDCT_CORE|Fracture of face bones|Fracture of face bones
C0159321|T037|IS|27477003|SNOMEDCT_CORE|Fracture of face bones, NOS|Fracture of face bones
C0159321|T037|SY|27477003|SNOMEDCT_CORE|Fracture of facial bone|Fracture of face bones
C0159321|T037|SY|27477003|SNOMEDCT_CORE|Fracture of facial bones|Fracture of face bones
C0159321|T037|IS|27477003|SNOMEDCT_CORE|Fracture of facial bones, NOS|Fracture of face bones
C0159322|T037|SY|81639003|SNOMEDCT_CORE|Closed fracture nasal bone|Closed fracture of nasal bones
C0159322|T037|SY|81639003|SNOMEDCT_CORE|Closed fracture nose|Closed fracture of nasal bones
C0159322|T037|PT|81639003|SNOMEDCT_CORE|Closed fracture of nasal bones|Closed fracture of nasal bones
C0159322|T037|FN|81639003|SNOMEDCT_CORE|Closed fracture of nasal bones|Closed fracture of nasal bones
C0159324|T037|SY|207753003|SNOMEDCT_CORE|Closed fracture of inferior maxilla|Fracture of mandible, closed
C0159324|T037|SY|207753003|SNOMEDCT_CORE|Closed fracture of lower jaw bone|Fracture of mandible, closed
C0159324|T037|SY|207753003|SNOMEDCT_CORE|Closed fracture of mandible|Fracture of mandible, closed
C0159324|T037|SY|207753003|SNOMEDCT_CORE|Fracture of lower jaw, closed|Fracture of mandible, closed
C0159324|T037|PT|207753003|SNOMEDCT_CORE|Fracture of mandible, closed|Fracture of mandible, closed
C0159324|T037|FN|207753003|SNOMEDCT_CORE|Fracture of mandible, closed|Fracture of mandible, closed
C0159553|T037|PT|207957008|SNOMEDCT_CORE|Closed fracture lumbar vertebra|Closed fracture lumbar vertebra
C0159553|T037|FN|207957008|SNOMEDCT_CORE|Closed fracture lumbar vertebra|Closed fracture lumbar vertebra
C0159618|T037|PT|45356009|SNOMEDCT_CORE|Closed fracture of one rib|Closed fracture of one rib
C0159618|T037|FN|45356009|SNOMEDCT_CORE|Closed fracture of one rib|Closed fracture of one rib
C0159619|T037|PT|3291007|SNOMEDCT_CORE|Closed fracture of two ribs|Closed fracture of two ribs
C0159619|T037|FN|3291007|SNOMEDCT_CORE|Closed fracture of two ribs|Closed fracture of two ribs
C0159620|T037|PT|79546008|SNOMEDCT_CORE|Closed fracture of three ribs|Closed fracture of three ribs
C0159620|T037|FN|79546008|SNOMEDCT_CORE|Closed fracture of three ribs|Closed fracture of three ribs
C0159621|T037|PT|39335003|SNOMEDCT_CORE|Closed fracture of four ribs|Closed fracture of four ribs
C0159621|T037|FN|39335003|SNOMEDCT_CORE|Closed fracture of four ribs|Closed fracture of four ribs
C0159626|T037|SY|12204004|SNOMEDCT_CORE|Closed fracture multiple ribs|Closed fracture of multiple ribs
C0159626|T037|PT|12204004|SNOMEDCT_CORE|Closed fracture of multiple ribs|Closed fracture of multiple ribs
C0159626|T037|FN|12204004|SNOMEDCT_CORE|Closed fracture of multiple ribs|Closed fracture of multiple ribs
C0159626|T037|IS|12204004|SNOMEDCT_CORE|Closed fracture of multiple ribs, NOS|Closed fracture of multiple ribs
C0159637|T037|PT|66112004|SNOMEDCT_CORE|Closed fracture of sternum|Closed fracture of sternum
C0159637|T037|FN|66112004|SNOMEDCT_CORE|Closed fracture of sternum|Closed fracture of sternum
C0159637|T037|SY|66112004|SNOMEDCT_CORE|Closed fracture sternum|Closed fracture of sternum
C0159641|T037|SY|33118001|SNOMEDCT_CORE|Closed fracture acetabulum|Closed fracture of acetabulum
C0159641|T037|PT|33118001|SNOMEDCT_CORE|Closed fracture of acetabulum|Closed fracture of acetabulum
C0159641|T037|FN|33118001|SNOMEDCT_CORE|Closed fracture of acetabulum|Closed fracture of acetabulum
C0159643|T037|SY|208164008|SNOMEDCT_CORE|Closed fracture of pubis|Closed fracture pubis
C0159643|T037|PT|208164008|SNOMEDCT_CORE|Closed fracture pubis|Closed fracture pubis
C0159643|T037|FN|208164008|SNOMEDCT_CORE|Closed fracture pubis|Closed fracture pubis
C0159658|T037|SY|58150001|SNOMEDCT_CORE|Collar bone fracture|Fracture of clavicle
C0159658|T037|PT|58150001|SNOMEDCT_CORE|Fracture of clavicle|Fracture of clavicle
C0159658|T037|FN|58150001|SNOMEDCT_CORE|Fracture of clavicle|Fracture of clavicle
C0159658|T037|IS|58150001|SNOMEDCT_CORE|Fracture of clavicle, NOS|Fracture of clavicle
C0159658|T037|SY|58150001|SNOMEDCT_CORE|Fracture of collar bone|Fracture of clavicle
C0159659|T037|PT|33173003|SNOMEDCT_CORE|Closed fracture of clavicle|Closed fracture of clavicle
C0159659|T037|FN|33173003|SNOMEDCT_CORE|Closed fracture of clavicle|Closed fracture of clavicle
C0159659|T037|IS|33173003|SNOMEDCT_CORE|Closed fracture of clavicle, NOS|Closed fracture of clavicle
C0159667|T037|PT|9682006|SNOMEDCT_CORE|Fracture of scapula|Fracture of scapula
C0159667|T037|FN|9682006|SNOMEDCT_CORE|Fracture of scapula|Fracture of scapula
C0159667|T037|IS|9682006|SNOMEDCT_CORE|Fracture of scapula, NOS|Fracture of scapula
C0159667|T037|SY|9682006|SNOMEDCT_CORE|Fracture of shoulder blade|Fracture of scapula
C0159667|T037|IS|9682006|SNOMEDCT_CORE|Fracture of shoulder blade, NOS|Fracture of scapula
C0159668|T037|PT|29749002|SNOMEDCT_CORE|Closed fracture of scapula|Closed fracture of scapula
C0159668|T037|FN|29749002|SNOMEDCT_CORE|Closed fracture of scapula|Closed fracture of scapula
C0159668|T037|IS|29749002|SNOMEDCT_CORE|Closed fracture of scapula, NOS|Closed fracture of scapula
C0159668|T037|SY|29749002|SNOMEDCT_CORE|Closed fracture of shoulder blade|Closed fracture of scapula
C0159668|T037|IS|29749002|SNOMEDCT_CORE|Closed fracture of shoulder blade, NOS|Closed fracture of scapula
C0159678|T037|SY|42636007|SNOMEDCT_CORE|Closed fracture of proximal end of humerus|Closed fracture of upper end of humerus
C0159678|T037|SY|42636007|SNOMEDCT_CORE|Closed fracture of the proximal humerus|Closed fracture of upper end of humerus
C0159678|T037|PT|42636007|SNOMEDCT_CORE|Closed fracture of upper end of humerus|Closed fracture of upper end of humerus
C0159678|T037|FN|42636007|SNOMEDCT_CORE|Closed fracture of upper end of humerus|Closed fracture of upper end of humerus
C0159678|T037|IS|42636007|SNOMEDCT_CORE|Closed fracture of upper end of humerus, NOS|Closed fracture of upper end of humerus
C0159680|T037|SY|73244003|SNOMEDCT_CORE|Closed fracture of neck of humerus|Closed fracture of surgical neck of humerus
C0159680|T037|IS|73244003|SNOMEDCT_CORE|Closed fracture of neck of humerus, NOS|Closed fracture of surgical neck of humerus
C0159680|T037|PT|73244003|SNOMEDCT_CORE|Closed fracture of surgical neck of humerus|Closed fracture of surgical neck of humerus
C0159680|T037|FN|73244003|SNOMEDCT_CORE|Closed fracture of surgical neck of humerus|Closed fracture of surgical neck of humerus
C0159692|T037|SY|90235006|SNOMEDCT_CORE|Closed fracture of humerus, shaft|Closed fracture of shaft of humerus
C0159692|T037|PT|90235006|SNOMEDCT_CORE|Closed fracture of shaft of humerus|Closed fracture of shaft of humerus
C0159692|T037|FN|90235006|SNOMEDCT_CORE|Closed fracture of shaft of humerus|Closed fracture of shaft of humerus
C0159710|T037|PT|75857000|SNOMEDCT_CORE|Fracture of radius AND ulna|Fracture of radius AND ulna
C0159710|T037|FN|75857000|SNOMEDCT_CORE|Fracture of radius AND ulna|Fracture of radius AND ulna
C0159710|T037|IS|75857000|SNOMEDCT_CORE|Fracture of radius and ulna, NOS|Fracture of radius AND ulna
C0159713|T037|PT|64902007|SNOMEDCT_CORE|Closed fracture of olecranon process of ulna|Closed fracture of olecranon process of ulna
C0159713|T037|FN|64902007|SNOMEDCT_CORE|Closed fracture of olecranon process of ulna|Closed fracture of olecranon process of ulna
C0159716|T037|PT|68854005|SNOMEDCT_CORE|Closed fracture of head of radius|Closed fracture of head of radius
C0159716|T037|FN|68854005|SNOMEDCT_CORE|Closed fracture of head of radius|Closed fracture of head of radius
C0159716|T037|SY|68854005|SNOMEDCT_CORE|Closed fracture radius, head|Closed fracture of head of radius
C0159730|T037|IS|28078000|SNOMEDCT_CORE|Closed fracture of radius and ulna, shaft|Closed fracture of radius and ulna, shaft
C0159730|T037|IS|28078000|SNOMEDCT_CORE|Closed fracture of shaft of radius AND ulna|Closed fracture of shaft of radius AND ulna
C0159738|T037|PT|33192001|SNOMEDCT_CORE|Closed fracture of lower end of radius AND ulna|Closed fracture of lower end of radius AND ulna
C0159738|T037|IS|33192001|SNOMEDCT_CORE|Closed fracture of lower end of radius and ulna|Closed fracture of lower end of radius AND ulna
C0159738|T037|FN|33192001|SNOMEDCT_CORE|Closed fracture of lower end of radius AND ulna|Closed fracture of lower end of radius AND ulna
C0159738|T037|SY|33192001|SNOMEDCT_CORE|Closed fracture of radius and ulna, lower end|Closed fracture of lower end of radius AND ulna
C0159738|T037|SY|33192001|SNOMEDCT_CORE|Closed fracture radius and ulna, distal|Closed fracture of lower end of radius AND ulna
C0159776|T037|OAP|91588005|SNOMEDCT_CORE|Closed fracture of metacarpal bone|Closed fracture of metacarpal bone
C0159776|T037|PT|208394006|SNOMEDCT_CORE|Closed fracture of metacarpal bone|Closed fracture of metacarpal bone
C0159776|T037|IS|208394006|SNOMEDCT_CORE|Closed fracture of metacarpal bone|Closed fracture of metacarpal bone
C0159776|T037|OAF|91588005|SNOMEDCT_CORE|Closed fracture of metacarpal bone|Closed fracture of metacarpal bone
C0159776|T037|FN|208394006|SNOMEDCT_CORE|Closed fracture of metacarpal bone|Closed fracture of metacarpal bone
C0159776|T037|OF|208394006|SNOMEDCT_CORE|Closed fracture of metacarpal bone|Closed fracture of metacarpal bone
C0159776|T037|IS|91588005|SNOMEDCT_CORE|Closed fracture of metacarpal bone, NOS|Closed fracture of metacarpal bone
C0159791|T037|PT|208430000|SNOMEDCT_CORE|Closed fracture of one or more phalanges of hand|Closed fracture of one or more phalanges of hand
C0159791|T037|FN|208430000|SNOMEDCT_CORE|Closed fracture of one or more phalanges of hand|Closed fracture of one or more phalanges of hand
C0159796|T037|PT|208463007|SNOMEDCT_CORE|Open fracture of one or more phalanges of hand|Open fracture of one or more phalanges of hand
C0159796|T037|FN|208463007|SNOMEDCT_CORE|Open fracture of one or more phalanges of hand|Open fracture of one or more phalanges of hand
C0159814|T037|PT|1705000|SNOMEDCT_CORE|Closed fracture of base of neck of femur|Closed fracture of base of neck of femur
C0159814|T037|FN|1705000|SNOMEDCT_CORE|Closed fracture of base of neck of femur|Closed fracture of base of neck of femur
C0159814|T037|SY|1705000|SNOMEDCT_CORE|Closed fracture of cervicotrochanteric section of femur|Closed fracture of base of neck of femur
C0159833|T037|PT|26442006|SNOMEDCT_CORE|Closed fracture of shaft of femur|Closed fracture of shaft of femur
C0159833|T037|FN|26442006|SNOMEDCT_CORE|Closed fracture of shaft of femur|Closed fracture of shaft of femur
C0159833|T037|SY|26442006|SNOMEDCT_CORE|Closed fracture shaft of femur|Closed fracture of shaft of femur
C0159837|T037|SY|263233008|SNOMEDCT_CORE|Closed fracture of distal end of femur|Closed fracture of femur, distal end
C0159837|T037|PT|263233008|SNOMEDCT_CORE|Closed fracture of femur, distal end|Closed fracture of femur, distal end
C0159837|T037|FN|263233008|SNOMEDCT_CORE|Closed fracture of femur, distal end|Closed fracture of femur, distal end
C0159837|T037|SY|263233008|SNOMEDCT_CORE|Closed fracture of lower end of femur|Closed fracture of femur, distal end
C0159849|T037|SY|51037009|SNOMEDCT_CORE|Fracture of knee-cap|Fracture of patella
C0159849|T037|PT|51037009|SNOMEDCT_CORE|Fracture of patella|Fracture of patella
C0159849|T037|FN|51037009|SNOMEDCT_CORE|Fracture of patella|Fracture of patella
C0159849|T037|IS|51037009|SNOMEDCT_CORE|Fracture of patella, NOS|Fracture of patella
C0159850|T037|PT|80756009|SNOMEDCT_CORE|Closed fracture of patella|Closed fracture of patella
C0159850|T037|FN|80756009|SNOMEDCT_CORE|Closed fracture of patella|Closed fracture of patella
C0159852|T037|PT|414293001|SNOMEDCT_CORE|Fracture of tibia AND fibula|Fracture of tibia AND fibula
C0159852|T037|FN|414293001|SNOMEDCT_CORE|Fracture of tibia AND fibula|Fracture of tibia AND fibula
C0159854|T037|PT|23900009|SNOMEDCT_CORE|Closed fracture of upper end of tibia|Closed fracture of upper end of tibia
C0159854|T037|FN|23900009|SNOMEDCT_CORE|Closed fracture of upper end of tibia|Closed fracture of upper end of tibia
C0159862|T037|PT|28012007|SNOMEDCT_CORE|Closed fracture of shaft of tibia|Closed fracture of shaft of tibia
C0159862|T037|FN|28012007|SNOMEDCT_CORE|Closed fracture of shaft of tibia|Closed fracture of shaft of tibia
C0159864|T037|PT|208629000|SNOMEDCT_CORE|Closed fracture of tibia and fibula, shaft|Closed fracture of tibia and fibula, shaft
C0159864|T037|FN|208629000|SNOMEDCT_CORE|Closed fracture of tibia and fibula, shaft|Closed fracture of tibia and fibula, shaft
C0159877|T037|SY|16114001|SNOMEDCT_CORE|Ankle fracture|Fracture of ankle
C0159877|T037|PT|16114001|SNOMEDCT_CORE|Fracture of ankle|Fracture of ankle
C0159877|T037|FN|16114001|SNOMEDCT_CORE|Fracture of ankle|Fracture of ankle
C0159877|T037|IS|16114001|SNOMEDCT_CORE|Fracture of ankle, NOS|Fracture of ankle
C0159877|T037|SY|16114001|SNOMEDCT_CORE|Fracture of distal end of tibia and fibula|Fracture of ankle
C0159883|T037|SY|6698000|SNOMEDCT_CORE|Closed fracture ankle, trimalleolar|Closed trimalleolar fracture
C0159883|T037|PT|6698000|SNOMEDCT_CORE|Closed trimalleolar fracture|Closed trimalleolar fracture
C0159883|T037|FN|6698000|SNOMEDCT_CORE|Closed trimalleolar fracture|Closed trimalleolar fracture
C0159888|T037|PT|64665009|SNOMEDCT_CORE|Closed fracture of calcaneus|Closed fracture of calcaneus
C0159888|T037|FN|64665009|SNOMEDCT_CORE|Closed fracture of calcaneus|Closed fracture of calcaneus
C0159888|T037|SY|64665009|SNOMEDCT_CORE|Closed fracture of heel bone|Closed fracture of calcaneus
C0159888|T037|SY|64665009|SNOMEDCT_CORE|Closed fracture of os calcis|Closed fracture of calcaneus
C0159917|T037|PT|34565006|SNOMEDCT_CORE|Closed anterior dislocation of humerus|Closed anterior dislocation of humerus
C0159917|T037|FN|34565006|SNOMEDCT_CORE|Closed anterior dislocation of humerus|Closed anterior dislocation of humerus
C0159920|T037|IS|208759001|SNOMEDCT_CORE|Closed dislocation of acromioclavicular joint|Closed traumatic dislocation acromioclavicular joint
C0159920|T037|PT|208759001|SNOMEDCT_CORE|Closed traumatic dislocation acromioclavicular joint|Closed traumatic dislocation acromioclavicular joint
C0159920|T037|FN|208759001|SNOMEDCT_CORE|Closed traumatic dislocation acromioclavicular joint|Closed traumatic dislocation acromioclavicular joint
C0159931|T037|PT|4273008|SNOMEDCT_CORE|Closed posterior dislocation of elbow|Closed posterior dislocation of elbow
C0159931|T037|FN|4273008|SNOMEDCT_CORE|Closed posterior dislocation of elbow|Closed posterior dislocation of elbow
C0159956|T037|OP|125619004|SNOMEDCT_CORE|Dislocation of finger|Traumatic dislocation of joint of finger
C0159956|T037|PT|125619004|SNOMEDCT_CORE|Traumatic dislocation of joint of finger|Traumatic dislocation of joint of finger
C0159956|T037|FN|125619004|SNOMEDCT_CORE|Traumatic dislocation of joint of finger|Traumatic dislocation of joint of finger
C0159957|T037|OP|75137002|SNOMEDCT_CORE|Closed dislocation of finger|Closed traumatic dislocation of joint of finger
C0159957|T037|IS|75137002|SNOMEDCT_CORE|Closed dislocation of finger, NOS|Closed traumatic dislocation of joint of finger
C0159957|T037|IS|75137002|SNOMEDCT_CORE|Closed dislocation of phalanx of hand|Closed traumatic dislocation of joint of finger
C0159957|T037|IS|75137002|SNOMEDCT_CORE|Closed dislocation of phalanx of hand, NOS|Closed traumatic dislocation of joint of finger
C0159957|T037|PT|75137002|SNOMEDCT_CORE|Closed traumatic dislocation of joint of finger|Closed traumatic dislocation of joint of finger
C0159957|T037|FN|75137002|SNOMEDCT_CORE|Closed traumatic dislocation of joint of finger|Closed traumatic dislocation of joint of finger
C0159970|T037|IS|58320001|SNOMEDCT_CORE|Dislocated knee|Traumatic dislocation of knee joint
C0159970|T037|OP|58320001|SNOMEDCT_CORE|Dislocation of knee|Traumatic dislocation of knee joint
C0159970|T037|IS|58320001|SNOMEDCT_CORE|Dislocation of knee, NOS|Traumatic dislocation of knee joint
C0159970|T037|IS|58320001|SNOMEDCT_CORE|Dislocation of tibiofemoral joint|Traumatic dislocation of knee joint
C0159970|T037|FN|58320001|SNOMEDCT_CORE|Traumatic dislocation of knee joint|Traumatic dislocation of knee joint
C0159970|T037|PT|58320001|SNOMEDCT_CORE|Traumatic dislocation of knee joint|Traumatic dislocation of knee joint
C0159971|T037|PT|302932006|SNOMEDCT_CORE|Tear of medial meniscus of knee|Tear of medial meniscus of knee
C0159971|T037|FN|302932006|SNOMEDCT_CORE|Tear of medial meniscus of knee|Tear of medial meniscus of knee
C0159971|T037|SY|302932006|SNOMEDCT_CORE|Tear of medial meniscus of knee joint|Tear of medial meniscus of knee
C0159971|T037|SY|302932006|SNOMEDCT_CORE|Torn medial meniscus|Tear of medial meniscus of knee
C0160063|T037|PT|70704007|SNOMEDCT_CORE|Sprain of wrist|Sprain of wrist
C0160063|T037|FN|70704007|SNOMEDCT_CORE|Sprain of wrist|Sprain of wrist
C0160063|T037|SY|70704007|SNOMEDCT_CORE|Sprain of wrist joint|Sprain of wrist
C0160063|T037|IS|70704007|SNOMEDCT_CORE|Sprain of wrist, NOS|Sprain of wrist
C0160063|T037|SY|70704007|SNOMEDCT_CORE|Wrist sprain|Sprain of wrist
C0160068|T037|SY|87778004|SNOMEDCT_CORE|Hand sprain|Sprain of hand
C0160068|T037|PT|87778004|SNOMEDCT_CORE|Sprain of hand|Sprain of hand
C0160068|T037|FN|87778004|SNOMEDCT_CORE|Sprain of hand|Sprain of hand
C0160068|T037|SY|87778004|SNOMEDCT_CORE|Sprain of hand joint|Sprain of hand
C0160068|T037|IS|87778004|SNOMEDCT_CORE|Sprain of hand, NOS|Sprain of hand
C0160068|T037|SY|87778004|SNOMEDCT_CORE|Sprain of joint of hand|Sprain of hand
C0160068|T037|SY|87778004|SNOMEDCT_CORE|Sprain of ligament of hand|Sprain of hand
C0160081|T037|PT|81902001|SNOMEDCT_CORE|Sprain of medial collateral ligament of knee|Sprain of medial collateral ligament of knee
C0160081|T037|FN|81902001|SNOMEDCT_CORE|Sprain of medial collateral ligament of knee|Sprain of medial collateral ligament of knee
C0160087|T037|SY|44465007|SNOMEDCT_CORE|Ankle sprain|Sprain of ankle
C0160087|T037|PT|44465007|SNOMEDCT_CORE|Sprain of ankle|Sprain of ankle
C0160087|T037|FN|44465007|SNOMEDCT_CORE|Sprain of ankle|Sprain of ankle
C0160087|T037|SY|44465007|SNOMEDCT_CORE|Sprain of ankle joint|Sprain of ankle
C0160087|T037|IS|44465007|SNOMEDCT_CORE|Sprain of ankle, NOS|Sprain of ankle
C0160087|T037|SY|44465007|SNOMEDCT_CORE|Sprain of ligament of ankle joint|Sprain of ankle
C0160093|T037|SY|49388007|SNOMEDCT_CORE|Foot sprain|Sprain of foot
C0160093|T037|SY|49388007|SNOMEDCT_CORE|FSPR - Foot sprain|Sprain of foot
C0160093|T037|PT|49388007|SNOMEDCT_CORE|Sprain of foot|Sprain of foot
C0160093|T037|FN|49388007|SNOMEDCT_CORE|Sprain of foot|Sprain of foot
C0160093|T037|IS|49388007|SNOMEDCT_CORE|Sprain of foot, NOS|Sprain of foot
C0160107|T037|PT|274162005|SNOMEDCT_CORE|Thoracic back sprain|Thoracic back sprain
C0160107|T037|FN|274162005|SNOMEDCT_CORE|Thoracic back sprain|Thoracic back sprain
C0160108|T037|SY|209565008|SNOMEDCT_CORE|Lumbar back sprain|Lumbar sprain
C0160108|T037|PT|209565008|SNOMEDCT_CORE|Lumbar sprain|Lumbar sprain
C0160108|T037|FN|209565008|SNOMEDCT_CORE|Lumbar sprain|Lumbar sprain
C0160111|T037|SY|281598004|SNOMEDCT_CORE|Back sprain|Back sprain
C0160121|T037|PT|62106007|SNOMEDCT_CORE|Concussion with no loss of consciousness|Concussion with no loss of consciousness
C0160121|T037|FN|62106007|SNOMEDCT_CORE|Concussion with no loss of consciousness|Concussion with no loss of consciousness
C0160122|T037|PT|209827006|SNOMEDCT_CORE|Concussion with less than 1 hour loss of consciousness|Concussion with less than 1 hour loss of consciousness
C0160122|T037|FN|209827006|SNOMEDCT_CORE|Concussion with less than 1 hour loss of consciousness|Concussion with less than 1 hour loss of consciousness
C0160126|T037|PT|62564004|SNOMEDCT_CORE|Concussion with loss of consciousness|Concussion with loss of consciousness
C0160126|T037|FN|62564004|SNOMEDCT_CORE|Concussion with loss of consciousness|Concussion with loss of consciousness
C0160126|T037|IS|62564004|SNOMEDCT_CORE|Concussion with loss of consciousness of unspecified duration|Concussion with loss of consciousness
C0160469|T037|PT|23293006|SNOMEDCT_CORE|Rupture of eye with partial loss of intraocular tissue|Rupture of eye with partial loss of intraocular tissue
C0160469|T037|FN|23293006|SNOMEDCT_CORE|Rupture of eye with partial loss of intraocular tissue|Rupture of eye with partial loss of intraocular tissue
C0160604|T037|PT|125649002|SNOMEDCT_CORE|Open wound of forearm|Open wound of forearm
C0160604|T037|FN|125649002|SNOMEDCT_CORE|Open wound of forearm|Open wound of forearm
C0160612|T037|PT|6154004|SNOMEDCT_CORE|Open wound of forearm with tendon involvement|Open wound of forearm with tendon involvement
C0160612|T037|FN|6154004|SNOMEDCT_CORE|Open wound of forearm with tendon involvement|Open wound of forearm with tendon involvement
C0160614|T037|PT|15550007|SNOMEDCT_CORE|Open wound of wrist with tendon involvement|Open wound of wrist with tendon involvement
C0160614|T037|FN|15550007|SNOMEDCT_CORE|Open wound of wrist with tendon involvement|Open wound of wrist with tendon involvement
C0160621|T037|PT|32348000|SNOMEDCT_CORE|Open wound of finger with complication|Open wound of finger with complication
C0160621|T037|FN|32348000|SNOMEDCT_CORE|Open wound of finger with complication|Open wound of finger with complication
C0160622|T037|PT|23777003|SNOMEDCT_CORE|Open wound of finger with tendon involvement|Open wound of finger with tendon involvement
C0160622|T037|FN|23777003|SNOMEDCT_CORE|Open wound of finger with tendon involvement|Open wound of finger with tendon involvement
C0160643|T037|SY|210661006|SNOMEDCT_CORE|Open wound of hip and thigh|Open wound of hip and/or thigh
C0160643|T037|OF|210661006|SNOMEDCT_CORE|Open wound of hip and thigh|Open wound of hip and/or thigh
C0160643|T037|PT|210661006|SNOMEDCT_CORE|Open wound of hip and/or thigh|Open wound of hip and/or thigh
C0160643|T037|FN|210661006|SNOMEDCT_CORE|Open wound of hip and/or thigh|Open wound of hip and/or thigh
C0160778|T046|PT|36758002|SNOMEDCT_CORE|Late effect of fracture of lower extremities|Late effect of fracture of lower extremities
C0160778|T046|FN|36758002|SNOMEDCT_CORE|Late effect of fracture of lower extremities|Late effect of fracture of lower extremities
C0160797|T046|PT|81642009|SNOMEDCT_CORE|Late effect of spinal cord injury|Late effect of spinal cord injury
C0160797|T046|FN|81642009|SNOMEDCT_CORE|Late effect of spinal cord injury|Late effect of spinal cord injury
C0160814|T046|SY|78523004|SNOMEDCT_CORE|Delayed effect of radiation|Late effect of radiation
C0160814|T046|PT|78523004|SNOMEDCT_CORE|Late effect of radiation|Late effect of radiation
C0160814|T046|FN|78523004|SNOMEDCT_CORE|Late effect of radiation|Late effect of radiation
C0160918|T037|SY|269214009|SNOMEDCT_CORE|Contusion face, scalp and neck, excluding eyes|Contusion of face, scalp and neck, excluding eye
C0160918|T037|PT|269214009|SNOMEDCT_CORE|Contusion of face, scalp and neck, excluding eye|Contusion of face, scalp and neck, excluding eye
C0160918|T037|FN|269214009|SNOMEDCT_CORE|Contusion of face, scalp and neck, excluding eye|Contusion of face, scalp and neck, excluding eye
C0160925|T037|PT|10050004|SNOMEDCT_CORE|Contusion of chest|Contusion of chest
C0160925|T037|FN|10050004|SNOMEDCT_CORE|Contusion of chest|Contusion of chest
C0160925|T037|SY|10050004|SNOMEDCT_CORE|Superficial bruising of chest wall|Contusion of chest
C0160926|T037|PT|37907001|SNOMEDCT_CORE|Contusion of abdominal wall|Contusion of abdominal wall
C0160926|T037|FN|37907001|SNOMEDCT_CORE|Contusion of abdominal wall|Contusion of abdominal wall
C0160926|T037|SY|37907001|SNOMEDCT_CORE|Superficial bruising of abdominal wall|Contusion of abdominal wall
C0160927|T037|PT|11437003|SNOMEDCT_CORE|Contusion of back|Contusion of back
C0160927|T037|FN|11437003|SNOMEDCT_CORE|Contusion of back|Contusion of back
C0160927|T037|SY|11437003|SNOMEDCT_CORE|Superficial bruising of back|Contusion of back
C0160931|T037|SY|68142008|SNOMEDCT_CORE|Arm bruise|Contusion of upper limb
C0160931|T037|SY|68142008|SNOMEDCT_CORE|Contusion of arm|Contusion of upper limb
C0160931|T037|IS|68142008|SNOMEDCT_CORE|Contusion of arm, NOS|Contusion of upper limb
C0160931|T037|PT|68142008|SNOMEDCT_CORE|Contusion of upper limb|Contusion of upper limb
C0160931|T037|FN|68142008|SNOMEDCT_CORE|Contusion of upper limb|Contusion of upper limb
C0160931|T037|IS|68142008|SNOMEDCT_CORE|Contusion of upper limb, NOS|Contusion of upper limb
C0160931|T037|SY|68142008|SNOMEDCT_CORE|Contusion, upper limb|Contusion of upper limb
C0160931|T037|SY|68142008|SNOMEDCT_CORE|Superficial bruising of arm|Contusion of upper limb
C0160931|T037|SY|68142008|SNOMEDCT_CORE|Superficial bruising of upper limb|Contusion of upper limb
C0160933|T037|PT|40257000|SNOMEDCT_CORE|Contusion of shoulder region|Contusion of shoulder region
C0160933|T037|FN|40257000|SNOMEDCT_CORE|Contusion of shoulder region|Contusion of shoulder region
C0160933|T037|SY|40257000|SNOMEDCT_CORE|Contusion, shoulder area|Contusion of shoulder region
C0160933|T037|SY|40257000|SNOMEDCT_CORE|Shoulder bruise|Contusion of shoulder region
C0160943|T037|PT|48123002|SNOMEDCT_CORE|Contusion of wrist|Contusion of wrist
C0160943|T037|FN|48123002|SNOMEDCT_CORE|Contusion of wrist|Contusion of wrist
C0160943|T037|SY|48123002|SNOMEDCT_CORE|Contusion, wrist|Contusion of wrist
C0160943|T037|SY|48123002|SNOMEDCT_CORE|Superficial bruising of wrist|Contusion of wrist
C0160949|T037|PT|84416003|SNOMEDCT_CORE|Contusion of thigh|Contusion of thigh
C0160949|T037|FN|84416003|SNOMEDCT_CORE|Contusion of thigh|Contusion of thigh
C0160949|T037|SY|84416003|SNOMEDCT_CORE|Contusion, thigh|Contusion of thigh
C0160949|T037|SY|84416003|SNOMEDCT_CORE|Superficial bruising of thigh|Contusion of thigh
C0160950|T037|PT|44801007|SNOMEDCT_CORE|Contusion of hip|Contusion of hip
C0160950|T037|FN|44801007|SNOMEDCT_CORE|Contusion of hip|Contusion of hip
C0160950|T037|SY|44801007|SNOMEDCT_CORE|Contusion, hip|Contusion of hip
C0160950|T037|SY|44801007|SNOMEDCT_CORE|Superficial bruising of hip|Contusion of hip
C0160952|T037|PT|45613006|SNOMEDCT_CORE|Contusion of lower leg|Contusion of lower leg
C0160952|T037|FN|45613006|SNOMEDCT_CORE|Contusion of lower leg|Contusion of lower leg
C0160952|T037|SY|45613006|SNOMEDCT_CORE|Contusion, lower leg|Contusion of lower leg
C0160952|T037|SY|45613006|SNOMEDCT_CORE|Leg bruise|Contusion of lower leg
C0160952|T037|SY|45613006|SNOMEDCT_CORE|Superficial bruising of leg|Contusion of lower leg
C0160952|T037|SY|45613006|SNOMEDCT_CORE|Superficial bruising of lower leg|Contusion of lower leg
C0160952|T037|SY|45613006|SNOMEDCT_CORE|Superficial bruising of lower limb|Contusion of lower leg
C0160953|T037|PT|22878006|SNOMEDCT_CORE|Contusion of knee|Contusion of knee
C0160953|T037|FN|22878006|SNOMEDCT_CORE|Contusion of knee|Contusion of knee
C0160953|T037|SY|22878006|SNOMEDCT_CORE|Contusion, knee|Contusion of knee
C0160953|T037|SY|22878006|SNOMEDCT_CORE|Superficial bruising of knee|Contusion of knee
C0160955|T033|PT|74814004|SNOMEDCT_CORE|Contusion of foot|Contusion of foot
C0160955|T033|FN|74814004|SNOMEDCT_CORE|Contusion of foot|Contusion of foot
C0160955|T033|SY|74814004|SNOMEDCT_CORE|Superficial bruising of foot|Contusion of foot
C0160956|T037|PT|55042009|SNOMEDCT_CORE|Contusion of ankle|Contusion of ankle
C0160956|T037|FN|55042009|SNOMEDCT_CORE|Contusion of ankle|Contusion of ankle
C0160956|T037|SY|55042009|SNOMEDCT_CORE|Contusion, ankle|Contusion of ankle
C0160956|T037|SY|55042009|SNOMEDCT_CORE|Superficial bruising of ankle|Contusion of ankle
C0160957|T037|SY|58075000|SNOMEDCT_CORE|Bruise of toe|Contusion of toe
C0160957|T037|PT|58075000|SNOMEDCT_CORE|Contusion of toe|Contusion of toe
C0160957|T037|FN|58075000|SNOMEDCT_CORE|Contusion of toe|Contusion of toe
C0160957|T037|SY|58075000|SNOMEDCT_CORE|Superficial bruising of toe|Contusion of toe
C0160993|T037|SY|43422002|SNOMEDCT_CORE|Crush injury of foot|Crushing injury of foot
C0160993|T037|SY|43422002|SNOMEDCT_CORE|Crush injury to foot|Crushing injury of foot
C0160993|T037|PT|43422002|SNOMEDCT_CORE|Crushing injury of foot|Crushing injury of foot
C0160993|T037|FN|43422002|SNOMEDCT_CORE|Crushing injury of foot|Crushing injury of foot
C0161002|T037|FN|37450000|SNOMEDCT_CORE|Corneal foreign body|Corneal foreign body
C0161002|T037|PT|37450000|SNOMEDCT_CORE|Corneal foreign body|Corneal foreign body
C0161003|T037|PT|52497002|SNOMEDCT_CORE|Foreign body in conjunctival sac|Foreign body in conjunctival sac
C0161003|T037|FN|52497002|SNOMEDCT_CORE|Foreign body in conjunctival sac|Foreign body in conjunctival sac
C0161003|T037|IS|52497002|SNOMEDCT_CORE|Foreign body in conjuntival sac|Foreign body in conjunctival sac
C0161007|T037|PT|75441006|SNOMEDCT_CORE|Foreign body in ear|Foreign body in ear
C0161007|T037|FN|75441006|SNOMEDCT_CORE|Foreign body in ear|Foreign body in ear
C0161008|T033|SY|74699008|SNOMEDCT_CORE|FB - Nasal foreign body|Foreign body in nose
C0161008|T033|PT|74699008|SNOMEDCT_CORE|Foreign body in nose|Foreign body in nose
C0161008|T033|FN|74699008|SNOMEDCT_CORE|Foreign body in nose|Foreign body in nose
C0161010|T037|PT|25479004|SNOMEDCT_CORE|Foreign body in pharynx|Foreign body in pharynx
C0161010|T037|FN|25479004|SNOMEDCT_CORE|Foreign body in pharynx|Foreign body in pharynx
C0161010|T037|SY|25479004|SNOMEDCT_CORE|Foreign body in throat|Foreign body in pharynx
C0161010|T037|IS|25479004|SNOMEDCT_CORE|Foreign body in throat, NOS|Foreign body in pharynx
C0161010|T037|SY|25479004|SNOMEDCT_CORE|Pharyngeal FB - foreign body|Foreign body in pharynx
C0161315|T037|PT|10132008|SNOMEDCT_CORE|Burns of multiple sites|Burns of multiple sites
C0161315|T037|FN|10132008|SNOMEDCT_CORE|Burns of multiple sites|Burns of multiple sites
C0161406|T037|SY|72556006|SNOMEDCT_CORE|Fifth cranial nerve injury|Injury of trigeminal nerve
C0161406|T037|SY|72556006|SNOMEDCT_CORE|Injury of fifth cranial nerve|Injury of trigeminal nerve
C0161406|T037|PT|72556006|SNOMEDCT_CORE|Injury of trigeminal nerve|Injury of trigeminal nerve
C0161406|T037|FN|72556006|SNOMEDCT_CORE|Injury of trigeminal nerve|Injury of trigeminal nerve
C0161406|T037|SY|72556006|SNOMEDCT_CORE|Injury to trigeminal nerve|Injury of trigeminal nerve
C0161406|T037|SY|72556006|SNOMEDCT_CORE|Trigeminal nerve injury|Injury of trigeminal nerve
C0161446|T037|SY|6836001|SNOMEDCT_CORE|Brachial plexus injury|Injury of brachial plexus
C0161446|T037|PT|6836001|SNOMEDCT_CORE|Injury of brachial plexus|Injury of brachial plexus
C0161446|T037|FN|6836001|SNOMEDCT_CORE|Injury of brachial plexus|Injury of brachial plexus
C0161446|T037|SY|6836001|SNOMEDCT_CORE|Traumatic brachial plexus lesion|Injury of brachial plexus
C0161458|T037|PT|62745008|SNOMEDCT_CORE|Injury of ulnar nerve|Injury of ulnar nerve
C0161458|T037|FN|62745008|SNOMEDCT_CORE|Injury of ulnar nerve|Injury of ulnar nerve
C0161470|T037|PT|25604001|SNOMEDCT_CORE|Traumatic injury of common peroneal nerve|Traumatic injury of common peroneal nerve
C0161470|T037|FN|25604001|SNOMEDCT_CORE|Traumatic injury of common peroneal nerve|Traumatic injury of common peroneal nerve
C0161530|T037|SY|67438002|SNOMEDCT_CORE|Anticoagulant poisoning|Poisoning by anticoagulant
C0161530|T037|PT|67438002|SNOMEDCT_CORE|Poisoning by anticoagulant|Poisoning by anticoagulant
C0161530|T037|OF|67438002|SNOMEDCT_CORE|Poisoning by anticoagulant|Poisoning by anticoagulant
C0161530|T037|IS|67438002|SNOMEDCT_CORE|Poisoning by anticoagulant, NOS|Poisoning by anticoagulant
C0161530|T037|FN|67438002|SNOMEDCT_CORE|Poisoning caused by anticoagulant|Poisoning by anticoagulant
C0161530|T037|SY|67438002|SNOMEDCT_CORE|Poisoning caused by anticoagulant|Poisoning by anticoagulant
C0161578|T037|PT|82276009|SNOMEDCT_CORE|Poisoning by antidepressant|Poisoning by antidepressant
C0161578|T037|OF|82276009|SNOMEDCT_CORE|Poisoning by antidepressant|Poisoning by antidepressant
C0161578|T037|SY|82276009|SNOMEDCT_CORE|Poisoning by antidepressant drug|Poisoning by antidepressant
C0161578|T037|IS|82276009|SNOMEDCT_CORE|Poisoning by antidepressant, NOS|Poisoning by antidepressant
C0161578|T037|SY|82276009|SNOMEDCT_CORE|Poisoning caused by antidepressant|Poisoning by antidepressant
C0161578|T037|FN|82276009|SNOMEDCT_CORE|Poisoning caused by antidepressant|Poisoning by antidepressant
C0161578|T037|SY|82276009|SNOMEDCT_CORE|Poisoning caused by antidepressant drug|Poisoning by antidepressant
C0161737|T037|PT|35195001|SNOMEDCT_CORE|Frostbite of foot|Frostbite of foot
C0161737|T037|FN|35195001|SNOMEDCT_CORE|Frostbite of foot|Frostbite of foot
C0161767|T046|PT|79315005|SNOMEDCT_CORE|Mechanical complication due to urethral indwelling catheter|Mechanical complication due to urethral indwelling catheter
C0161767|T046|FN|79315005|SNOMEDCT_CORE|Mechanical complication due to urethral indwelling catheter|Mechanical complication due to urethral indwelling catheter
C0161803|T046|PT|79369007|SNOMEDCT_CORE|Complication of transplanted pancreas|Complication of transplanted pancreas
C0161803|T046|FN|79369007|SNOMEDCT_CORE|Complication of transplanted pancreas|Complication of transplanted pancreas
C0161836|T046|PT|35688006|SNOMEDCT_CORE|Complication of medical care|Complication of medical care
C0161836|T046|FN|35688006|SNOMEDCT_CORE|Complication of medical care|Complication of medical care
C0161836|T046|IS|35688006|SNOMEDCT_CORE|Complication of medical care, NOS|Complication of medical care
C0161836|T046|SY|35688006|SNOMEDCT_CORE|Medical care complication|Complication of medical care
C0162164|T019|PT|67278007|SNOMEDCT_CORE|Congenital stenosis of pulmonary valve|Congenital stenosis of pulmonary valve
C0162164|T019|FN|67278007|SNOMEDCT_CORE|Congenital stenosis of pulmonary valve|Congenital stenosis of pulmonary valve
C0162164|T019|SY|67278007|SNOMEDCT_CORE|Congenital valvular pulmonic stenosis|Congenital stenosis of pulmonary valve
C0162164|T019|SY|67278007|SNOMEDCT_CORE|PV - Congenital pulmonary valve stenosis|Congenital stenosis of pulmonary valve
C0162285|T046|IS|89091004|SNOMEDCT_CORE|Blepharoedema|Edema of eyelid
C0162285|T046|PT|89091004|SNOMEDCT_CORE|Edema of eyelid|Edema of eyelid
C0162285|T046|FN|89091004|SNOMEDCT_CORE|Edema of eyelid|Edema of eyelid
C0162285|T046|SY|89091004|SNOMEDCT_CORE|Hydroblepharon|Edema of eyelid
C0162285|T046|PTGB|89091004|SNOMEDCT_CORE|Oedema of eyelid|Edema of eyelid
C0162296|T047|SY|35678005|SNOMEDCT_CORE|Arthralgia of multiple joints|Multiple joint pain
C0162296|T047|PT|35678005|SNOMEDCT_CORE|Multiple joint pain|Multiple joint pain
C0162296|T047|FN|35678005|SNOMEDCT_CORE|Multiple joint pain|Multiple joint pain
C0162296|T047|SY|35678005|SNOMEDCT_CORE|Polyarthralgia|Multiple joint pain
C0162297|T046|PT|87317003|SNOMEDCT_CORE|Respiratory arrest|Respiratory arrest
C0162297|T046|FN|87317003|SNOMEDCT_CORE|Respiratory arrest|Respiratory arrest
C0162299|T047|PT|72325004|SNOMEDCT_CORE|Cyst of thyroid|Cyst of thyroid
C0162299|T047|FN|72325004|SNOMEDCT_CORE|Cyst of thyroid|Cyst of thyroid
C0162301|T047|PT|20342001|SNOMEDCT_CORE|Calculus in urethra|Calculus in urethra
C0162301|T047|FN|20342001|SNOMEDCT_CORE|Calculus in urethra|Calculus in urethra
C0162301|T047|SY|20342001|SNOMEDCT_CORE|Urethral calculus|Calculus in urethra
C0162301|T047|SY|20342001|SNOMEDCT_CORE|Urethral stone|Calculus in urethra
C0162316|T047|SYGB|87522002|SNOMEDCT_CORE|IDA - Iron deficiency anaemia|Iron deficiency anemia
C0162316|T047|SY|87522002|SNOMEDCT_CORE|IDA - Iron deficiency anemia|Iron deficiency anemia
C0162316|T047|PTGB|87522002|SNOMEDCT_CORE|Iron deficiency anaemia|Iron deficiency anemia
C0162316|T047|SYGB|87522002|SNOMEDCT_CORE|Iron deficiency anaemia syndrome|Iron deficiency anemia
C0162316|T047|PT|87522002|SNOMEDCT_CORE|Iron deficiency anemia|Iron deficiency anemia
C0162316|T047|FN|87522002|SNOMEDCT_CORE|Iron deficiency anemia|Iron deficiency anemia
C0162316|T047|SY|87522002|SNOMEDCT_CORE|Iron deficiency anemia syndrome|Iron deficiency anemia
C0162316|T047|IS|87522002|SNOMEDCT_CORE|Iron deficiency anemia, NOS|Iron deficiency anemia
C0162316|T047|SYGB|87522002|SNOMEDCT_CORE|Sideropenic anaemia|Iron deficiency anemia
C0162316|T047|SY|87522002|SNOMEDCT_CORE|Sideropenic anemia|Iron deficiency anemia
C0162323|T047|SY|417373000|SNOMEDCT_CORE|Inflammatory arthritis of multiple joints|Inflammatory polyarthropathy
C0162323|T047|PT|417373000|SNOMEDCT_CORE|Inflammatory polyarthropathy|Inflammatory polyarthropathy
C0162323|T047|FN|417373000|SNOMEDCT_CORE|Inflammatory polyarthropathy|Inflammatory polyarthropathy
C0162323|T047|SY|416956002|SNOMEDCT_CORE|Polyarthritis|Inflammatory polyarthropathy
C0162351|T046|PT|29268000|SNOMEDCT_CORE|Contact hypersensitivity|Contact hypersensitivity
C0162351|T046|FN|29268000|SNOMEDCT_CORE|Contact hypersensitivity|Contact hypersensitivity
C0162385|T037|PT|127287001|SNOMEDCT_CORE|Intertrochanteric fracture|Intertrochanteric fracture
C0162385|T037|FN|127287001|SNOMEDCT_CORE|Intertrochanteric fracture|Intertrochanteric fracture
C0162385|T037|SY|127287001|SNOMEDCT_CORE|Intertrochanteric fracture of femur|Intertrochanteric fracture
C0162386|T037|SY|263229001|SNOMEDCT_CORE|Subtrochanteric fracture|Subtrochanteric fracture of femur
C0162386|T037|PT|263229001|SNOMEDCT_CORE|Subtrochanteric fracture of femur|Subtrochanteric fracture of femur
C0162386|T037|FN|263229001|SNOMEDCT_CORE|Subtrochanteric fracture of femur|Subtrochanteric fracture of femur
C0162423|T047|SY|72658003|SNOMEDCT_CORE|Heat rash|Prickly heat
C0162423|T047|SY|72658003|SNOMEDCT_CORE|Miliaria rubra|Prickly heat
C0162423|T047|SY|72658003|SNOMEDCT_CORE|Miliaria tropicalis|Prickly heat
C0162423|T047|PT|72658003|SNOMEDCT_CORE|Prickly heat|Prickly heat
C0162423|T047|FN|72658003|SNOMEDCT_CORE|Prickly heat|Prickly heat
C0162429|T047|SY|2492009|SNOMEDCT_CORE|Malnutrition|Malnutrition
C0162429|T047|IS|70241007|SNOMEDCT_CORE|Undernutrition|Malnutrition
C0162451|T047|SY|200823002|SNOMEDCT_CORE|Allergic dermatitis caused by poison ivy|Contact dermatitis due to poison ivy
C0162451|T047|SY|200823002|SNOMEDCT_CORE|Allergic dermatitis caused by Rhus toxicodendron|Contact dermatitis due to poison ivy
C0162451|T047|SY|200823002|SNOMEDCT_CORE|Allergic dermatitis due to poison ivy|Contact dermatitis due to poison ivy
C0162451|T047|SY|200823002|SNOMEDCT_CORE|Allergic dermatitis due to Rhus toxicodendron|Contact dermatitis due to poison ivy
C0162451|T047|SY|200823002|SNOMEDCT_CORE|Contact dermatitis caused by poison ivy|Contact dermatitis due to poison ivy
C0162451|T047|FN|200823002|SNOMEDCT_CORE|Contact dermatitis caused by poison ivy|Contact dermatitis due to poison ivy
C0162451|T047|SY|200823002|SNOMEDCT_CORE|Contact dermatitis caused by poison-ivy|Contact dermatitis due to poison ivy
C0162451|T047|SY|200823002|SNOMEDCT_CORE|Contact dermatitis caused by Rhus toxicodendron|Contact dermatitis due to poison ivy
C0162451|T047|PT|200823002|SNOMEDCT_CORE|Contact dermatitis due to poison ivy|Contact dermatitis due to poison ivy
C0162451|T047|OF|200823002|SNOMEDCT_CORE|Contact dermatitis due to poison ivy|Contact dermatitis due to poison ivy
C0162451|T047|SY|200823002|SNOMEDCT_CORE|Contact dermatitis due to poison-ivy|Contact dermatitis due to poison ivy
C0162451|T047|OF|200823002|SNOMEDCT_CORE|Contact dermatitis due to poison-ivy|Contact dermatitis due to poison ivy
C0162451|T047|SY|200823002|SNOMEDCT_CORE|Contact dermatitis due to Rhus toxicodendron|Contact dermatitis due to poison ivy
C0162529|T047|SYGB|30588004|SNOMEDCT_CORE|Colonic ischaemia|Ischemic colitis
C0162529|T047|SY|30588004|SNOMEDCT_CORE|Colonic ischemia|Ischemic colitis
C0162529|T047|PTGB|30588004|SNOMEDCT_CORE|Ischaemic colitis|Ischemic colitis
C0162529|T047|IS|30588004|SNOMEDCT_CORE|Ischaemic colitis, NOS|Ischemic colitis
C0162529|T047|PT|30588004|SNOMEDCT_CORE|Ischemic colitis|Ischemic colitis
C0162529|T047|FN|30588004|SNOMEDCT_CORE|Ischemic colitis|Ischemic colitis
C0162529|T047|IS|30588004|SNOMEDCT_CORE|Ischemic colitis, NOS|Ischemic colitis
C0162538|T047|SY|29260007|SNOMEDCT_CORE|IgA deficiency|Immunoglobulin A deficiency
C0162538|T047|FN|29260007|SNOMEDCT_CORE|Immunoglobulin A deficiency|Immunoglobulin A deficiency
C0162538|T047|PT|29260007|SNOMEDCT_CORE|Immunoglobulin A deficiency|Immunoglobulin A deficiency
C0162557|T047|PT|197270009|SNOMEDCT_CORE|Acute hepatic failure|Acute hepatic failure
C0162557|T047|FN|197270009|SNOMEDCT_CORE|Acute hepatic failure|Acute hepatic failure
C0162557|T047|SY|197270009|SNOMEDCT_CORE|Acute liver failure|Acute hepatic failure
C0162557|T047|SY|197270009|SNOMEDCT_CORE|ALF - Acute liver failure|Acute hepatic failure
C0162670|T047|PT|16851005|SNOMEDCT_CORE|Mitochondrial myopathy|Mitochondrial myopathy
C0162670|T047|FN|16851005|SNOMEDCT_CORE|Mitochondrial myopathy|Mitochondrial myopathy
C0162670|T047|SY|16851005|SNOMEDCT_CORE|Ragged red myopathy|Mitochondrial myopathy
C0162678|T191|SY|19133005|SNOMEDCT_CORE|Clinical neurofibromatosis|Neurofibromatosis syndrome
C0162678|T191|PT|19133005|SNOMEDCT_CORE|Neurofibromatosis syndrome|Neurofibromatosis syndrome
C0162678|T191|FN|19133005|SNOMEDCT_CORE|Neurofibromatosis syndrome|Neurofibromatosis syndrome
C0162678|T191|SY|19133005|SNOMEDCT_CORE|NF - Neurofibromatosis|Neurofibromatosis syndrome
C0162809|T047|IS|33927004|SNOMEDCT_CORE|Anosmia eunuchoidism|Olfactogenital dysplasia
C0162809|T047|IS|33927004|SNOMEDCT_CORE|Dysplasia olfactogenitalis of de Morsier|Olfactogenital dysplasia
C0162809|T047|IS|33927004|SNOMEDCT_CORE|Kallman syndrome|Olfactogenital dysplasia
C0162809|T047|IS|33927004|SNOMEDCT_CORE|Olfactogenital dysplasia|Olfactogenital dysplasia
C0162810|T020|OAP|267821008|SNOMEDCT_CORE|Hypertrophic cicatrix|Hypertrophic scar
C0162810|T020|SY|19843006|SNOMEDCT_CORE|Hypertrophic cicatrix|Hypertrophic scar
C0162810|T020|OAF|267821008|SNOMEDCT_CORE|Hypertrophic cicatrix|Hypertrophic scar
C0162810|T020|PT|19843006|SNOMEDCT_CORE|Hypertrophic scar|Hypertrophic scar
C0162810|T020|FN|19843006|SNOMEDCT_CORE|Hypertrophic scar|Hypertrophic scar
C0162810|T020|IS|19843006|SNOMEDCT_CORE|Hypertrophic scar of skin|Hypertrophic scar
C0162820|T047|SY|238575004|SNOMEDCT_CORE|ACD - Allergic contact dermatitis|Allergic contact dermatitis
C0162820|T047|PT|238575004|SNOMEDCT_CORE|Allergic contact dermatitis|Allergic contact dermatitis
C0162820|T047|FN|238575004|SNOMEDCT_CORE|Allergic contact dermatitis|Allergic contact dermatitis
C0162823|T047|SY|110979008|SNOMEDCT_CORE|ICD - Irritant contact dermatitis|Irritant contact dermatitis
C0162823|T047|PT|110979008|SNOMEDCT_CORE|Irritant contact dermatitis|Irritant contact dermatitis
C0162823|T047|FN|110979008|SNOMEDCT_CORE|Irritant contact dermatitis|Irritant contact dermatitis
C0162823|T047|SY|110979008|SNOMEDCT_CORE|Non-allergic contact dermatitis|Irritant contact dermatitis
C0162823|T047|SY|110979008|SNOMEDCT_CORE|Primary irritant dermatitis|Irritant contact dermatitis
C0162823|T047|OF|110979008|SNOMEDCT_CORE|Primary irritant dermatitis|Irritant contact dermatitis
C0162834|T046|SY|49765009|SNOMEDCT_CORE|Hyperpigmentation|Hyperpigmentation of skin
C0162834|T046|SY|49765009|SNOMEDCT_CORE|Hyperpigmentation disorder|Hyperpigmentation of skin
C0162834|T046|PT|49765009|SNOMEDCT_CORE|Hyperpigmentation of skin|Hyperpigmentation of skin
C0162834|T046|FN|49765009|SNOMEDCT_CORE|Hyperpigmentation of skin|Hyperpigmentation of skin
C0162834|T046|IS|49765009|SNOMEDCT_CORE|Hyperpigmentation of skin, NOS|Hyperpigmentation of skin
C0162836|T047|SY|59393003|SNOMEDCT_CORE|Apocrine acne|Hidradenitis suppurativa
C0162836|T047|SY|59393003|SNOMEDCT_CORE|Hidradenitis axillaris|Hidradenitis suppurativa
C0162836|T047|PT|59393003|SNOMEDCT_CORE|Hidradenitis suppurativa|Hidradenitis suppurativa
C0162836|T047|FN|59393003|SNOMEDCT_CORE|Hidradenitis suppurativa|Hidradenitis suppurativa
C0162836|T047|SY|59393003|SNOMEDCT_CORE|Suppurative hidradenitis|Hidradenitis suppurativa
C0162836|T047|SY|59393003|SNOMEDCT_CORE|Verneuil's disease|Hidradenitis suppurativa
C0162870|T190|PT|13290008|SNOMEDCT_CORE|Aneurysm of iliac artery|Aneurysm of iliac artery
C0162870|T190|FN|13290008|SNOMEDCT_CORE|Aneurysm of iliac artery|Aneurysm of iliac artery
C0162871|T047|SY|233985008|SNOMEDCT_CORE|AAA - Abdominal aortic aneurysm|Abdominal aortic aneurysm
C0162871|T047|PT|233985008|SNOMEDCT_CORE|Abdominal aortic aneurysm|Abdominal aortic aneurysm
C0162871|T047|FN|233985008|SNOMEDCT_CORE|Abdominal aortic aneurysm|Abdominal aortic aneurysm
C0162872|T047|PT|433068007|SNOMEDCT_CORE|Aneurysm of thoracic aorta|Aneurysm of thoracic aorta
C0162872|T047|FN|433068007|SNOMEDCT_CORE|Aneurysm of thoracic aorta|Aneurysm of thoracic aorta
C0175708|T047|SY|87648004|SNOMEDCT_CORE|Chronic rheumatic carditis|Chronic rheumatic heart disease
C0175708|T047|PT|87648004|SNOMEDCT_CORE|Chronic rheumatic heart disease|Chronic rheumatic heart disease
C0175708|T047|FN|87648004|SNOMEDCT_CORE|Chronic rheumatic heart disease|Chronic rheumatic heart disease
C0176005|T033|PT|218246003|SNOMEDCT_CORE|Late effect of accidental injury|Late effect of accidental injury
C0176005|T033|FN|218246003|SNOMEDCT_CORE|Late effect of accidental injury|Late effect of accidental injury
C0176005|T033|IS|218246003|SNOMEDCT_CORE|Late effects of accidental injury|Late effect of accidental injury
C0176005|T033|OF|218246003|SNOMEDCT_CORE|Late effects of accidental injury|Late effect of accidental injury
C0178274|T047|OAP|266259002|SNOMEDCT_CORE|Arterial, arteriole and capillary disease|Arterial, arteriole and capillary disease
C0178274|T047|OAF|266259002|SNOMEDCT_CORE|Arterial, arteriole and capillary disease|Arterial, arteriole and capillary disease
C0178282|T190|SY|52515009|SNOMEDCT_CORE|Abdominal hernia|Hernia of abdominal cavity
C0178282|T190|PT|52515009|SNOMEDCT_CORE|Hernia of abdominal cavity|Hernia of abdominal cavity
C0178282|T190|FN|52515009|SNOMEDCT_CORE|Hernia of abdominal cavity|Hernia of abdominal cavity
C0178282|T190|IS|52515009|SNOMEDCT_CORE|Hernia of abdominal cavity, NOS|Hernia of abdominal cavity
C0178283|T047|PT|307418008|SNOMEDCT_CORE|Non-infective enteritis and colitis|Non-infective enteritis and colitis
C0178283|T047|FN|307418008|SNOMEDCT_CORE|Non-infective enteritis and colitis|Non-infective enteritis and colitis
C0178298|T047|IS|80659006|SNOMEDCT_CORE|Disease of skin and subcutaneous tissue, NOS|Disorder of skin and/or subcutaneous tissue
C0178298|T047|OF|80659006|SNOMEDCT_CORE|Disease of skin AND/OR subcutaneous tissue|Disorder of skin and/or subcutaneous tissue
C0178298|T047|IS|80659006|SNOMEDCT_CORE|Disease of skin AND/OR subcutaneous tissue|Disorder of skin and/or subcutaneous tissue
C0178298|T047|SY|80659006|SNOMEDCT_CORE|Disorder of skin and subcutaneous tissue|Disorder of skin and/or subcutaneous tissue
C0178298|T047|FN|80659006|SNOMEDCT_CORE|Disorder of skin and/or subcutaneous tissue|Disorder of skin and/or subcutaneous tissue
C0178298|T047|OF|80659006|SNOMEDCT_CORE|Disorder of skin AND/OR subcutaneous tissue|Disorder of skin and/or subcutaneous tissue
C0178298|T047|PT|80659006|SNOMEDCT_CORE|Disorder of skin and/or subcutaneous tissue|Disorder of skin and/or subcutaneous tissue
C0178298|T047|OP|80659006|SNOMEDCT_CORE|Disorder of skin AND/OR subcutaneous tissue|Disorder of skin and/or subcutaneous tissue
C0178298|T047|SY|80659006|SNOMEDCT_CORE|Disorder of the dermis and subcutaneous tissue|Disorder of skin and/or subcutaneous tissue
C0178298|T047|SY|80659006|SNOMEDCT_CORE|Skin and subcutaneous tissue disease|Disorder of skin and/or subcutaneous tissue
C0178316|T037|SY|23406007|SNOMEDCT_CORE|Arm fracture|Fracture of upper limb
C0178316|T037|SY|23406007|SNOMEDCT_CORE|Fracture of arm|Fracture of upper limb
C0178316|T037|IS|23406007|SNOMEDCT_CORE|Fracture of arm, NOS|Fracture of upper limb
C0178316|T037|SY|23406007|SNOMEDCT_CORE|Fracture of bone of upper limb|Fracture of upper limb
C0178316|T037|PT|23406007|SNOMEDCT_CORE|Fracture of upper limb|Fracture of upper limb
C0178316|T037|FN|23406007|SNOMEDCT_CORE|Fracture of upper limb|Fracture of upper limb
C0178316|T037|IS|23406007|SNOMEDCT_CORE|Fracture of upper limb, NOS|Fracture of upper limb
C0178323|T037|PT|26947005|SNOMEDCT_CORE|Open wound of lower limb|Open wound of lower limb
C0178323|T037|FN|26947005|SNOMEDCT_CORE|Open wound of lower limb|Open wound of lower limb
C0178323|T037|IS|26947005|SNOMEDCT_CORE|Open wound of lower limb, NOS|Open wound of lower limb
C0178405|T033|PT|129903002|SNOMEDCT_CORE|Ineffective infant feeding pattern|Ineffective infant feeding pattern
C0178405|T033|FN|129903002|SNOMEDCT_CORE|Ineffective infant feeding pattern|Ineffective infant feeding pattern
C0178415|T033|SY|396152005|SNOMEDCT_CORE|Elevated PSA|Raised prostate specific antigen
C0178415|T033|PT|396152005|SNOMEDCT_CORE|Raised prostate specific antigen|Raised prostate specific antigen
C0178415|T033|FN|396152005|SNOMEDCT_CORE|Raised prostate specific antigen|Raised prostate specific antigen
C0178415|T033|SY|396152005|SNOMEDCT_CORE|Raised PSA|Raised prostate specific antigen
C0178421|T191|SY|254845004|SNOMEDCT_CORE|Breast mouse|Fibroadenoma of breast
C0178421|T191|PT|254845004|SNOMEDCT_CORE|Fibroadenoma of breast|Fibroadenoma of breast
C0178421|T191|FN|254845004|SNOMEDCT_CORE|Fibroadenoma of breast|Fibroadenoma of breast
C0178671|T037|PT|282749008|SNOMEDCT_CORE|Head and neck injury|Head and neck injury
C0178671|T037|FN|282749008|SNOMEDCT_CORE|Head and neck injury|Head and neck injury
C0178879|T047|SY|7163005|SNOMEDCT_CORE|Obstructive uropathy|Urinary tract obstruction
C0178879|T047|IS|7163005|SNOMEDCT_CORE|Obstructive uropathy, NOS|Urinary tract obstruction
C0178879|T047|PT|7163005|SNOMEDCT_CORE|Urinary tract obstruction|Urinary tract obstruction
C0178879|T047|FN|7163005|SNOMEDCT_CORE|Urinary tract obstruction|Urinary tract obstruction
C0178879|T047|IS|7163005|SNOMEDCT_CORE|Urinary tract obstruction, NOS|Urinary tract obstruction
C0184543|T033|SY|129836000|SNOMEDCT_CORE|Nonadherence with therapeutic regimen|Noncompliance with therapeutic regimen
C0184543|T033|PT|129836000|SNOMEDCT_CORE|Noncompliance with therapeutic regimen|Noncompliance with therapeutic regimen
C0184543|T033|FN|129836000|SNOMEDCT_CORE|Noncompliance with therapeutic regimen|Noncompliance with therapeutic regimen
C0184543|T033|SY|129836000|SNOMEDCT_CORE|Noncompliance: therapeutic regimen|Noncompliance with therapeutic regimen
C0184567|T184|PT|274663001|SNOMEDCT_CORE|Acute pain|Acute pain
C0184567|T184|FN|274663001|SNOMEDCT_CORE|Acute pain|Acute pain
C0205642|T191|SY|57596004|SNOMEDCT_CORE|Follicular carcinoma, oxyphilic cell|Oxyphilic adenocarcinoma
C0205642|T191|SY|57596004|SNOMEDCT_CORE|Hurthle cell adenocarcinoma|Oxyphilic adenocarcinoma
C0205642|T191|SY|57596004|SNOMEDCT_CORE|Hurthle cell carcinoma|Oxyphilic adenocarcinoma
C0205642|T191|SY|57596004|SNOMEDCT_CORE|Oncocytic adenocarcinoma|Oxyphilic adenocarcinoma
C0205642|T191|SY|57596004|SNOMEDCT_CORE|Oncocytic carcinoma|Oxyphilic adenocarcinoma
C0205642|T191|PT|443261008|SNOMEDCT_CORE|Oxyphilic adenocarcinoma|Oxyphilic adenocarcinoma
C0205642|T191|PT|57596004|SNOMEDCT_CORE|Oxyphilic adenocarcinoma|Oxyphilic adenocarcinoma
C0205642|T191|FN|57596004|SNOMEDCT_CORE|Oxyphilic adenocarcinoma|Oxyphilic adenocarcinoma
C0205642|T191|FN|443261008|SNOMEDCT_CORE|Oxyphilic adenocarcinoma|Oxyphilic adenocarcinoma
C0205699|T191|PT|307593001|SNOMEDCT_CORE|Carcinomatosis|Carcinomatosis
C0205699|T191|FN|307593001|SNOMEDCT_CORE|Carcinomatosis|Carcinomatosis
C0205699|T191|SY|307593001|SNOMEDCT_CORE|Disseminated carcinomatosis|Carcinomatosis
C0205748|T191|SYGB|254818000|SNOMEDCT_CORE|Atypical naevus of skin|Dysplastic nevus of skin
C0205748|T191|SY|254818000|SNOMEDCT_CORE|Atypical nevus of skin|Dysplastic nevus of skin
C0205748|T191|PTGB|254818000|SNOMEDCT_CORE|Dysplastic naevus of skin|Dysplastic nevus of skin
C0205748|T191|PT|254818000|SNOMEDCT_CORE|Dysplastic nevus of skin|Dysplastic nevus of skin
C0205748|T191|FN|254818000|SNOMEDCT_CORE|Dysplastic nevus of skin|Dysplastic nevus of skin
C0205765|T047|SY|27431007|SNOMEDCT_CORE|Chronic cystic mastitis|Chronic cystic mastitis
C0205792|T190|SY|398061002|SNOMEDCT_CORE|Enterocele|Vaginal enterocele
C0205792|T190|SY|398061002|SNOMEDCT_CORE|Hernia into pouch of Douglas|Vaginal enterocele
C0205792|T190|SY|398061002|SNOMEDCT_CORE|Posterior vaginal hernia|Vaginal enterocele
C0205792|T190|SY|398061002|SNOMEDCT_CORE|Pouch of Douglas hernia|Vaginal enterocele
C0205792|T190|PT|398061002|SNOMEDCT_CORE|Vaginal enterocele|Vaginal enterocele
C0205792|T190|FN|398061002|SNOMEDCT_CORE|Vaginal enterocele|Vaginal enterocele
C0205851|T191|SY|402878003|SNOMEDCT_CORE|Germ cell neoplasm|Germ cell tumor
C0205851|T191|PT|402878003|SNOMEDCT_CORE|Germ cell tumor|Germ cell tumor
C0205851|T191|FN|402878003|SNOMEDCT_CORE|Germ cell tumor|Germ cell tumor
C0205851|T191|PTGB|402878003|SNOMEDCT_CORE|Germ cell tumour|Germ cell tumor
C0205929|T020|IS|72779005|SNOMEDCT_CORE|Fistula in ano|Fistula-in-ano
C0205929|T020|IS|72779005|SNOMEDCT_CORE|Fistula-in-ano|Fistula-in-ano
C0205969|T191|SY|128717008|SNOMEDCT_CORE|Thymic carcinoma|Thymoma, type C
C0205969|T191|FN|128717008|SNOMEDCT_CORE|Thymoma, type C|Thymoma, type C
C0205969|T191|PT|128717008|SNOMEDCT_CORE|Thymoma, type C|Thymoma, type C
C0205969|T191|PT|444374006|SNOMEDCT_CORE|Type C thymoma|Thymoma, type C
C0205969|T191|FN|444374006|SNOMEDCT_CORE|Type C thymoma|Thymoma, type C
C0205990|T020|PT|398022005|SNOMEDCT_CORE|Vaginal wall prolapse|Vaginal wall prolapse
C0205990|T020|FN|398022005|SNOMEDCT_CORE|Vaginal wall prolapse|Vaginal wall prolapse
C0206051|T047|IS|90128006|SNOMEDCT_CORE|Photoallergy|Photoallergy
C0206061|T047|PT|64667001|SNOMEDCT_CORE|Interstitial pneumonia|Interstitial pneumonia
C0206061|T047|FN|64667001|SNOMEDCT_CORE|Interstitial pneumonia|Interstitial pneumonia
C0206061|T047|SY|64667001|SNOMEDCT_CORE|Interstitial pneumonitis|Interstitial pneumonia
C0206062|T047|SY|233703007|SNOMEDCT_CORE|Diffuse parenchymal lung disease|Interstitial lung disease
C0206062|T047|SY|233703007|SNOMEDCT_CORE|ILD - Interstitial lung disease|Interstitial lung disease
C0206062|T047|IS|64667001|SNOMEDCT_CORE|Interstitial lung disease|Interstitial lung disease
C0206062|T047|PT|233703007|SNOMEDCT_CORE|Interstitial lung disease|Interstitial lung disease
C0206062|T047|FN|233703007|SNOMEDCT_CORE|Interstitial lung disease|Interstitial lung disease
C0206064|T047|PT|233845001|SNOMEDCT_CORE|Cardiac syndrome X|Cardiac syndrome X
C0206064|T047|FN|233845001|SNOMEDCT_CORE|Cardiac syndrome X|Cardiac syndrome X
C0206064|T047|SY|233845001|SNOMEDCT_CORE|Chest pain with normal coronary angiography|Cardiac syndrome X
C0206064|T047|SY|233845001|SNOMEDCT_CORE|Coronary microvascular disease|Cardiac syndrome X
C0206064|T047|SY|233845001|SNOMEDCT_CORE|Coronary small artery disease|Cardiac syndrome X
C0206064|T047|SY|233845001|SNOMEDCT_CORE|Microvascular angina|Cardiac syndrome X
C0206073|T048|PT|404189009|SNOMEDCT_CORE|Domestic violence|Domestic violence
C0206073|T048|OF|404189009|SNOMEDCT_CORE|Domestic violence|Domestic violence
C0206073|T048|FN|404189009|SNOMEDCT_CORE|Domestic violence|Domestic violence
C0206139|T047|SY|235049008|SNOMEDCT_CORE|OLP - Oral lichen planus|Oral lichen planus
C0206139|T047|PT|235049008|SNOMEDCT_CORE|Oral lichen planus|Oral lichen planus
C0206139|T047|FN|235049008|SNOMEDCT_CORE|Oral lichen planus|Oral lichen planus
C0206141|T047|IS|423294001|SNOMEDCT_CORE|HES|Idiopathic hypereosinophilic syndrome
C0206141|T047|IS|423294001|SNOMEDCT_CORE|Hypereosinophilic syndrome|Idiopathic hypereosinophilic syndrome
C0206141|T047|PT|423294001|SNOMEDCT_CORE|Idiopathic hypereosinophilic syndrome|Idiopathic hypereosinophilic syndrome
C0206141|T047|FN|423294001|SNOMEDCT_CORE|Idiopathic hypereosinophilic syndrome|Idiopathic hypereosinophilic syndrome
C0206141|T047|SY|423294001|SNOMEDCT_CORE|Idiopathic hypereosinophilic syndrome|Idiopathic hypereosinophilic syndrome
C0206180|T191|PT|277637000|SNOMEDCT_CORE|Large cell anaplastic lymphoma|Large cell anaplastic lymphoma
C0206180|T191|FN|277637000|SNOMEDCT_CORE|Large cell anaplastic lymphoma|Large cell anaplastic lymphoma
C0206239|T037|PT|56177003|SNOMEDCT_CORE|Cubital tunnel syndrome|Cubital tunnel syndrome
C0206239|T037|FN|56177003|SNOMEDCT_CORE|Cubital tunnel syndrome|Cubital tunnel syndrome
C0206368|T047|SY|111514006|SNOMEDCT_CORE|Glaucoma capsulare|Pseudoexfoliation glaucoma
C0206368|T047|PT|111514006|SNOMEDCT_CORE|Pseudoexfoliation glaucoma|Pseudoexfoliation glaucoma
C0206368|T047|FN|111514006|SNOMEDCT_CORE|Pseudoexfoliation glaucoma|Pseudoexfoliation glaucoma
C0206368|T047|SY|44219007|SNOMEDCT_CORE|Pseudoexfoliation syndrome|Pseudoexfoliation glaucoma
C0206368|T047|SY|111514006|SNOMEDCT_CORE|Secondary open-angle glaucoma with pseudoexfoliation|Pseudoexfoliation glaucoma
C0206504|T037|SY|60442001|SNOMEDCT_CORE|Perforated eardrum|Perforation of tympanic membrane
C0206504|T037|SY|60442001|SNOMEDCT_CORE|Perforation of ear drum|Perforation of tympanic membrane
C0206504|T037|IS|60442001|SNOMEDCT_CORE|Perforation of ear drum, NOS|Perforation of tympanic membrane
C0206504|T037|SY|60442001|SNOMEDCT_CORE|Perforation of eardrum|Perforation of tympanic membrane
C0206504|T037|PT|60442001|SNOMEDCT_CORE|Perforation of tympanic membrane|Perforation of tympanic membrane
C0206504|T037|FN|60442001|SNOMEDCT_CORE|Perforation of tympanic membrane|Perforation of tympanic membrane
C0206504|T037|IS|60442001|SNOMEDCT_CORE|Perforation of tympanic membrane, NOS|Perforation of tympanic membrane
C0206504|T037|SY|60442001|SNOMEDCT_CORE|Perforation tympanic membrane|Perforation of tympanic membrane
C0206586|T047|PT|9794007|SNOMEDCT_CORE|Endolymphatic hydrops|Endolymphatic hydrops
C0206586|T047|FN|9794007|SNOMEDCT_CORE|Endolymphatic hydrops|Endolymphatic hydrops
C0206624|T191|PT|109843000|SNOMEDCT_CORE|Hepatoblastoma|Hepatoblastoma
C0206624|T191|OP|109843000|SNOMEDCT_CORE|Hepatoblastoma|Hepatoblastoma
C0206624|T191|FN|109843000|SNOMEDCT_CORE|Hepatoblastoma|Hepatoblastoma
C0206624|T191|SY|109843000|SNOMEDCT_CORE|Hepatoblastoma of liver|Hepatoblastoma
C0206646|T191|SY|400153009|SNOMEDCT_CORE|Abdominal desmoid tumor|Abdominal fibromatosis
C0206646|T191|SYGB|400153009|SNOMEDCT_CORE|Abdominal desmoid tumour|Abdominal fibromatosis
C0206646|T191|PT|400153009|SNOMEDCT_CORE|Abdominal fibromatosis|Abdominal fibromatosis
C0206646|T191|FN|400153009|SNOMEDCT_CORE|Abdominal fibromatosis|Abdominal fibromatosis
C0206667|T191|PT|302826002|SNOMEDCT_CORE|Adrenal cortical adenoma|Adrenal cortical adenoma
C0206667|T191|FN|302826002|SNOMEDCT_CORE|Adrenal cortical adenoma|Adrenal cortical adenoma
C0206682|T191|PT|255028004|SNOMEDCT_CORE|Follicular thyroid carcinoma|Follicular thyroid carcinoma
C0206682|T191|FN|255028004|SNOMEDCT_CORE|Follicular thyroid carcinoma|Follicular thyroid carcinoma
C0206682|T191|SY|255028004|SNOMEDCT_CORE|FTC - follicular thyroid carcinoma|Follicular thyroid carcinoma
C0206682|T191|IS|255028004|SNOMEDCT_CORE|FTC - Follicular thyroid carcinoma|Follicular thyroid carcinoma
C0206686|T191|PT|255035007|SNOMEDCT_CORE|Adrenal carcinoma|Adrenal carcinoma
C0206686|T191|FN|255035007|SNOMEDCT_CORE|Adrenal carcinoma|Adrenal carcinoma
C0206686|T191|SY|255035007|SNOMEDCT_CORE|Adrenal cortical adenocarcinoma|Adrenal carcinoma
C0206698|T191|PT|312104005|SNOMEDCT_CORE|Cholangiocarcinoma of biliary tract|Cholangiocarcinoma of biliary tract
C0206698|T191|FN|312104005|SNOMEDCT_CORE|Cholangiocarcinoma of biliary tract|Cholangiocarcinoma of biliary tract
C0206708|T191|PT|285636001|SNOMEDCT_CORE|Cervical intraepithelial neoplasia|Cervical intraepithelial neoplasia
C0206708|T191|FN|285636001|SNOMEDCT_CORE|Cervical intraepithelial neoplasia|Cervical intraepithelial neoplasia
C0206708|T191|SY|285636001|SNOMEDCT_CORE|CIN - Cervical intraepithelial neoplasia|Cervical intraepithelial neoplasia
C0206717|T191|SYGB|422886007|SNOMEDCT_CORE|Aesthesioneuroblastoma|Olfactory neuroblastoma
C0206717|T191|SY|422886007|SNOMEDCT_CORE|Esthesioneuroblastoma|Olfactory neuroblastoma
C0206717|T191|PT|422886007|SNOMEDCT_CORE|Olfactory neuroblastoma|Olfactory neuroblastoma
C0206717|T191|FN|422886007|SNOMEDCT_CORE|Olfactory neuroblastoma|Olfactory neuroblastoma
C0206733|T191|SY|195382003|SNOMEDCT_CORE|Capillary angioma|Capillary angioma
C0206737|T191|SYGB|302838006|SNOMEDCT_CORE|Cellular naevus|Dermal cellular nevus
C0206737|T191|SY|302838006|SNOMEDCT_CORE|Cellular nevus|Dermal cellular nevus
C0206737|T191|PTGB|302838006|SNOMEDCT_CORE|Dermal cellular naevus|Dermal cellular nevus
C0206737|T191|PT|302838006|SNOMEDCT_CORE|Dermal cellular nevus|Dermal cellular nevus
C0206737|T191|FN|302838006|SNOMEDCT_CORE|Dermal cellular nevus|Dermal cellular nevus
C0206737|T191|SYGB|302838006|SNOMEDCT_CORE|Dermal naevus|Dermal cellular nevus
C0206737|T191|SY|302838006|SNOMEDCT_CORE|Dermal nevus|Dermal cellular nevus
C0206737|T191|SYGB|302838006|SNOMEDCT_CORE|IDN - Intradermal naevus|Dermal cellular nevus
C0206737|T191|SY|302838006|SNOMEDCT_CORE|IDN - Intradermal nevus|Dermal cellular nevus
C0206737|T191|SYGB|302838006|SNOMEDCT_CORE|Intradermal melanocytic naevus|Dermal cellular nevus
C0206737|T191|SY|302838006|SNOMEDCT_CORE|Intradermal melanocytic nevus|Dermal cellular nevus
C0220636|T191|SY|255072001|SNOMEDCT_CORE|CA - Cancer of salivary gland|Malignant tumor of salivary gland
C0220636|T191|SY|255072001|SNOMEDCT_CORE|Cancer of salivary gland|Malignant tumor of salivary gland
C0220636|T191|PT|255072001|SNOMEDCT_CORE|Malignant tumor of salivary gland|Malignant tumor of salivary gland
C0220636|T191|FN|255072001|SNOMEDCT_CORE|Malignant tumor of salivary gland|Malignant tumor of salivary gland
C0220636|T191|PTGB|255072001|SNOMEDCT_CORE|Malignant tumour of salivary gland|Malignant tumor of salivary gland
C0220636|T191|SY|255072001|SNOMEDCT_CORE|Salivary gland cancer|Malignant tumor of salivary gland
C0220650|T191|SY|94225005|SNOMEDCT_CORE|Cancer metastatic to brain|Secondary malignant neoplasm of brain
C0220650|T191|SY|94225005|SNOMEDCT_CORE|Metastasis to brain|Secondary malignant neoplasm of brain
C0220650|T191|SY|94225005|SNOMEDCT_CORE|Metastatic malignant neoplasm to brain|Secondary malignant neoplasm of brain
C0220650|T191|IS|94225005|SNOMEDCT_CORE|Metastatic malignant neoplasm to brain, NOS|Secondary malignant neoplasm of brain
C0220650|T191|SY|94225005|SNOMEDCT_CORE|Secondary cancer of brain|Secondary malignant neoplasm of brain
C0220650|T191|PT|94225005|SNOMEDCT_CORE|Secondary malignant neoplasm of brain|Secondary malignant neoplasm of brain
C0220650|T191|FN|94225005|SNOMEDCT_CORE|Secondary malignant neoplasm of brain|Secondary malignant neoplasm of brain
C0220650|T191|IS|94225005|SNOMEDCT_CORE|Secondary malignant neoplasm of brain, NOS|Secondary malignant neoplasm of brain
C0220654|T191|SY|230156002|SNOMEDCT_CORE|Carcinomatous meningitis|Malignant meningitis
C0220654|T191|PT|230156002|SNOMEDCT_CORE|Malignant meningitis|Malignant meningitis
C0220654|T191|FN|230156002|SNOMEDCT_CORE|Malignant meningitis|Malignant meningitis
C0220654|T191|SY|230156002|SNOMEDCT_CORE|Meningeal carcinomatosis|Malignant meningitis
C0220656|T191|PT|236005001|SNOMEDCT_CORE|Malignant ascites|Malignant ascites
C0220656|T191|FN|236005001|SNOMEDCT_CORE|Malignant ascites|Malignant ascites
C0220870|T184|SY|386705008|SNOMEDCT_CORE|Dizziness - light-headed|Lightheadedness
C0220870|T184|SY|386705008|SNOMEDCT_CORE|Feels light headed|Lightheadedness
C0220870|T184|SY|386705008|SNOMEDCT_CORE|Light-headedness|Lightheadedness
C0220870|T184|SY|386705008|SNOMEDCT_CORE|Lightheaded|Lightheadedness
C0220870|T184|PT|386705008|SNOMEDCT_CORE|Lightheadedness|Lightheadedness
C0220870|T184|FN|386705008|SNOMEDCT_CORE|Lightheadedness|Lightheadedness
C0220981|T046|PT|59455009|SNOMEDCT_CORE|Metabolic acidosis|Metabolic acidosis
C0220981|T046|FN|59455009|SNOMEDCT_CORE|Metabolic acidosis|Metabolic acidosis
C0220981|T046|IS|59455009|SNOMEDCT_CORE|Metabolic acidosis, NOS|Metabolic acidosis
C0221002|T047|PT|36348003|SNOMEDCT_CORE|Primary hyperparathyroidism|Primary hyperparathyroidism
C0221002|T047|FN|36348003|SNOMEDCT_CORE|Primary hyperparathyroidism|Primary hyperparathyroidism
C0221013|T191|SY|397016004|SNOMEDCT_CORE|SMCD - systemic mast cell disease|Systemic mast cell disease
C0221013|T191|PT|397016004|SNOMEDCT_CORE|Systemic mast cell disease|Systemic mast cell disease
C0221013|T191|FN|397016004|SNOMEDCT_CORE|Systemic mast cell disease|Systemic mast cell disease
C0221013|T191|SY|397016004|SNOMEDCT_CORE|Systemic mastocytosis|Systemic mast cell disease
C0221047|T047|SY|74615001|SNOMEDCT_CORE|Brady-tachy syndrome|Tachycardia-bradycardia
C0221047|T047|SY|74615001|SNOMEDCT_CORE|Bradycardia-tachycardia syndrome|Tachycardia-bradycardia
C0221047|T047|SY|74615001|SNOMEDCT_CORE|Tachycardia bradycardia syndrome|Tachycardia-bradycardia
C0221047|T047|PT|74615001|SNOMEDCT_CORE|Tachycardia-bradycardia|Tachycardia-bradycardia
C0221047|T047|FN|74615001|SNOMEDCT_CORE|Tachycardia-bradycardia|Tachycardia-bradycardia
C0221069|T047|PT|282785008|SNOMEDCT_CORE|Anterior cord syndrome|Anterior cord syndrome
C0221069|T047|FN|282785008|SNOMEDCT_CORE|Anterior cord syndrome|Anterior cord syndrome
C0221069|T047|OAP|2972007|SNOMEDCT_CORE|Anterior spinal artery occlusion syndrome|Anterior cord syndrome
C0221069|T047|SY|282785008|SNOMEDCT_CORE|Anterior spinal artery occlusion syndrome|Anterior cord syndrome
C0221069|T047|OAF|2972007|SNOMEDCT_CORE|Anterior spinal artery occlusion syndrome|Anterior cord syndrome
C0221069|T047|SY|282785008|SNOMEDCT_CORE|Anterior spinal artery syndrome|Anterior cord syndrome
C0221069|T047|OAS|2972007|SNOMEDCT_CORE|Beck's syndrome|Anterior cord syndrome
C0221069|T047|SY|282785008|SNOMEDCT_CORE|Beck's syndrome|Anterior cord syndrome
C0221069|T047|OAS|2972007|SNOMEDCT_CORE|Occlusion of anterior spinal artery|Anterior cord syndrome
C0221069|T047|IS|2972007|SNOMEDCT_CORE|Ventral medullary syndrome|Anterior cord syndrome
C0221074|T048|PT|58703003|SNOMEDCT_CORE|Postpartum depression|Postpartum depression
C0221074|T048|FN|58703003|SNOMEDCT_CORE|Postpartum depression|Postpartum depression
C0221074|T048|SY|58703003|SNOMEDCT_CORE|Puerperal depression|Postpartum depression
C0221098|T184|IS|9991008|SNOMEDCT_CORE|Acute abdominal complaint|Acute abdominal complaint
C0221150|T184|SY|30233002|SNOMEDCT_CORE|Odynophagia|Swallowing painful
C0221150|T184|SY|30233002|SNOMEDCT_CORE|Pain on swallowing|Swallowing painful
C0221150|T184|SY|30233002|SNOMEDCT_CORE|Painful swallowing|Swallowing painful
C0221150|T184|PT|30233002|SNOMEDCT_CORE|Swallowing painful|Swallowing painful
C0221150|T184|FN|30233002|SNOMEDCT_CORE|Swallowing painful|Swallowing painful
C0221155|T047|PT|56218007|SNOMEDCT_CORE|Systolic hypertension|Systolic hypertension
C0221155|T047|FN|56218007|SNOMEDCT_CORE|Systolic hypertension|Systolic hypertension
C0221184|T033|PT|61917005|SNOMEDCT_CORE|Bitemporal hemianopia|Bitemporal hemianopia
C0221184|T033|FN|61917005|SNOMEDCT_CORE|Bitemporal hemianopia|Bitemporal hemianopia
C0221184|T033|IS|61917005|SNOMEDCT_CORE|Bitemporal hemianopsia|Bitemporal hemianopia
C0221201|T184|PT|271756005|SNOMEDCT_CORE|Macular eruption|Macular eruption
C0221201|T184|FN|271756005|SNOMEDCT_CORE|Macular eruption|Macular eruption
C0221201|T184|SY|271756005|SNOMEDCT_CORE|Macular rash|Macular eruption
C0221228|T047|PT|247467008|SNOMEDCT_CORE|Comedone|Comedone
C0221228|T047|FN|247467008|SNOMEDCT_CORE|Comedone|Comedone
C0221244|T047|SY|156329007|SNOMEDCT_CORE|Seborrhea capitis|Seborrheic dermatitis of scalp
C0221244|T047|PT|156329007|SNOMEDCT_CORE|Seborrheic dermatitis of scalp|Seborrheic dermatitis of scalp
C0221244|T047|FN|156329007|SNOMEDCT_CORE|Seborrheic dermatitis of scalp|Seborrheic dermatitis of scalp
C0221244|T047|SY|156329007|SNOMEDCT_CORE|Seborrheic eczema of scalp|Seborrheic dermatitis of scalp
C0221244|T047|SYGB|156329007|SNOMEDCT_CORE|Seborrhoea capitis|Seborrheic dermatitis of scalp
C0221244|T047|OF|156329007|SNOMEDCT_CORE|Seborrhoeic dermatitis of scalp|Seborrheic dermatitis of scalp
C0221244|T047|PTGB|156329007|SNOMEDCT_CORE|Seborrhoeic dermatitis of scalp|Seborrheic dermatitis of scalp
C0221244|T047|SYGB|156329007|SNOMEDCT_CORE|Seborrhoeic eczema of scalp|Seborrheic dermatitis of scalp
C0221248|T020|PT|240042004|SNOMEDCT_CORE|Tophus|Tophus
C0221248|T020|FN|240042004|SNOMEDCT_CORE|Tophus|Tophus
C0221258|T047|OAF|76226003|SNOMEDCT_CORE|Tattoo|Tattoo
C0221258|T047|OAP|76226003|SNOMEDCT_CORE|Tattoo|Tattoo
C0221259|T047|PT|60332004|SNOMEDCT_CORE|Malposition of eyelashes|Malposition of eyelashes
C0221259|T047|SY|60332004|SNOMEDCT_CORE|Trichiasis|Malposition of eyelashes
C0221259|T047|FN|60332004|SNOMEDCT_CORE|Trichiasis|Malposition of eyelashes
C0221259|T047|IS|60332004|SNOMEDCT_CORE|Trichiasis, NOS|Malposition of eyelashes
C0221260|T047|PT|87065009|SNOMEDCT_CORE|Dystrophia unguium|Dystrophia unguium
C0221260|T047|FN|87065009|SNOMEDCT_CORE|Dystrophia unguium|Dystrophia unguium
C0221260|T047|SY|87065009|SNOMEDCT_CORE|Dystrophic nail|Dystrophia unguium
C0221260|T047|SY|87065009|SNOMEDCT_CORE|Nail dystrophy|Dystrophia unguium
C0221260|T047|SY|87065009|SNOMEDCT_CORE|Onychodystrophy|Dystrophia unguium
C0221263|T033|SY|201281002|SNOMEDCT_CORE|Café au lait spot|Café au lait spots
C0221263|T033|FN|201281002|SNOMEDCT_CORE|Café au lait spot|Café au lait spots
C0221263|T033|PT|201281002|SNOMEDCT_CORE|Café au lait spots|Café au lait spots
C0221263|T033|SY|201281002|SNOMEDCT_CORE|Cafe au lait spots|Café au lait spots
C0221263|T033|SY|201281002|SNOMEDCT_CORE|Cafe-au-lait spots|Café au lait spots
C0221263|T033|OF|201281002|SNOMEDCT_CORE|Cafe-au-lait spots|Café au lait spots
C0221265|T033|PT|165474009|SNOMEDCT_CORE|Microcytosis|Microcytosis
C0221265|T033|OF|165474009|SNOMEDCT_CORE|Microcytosis|Microcytosis
C0221265|T033|FN|165474009|SNOMEDCT_CORE|Microcytosis, red cells|Microcytosis
C0221265|T033|SY|165474009|SNOMEDCT_CORE|Microcytosis, red cells|Microcytosis
C0221276|T047|IS|44865000|SNOMEDCT_CORE|Spurious polycythaemia|Spurious polycythemia
C0221276|T047|IS|44865000|SNOMEDCT_CORE|Spurious polycythemia|Spurious polycythemia
C0221355|T019|SY|19410003|SNOMEDCT_CORE|Macrocephalus|Macrocephaly
C0221355|T019|PT|19410003|SNOMEDCT_CORE|Macrocephaly|Macrocephaly
C0221355|T019|FN|19410003|SNOMEDCT_CORE|Macrocephaly|Macrocephaly
C0221376|T047|PT|21711003|SNOMEDCT_CORE|Hydrosalpinx|Hydrosalpinx
C0221376|T047|FN|21711003|SNOMEDCT_CORE|Hydrosalpinx|Hydrosalpinx
C0221388|T047|PT|79720007|SNOMEDCT_CORE|Chronic nonalcoholic liver disease|Chronic nonalcoholic liver disease
C0221388|T047|FN|79720007|SNOMEDCT_CORE|Chronic nonalcoholic liver disease|Chronic nonalcoholic liver disease
C0221388|T047|IS|79720007|SNOMEDCT_CORE|Chronic nonalcoholic liver disease, NOS|Chronic nonalcoholic liver disease
C0221388|T047|SY|79720007|SNOMEDCT_CORE|Fatty metamorphosis of liver|Chronic nonalcoholic liver disease
C0221392|T047|PT|52441000|SNOMEDCT_CORE|Atrophic vaginitis|Atrophic vaginitis
C0221392|T047|FN|52441000|SNOMEDCT_CORE|Atrophic vaginitis|Atrophic vaginitis
C0221406|T047|SY|190502001|SNOMEDCT_CORE|Cushing basophilism|Pituitary dependent hypercortisolism
C0221406|T047|SY|190502001|SNOMEDCT_CORE|Cushing disease|Pituitary dependent hypercortisolism
C0221406|T047|SY|190502001|SNOMEDCT_CORE|Cushing's disease|Pituitary dependent hypercortisolism
C0221406|T047|SY|190502001|SNOMEDCT_CORE|Pituitary Cushing syndrome|Pituitary dependent hypercortisolism
C0221406|T047|SY|190502001|SNOMEDCT_CORE|Pituitary dependent Cushing disease|Pituitary dependent hypercortisolism
C0221406|T047|PT|190502001|SNOMEDCT_CORE|Pituitary dependent hypercortisolism|Pituitary dependent hypercortisolism
C0221406|T047|SY|190502001|SNOMEDCT_CORE|Pituitary hyperadrenal corticism|Pituitary dependent hypercortisolism
C0221406|T047|SY|190502001|SNOMEDCT_CORE|Pituitary-dependent Cushing's disease|Pituitary dependent hypercortisolism
C0221406|T047|FN|190502001|SNOMEDCT_CORE|Pituitary-dependent Cushing's disease|Pituitary dependent hypercortisolism
C0221480|T048|PT|191616006|SNOMEDCT_CORE|Recurrent depression|Recurrent depression
C0221480|T048|FN|191616006|SNOMEDCT_CORE|Recurrent depression|Recurrent depression
C0221505|T047|PT|301766008|SNOMEDCT_CORE|Lesion of brain|Lesion of brain
C0221505|T047|FN|301766008|SNOMEDCT_CORE|Lesion of brain|Lesion of brain
C0221508|T048|IS|78667006|SNOMEDCT_CORE|Nervous breakdown|Nervous breakdown
C0221520|T048|SY|191527001|SNOMEDCT_CORE|Schizophrenia simplex|Simple schizophrenia
C0221520|T048|PT|191527001|SNOMEDCT_CORE|Simple schizophrenia|Simple schizophrenia
C0221520|T048|FN|191527001|SNOMEDCT_CORE|Simple schizophrenia|Simple schizophrenia
C0221628|T033|PT|371434005|SNOMEDCT_CORE|History of alcohol abuse|History of alcohol abuse
C0221628|T033|OF|371434005|SNOMEDCT_CORE|History of alcohol abuse|History of alcohol abuse
C0221628|T033|FN|371434005|SNOMEDCT_CORE|History of alcohol abuse|History of alcohol abuse
C0221629|T033|PT|249939004|SNOMEDCT_CORE|Proximal muscle weakness|Proximal muscle weakness
C0221629|T033|FN|249939004|SNOMEDCT_CORE|Proximal muscle weakness|Proximal muscle weakness
C0221755|T184|PT|249590007|SNOMEDCT_CORE|Abdominal bruit|Abdominal bruit
C0221755|T184|FN|249590007|SNOMEDCT_CORE|Abdominal bruit|Abdominal bruit
C0221757|T047|IS|30188007|SNOMEDCT_CORE|alpha-1-Antitrypsin deficiency|Alpha-1-antitrypsin deficiency
C0221757|T047|PT|30188007|SNOMEDCT_CORE|Alpha-1-antitrypsin deficiency|Alpha-1-antitrypsin deficiency
C0221757|T047|FN|30188007|SNOMEDCT_CORE|Alpha-1-antitrypsin deficiency|Alpha-1-antitrypsin deficiency
C0221757|T047|OF|30188007|SNOMEDCT_CORE|alpha-1-Antitrypsin deficiency|Alpha-1-antitrypsin deficiency
C0221757|T047|SY|30188007|SNOMEDCT_CORE|alpha-1-Proteinase inhibitor deficiency|Alpha-1-antitrypsin deficiency
C0221759|T047|IS|3548001|SNOMEDCT_CORE|Brachial neuritis|Brachial neuritis
C0221759|T047|PT|72893007|SNOMEDCT_CORE|Brachial neuritis|Brachial neuritis
C0221759|T047|FN|72893007|SNOMEDCT_CORE|Brachial neuritis|Brachial neuritis
C0221759|T047|IS|72893007|SNOMEDCT_CORE|Brachial neuritis, NOS|Brachial neuritis
C0221776|T184|SY|102616008|SNOMEDCT_CORE|Oral cavity pain|Painful mouth
C0221776|T184|SY|102616008|SNOMEDCT_CORE|Oral pain|Painful mouth
C0221776|T184|IS|102616008|SNOMEDCT_CORE|Pain in oral cavity|Painful mouth
C0221776|T184|PT|102616008|SNOMEDCT_CORE|Painful mouth|Painful mouth
C0221776|T184|FN|102616008|SNOMEDCT_CORE|Painful mouth|Painful mouth
C0221777|T047|SY|267369002|SNOMEDCT_CORE|Non-toxic goiter|Non-toxic simple goiter
C0221777|T047|SYGB|267369002|SNOMEDCT_CORE|Non-toxic goitre|Non-toxic simple goiter
C0221777|T047|SY|267369002|SNOMEDCT_CORE|Non-toxic simple goiter|Non-toxic simple goiter
C0221777|T047|SYGB|267369002|SNOMEDCT_CORE|Non-toxic simple goitre|Non-toxic simple goiter
C0221784|T033|PT|289474006|SNOMEDCT_CORE|Lesion of vulva|Lesion of vulva
C0221784|T033|FN|289474006|SNOMEDCT_CORE|Lesion of vulva|Lesion of vulva
C0221785|T184|SY|202482009|SNOMEDCT_CORE|Arthralgia of wrist|Pain in wrist
C0221785|T184|PT|56608008|SNOMEDCT_CORE|Pain in wrist|Pain in wrist
C0221785|T184|FN|56608008|SNOMEDCT_CORE|Pain in wrist|Pain in wrist
C0221785|T184|PT|202482009|SNOMEDCT_CORE|Wrist joint pain|Pain in wrist
C0221785|T184|FN|202482009|SNOMEDCT_CORE|Wrist joint pain|Pain in wrist
C0221785|T184|SY|56608008|SNOMEDCT_CORE|Wrist pain|Pain in wrist
C0227791|T033|PT|271939006|SNOMEDCT_CORE|Vaginal discharge|Vaginal discharge
C0227791|T033|FN|271939006|SNOMEDCT_CORE|Vaginal discharge|Vaginal discharge
C0231218|T184|SY|367391008|SNOMEDCT_CORE|Does not feel right|Malaise
C0231218|T184|SY|367391008|SNOMEDCT_CORE|Feels off-color|Malaise
C0231218|T184|SYGB|367391008|SNOMEDCT_CORE|Feels off-colour|Malaise
C0231218|T184|SY|367391008|SNOMEDCT_CORE|Feels poorly|Malaise
C0231218|T184|SY|367391008|SNOMEDCT_CORE|Feels unwell|Malaise
C0231218|T184|SY|367391008|SNOMEDCT_CORE|Ill-defined experience|Malaise
C0231218|T184|PT|367391008|SNOMEDCT_CORE|Malaise|Malaise
C0231218|T184|FN|367391008|SNOMEDCT_CORE|Malaise|Malaise
C0231218|T184|SY|367391008|SNOMEDCT_CORE|Not feeling great|Malaise
C0231218|T184|SY|367391008|SNOMEDCT_CORE|Not feeling well|Malaise
C0231218|T184|SY|367391008|SNOMEDCT_CORE|Vague bodily discomfort|Malaise
C0231246|T033|PT|36440009|SNOMEDCT_CORE|Failure to gain weight|Failure to gain weight
C0231246|T033|FN|36440009|SNOMEDCT_CORE|Failure to gain weight|Failure to gain weight
C0231246|T033|SY|36440009|SNOMEDCT_CORE|Not gaining weight|Failure to gain weight
C0231246|T033|SY|36440009|SNOMEDCT_CORE|Not putting on weight|Failure to gain weight
C0231246|T033|SY|36440009|SNOMEDCT_CORE|Poor weight gain|Failure to gain weight
C0231246|T033|SY|36440009|SNOMEDCT_CORE|Unable to gain weight|Failure to gain weight
C0231274|T046|SY|69215007|SNOMEDCT_CORE|Gets overheated|Intolerant of heat
C0231274|T046|IS|69215007|SNOMEDCT_CORE|Heat intolerance|Intolerant of heat
C0231274|T046|PT|69215007|SNOMEDCT_CORE|Intolerant of heat|Intolerant of heat
C0231274|T046|FN|69215007|SNOMEDCT_CORE|Intolerant of heat|Intolerant of heat
C0231274|T046|SY|69215007|SNOMEDCT_CORE|Sensitive to heat|Intolerant of heat
C0231347|T033|PT|45704003|SNOMEDCT_CORE|At risk for noncompliance|At risk for noncompliance
C0231347|T033|FN|45704003|SNOMEDCT_CORE|At risk for noncompliance|At risk for noncompliance
C0231347|T033|IS|45704003|SNOMEDCT_CORE|Potential noncompliance|At risk for noncompliance
C0231347|T033|SY|45704003|SNOMEDCT_CORE|Potential noncompliance|At risk for noncompliance
C0231353|T033|PT|88202002|SNOMEDCT_CORE|Alteration in nutrition: less than body requirements|Alteration in nutrition: less than body requirements
C0231353|T033|FN|88202002|SNOMEDCT_CORE|Alteration in nutrition: less than body requirements|Alteration in nutrition: less than body requirements
C0231353|T033|IS|88202002|SNOMEDCT_CORE|Alteration in nutrition: less than body requirements.|Alteration in nutrition: less than body requirements
C0231353|T033|SY|88202002|SNOMEDCT_CORE|Body nutrition deficit|Alteration in nutrition: less than body requirements
C0231353|T033|SY|88202002|SNOMEDCT_CORE|Imbalanced nutrition: Less than body requirements|Alteration in nutrition: less than body requirements
C0231353|T033|IS|88202002|SNOMEDCT_CORE|Nutritional deficit|Alteration in nutrition: less than body requirements
C0231357|T033|PT|70693003|SNOMEDCT_CORE|At risk for impaired skin integrity|At risk for impaired skin integrity
C0231357|T033|FN|70693003|SNOMEDCT_CORE|At risk for impaired skin integrity|At risk for impaired skin integrity
C0231357|T033|SY|70693003|SNOMEDCT_CORE|At risk for skin ulceration|At risk for impaired skin integrity
C0231357|T033|IS|70693003|SNOMEDCT_CORE|At risk to skin ulceration|At risk for impaired skin integrity
C0231357|T033|IS|70693003|SNOMEDCT_CORE|Potential for skin breakdown|At risk for impaired skin integrity
C0231357|T033|IS|70693003|SNOMEDCT_CORE|Potential impairment of skin integrity|At risk for impaired skin integrity
C0231357|T033|SY|70693003|SNOMEDCT_CORE|Potential skin breakdown|At risk for impaired skin integrity
C0231357|T033|SY|70693003|SNOMEDCT_CORE|Skin at risk of breakdown|At risk for impaired skin integrity
C0231357|T033|SY|70693003|SNOMEDCT_CORE|Skin integrity at risk|At risk for impaired skin integrity
C0231357|T033|SY|70693003|SNOMEDCT_CORE|Skin integrity impairment risk|At risk for impaired skin integrity
C0231357|T033|SY|70693003|SNOMEDCT_CORE|Vulnerable to skin tissue breakdown|At risk for impaired skin integrity
C0231367|T033|PT|77427003|SNOMEDCT_CORE|Activity intolerance|Activity intolerance
C0231367|T033|IS|77427003|SNOMEDCT_CORE|Activity intolerance|Activity intolerance
C0231367|T033|FN|77427003|SNOMEDCT_CORE|Activity intolerance|Activity intolerance
C0231417|T033|PT|406161008|SNOMEDCT_CORE|Alteration in parenting|Alteration in parenting
C0231417|T033|FN|406161008|SNOMEDCT_CORE|Alteration in parenting|Alteration in parenting
C0231417|T033|SY|406161008|SNOMEDCT_CORE|Parenting alteration|Alteration in parenting
C0231471|T033|SY|43029002|SNOMEDCT_CORE|Abnormal body position|Abnormal posture
C0231471|T033|PT|43029002|SNOMEDCT_CORE|Abnormal posture|Abnormal posture
C0231471|T033|FN|43029002|SNOMEDCT_CORE|Abnormal posture|Abnormal posture
C0231513|T033|PT|90392009|SNOMEDCT_CORE|Nocturnal muscle spasm|Nocturnal muscle spasm
C0231513|T033|FN|90392009|SNOMEDCT_CORE|Nocturnal muscle spasm|Nocturnal muscle spasm
C0231528|T184|SY|68962001|SNOMEDCT_CORE|Aching muscles|Muscle pain
C0231528|T184|SY|68962001|SNOMEDCT_CORE|Muscle ache|Muscle pain
C0231528|T184|PT|68962001|SNOMEDCT_CORE|Muscle pain|Muscle pain
C0231528|T184|FN|68962001|SNOMEDCT_CORE|Muscle pain|Muscle pain
C0231528|T184|SY|68962001|SNOMEDCT_CORE|Myalgia|Muscle pain
C0231528|T184|SY|68962001|SNOMEDCT_CORE|Myodynia|Muscle pain
C0231528|T184|SY|68962001|SNOMEDCT_CORE|Myoneuralgia|Muscle pain
C0231528|T184|SY|68962001|SNOMEDCT_CORE|Myosalgia|Muscle pain
C0231613|T184|PT|330007|SNOMEDCT_CORE|Occipital headache|Occipital headache
C0231613|T184|FN|330007|SNOMEDCT_CORE|Occipital headache|Occipital headache
C0231655|T184|SY|20793008|SNOMEDCT_CORE|Pain in scapula|Scapulalgia
C0231655|T184|PT|20793008|SNOMEDCT_CORE|Scapulalgia|Scapulalgia
C0231655|T184|FN|20793008|SNOMEDCT_CORE|Scapulalgia|Scapulalgia
C0231655|T184|SY|20793008|SNOMEDCT_CORE|Scapulodynia|Scapulalgia
C0231655|T184|SY|20793008|SNOMEDCT_CORE|Shoulder blade pain|Scapulalgia
C0231686|T033|SY|22631008|SNOMEDCT_CORE|Disequilibrium when walking|Unsteady when walking
C0231686|T033|OAS|394616008|SNOMEDCT_CORE|Instability of gait|Unsteady when walking
C0231686|T033|SY|22631008|SNOMEDCT_CORE|Instability of gait|Unsteady when walking
C0231686|T033|SY|22631008|SNOMEDCT_CORE|Unstable when walking|Unsteady when walking
C0231686|T033|OAP|394616008|SNOMEDCT_CORE|Unsteady gait|Unsteady when walking
C0231686|T033|SY|22631008|SNOMEDCT_CORE|Unsteady gait|Unsteady when walking
C0231686|T033|OAF|394616008|SNOMEDCT_CORE|Unsteady gait|Unsteady when walking
C0231686|T033|PT|22631008|SNOMEDCT_CORE|Unsteady when walking|Unsteady when walking
C0231686|T033|FN|22631008|SNOMEDCT_CORE|Unsteady when walking|Unsteady when walking
C0231710|T184|SY|279043006|SNOMEDCT_CORE|Buttock pain|Pain in buttock
C0231710|T184|PT|279043006|SNOMEDCT_CORE|Pain in buttock|Pain in buttock
C0231710|T184|FN|279043006|SNOMEDCT_CORE|Pain in buttock|Pain in buttock
C0231710|T184|SY|279043006|SNOMEDCT_CORE|Pygalgia|Pain in buttock
C0231749|T184|SY|30989003|SNOMEDCT_CORE|Arthralgia of knee|Knee pain
C0231749|T184|SY|30989003|SNOMEDCT_CORE|Gonalgia|Knee pain
C0231749|T184|SY|30989003|SNOMEDCT_CORE|Knee joint pain|Knee pain
C0231749|T184|PT|30989003|SNOMEDCT_CORE|Knee pain|Knee pain
C0231749|T184|FN|30989003|SNOMEDCT_CORE|Knee pain|Knee pain
C0231780|T184|PT|2733002|SNOMEDCT_CORE|Heel pain|Heel pain
C0231780|T184|FN|2733002|SNOMEDCT_CORE|Heel pain|Heel pain
C0231780|T184|SY|2733002|SNOMEDCT_CORE|Talalgia|Heel pain
C0231807|T184|SY|60845006|SNOMEDCT_CORE|Breathlessness on exertion|Dyspnea on exertion
C0231807|T184|SY|60845006|SNOMEDCT_CORE|Dyspnea on effort|Dyspnea on exertion
C0231807|T184|PT|60845006|SNOMEDCT_CORE|Dyspnea on exertion|Dyspnea on exertion
C0231807|T184|FN|60845006|SNOMEDCT_CORE|Dyspnea on exertion|Dyspnea on exertion
C0231807|T184|SYGB|60845006|SNOMEDCT_CORE|Dyspnoea on effort|Dyspnea on exertion
C0231807|T184|PTGB|60845006|SNOMEDCT_CORE|Dyspnoea on exertion|Dyspnea on exertion
C0231807|T184|SY|60845006|SNOMEDCT_CORE|Exertional dyspnea|Dyspnea on exertion
C0231807|T184|SYGB|60845006|SNOMEDCT_CORE|Exertional dyspnoea|Dyspnea on exertion
C0231807|T184|SY|60845006|SNOMEDCT_CORE|Short of breath on exertion|Dyspnea on exertion
C0231807|T184|SY|60845006|SNOMEDCT_CORE|SOBOE - Shortness of breath on exertion|Dyspnea on exertion
C0231835|T033|SY|271823003|SNOMEDCT_CORE|Rapid breathing|Tachypnea
C0231835|T033|SY|271823003|SNOMEDCT_CORE|Rapid respiration|Tachypnea
C0231835|T033|PT|271823003|SNOMEDCT_CORE|Tachypnea|Tachypnea
C0231835|T033|FN|271823003|SNOMEDCT_CORE|Tachypnea|Tachypnea
C0231835|T033|SY|271823003|SNOMEDCT_CORE|Tachypneic|Tachypnea
C0231835|T033|PTGB|271823003|SNOMEDCT_CORE|Tachypnoea|Tachypnea
C0231835|T033|SYGB|271823003|SNOMEDCT_CORE|Tachypnoeic|Tachypnea
C0232058|T047|PT|13094009|SNOMEDCT_CORE|Apnea in the newborn|Apnea in the newborn
C0232058|T047|FN|13094009|SNOMEDCT_CORE|Apnea in the newborn|Apnea in the newborn
C0232058|T047|SY|13094009|SNOMEDCT_CORE|Apnea neonatorum|Apnea in the newborn
C0232058|T047|SY|13094009|SNOMEDCT_CORE|Apnea of newborn|Apnea in the newborn
C0232058|T047|PTGB|13094009|SNOMEDCT_CORE|Apnoea in the newborn|Apnea in the newborn
C0232058|T047|SYGB|13094009|SNOMEDCT_CORE|Apnoea neonatorum|Apnea in the newborn
C0232058|T047|SYGB|13094009|SNOMEDCT_CORE|Apnoea of newborn|Apnea in the newborn
C0232058|T047|SY|13094009|SNOMEDCT_CORE|Neonatal apnea|Apnea in the newborn
C0232058|T047|SYGB|13094009|SNOMEDCT_CORE|Neonatal apnoea|Apnea in the newborn
C0232071|T037|PT|58849003|SNOMEDCT_CORE|Aspiration of food|Aspiration of food
C0232071|T037|FN|58849003|SNOMEDCT_CORE|Aspiration of food|Aspiration of food
C0232071|T037|IS|58849003|SNOMEDCT_CORE|Aspiration of food material|Aspiration of food
C0232255|T033|SY|59935001|SNOMEDCT_CORE|Functional cardiac murmur|Functional heart murmur
C0232255|T033|SY|59935001|SNOMEDCT_CORE|Functional flow murmur|Functional heart murmur
C0232255|T033|PT|59935001|SNOMEDCT_CORE|Functional heart murmur|Functional heart murmur
C0232255|T033|FN|59935001|SNOMEDCT_CORE|Functional heart murmur|Functional heart murmur
C0232255|T033|SY|59935001|SNOMEDCT_CORE|Innocent heart murmur|Functional heart murmur
C0232257|T033|SY|31574009|SNOMEDCT_CORE|SM - Systolic murmur|Systolic murmur
C0232257|T033|PT|31574009|SNOMEDCT_CORE|Systolic murmur|Systolic murmur
C0232257|T033|FN|31574009|SNOMEDCT_CORE|Systolic murmur|Systolic murmur
C0232257|T033|IS|31574009|SNOMEDCT_CORE|Systolic murmur, NOS|Systolic murmur
C0232286|T184|IS|71884009|SNOMEDCT_CORE|Precordial chest pain|Precordial pain
C0232286|T184|PT|71884009|SNOMEDCT_CORE|Precordial pain|Precordial pain
C0232286|T184|FN|71884009|SNOMEDCT_CORE|Precordial pain|Precordial pain
C0232288|T184|PT|81953000|SNOMEDCT_CORE|Chest pain on exertion|Chest pain on exertion
C0232288|T184|FN|81953000|SNOMEDCT_CORE|Chest pain on exertion|Chest pain on exertion
C0232288|T184|IS|81953000|SNOMEDCT_CORE|Exertional chest pain|Chest pain on exertion
C0232292|T184|SY|23924001|SNOMEDCT_CORE|Chest tightness|Tight chest
C0232292|T184|IS|23924001|SNOMEDCT_CORE|Feeling of chest tightness|Tight chest
C0232292|T184|PT|23924001|SNOMEDCT_CORE|Tight chest|Tight chest
C0232292|T184|FN|23924001|SNOMEDCT_CORE|Tight chest|Tight chest
C0232466|T033|PT|78164000|SNOMEDCT_CORE|Feeding problem|Feeding problem
C0232466|T033|FN|78164000|SNOMEDCT_CORE|Feeding problem|Feeding problem
C0232483|T046|OAP|47268002|SNOMEDCT_CORE|Reflux|Reflux
C0232483|T046|OAF|47268002|SNOMEDCT_CORE|Reflux|Reflux
C0232483|T046|IS|47268002|SNOMEDCT_CORE|Reflux, NOS|Reflux
C0232487|T184|PT|43364001|SNOMEDCT_CORE|Abdominal discomfort|Abdominal discomfort
C0232487|T184|FN|43364001|SNOMEDCT_CORE|Abdominal discomfort|Abdominal discomfort
C0232488|T033|PT|9991008|SNOMEDCT_CORE|Abdominal colic|Abdominal colic
C0232488|T033|FN|9991008|SNOMEDCT_CORE|Abdominal colic|Abdominal colic
C0232488|T033|SY|9991008|SNOMEDCT_CORE|Colic|Abdominal colic
C0232488|T033|SY|9991008|SNOMEDCT_CORE|Colicky abdominal pain|Abdominal colic
C0232488|T033|SY|9991008|SNOMEDCT_CORE|Spasmodic abdominal pain|Abdominal colic
C0232490|T047|IS|9991008|SNOMEDCT_CORE|Abdominal crisis|Abdominal crisis
C0232491|T184|PT|111985007|SNOMEDCT_CORE|Chronic abdominal pain|Chronic abdominal pain
C0232491|T184|FN|111985007|SNOMEDCT_CORE|Chronic abdominal pain|Chronic abdominal pain
C0232492|T184|PT|83132003|SNOMEDCT_CORE|Upper abdominal pain|Upper abdominal pain
C0232492|T184|FN|83132003|SNOMEDCT_CORE|Upper abdominal pain|Upper abdominal pain
C0232493|T184|PT|79922009|SNOMEDCT_CORE|Epigastric pain|Epigastric pain
C0232493|T184|FN|79922009|SNOMEDCT_CORE|Epigastric pain|Epigastric pain
C0232495|T184|PT|54586004|SNOMEDCT_CORE|Lower abdominal pain|Lower abdominal pain
C0232495|T184|FN|54586004|SNOMEDCT_CORE|Lower abdominal pain|Lower abdominal pain
C0232502|T184|PT|35745008|SNOMEDCT_CORE|Umbilical discharge|Umbilical discharge
C0232502|T184|FN|35745008|SNOMEDCT_CORE|Umbilical discharge|Umbilical discharge
C0232519|T046|PT|47717004|SNOMEDCT_CORE|Abnormal deglutition|Abnormal deglutition
C0232519|T046|FN|47717004|SNOMEDCT_CORE|Abnormal deglutition|Abnormal deglutition
C0232519|T046|SY|47717004|SNOMEDCT_CORE|Abnormal swallowing|Abnormal deglutition
C0232598|T184|PT|63722008|SNOMEDCT_CORE|Chronic vomiting|Chronic vomiting
C0232598|T184|FN|63722008|SNOMEDCT_CORE|Chronic vomiting|Chronic vomiting
C0232698|T184|PTGB|179950008|SNOMEDCT_CORE|Abnormal defaecation|Abnormal defecation
C0232698|T184|PT|179950008|SNOMEDCT_CORE|Abnormal defecation|Abnormal defecation
C0232698|T184|FN|179950008|SNOMEDCT_CORE|Abnormal defecation|Abnormal defecation
C0232808|T047|PT|112066009|SNOMEDCT_CORE|Absent renal function|Absent renal function
C0232808|T047|OF|112066009|SNOMEDCT_CORE|Absent renal function|Absent renal function
C0232808|T047|FN|112066009|SNOMEDCT_CORE|Absent renal function|Absent renal function
C0232808|T047|IS|112066009|SNOMEDCT_CORE|NFK - Non-functioning kidney|Absent renal function
C0232808|T047|IS|112066009|SNOMEDCT_CORE|Non-functioning kidney|Absent renal function
C0232841|T046|PT|40492006|SNOMEDCT_CORE|Bladder dysfunction|Bladder dysfunction
C0232841|T046|FN|40492006|SNOMEDCT_CORE|Bladder dysfunction|Bladder dysfunction
C0232841|T046|IS|40492006|SNOMEDCT_CORE|Bladder dysfunction, NOS|Bladder dysfunction
C0232849|T184|PT|15803009|SNOMEDCT_CORE|Bladder pain|Bladder pain
C0232849|T184|FN|15803009|SNOMEDCT_CORE|Bladder pain|Bladder pain
C0232849|T184|SY|15803009|SNOMEDCT_CORE|Urinary bladder pain|Bladder pain
C0232849|T184|SY|15803009|SNOMEDCT_CORE|Vesical pain|Bladder pain
C0232854|T184|PT|84471002|SNOMEDCT_CORE|Slowing of urinary stream|Slowing of urinary stream
C0232854|T184|FN|84471002|SNOMEDCT_CORE|Slowing of urinary stream|Slowing of urinary stream
C0232861|T184|PT|2910007|SNOMEDCT_CORE|Discharge from penis|Discharge from penis
C0232861|T184|FN|2910007|SNOMEDCT_CORE|Discharge from penis|Discharge from penis
C0232861|T184|IS|2910007|SNOMEDCT_CORE|Penile discharge|Discharge from penis
C0232940|T047|IS|86030004|SNOMEDCT_CORE|Loss of menstrual period|Secondary physiologic amenorrhea
C0232940|T047|IS|86030004|SNOMEDCT_CORE|Secondary amenorrhea|Secondary physiologic amenorrhea
C0232940|T047|IS|86030004|SNOMEDCT_CORE|Secondary amenorrhoea|Secondary physiologic amenorrhea
C0232940|T047|PT|86030004|SNOMEDCT_CORE|Secondary physiologic amenorrhea|Secondary physiologic amenorrhea
C0232940|T047|FN|86030004|SNOMEDCT_CORE|Secondary physiologic amenorrhea|Secondary physiologic amenorrhea
C0232940|T047|PTGB|86030004|SNOMEDCT_CORE|Secondary physiologic amenorrhoea|Secondary physiologic amenorrhea
C0232943|T184|PT|314631008|SNOMEDCT_CORE|Menometrorrhagia|Menometrorrhagia
C0232943|T184|FN|314631008|SNOMEDCT_CORE|Menometrorrhagia|Menometrorrhagia
C0232943|T184|SY|314631008|SNOMEDCT_CORE|Metromenorrhagia|Menometrorrhagia
C0232968|T184|PT|68811000|SNOMEDCT_CORE|Menopausal problem|Menopausal problem
C0232968|T184|FN|68811000|SNOMEDCT_CORE|Menopausal problem|Menopausal problem
C0232968|T184|IS|68811000|SNOMEDCT_CORE|Menopausal problem, NOS|Menopausal problem
C0232970|T033|SY|76498008|SNOMEDCT_CORE|Postmenopausal|Postmenopausal state
C0232970|T033|PT|76498008|SNOMEDCT_CORE|Postmenopausal state|Postmenopausal state
C0232970|T033|FN|76498008|SNOMEDCT_CORE|Postmenopausal state|Postmenopausal state
C0232989|T033|PT|72892002|SNOMEDCT_CORE|Normal pregnancy|Normal pregnancy
C0232989|T033|FN|72892002|SNOMEDCT_CORE|Normal pregnancy|Normal pregnancy
C0233105|T046|OAP|69124005|SNOMEDCT_CORE|Complete abortion|Complete abortion
C0233105|T046|OAF|69124005|SNOMEDCT_CORE|Complete abortion|Complete abortion
C0233214|T033|PT|28701003|SNOMEDCT_CORE|Low maternal weight gain|Low maternal weight gain
C0233214|T033|FN|28701003|SNOMEDCT_CORE|Low maternal weight gain|Low maternal weight gain
C0233308|T033|PT|169734005|SNOMEDCT_CORE|Spontaneous rupture of fetal membranes|Spontaneous rupture of fetal membranes
C0233308|T033|SYGB|169734005|SNOMEDCT_CORE|Spontaneous rupture of foetal membranes|Spontaneous rupture of fetal membranes
C0233308|T033|SY|169734005|SNOMEDCT_CORE|Spontaneous rupture of membranes|Spontaneous rupture of fetal membranes
C0233308|T033|FN|169734005|SNOMEDCT_CORE|Spontaneous rupture of membranes|Spontaneous rupture of fetal membranes
C0233308|T033|SY|169734005|SNOMEDCT_CORE|SRM - Spontaneous rupture of membranes|Spontaneous rupture of fetal membranes
C0233308|T033|SY|169734005|SNOMEDCT_CORE|SROM - Spontaneous rupture of membranes|Spontaneous rupture of fetal membranes
C0233315|T033|PT|367494004|SNOMEDCT_CORE|Premature birth of newborn|Premature birth of newborn
C0233315|T033|FN|367494004|SNOMEDCT_CORE|Premature birth of newborn|Premature birth of newborn
C0233403|T048|SY|81302005|SNOMEDCT_CORE|Physically well but worried|Worried well
C0233403|T048|SY|81302005|SNOMEDCT_CORE|Psyche disturbed with normal general body function|Worried well
C0233403|T048|PT|81302005|SNOMEDCT_CORE|Worried well|Worried well
C0233403|T048|FN|81302005|SNOMEDCT_CORE|Worried well|Worried well
C0233439|T048|PT|386822001|SNOMEDCT_CORE|Adjustment reaction of adolescence|Adjustment reaction of adolescence
C0233439|T048|FN|386822001|SNOMEDCT_CORE|Adjustment reaction of adolescence|Adjustment reaction of adolescence
C0233439|T048|SY|386822001|SNOMEDCT_CORE|Adolescent situation reaction|Adjustment reaction of adolescence
C0233439|T048|SY|386822001|SNOMEDCT_CORE|Adolescent turmoil|Adjustment reaction of adolescence
C0233514|T048|SY|277843001|SNOMEDCT_CORE|Behavioral concern|Problem behavior
C0233514|T048|SY|277843001|SNOMEDCT_CORE|Behavioral problem|Problem behavior
C0233514|T048|SYGB|277843001|SNOMEDCT_CORE|Behavioural concern|Problem behavior
C0233514|T048|SYGB|277843001|SNOMEDCT_CORE|Behavioural problem|Problem behavior
C0233514|T048|PT|277843001|SNOMEDCT_CORE|Problem behavior|Problem behavior
C0233514|T048|FN|277843001|SNOMEDCT_CORE|Problem behavior|Problem behavior
C0233514|T048|PTGB|277843001|SNOMEDCT_CORE|Problem behaviour|Problem behavior
C0233530|T048|PTGB|82096005|SNOMEDCT_CORE|Aggressive type unsocialised behaviour disorder|Aggressive type unsocialized behavior disorder
C0233530|T048|IS|82096005|SNOMEDCT_CORE|Aggressive type unsocialised conduct disorder|Aggressive type unsocialized behavior disorder
C0233530|T048|PT|82096005|SNOMEDCT_CORE|Aggressive type unsocialized behavior disorder|Aggressive type unsocialized behavior disorder
C0233530|T048|FN|82096005|SNOMEDCT_CORE|Aggressive type unsocialized behavior disorder|Aggressive type unsocialized behavior disorder
C0233530|T048|OF|82096005|SNOMEDCT_CORE|Aggressive type unsocialized behavior disorder|Aggressive type unsocialized behavior disorder
C0233530|T048|IS|82096005|SNOMEDCT_CORE|Aggressive type unsocialized conduct disorder|Aggressive type unsocialized behavior disorder
C0233715|T033|PT|29164008|SNOMEDCT_CORE|Disturbance in speech|Disturbance in speech
C0233715|T033|FN|29164008|SNOMEDCT_CORE|Disturbance in speech|Disturbance in speech
C0233715|T033|IS|29164008|SNOMEDCT_CORE|Disturbance in speech, NOS|Disturbance in speech
C0233715|T033|SY|29164008|SNOMEDCT_CORE|Speech abnormality|Disturbance in speech
C0233715|T033|IS|29164008|SNOMEDCT_CORE|Speech abnormality, NOS|Disturbance in speech
C0233715|T033|SY|29164008|SNOMEDCT_CORE|Speech impairment|Disturbance in speech
C0233794|T048|SY|386807006|SNOMEDCT_CORE|Bad memory|Memory impairment
C0233794|T048|SY|386807006|SNOMEDCT_CORE|Disturbance of memory|Memory impairment
C0233794|T048|SY|386807006|SNOMEDCT_CORE|Impaired memory|Memory impairment
C0233794|T048|SY|386807006|SNOMEDCT_CORE|Memory deficit|Memory impairment
C0233794|T048|PT|386807006|SNOMEDCT_CORE|Memory impairment|Memory impairment
C0233794|T048|FN|386807006|SNOMEDCT_CORE|Memory impairment|Memory impairment
C0233794|T048|SY|386807006|SNOMEDCT_CORE|Memory problem|Memory impairment
C0233794|T048|SY|386807006|SNOMEDCT_CORE|Poor memory|Memory impairment
C0234016|T048|PT|73491007|SNOMEDCT_CORE|Psychogenic impotence|Psychogenic impotence
C0234016|T048|OF|73491007|SNOMEDCT_CORE|Psychogenic impotence|Psychogenic impotence
C0234016|T048|FN|73491007|SNOMEDCT_CORE|Psychogenic impotence|Psychogenic impotence
C0234233|T184|SY|247348008|SNOMEDCT_CORE|Sore to touch|Tenderness
C0234233|T184|SY|247348008|SNOMEDCT_CORE|Tender pain|Tenderness
C0234233|T184|PT|247348008|SNOMEDCT_CORE|Tenderness|Tenderness
C0234233|T184|FN|247348008|SNOMEDCT_CORE|Tenderness|Tenderness
C0234369|T184|SY|26079004|SNOMEDCT_CORE|Involuntary trembling|Trembling
C0234369|T184|SY|26079004|SNOMEDCT_CORE|Trembling|Trembling
C0234376|T184|SY|30721006|SNOMEDCT_CORE|Action tremor|Action tremor
C0234379|T184|IS|25082004|SNOMEDCT_CORE|Rest tremor|Resting tremor
C0234379|T184|PT|25082004|SNOMEDCT_CORE|Resting tremor|Resting tremor
C0234379|T184|FN|25082004|SNOMEDCT_CORE|Resting tremor|Resting tremor
C0234632|T033|PT|13164000|SNOMEDCT_CORE|Reduced visual acuity|Reduced visual acuity
C0234632|T033|FN|13164000|SNOMEDCT_CORE|Reduced visual acuity|Reduced visual acuity
C0234655|T184|PT|2070002|SNOMEDCT_CORE|Burning sensation in eye|Burning sensation in eye
C0234655|T184|FN|2070002|SNOMEDCT_CORE|Burning sensation in eye|Burning sensation in eye
C0234665|T033|PT|43854003|SNOMEDCT_CORE|Retraction of eyelid|Retraction of eyelid
C0234665|T033|FN|43854003|SNOMEDCT_CORE|Retraction of eyelid|Retraction of eyelid
C0234665|T033|IS|43854003|SNOMEDCT_CORE|Retraction of eyelid, NOS|Retraction of eyelid
C0234927|T046|SY|86708008|SNOMEDCT_CORE|Hypersteatosis|Sebaceous gland overactivity
C0234927|T046|SY|86708008|SNOMEDCT_CORE|Sebaceous gland overactivity|Sebaceous gland overactivity
C0234935|T047|PT|402408009|SNOMEDCT_CORE|Acute urticaria|Acute urticaria
C0234935|T047|FN|402408009|SNOMEDCT_CORE|Acute urticaria|Acute urticaria
C0234974|T047|PT|79348005|SNOMEDCT_CORE|Simple partial seizure, consciousness not impaired|Simple partial seizure, consciousness not impaired
C0234974|T047|OF|79348005|SNOMEDCT_CORE|Simple partial seizure, consciousness not impaired|Simple partial seizure, consciousness not impaired
C0234974|T047|FN|79348005|SNOMEDCT_CORE|Simple partial seizure, consciousness not impaired|Simple partial seizure, consciousness not impaired
C0234974|T047|IS|79348005|SNOMEDCT_CORE|Simple partial seizures with consciousness preserved|Simple partial seizure, consciousness not impaired
C0235025|T047|SY|95663000|SNOMEDCT_CORE|Motor neuritis|Peripheral motor neuropathy
C0235025|T047|IS|95663000|SNOMEDCT_CORE|Motor neuropathy|Peripheral motor neuropathy
C0235025|T047|SY|95663000|SNOMEDCT_CORE|Motor peripheral neuropathy|Peripheral motor neuropathy
C0235025|T047|PT|95663000|SNOMEDCT_CORE|Peripheral motor neuropathy|Peripheral motor neuropathy
C0235025|T047|FN|95663000|SNOMEDCT_CORE|Peripheral motor neuropathy|Peripheral motor neuropathy
C0235136|T048|PT|83458005|SNOMEDCT_CORE|Agitated depression|Agitated depression
C0235136|T048|FN|83458005|SNOMEDCT_CORE|Agitated depression|Agitated depression
C0235162|T184|PT|301345002|SNOMEDCT_CORE|Difficulty sleeping|Difficulty sleeping
C0235162|T184|FN|301345002|SNOMEDCT_CORE|Difficulty sleeping|Difficulty sleeping
C0235162|T184|SY|301345002|SNOMEDCT_CORE|Poor sleep|Difficulty sleeping
C0235198|T033|SY|60032008|SNOMEDCT_CORE|Concentration impairment|Unable to concentrate
C0235198|T033|IS|60032008|SNOMEDCT_CORE|Lack of concentration|Unable to concentrate
C0235198|T033|PT|60032008|SNOMEDCT_CORE|Unable to concentrate|Unable to concentrate
C0235198|T033|FN|60032008|SNOMEDCT_CORE|Unable to concentrate|Unable to concentrate
C0235222|T047|PT|48146000|SNOMEDCT_CORE|Diastolic hypertension|Diastolic hypertension
C0235222|T047|FN|48146000|SNOMEDCT_CORE|Diastolic hypertension|Diastolic hypertension
C0235222|T047|IS|48146000|SNOMEDCT_CORE|Diastolic hypertension, NOS|Diastolic hypertension
C0235259|T020|PT|95723009|SNOMEDCT_CORE|Subcapsular cataract|Subcapsular cataract
C0235259|T020|FN|95723009|SNOMEDCT_CORE|Subcapsular cataract|Subcapsular cataract
C0235259|T020|IS|95723009|SNOMEDCT_CORE|Subcapsular cataract, NOS|Subcapsular cataract
C0235267|T184|PT|75705005|SNOMEDCT_CORE|Red eye|Red eye
C0235267|T184|FN|75705005|SNOMEDCT_CORE|Red eye|Red eye
C0235267|T184|IS|75705005|SNOMEDCT_CORE|Redness of eye|Red eye
C0235299|T184|PT|301717006|SNOMEDCT_CORE|Right upper quadrant pain|Right upper quadrant pain
C0235299|T184|FN|301717006|SNOMEDCT_CORE|Right upper quadrant pain|Right upper quadrant pain
C0235325|T046|SY|61401005|SNOMEDCT_CORE|Gastric bleeding|Gastric hemorrhage
C0235325|T046|IS|61401005|SNOMEDCT_CORE|Gastric bleeding, NOS|Gastric hemorrhage
C0235325|T046|PTGB|61401005|SNOMEDCT_CORE|Gastric haemorrhage|Gastric hemorrhage
C0235325|T046|PT|61401005|SNOMEDCT_CORE|Gastric hemorrhage|Gastric hemorrhage
C0235325|T046|FN|61401005|SNOMEDCT_CORE|Gastric hemorrhage|Gastric hemorrhage
C0235325|T046|IS|61401005|SNOMEDCT_CORE|Gastric hemorrhage, NOS|Gastric hemorrhage
C0235325|T046|SY|61401005|SNOMEDCT_CORE|Gastrorrhagia|Gastric hemorrhage
C0235326|T047|PTGB|75955007|SNOMEDCT_CORE|Thrombosed haemorrhoids|Thrombosed hemorrhoids
C0235326|T047|PT|75955007|SNOMEDCT_CORE|Thrombosed hemorrhoids|Thrombosed hemorrhoids
C0235326|T047|FN|75955007|SNOMEDCT_CORE|Thrombosed hemorrhoids|Thrombosed hemorrhoids
C0235326|T047|IS|75955007|SNOMEDCT_CORE|Thrombosed hemorrhoids, NOS|Thrombosed hemorrhoids
C0235327|T047|PT|235849009|SNOMEDCT_CORE|Small intestinal gangrene|Small intestinal gangrene
C0235327|T047|FN|235849009|SNOMEDCT_CORE|Small intestinal gangrene|Small intestinal gangrene
C0235328|T047|PT|40650009|SNOMEDCT_CORE|Obstruction of colon|Obstruction of colon
C0235328|T047|FN|40650009|SNOMEDCT_CORE|Obstruction of colon|Obstruction of colon
C0235328|T047|IS|40650009|SNOMEDCT_CORE|Occlusion of colon|Obstruction of colon
C0235329|T047|SY|281255004|SNOMEDCT_CORE|SBO - Small bowel obstruction|Small bowel obstruction
C0235329|T047|PT|281255004|SNOMEDCT_CORE|Small bowel obstruction|Small bowel obstruction
C0235329|T047|FN|281255004|SNOMEDCT_CORE|Small bowel obstruction|Small bowel obstruction
C0235351|T047|SY|66123000|SNOMEDCT_CORE|Tongue ulceration|Ulcer on tongue
C0235351|T047|IS|66123000|SNOMEDCT_CORE|Tongue ulceration, NOS|Ulcer on tongue
C0235351|T047|IS|66123000|SNOMEDCT_CORE|Ulcer of tongue|Ulcer on tongue
C0235351|T047|IS|66123000|SNOMEDCT_CORE|Ulcer of tongue, NOS|Ulcer on tongue
C0235351|T047|PT|66123000|SNOMEDCT_CORE|Ulcer on tongue|Ulcer on tongue
C0235351|T047|FN|66123000|SNOMEDCT_CORE|Ulcer on tongue|Ulcer on tongue
C0235439|T046|FN|26237000|SNOMEDCT_CORE|Ankle edema|Ankle edema
C0235439|T046|PT|26237000|SNOMEDCT_CORE|Ankle edema|Ankle edema
C0235439|T046|PTGB|26237000|SNOMEDCT_CORE|Ankle oedema|Ankle edema
C0235439|T046|SY|26237000|SNOMEDCT_CORE|Swollen ankle - edema|Ankle edema
C0235439|T046|SYGB|26237000|SNOMEDCT_CORE|Swollen ankle - oedema|Ankle edema
C0235470|T033|SY|23687008|SNOMEDCT_CORE|Angina pectoris with documented spasm|Angina pectoris with documented spasm
C0235480|T047|SY|282825002|SNOMEDCT_CORE|AF - Paroxysmal atrial fibrillation|Paroxysmal atrial fibrillation
C0235480|T047|SY|282825002|SNOMEDCT_CORE|Intermittent atrial fibrillation|Paroxysmal atrial fibrillation
C0235480|T047|SY|282825002|SNOMEDCT_CORE|PAF - Paroxysmal atrial fibrillation|Paroxysmal atrial fibrillation
C0235480|T047|PT|282825002|SNOMEDCT_CORE|Paroxysmal atrial fibrillation|Paroxysmal atrial fibrillation
C0235480|T047|FN|282825002|SNOMEDCT_CORE|Paroxysmal atrial fibrillation|Paroxysmal atrial fibrillation
C0235501|T047|SY|95451004|SNOMEDCT_CORE|Superficial thrombophlebitis of arm|Thrombophlebitis of superficial veins of upper extremities
C0235501|T047|PT|95451004|SNOMEDCT_CORE|Thrombophlebitis of superficial veins of upper extremities|Thrombophlebitis of superficial veins of upper extremities
C0235501|T047|FN|95451004|SNOMEDCT_CORE|Thrombophlebitis of superficial veins of upper extremities|Thrombophlebitis of superficial veins of upper extremities
C0235511|T046|PT|275517008|SNOMEDCT_CORE|Superficial vein thrombosis|Superficial vein thrombosis
C0235511|T046|FN|275517008|SNOMEDCT_CORE|Superficial vein thrombosis|Superficial vein thrombosis
C0235527|T047|OAP|128404006|SNOMEDCT_CORE|Right heart failure|Right heart failure
C0235527|T047|OAF|128404006|SNOMEDCT_CORE|Right heart failure|Right heart failure
C0235592|T047|PT|127086001|SNOMEDCT_CORE|Cervical lymphadenopathy|Cervical lymphadenopathy
C0235592|T047|FN|127086001|SNOMEDCT_CORE|Cervical lymphadenopathy|Cervical lymphadenopathy
C0235632|T184|PT|271857006|SNOMEDCT_CORE|Loin pain|Loin pain
C0235632|T184|FN|271857006|SNOMEDCT_CORE|Loin pain|Loin pain
C0235639|T033|PT|102866000|SNOMEDCT_CORE|Abnormal urine|Abnormal urine
C0235639|T033|FN|102866000|SNOMEDCT_CORE|Abnormal urine|Abnormal urine
C0235639|T033|IS|102866000|SNOMEDCT_CORE|Abnormal urine, NOS|Abnormal urine
C0235653|T191|SY|372064008|SNOMEDCT_CORE|Cancer of female breast|Malignant neoplasm of female breast
C0235653|T191|SY|372064008|SNOMEDCT_CORE|Female breast cancer|Malignant neoplasm of female breast
C0235653|T191|PT|372064008|SNOMEDCT_CORE|Malignant neoplasm of female breast|Malignant neoplasm of female breast
C0235653|T191|FN|372064008|SNOMEDCT_CORE|Malignant neoplasm of female breast|Malignant neoplasm of female breast
C0235656|T046|PT|289794001|SNOMEDCT_CORE|Lesion of cervix|Lesion of cervix
C0235656|T046|FN|289794001|SNOMEDCT_CORE|Lesion of cervix|Lesion of cervix
C0235659|T033|SY|276369006|SNOMEDCT_CORE|Baby kicking less|Reduced fetal movement
C0235659|T033|SY|276369006|SNOMEDCT_CORE|Baby moving less|Reduced fetal movement
C0235659|T033|SY|276369006|SNOMEDCT_CORE|Low fetal movement|Reduced fetal movement
C0235659|T033|SYGB|276369006|SNOMEDCT_CORE|Low foetal movement|Reduced fetal movement
C0235659|T033|PT|276369006|SNOMEDCT_CORE|Reduced fetal movement|Reduced fetal movement
C0235659|T033|FN|276369006|SNOMEDCT_CORE|Reduced fetal movement|Reduced fetal movement
C0235659|T033|PTGB|276369006|SNOMEDCT_CORE|Reduced foetal movement|Reduced fetal movement
C0235660|T047|IS|78622004|SNOMEDCT_CORE|Galactorrhea|Galactorrhea not associated with childbirth
C0235660|T047|PT|78622004|SNOMEDCT_CORE|Galactorrhea not associated with childbirth|Galactorrhea not associated with childbirth
C0235660|T047|FN|78622004|SNOMEDCT_CORE|Galactorrhea not associated with childbirth|Galactorrhea not associated with childbirth
C0235660|T047|IS|78622004|SNOMEDCT_CORE|Galactorrhea, NOS|Galactorrhea not associated with childbirth
C0235660|T047|IS|78622004|SNOMEDCT_CORE|Galactorrhoea|Galactorrhea not associated with childbirth
C0235660|T047|PTGB|78622004|SNOMEDCT_CORE|Galactorrhoea not associated with childbirth|Galactorrhea not associated with childbirth
C0235660|T047|SY|78622004|SNOMEDCT_CORE|Inappropriate lactation|Galactorrhea not associated with childbirth
C0235660|T047|SY|78622004|SNOMEDCT_CORE|Inappropriate production of milk|Galactorrhea not associated with childbirth
C0235660|T047|SY|78622004|SNOMEDCT_CORE|Milk from non-pregnant breast|Galactorrhea not associated with childbirth
C0235710|T184|PT|279084009|SNOMEDCT_CORE|Chest discomfort|Chest discomfort
C0235710|T184|FN|279084009|SNOMEDCT_CORE|Chest discomfort|Chest discomfort
C0235752|T019|SYGB|416377005|SNOMEDCT_CORE|Naevus flammeus|Port-wine stain of skin
C0235752|T019|SY|416377005|SNOMEDCT_CORE|Nevus flammeus|Port-wine stain of skin
C0235752|T019|SY|416377005|SNOMEDCT_CORE|Port wine stain of skin|Port-wine stain of skin
C0235752|T019|SY|416377005|SNOMEDCT_CORE|Port-wine birthmark|Port-wine stain of skin
C0235752|T019|SYGB|416377005|SNOMEDCT_CORE|Port-wine naevus|Port-wine stain of skin
C0235752|T019|SY|416377005|SNOMEDCT_CORE|Port-wine nevus|Port-wine stain of skin
C0235752|T019|SY|416377005|SNOMEDCT_CORE|Port-wine stain|Port-wine stain of skin
C0235752|T019|PT|416377005|SNOMEDCT_CORE|Port-wine stain of skin|Port-wine stain of skin
C0235752|T019|FN|416377005|SNOMEDCT_CORE|Port-wine stain of skin|Port-wine stain of skin
C0235752|T019|SYGB|416377005|SNOMEDCT_CORE|Portwine naevus|Port-wine stain of skin
C0235752|T019|SY|416377005|SNOMEDCT_CORE|Portwine nevus|Port-wine stain of skin
C0235752|T019|SY|416377005|SNOMEDCT_CORE|PWS - Port-wine stain|Port-wine stain of skin
C0235761|T190|SY|80142000|SNOMEDCT_CORE|Nasal septal perforation|Perforation of nasal septum
C0235761|T190|SY|80142000|SNOMEDCT_CORE|Perforated nasal septum|Perforation of nasal septum
C0235761|T190|PT|80142000|SNOMEDCT_CORE|Perforation of nasal septum|Perforation of nasal septum
C0235761|T190|FN|80142000|SNOMEDCT_CORE|Perforation of nasal septum|Perforation of nasal septum
C0235777|T184|PT|95617006|SNOMEDCT_CORE|Neonatal cyanosis|Neonatal cyanosis
C0235777|T184|FN|95617006|SNOMEDCT_CORE|Neonatal cyanosis|Neonatal cyanosis
C0235777|T184|IS|95617006|SNOMEDCT_CORE|Neonatal cyanosis, NOS|Neonatal cyanosis
C0235782|T191|PT|372140005|SNOMEDCT_CORE|Carcinoma of gallbladder|Carcinoma of gallbladder
C0235782|T191|FN|372140005|SNOMEDCT_CORE|Carcinoma of gallbladder|Carcinoma of gallbladder
C0235808|T184|SY|430968008|SNOMEDCT_CORE|Male perineal pain|Pain in male perineum
C0235808|T184|PT|430968008|SNOMEDCT_CORE|Pain in male perineum|Pain in male perineum
C0235808|T184|FN|430968008|SNOMEDCT_CORE|Pain in male perineum|Pain in male perineum
C0235880|T047|PT|32595002|SNOMEDCT_CORE|Mononeuritis|Mononeuritis
C0235880|T047|FN|32595002|SNOMEDCT_CORE|Mononeuritis|Mononeuritis
C0235880|T047|IS|32595002|SNOMEDCT_CORE|Mononeuritis, NOS|Mononeuritis
C0235886|T046|OAP|102574007|SNOMEDCT_CORE|Edema of leg|Leg edema
C0235886|T046|OAF|102574007|SNOMEDCT_CORE|Edema of leg|Leg edema
C0235886|T046|OAS|102574007|SNOMEDCT_CORE|Leg edema|Leg edema
C0235886|T046|OAS|102574007|SNOMEDCT_CORE|Leg oedema|Leg edema
C0235886|T046|OAP|102574007|SNOMEDCT_CORE|Oedema of leg|Leg edema
C0235895|T046|PT|19220005|SNOMEDCT_CORE|Complication of implant|Complication of implant
C0235895|T046|FN|19220005|SNOMEDCT_CORE|Complication of implant|Complication of implant
C0235922|T191|PT|92102001|SNOMEDCT_CORE|Benign neoplasm of female breast|Benign neoplasm of female breast
C0235922|T191|FN|92102001|SNOMEDCT_CORE|Benign neoplasm of female breast|Benign neoplasm of female breast
C0235922|T191|IS|92102001|SNOMEDCT_CORE|Benign neoplasm of female breast, NOS|Benign neoplasm of female breast
C0235972|T020|PT|95689000|SNOMEDCT_CORE|Retinal deposits|Retinal deposits
C0235972|T020|FN|95689000|SNOMEDCT_CORE|Retinal deposits|Retinal deposits
C0235974|T191|PT|372142002|SNOMEDCT_CORE|Carcinoma of pancreas|Carcinoma of pancreas
C0235974|T191|FN|372142002|SNOMEDCT_CORE|Carcinoma of pancreas|Carcinoma of pancreas
C0235982|T047|PT|43797002|SNOMEDCT_CORE|Stricture of bile duct|Stricture of bile duct
C0235982|T047|FN|43797002|SNOMEDCT_CORE|Stricture of bile duct|Stricture of bile duct
C0236000|T184|PT|274667000|SNOMEDCT_CORE|Jaw pain|Jaw pain
C0236000|T184|FN|274667000|SNOMEDCT_CORE|Jaw pain|Jaw pain
C0236000|T184|SY|274667000|SNOMEDCT_CORE|Pain of jaw|Jaw pain
C0236038|T047|PT|95827002|SNOMEDCT_CORE|Congenital hearing disorder|Congenital hearing disorder
C0236038|T047|FN|95827002|SNOMEDCT_CORE|Congenital hearing disorder|Congenital hearing disorder
C0236038|T047|IS|95827002|SNOMEDCT_CORE|Congenital hearing disorder, NOS|Congenital hearing disorder
C0236040|T184|SY|300954003|SNOMEDCT_CORE|Calf pain|Pain in calf
C0236040|T184|PT|300954003|SNOMEDCT_CORE|Pain in calf|Pain in calf
C0236040|T184|FN|300954003|SNOMEDCT_CORE|Pain in calf|Pain in calf
C0236048|T047|PT|78809005|SNOMEDCT_CORE|Gastric polyp|Gastric polyp
C0236048|T047|FN|78809005|SNOMEDCT_CORE|Gastric polyp|Gastric polyp
C0236048|T047|IS|78809005|SNOMEDCT_CORE|Gastric polyp, NOS|Gastric polyp
C0236048|T047|SY|78809005|SNOMEDCT_CORE|Polyp of stomach|Gastric polyp
C0236075|T184|PT|21801002|SNOMEDCT_CORE|Menopausal symptom|Menopausal symptom
C0236075|T184|FN|21801002|SNOMEDCT_CORE|Menopausal symptom|Menopausal symptom
C0236075|T184|IS|21801002|SNOMEDCT_CORE|Menopausal symptom, NOS|Menopausal symptom
C0236078|T184|PT|20502007|SNOMEDCT_CORE|Pain in scrotum|Pain in scrotum
C0236078|T184|FN|20502007|SNOMEDCT_CORE|Pain in scrotum|Pain in scrotum
C0236078|T184|SY|20502007|SNOMEDCT_CORE|Pain of scrotum|Pain in scrotum
C0236078|T184|SY|20502007|SNOMEDCT_CORE|Scrotal pain|Pain in scrotum
C0236082|T184|SY|38343000|SNOMEDCT_CORE|Pain in vagina|Vaginal pain
C0236082|T184|PT|38343000|SNOMEDCT_CORE|Vaginal pain|Vaginal pain
C0236082|T184|FN|38343000|SNOMEDCT_CORE|Vaginal pain|Vaginal pain
C0236127|T047|SY|57748001|SNOMEDCT_CORE|Bleeding esophageal ulcer|Bleeding ulcer of esophagus
C0236127|T047|SYGB|57748001|SNOMEDCT_CORE|Bleeding oesophageal ulcer|Bleeding ulcer of esophagus
C0236127|T047|PT|57748001|SNOMEDCT_CORE|Bleeding ulcer of esophagus|Bleeding ulcer of esophagus
C0236127|T047|FN|57748001|SNOMEDCT_CORE|Bleeding ulcer of esophagus|Bleeding ulcer of esophagus
C0236127|T047|PTGB|57748001|SNOMEDCT_CORE|Bleeding ulcer of oesophagus|Bleeding ulcer of esophagus
C0236127|T047|SYGB|57748001|SNOMEDCT_CORE|Haemorrhagic ulcer of oesophagus|Bleeding ulcer of esophagus
C0236127|T047|SY|57748001|SNOMEDCT_CORE|Hemorrhagic ulcer of esophagus|Bleeding ulcer of esophagus
C0236151|T033|SY|167180005|SNOMEDCT_CORE|Abnormal results of kidney function studies|Renal function tests abnormal
C0236151|T033|PT|167180005|SNOMEDCT_CORE|Renal function tests abnormal|Renal function tests abnormal
C0236151|T033|FN|167180005|SNOMEDCT_CORE|Renal function tests abnormal|Renal function tests abnormal
C0236640|T048|SY|66108005|SNOMEDCT_CORE|Dementia of the Alzheimer's type, with late onset, uncomplicated|Primary degenerative dementia of the Alzheimer type, senile onset, uncomplicated
C0236640|T048|PT|66108005|SNOMEDCT_CORE|Primary degenerative dementia of the Alzheimer type, senile onset, uncomplicated|Primary degenerative dementia of the Alzheimer type, senile onset, uncomplicated
C0236640|T048|FN|66108005|SNOMEDCT_CORE|Primary degenerative dementia of the Alzheimer type, senile onset, uncomplicated|Primary degenerative dementia of the Alzheimer type, senile onset, uncomplicated
C0236650|T048|SY|70936005|SNOMEDCT_CORE|Multi infarct dementia, uncomplicated|Multi-infarct dementia, uncomplicated
C0236650|T048|PT|70936005|SNOMEDCT_CORE|Multi-infarct dementia, uncomplicated|Multi-infarct dementia, uncomplicated
C0236650|T048|FN|70936005|SNOMEDCT_CORE|Multi-infarct dementia, uncomplicated|Multi-infarct dementia, uncomplicated
C0236650|T048|SY|70936005|SNOMEDCT_CORE|Vascular dementia, uncomplicated|Multi-infarct dementia, uncomplicated
C0236653|T048|PT|14070001|SNOMEDCT_CORE|Multi-infarct dementia with depression|Multi-infarct dementia with depression
C0236653|T048|FN|14070001|SNOMEDCT_CORE|Multi-infarct dementia with depression|Multi-infarct dementia with depression
C0236653|T048|SY|14070001|SNOMEDCT_CORE|Vascular dementia, with depressive mood|Multi-infarct dementia with depression
C0236654|T048|PT|18653004|SNOMEDCT_CORE|Alcohol intoxication delirium|Alcohol intoxication delirium
C0236654|T048|FN|18653004|SNOMEDCT_CORE|Alcohol intoxication delirium|Alcohol intoxication delirium
C0236656|T048|SY|281004|SNOMEDCT_CORE|Alcohol-induced persisting dementia|Dementia associated with alcoholism
C0236656|T048|SY|281004|SNOMEDCT_CORE|Alcoholic dementia|Dementia associated with alcoholism
C0236656|T048|PT|281004|SNOMEDCT_CORE|Dementia associated with alcoholism|Dementia associated with alcoholism
C0236656|T048|FN|281004|SNOMEDCT_CORE|Dementia associated with alcoholism|Dementia associated with alcoholism
C0236660|T048|SY|53936005|SNOMEDCT_CORE|Alcohol induced mood disorder|Alcohol-induced mood disorder
C0236660|T048|PT|53936005|SNOMEDCT_CORE|Alcohol-induced mood disorder|Alcohol-induced mood disorder
C0236660|T048|FN|53936005|SNOMEDCT_CORE|Alcohol-induced mood disorder|Alcohol-induced mood disorder
C0236663|T047|PT|191480000|SNOMEDCT_CORE|Alcohol withdrawal syndrome|Alcohol withdrawal syndrome
C0236663|T047|FN|191480000|SNOMEDCT_CORE|Alcohol withdrawal syndrome|Alcohol withdrawal syndrome
C0236734|T048|PT|308374001|SNOMEDCT_CORE|Caffeine-related disorder|Caffeine-related disorder
C0236734|T048|FN|308374001|SNOMEDCT_CORE|Caffeine-related disorder|Caffeine-related disorder
C0236736|T048|SY|46975003|SNOMEDCT_CORE|Cocaine induced mental disorder|Cocaine-induced organic mental disorder
C0236736|T048|PT|46975003|SNOMEDCT_CORE|Cocaine-induced organic mental disorder|Cocaine-induced organic mental disorder
C0236736|T048|FN|46975003|SNOMEDCT_CORE|Cocaine-induced organic mental disorder|Cocaine-induced organic mental disorder
C0236736|T048|IS|46975003|SNOMEDCT_CORE|Cocaine-induced organic mental disorder, NOS|Cocaine-induced organic mental disorder
C0236736|T048|SY|46975003|SNOMEDCT_CORE|Cocaine-related disorder|Cocaine-induced organic mental disorder
C0236736|T048|IS|46975003|SNOMEDCT_CORE|Cocaine-related disorder, NOS|Cocaine-induced organic mental disorder
C0236747|T048|PT|37739004|SNOMEDCT_CORE|Mood disorder due to a general medical condition|Mood disorder due to a general medical condition
C0236747|T048|FN|37739004|SNOMEDCT_CORE|Mood disorder due to a general medical condition|Mood disorder due to a general medical condition
C0236748|T048|PT|52910006|SNOMEDCT_CORE|Anxiety disorder due to a general medical condition|Anxiety disorder due to a general medical condition
C0236748|T048|FN|52910006|SNOMEDCT_CORE|Anxiety disorder due to a general medical condition|Anxiety disorder due to a general medical condition
C0236748|T048|SY|52910006|SNOMEDCT_CORE|Anxiety disorder due to general medical condition|Anxiety disorder due to a general medical condition
C0236748|T048|SY|52910006|SNOMEDCT_CORE|Anxiety disorder due to medical disorder|Anxiety disorder due to a general medical condition
C0236758|T048|PT|28884001|SNOMEDCT_CORE|Moderate bipolar I disorder, single manic episode|Moderate bipolar I disorder, single manic episode
C0236758|T048|FN|28884001|SNOMEDCT_CORE|Moderate bipolar I disorder, single manic episode|Moderate bipolar I disorder, single manic episode
C0236761|T048|SY|78269000|SNOMEDCT_CORE|Bipolar 1 disorder, single manic episode, in partial remission|Bipolar I disorder, single manic episode, in partial remission
C0236761|T048|PT|78269000|SNOMEDCT_CORE|Bipolar I disorder, single manic episode, in partial remission|Bipolar I disorder, single manic episode, in partial remission
C0236761|T048|FN|78269000|SNOMEDCT_CORE|Bipolar I disorder, single manic episode, in partial remission|Bipolar I disorder, single manic episode, in partial remission
C0236763|T048|PT|70747007|SNOMEDCT_CORE|Major depression single episode, in partial remission|Major depression single episode, in partial remission
C0236763|T048|FN|70747007|SNOMEDCT_CORE|Major depression single episode, in partial remission|Major depression single episode, in partial remission
C0236763|T048|SY|70747007|SNOMEDCT_CORE|Major depression, single episode, in partial remission|Major depression single episode, in partial remission
C0236764|T048|PT|33135002|SNOMEDCT_CORE|Recurrent major depression in partial remission|Recurrent major depression in partial remission
C0236764|T048|FN|33135002|SNOMEDCT_CORE|Recurrent major depression in partial remission|Recurrent major depression in partial remission
C0236765|T048|SY|31446002|SNOMEDCT_CORE|Bipolar affective disorder, current episode hypomanic|Bipolar I disorder, most recent episode hypomanic
C0236765|T048|PT|31446002|SNOMEDCT_CORE|Bipolar I disorder, most recent episode hypomanic|Bipolar I disorder, most recent episode hypomanic
C0236765|T048|FN|31446002|SNOMEDCT_CORE|Bipolar I disorder, most recent episode hypomanic|Bipolar I disorder, most recent episode hypomanic
C0236767|T048|SY|71984005|SNOMEDCT_CORE|Mild bipolar I disorder, most recent episode manic|Mild manic bipolar I disorder
C0236767|T048|IS|71984005|SNOMEDCT_CORE|Mild manic bipolar disorder|Mild manic bipolar I disorder
C0236767|T048|PT|71984005|SNOMEDCT_CORE|Mild manic bipolar I disorder|Mild manic bipolar I disorder
C0236767|T048|FN|71984005|SNOMEDCT_CORE|Mild manic bipolar I disorder|Mild manic bipolar I disorder
C0236768|T048|SY|82998009|SNOMEDCT_CORE|Moderate bipolar I disorder, most recent episode manic|Moderate manic bipolar I disorder
C0236768|T048|IS|82998009|SNOMEDCT_CORE|Moderate manic bipolar disorder|Moderate manic bipolar I disorder
C0236768|T048|PT|82998009|SNOMEDCT_CORE|Moderate manic bipolar I disorder|Moderate manic bipolar I disorder
C0236768|T048|FN|82998009|SNOMEDCT_CORE|Moderate manic bipolar I disorder|Moderate manic bipolar I disorder
C0236770|T048|SY|28663008|SNOMEDCT_CORE|Severe bipolar I disorder, most recent episode manic, with psychotic features|Severe manic bipolar I disorder with psychotic features
C0236770|T048|IS|28663008|SNOMEDCT_CORE|Severe manic bipolar disorder with psychotic features|Severe manic bipolar I disorder with psychotic features
C0236770|T048|PT|28663008|SNOMEDCT_CORE|Severe manic bipolar I disorder with psychotic features|Severe manic bipolar I disorder with psychotic features
C0236770|T048|FN|28663008|SNOMEDCT_CORE|Severe manic bipolar I disorder with psychotic features|Severe manic bipolar I disorder with psychotic features
C0236771|T048|SY|63249007|SNOMEDCT_CORE|Bipolar I disorder, most recent episode manic, in partial remission|Manic bipolar I disorder in partial remission
C0236771|T048|IS|63249007|SNOMEDCT_CORE|Manic bipolar disorder in partial remission|Manic bipolar I disorder in partial remission
C0236771|T048|PT|63249007|SNOMEDCT_CORE|Manic bipolar I disorder in partial remission|Manic bipolar I disorder in partial remission
C0236771|T048|FN|63249007|SNOMEDCT_CORE|Manic bipolar I disorder in partial remission|Manic bipolar I disorder in partial remission
C0236772|T048|SY|30935000|SNOMEDCT_CORE|Bipolar I disorder, most recent episode manic, in full remission|Manic bipolar I disorder in full remission
C0236772|T048|IS|30935000|SNOMEDCT_CORE|Manic bipolar disorder in full remission|Manic bipolar I disorder in full remission
C0236772|T048|PT|30935000|SNOMEDCT_CORE|Manic bipolar I disorder in full remission|Manic bipolar I disorder in full remission
C0236772|T048|FN|30935000|SNOMEDCT_CORE|Manic bipolar I disorder in full remission|Manic bipolar I disorder in full remission
C0236773|T048|IS|49468007|SNOMEDCT_CORE|Bipolar I disorder, most recent episode depressed|Depressed bipolar I disorder
C0236773|T048|IS|49468007|SNOMEDCT_CORE|Depressed bipolar disorder, NOS|Depressed bipolar I disorder
C0236773|T048|PT|49468007|SNOMEDCT_CORE|Depressed bipolar I disorder|Depressed bipolar I disorder
C0236773|T048|FN|49468007|SNOMEDCT_CORE|Depressed bipolar I disorder|Depressed bipolar I disorder
C0236773|T048|IS|49468007|SNOMEDCT_CORE|Depressed bipolar I disorder, NOS|Depressed bipolar I disorder
C0236774|T048|SY|74686005|SNOMEDCT_CORE|Mild bipolar I disorder, most recent episode depressed|Mild depressed bipolar I disorder
C0236774|T048|IS|74686005|SNOMEDCT_CORE|Mild depressed bipolar disorder|Mild depressed bipolar I disorder
C0236774|T048|PT|74686005|SNOMEDCT_CORE|Mild depressed bipolar I disorder|Mild depressed bipolar I disorder
C0236774|T048|FN|74686005|SNOMEDCT_CORE|Mild depressed bipolar I disorder|Mild depressed bipolar I disorder
C0236775|T048|SY|66631006|SNOMEDCT_CORE|Moderate bipolar I disorder, most recent episode depressed|Moderate depressed bipolar I disorder
C0236775|T048|IS|66631006|SNOMEDCT_CORE|Moderate depressed bipolar disorder|Moderate depressed bipolar I disorder
C0236775|T048|PT|66631006|SNOMEDCT_CORE|Moderate depressed bipolar I disorder|Moderate depressed bipolar I disorder
C0236775|T048|FN|66631006|SNOMEDCT_CORE|Moderate depressed bipolar I disorder|Moderate depressed bipolar I disorder
C0236776|T048|SY|61403008|SNOMEDCT_CORE|Severe bipolar I disorder, most recent episode depressed without psychotic features|Severe depressed bipolar I disorder without psychotic features
C0236776|T048|IS|61403008|SNOMEDCT_CORE|Severe depressed bipolar disorder without psychotic features|Severe depressed bipolar I disorder without psychotic features
C0236776|T048|PT|61403008|SNOMEDCT_CORE|Severe depressed bipolar I disorder without psychotic features|Severe depressed bipolar I disorder without psychotic features
C0236776|T048|FN|61403008|SNOMEDCT_CORE|Severe depressed bipolar I disorder without psychotic features|Severe depressed bipolar I disorder without psychotic features
C0236777|T048|SY|59617007|SNOMEDCT_CORE|Severe bipolar I disorder, most recent episode depressed with psychotic features|Severe depressed bipolar I disorder with psychotic features
C0236777|T048|IS|59617007|SNOMEDCT_CORE|Severe depressed bipolar disorder with psychotic features|Severe depressed bipolar I disorder with psychotic features
C0236777|T048|PT|59617007|SNOMEDCT_CORE|Severe depressed bipolar I disorder with psychotic features|Severe depressed bipolar I disorder with psychotic features
C0236777|T048|FN|59617007|SNOMEDCT_CORE|Severe depressed bipolar I disorder with psychotic features|Severe depressed bipolar I disorder with psychotic features
C0236778|T048|SY|49512000|SNOMEDCT_CORE|Bipolar I disorder, most recent episode depressed, in partial remission|Depressed bipolar I disorder in partial remission
C0236778|T048|IS|49512000|SNOMEDCT_CORE|Depressed bipolar disorder in partial remission|Depressed bipolar I disorder in partial remission
C0236778|T048|PT|49512000|SNOMEDCT_CORE|Depressed bipolar I disorder in partial remission|Depressed bipolar I disorder in partial remission
C0236778|T048|FN|49512000|SNOMEDCT_CORE|Depressed bipolar I disorder in partial remission|Depressed bipolar I disorder in partial remission
C0236779|T048|SY|22121000|SNOMEDCT_CORE|Bipolar I disorder, most recent episode depressed, in full remission|Depressed bipolar I disorder in full remission
C0236779|T048|IS|22121000|SNOMEDCT_CORE|Depressed bipolar disorder in full remission|Depressed bipolar I disorder in full remission
C0236779|T048|PT|22121000|SNOMEDCT_CORE|Depressed bipolar I disorder in full remission|Depressed bipolar I disorder in full remission
C0236779|T048|FN|22121000|SNOMEDCT_CORE|Depressed bipolar I disorder in full remission|Depressed bipolar I disorder in full remission
C0236780|T048|SY|16506000|SNOMEDCT_CORE|Bipolar I disorder, most recent episode mixed|Mixed bipolar I disorder
C0236780|T048|IS|16506000|SNOMEDCT_CORE|Mixed bipolar disorder, NOS|Mixed bipolar I disorder
C0236780|T048|PT|16506000|SNOMEDCT_CORE|Mixed bipolar I disorder|Mixed bipolar I disorder
C0236780|T048|FN|16506000|SNOMEDCT_CORE|Mixed bipolar I disorder|Mixed bipolar I disorder
C0236780|T048|IS|16506000|SNOMEDCT_CORE|Mixed bipolar I disorder, NOS|Mixed bipolar I disorder
C0236781|T048|SY|43769008|SNOMEDCT_CORE|Mild bipolar I disorder, most recent episode mixed|Mild mixed bipolar I disorder
C0236781|T048|IS|43769008|SNOMEDCT_CORE|Mild mixed bipolar disorder|Mild mixed bipolar I disorder
C0236781|T048|PT|43769008|SNOMEDCT_CORE|Mild mixed bipolar I disorder|Mild mixed bipolar I disorder
C0236781|T048|FN|43769008|SNOMEDCT_CORE|Mild mixed bipolar I disorder|Mild mixed bipolar I disorder
C0236782|T048|SY|40926005|SNOMEDCT_CORE|Moderate bipolar I disorder, most recent episode mixed|Moderate mixed bipolar I disorder
C0236782|T048|IS|40926005|SNOMEDCT_CORE|Moderate mixed bipolar disorder|Moderate mixed bipolar I disorder
C0236782|T048|FN|40926005|SNOMEDCT_CORE|Moderate mixed bipolar I disorder|Moderate mixed bipolar I disorder
C0236782|T048|PT|40926005|SNOMEDCT_CORE|Moderate mixed bipolar I disorder|Moderate mixed bipolar I disorder
C0236783|T048|SY|46229002|SNOMEDCT_CORE|Severe bipolar I disorder, most recent episode mixed, without psychotic features|Severe mixed bipolar I disorder without psychotic features
C0236783|T048|IS|46229002|SNOMEDCT_CORE|Severe mixed bipolar disorder without psychotic features|Severe mixed bipolar I disorder without psychotic features
C0236783|T048|PT|46229002|SNOMEDCT_CORE|Severe mixed bipolar I disorder without psychotic features|Severe mixed bipolar I disorder without psychotic features
C0236783|T048|FN|46229002|SNOMEDCT_CORE|Severe mixed bipolar I disorder without psychotic features|Severe mixed bipolar I disorder without psychotic features
C0236784|T048|SY|10981006|SNOMEDCT_CORE|Severe bipolar I disorder, most recent episode mixed, with psychotic features|Severe mixed bipolar I disorder with psychotic features
C0236784|T048|IS|10981006|SNOMEDCT_CORE|Severe mixed bipolar disorder with psychotic features|Severe mixed bipolar I disorder with psychotic features
C0236784|T048|PT|10981006|SNOMEDCT_CORE|Severe mixed bipolar I disorder with psychotic features|Severe mixed bipolar I disorder with psychotic features
C0236784|T048|FN|10981006|SNOMEDCT_CORE|Severe mixed bipolar I disorder with psychotic features|Severe mixed bipolar I disorder with psychotic features
C0236785|T048|SY|36583000|SNOMEDCT_CORE|Bipolar I disorder, most recent episode mixed, in partial remission|Mixed bipolar I disorder in partial remission
C0236785|T048|IS|36583000|SNOMEDCT_CORE|Mixed bipolar disorder in partial remission|Mixed bipolar I disorder in partial remission
C0236785|T048|PT|36583000|SNOMEDCT_CORE|Mixed bipolar I disorder in partial remission|Mixed bipolar I disorder in partial remission
C0236785|T048|FN|36583000|SNOMEDCT_CORE|Mixed bipolar I disorder in partial remission|Mixed bipolar I disorder in partial remission
C0236786|T048|SY|111485001|SNOMEDCT_CORE|Bipolar I disorder, most recent episode mixed, in full remission|Mixed bipolar I disorder in full remission
C0236786|T048|IS|111485001|SNOMEDCT_CORE|Mixed bipolar disorder in full remission|Mixed bipolar I disorder in full remission
C0236786|T048|PT|111485001|SNOMEDCT_CORE|Mixed bipolar I disorder in full remission|Mixed bipolar I disorder in full remission
C0236786|T048|FN|111485001|SNOMEDCT_CORE|Mixed bipolar I disorder in full remission|Mixed bipolar I disorder in full remission
C0236788|T048|SY|83225003|SNOMEDCT_CORE|Bipolar 2 disorder|Bipolar II disorder
C0236788|T048|PT|83225003|SNOMEDCT_CORE|Bipolar II disorder|Bipolar II disorder
C0236788|T048|FN|83225003|SNOMEDCT_CORE|Bipolar II disorder|Bipolar II disorder
C0236788|T048|IS|83225003|SNOMEDCT_CORE|Bipolar II disorder, NOS|Bipolar II disorder
C0236792|T048|SY|23560001|SNOMEDCT_CORE|Asperger disorder|Asperger's disorder
C0236792|T048|PT|23560001|SNOMEDCT_CORE|Asperger's disorder|Asperger's disorder
C0236792|T048|FN|23560001|SNOMEDCT_CORE|Asperger's disorder|Asperger's disorder
C0236792|T048|SY|23560001|SNOMEDCT_CORE|Asperger's syndrome|Asperger's disorder
C0236792|T048|SY|23560001|SNOMEDCT_CORE|Aspergers disorder|Asperger's disorder
C0236794|T048|PT|56576003|SNOMEDCT_CORE|Panic disorder without agoraphobia|Panic disorder without agoraphobia
C0236794|T048|FN|56576003|SNOMEDCT_CORE|Panic disorder without agoraphobia|Panic disorder without agoraphobia
C0236794|T048|IS|56576003|SNOMEDCT_CORE|Panic disorder without agoraphobia, NOS|Panic disorder without agoraphobia
C0236800|T048|PT|35607004|SNOMEDCT_CORE|Panic disorder with agoraphobia|Panic disorder with agoraphobia
C0236800|T048|FN|35607004|SNOMEDCT_CORE|Panic disorder with agoraphobia|Panic disorder with agoraphobia
C0236800|T048|IS|35607004|SNOMEDCT_CORE|Panic disorder with agoraphobia, NOS|Panic disorder with agoraphobia
C0236801|T048|SY|54587008|SNOMEDCT_CORE|Isolated phobia|Simple phobia
C0236801|T048|PT|54587008|SNOMEDCT_CORE|Simple phobia|Simple phobia
C0236801|T048|FN|54587008|SNOMEDCT_CORE|Simple phobia|Simple phobia
C0236801|T048|SY|54587008|SNOMEDCT_CORE|Specific phobia|Simple phobia
C0236804|T048|SY|21647008|SNOMEDCT_CORE|Amfetamine dependence|Amphetamine dependence
C0236804|T048|PT|21647008|SNOMEDCT_CORE|Amphetamine dependence|Amphetamine dependence
C0236804|T048|FN|21647008|SNOMEDCT_CORE|Amphetamine dependence|Amphetamine dependence
C0236807|T048|SY|84758004|SNOMEDCT_CORE|Amfetamine abuse|Amphetamine abuse
C0236807|T048|PT|84758004|SNOMEDCT_CORE|Amphetamine abuse|Amphetamine abuse
C0236807|T048|FN|84758004|SNOMEDCT_CORE|Amphetamine abuse|Amphetamine abuse
C0236807|T048|SY|84758004|SNOMEDCT_CORE|Drug abuse using speed|Amphetamine abuse
C0236812|T048|PT|74142004|SNOMEDCT_CORE|Feeding disorder of infancy OR early childhood|Feeding disorder of infancy OR early childhood
C0236812|T048|IS|74142004|SNOMEDCT_CORE|Feeding disorder of infancy or early childhood|Feeding disorder of infancy OR early childhood
C0236812|T048|FN|74142004|SNOMEDCT_CORE|Feeding disorder of infancy OR early childhood|Feeding disorder of infancy OR early childhood
C0236812|T048|SY|74142004|SNOMEDCT_CORE|Feeding disorder, infancy or early childhood|Feeding disorder of infancy OR early childhood
C0236816|T048|SY|67195008|SNOMEDCT_CORE|Acute crisis reaction|Acute stress disorder
C0236816|T048|SY|67195008|SNOMEDCT_CORE|Acute reaction to stress|Acute stress disorder
C0236816|T048|PT|67195008|SNOMEDCT_CORE|Acute stress disorder|Acute stress disorder
C0236816|T048|FN|67195008|SNOMEDCT_CORE|Acute stress disorder|Acute stress disorder
C0236816|T048|SY|67195008|SNOMEDCT_CORE|Acute stress reaction|Acute stress disorder
C0236816|T048|SY|67195008|SNOMEDCT_CORE|Gross stress reaction|Acute stress disorder
C0236816|T048|IS|67195008|SNOMEDCT_CORE|Gross stress reaction, NOS|Acute stress disorder
C0236816|T048|SY|67195008|SNOMEDCT_CORE|Psychic shock|Acute stress disorder
C0236826|T048|PT|229733002|SNOMEDCT_CORE|Expressive language disorder|Expressive language disorder
C0236826|T048|FN|229733002|SNOMEDCT_CORE|Expressive language disorder|Expressive language disorder
C0236827|T048|PT|25766007|SNOMEDCT_CORE|Mixed receptive-expressive language disorder|Mixed receptive-expressive language disorder
C0236827|T048|FN|25766007|SNOMEDCT_CORE|Mixed receptive-expressive language disorder|Mixed receptive-expressive language disorder
C0236828|T048|PT|386701004|SNOMEDCT_CORE|Developmental articulation disorder|Developmental articulation disorder
C0236828|T048|FN|386701004|SNOMEDCT_CORE|Developmental articulation disorder|Developmental articulation disorder
C0236828|T048|SY|386701004|SNOMEDCT_CORE|Developmental speech articulation disorder|Developmental articulation disorder
C0236828|T048|IS|386701004|SNOMEDCT_CORE|Developmental speech articulation disorder|Developmental articulation disorder
C0236845|T047|PT|111489007|SNOMEDCT_CORE|Breathing-related sleep disorder|Breathing-related sleep disorder
C0236845|T047|FN|111489007|SNOMEDCT_CORE|Breathing-related sleep disorder|Breathing-related sleep disorder
C0236845|T047|IS|111489007|SNOMEDCT_CORE|Breathing-related sleep disorder, NOS|Breathing-related sleep disorder
C0236848|T048|PT|102891000|SNOMEDCT_CORE|Age-related cognitive decline|Age-related cognitive decline
C0236848|T048|FN|102891000|SNOMEDCT_CORE|Age-related cognitive decline|Age-related cognitive decline
C0236849|T048|PT|73149003|SNOMEDCT_CORE|Encopresis with constipation AND overflow incontinence|Encopresis with constipation AND overflow incontinence
C0236849|T048|IS|73149003|SNOMEDCT_CORE|Encopresis with constipation and overflow incontinence|Encopresis with constipation AND overflow incontinence
C0236849|T048|OF|73149003|SNOMEDCT_CORE|Encopresis with constipation AND overflow incontinence|Encopresis with constipation AND overflow incontinence
C0236849|T048|FN|73149003|SNOMEDCT_CORE|Encopresis with constipation AND overflow incontinence|Encopresis with constipation AND overflow incontinence
C0236861|T033|SY|371779005|SNOMEDCT_CORE|Physical abuse of child|Physical child abuse
C0236861|T033|PT|371779005|SNOMEDCT_CORE|Physical child abuse|Physical child abuse
C0236861|T033|OF|371779005|SNOMEDCT_CORE|Physical child abuse|Physical child abuse
C0236861|T033|FN|371779005|SNOMEDCT_CORE|Physical child abuse|Physical child abuse
C0237020|T191|OAS|119424003|SNOMEDCT_CORE|Benign cystic ovarian teratoma|Dermoid cyst of ovary
C0237020|T191|OAP|119424003|SNOMEDCT_CORE|Dermoid cyst of ovary|Dermoid cyst of ovary
C0237020|T191|OF|119424003|SNOMEDCT_CORE|Dermoid cyst of ovary|Dermoid cyst of ovary
C0237020|T191|OAS|119424003|SNOMEDCT_CORE|Mature cystic teratoma of ovary|Dermoid cyst of ovary
C0237020|T191|OAF|119424003|SNOMEDCT_CORE|Mature cystic teratoma of ovary|Dermoid cyst of ovary
C0237154|T033|PT|32911000|SNOMEDCT_CORE|Homeless|Homeless
C0237154|T033|FN|32911000|SNOMEDCT_CORE|Homeless|Homeless
C0237154|T033|PT|266935003|SNOMEDCT_CORE|Housing lack|Homeless
C0237154|T033|FN|266935003|SNOMEDCT_CORE|Housing lack|Homeless
C0237154|T033|SY|32911000|SNOMEDCT_CORE|Living on the street|Homeless
C0237236|T048|PT|248110007|SNOMEDCT_CORE|Sexual assault|Sexual assault
C0237236|T048|OAP|422608009|SNOMEDCT_CORE|Sexual assault|Sexual assault
C0237236|T048|OF|248110007|SNOMEDCT_CORE|Sexual assault|Sexual assault
C0237236|T048|OAF|422608009|SNOMEDCT_CORE|Sexual assault|Sexual assault
C0237236|T048|FN|248110007|SNOMEDCT_CORE|Sexual assault|Sexual assault
C0237284|T033|PT|422768004|SNOMEDCT_CORE|Unresponsive|Unresponsive
C0237284|T033|FN|422768004|SNOMEDCT_CORE|Unresponsive|Unresponsive
C0237314|T033|OAS|248650006|SNOMEDCT_CORE|Heart beats irregular|Irregular heart beat
C0237314|T033|OAP|248650006|SNOMEDCT_CORE|Heart irregular|Irregular heart beat
C0237314|T033|OAF|248650006|SNOMEDCT_CORE|Heart irregular|Irregular heart beat
C0237314|T033|PT|361137007|SNOMEDCT_CORE|Irregular heart beat|Irregular heart beat
C0237314|T033|FN|361137007|SNOMEDCT_CORE|Irregular heart beat|Irregular heart beat
C0237314|T033|OAS|248650006|SNOMEDCT_CORE|Palpitations - irregular|Irregular heart beat
C0237349|T033|PT|424890008|SNOMEDCT_CORE|Unbalanced diet|Unbalanced diet
C0237349|T033|FN|424890008|SNOMEDCT_CORE|Unbalanced diet|Unbalanced diet
C0238015|T047|PT|129618003|SNOMEDCT_CORE|Autonomic dysreflexia|Autonomic dysreflexia
C0238015|T047|FN|129618003|SNOMEDCT_CORE|Autonomic dysreflexia|Autonomic dysreflexia
C0238015|T047|SY|129618003|SNOMEDCT_CORE|Dysreflexia|Autonomic dysreflexia
C0238033|T191|PT|372096000|SNOMEDCT_CORE|Carcinoma of male breast|Carcinoma of male breast
C0238033|T191|FN|372096000|SNOMEDCT_CORE|Carcinoma of male breast|Carcinoma of male breast
C0238051|T047|PT|427020007|SNOMEDCT_CORE|Cerebral vasculitis|Cerebral vasculitis
C0238051|T047|FN|427020007|SNOMEDCT_CORE|Cerebral vasculitis|Cerebral vasculitis
C0238067|T047|SY|19311003|SNOMEDCT_CORE|CC - Collagenous colitis|Collagenous colitis
C0238067|T047|PT|19311003|SNOMEDCT_CORE|Collagenous colitis|Collagenous colitis
C0238067|T047|FN|19311003|SNOMEDCT_CORE|Collagenous colitis|Collagenous colitis
C0238074|T047|SY|87837008|SNOMEDCT_CORE|Chronic cardiopulmonary disease|Chronic pulmonary heart disease
C0238074|T047|PT|87837008|SNOMEDCT_CORE|Chronic pulmonary heart disease|Chronic pulmonary heart disease
C0238074|T047|FN|87837008|SNOMEDCT_CORE|Chronic pulmonary heart disease|Chronic pulmonary heart disease
C0238074|T047|IS|87837008|SNOMEDCT_CORE|Chronic pulmonary heart disease, NOS|Chronic pulmonary heart disease
C0238106|T047|PT|423590009|SNOMEDCT_CORE|Clostridium difficile colitis|Clostridium difficile colitis
C0238106|T047|FN|423590009|SNOMEDCT_CORE|Clostridium difficile colitis|Clostridium difficile colitis
C0238106|T047|SY|423590009|SNOMEDCT_CORE|Pseudomembranous colitis|Clostridium difficile colitis
C0238106|T047|SY|423590009|SNOMEDCT_CORE|Pseudomembranous enterocolitis|Clostridium difficile colitis
C0238122|T191|PT|276870001|SNOMEDCT_CORE|Carcinoma of fallopian tube|Carcinoma of fallopian tube
C0238122|T191|FN|276870001|SNOMEDCT_CORE|Carcinoma of fallopian tube|Carcinoma of fallopian tube
C0238124|T047|SYGB|52486002|SNOMEDCT_CORE|Necrotising cellulitis|Necrotizing fasciitis
C0238124|T047|IS|52486002|SNOMEDCT_CORE|Necrotising erysipelas|Necrotizing fasciitis
C0238124|T047|PTGB|52486002|SNOMEDCT_CORE|Necrotising fasciitis|Necrotizing fasciitis
C0238124|T047|SYGB|52486002|SNOMEDCT_CORE|Necrotising myositis|Necrotizing fasciitis
C0238124|T047|SY|52486002|SNOMEDCT_CORE|Necrotizing cellulitis|Necrotizing fasciitis
C0238124|T047|IS|52486002|SNOMEDCT_CORE|Necrotizing erysipelas|Necrotizing fasciitis
C0238124|T047|PT|52486002|SNOMEDCT_CORE|Necrotizing fasciitis|Necrotizing fasciitis
C0238124|T047|FN|52486002|SNOMEDCT_CORE|Necrotizing fasciitis|Necrotizing fasciitis
C0238124|T047|SY|52486002|SNOMEDCT_CORE|Necrotizing myositis|Necrotizing fasciitis
C0238124|T047|IS|52486002|SNOMEDCT_CORE|Streptococcal gangrene|Necrotizing fasciitis
C0238190|T047|SY|72315009|SNOMEDCT_CORE|IBM - Inclusion body myositis|Inclusion body myositis
C0238190|T047|FN|72315009|SNOMEDCT_CORE|Inclusion body myositis|Inclusion body myositis
C0238190|T047|PT|72315009|SNOMEDCT_CORE|Inclusion body myositis|Inclusion body myositis
C0238198|T191|PT|420120006|SNOMEDCT_CORE|Gastrointestinal stromal tumor|Gastrointestinal stromal tumor
C0238198|T191|FN|420120006|SNOMEDCT_CORE|Gastrointestinal stromal tumor|Gastrointestinal stromal tumor
C0238198|T191|PTGB|420120006|SNOMEDCT_CORE|Gastrointestinal stromal tumour|Gastrointestinal stromal tumor
C0238198|T191|SY|420120006|SNOMEDCT_CORE|GIST - Gastrointestinal stromal tumor|Gastrointestinal stromal tumor
C0238198|T191|SYGB|420120006|SNOMEDCT_CORE|GIST - Gastrointestinal stromal tumour|Gastrointestinal stromal tumor
C0238217|T046|PT|236570004|SNOMEDCT_CORE|Renal transplant rejection|Renal transplant rejection
C0238217|T046|FN|236570004|SNOMEDCT_CORE|Renal transplant rejection|Renal transplant rejection
C0238218|T037|SY|239720000|SNOMEDCT_CORE|Tear of cartilage of knee|Tear of meniscus of knee
C0238218|T037|PT|239720000|SNOMEDCT_CORE|Tear of meniscus of knee|Tear of meniscus of knee
C0238218|T037|FN|239720000|SNOMEDCT_CORE|Tear of meniscus of knee|Tear of meniscus of knee
C0238218|T037|IS|239720000|SNOMEDCT_CORE|Torn cartilage|Tear of meniscus of knee
C0238218|T037|SY|239720000|SNOMEDCT_CORE|Torn meniscus|Tear of meniscus of knee
C0238246|T191|PTGB|93469006|SNOMEDCT_CORE|Haemangioma of liver|Hemangioma of liver
C0238246|T191|PT|93469006|SNOMEDCT_CORE|Hemangioma of liver|Hemangioma of liver
C0238246|T191|FN|93469006|SNOMEDCT_CORE|Hemangioma of liver|Hemangioma of liver
C0238246|T191|SY|93469006|SNOMEDCT_CORE|Hepatic angioma|Hemangioma of liver
C0238246|T191|SYGB|93469006|SNOMEDCT_CORE|Hepatic haemangioma|Hemangioma of liver
C0238246|T191|SY|93469006|SNOMEDCT_CORE|Hepatic hemangioma|Hemangioma of liver
C0238300|T033|PT|231841004|SNOMEDCT_CORE|Stenosis of nasolacrimal duct|Stenosis of nasolacrimal duct
C0238300|T033|FN|231841004|SNOMEDCT_CORE|Stenosis of nasolacrimal duct|Stenosis of nasolacrimal duct
C0238301|T191|SY|187692001|SNOMEDCT_CORE|CA - Cancer of nasopharynx|CA - Cancer of nasopharynx
C0238301|T191|SY|187692001|SNOMEDCT_CORE|Cancer of nasopharynx|CA - Cancer of nasopharynx
C0238358|T047|OAS|240093008|SNOMEDCT_CORE|Familial hypokalaemic periodic paralysis|Familial hypokalemic periodic paralysis
C0238358|T047|PTGB|82732003|SNOMEDCT_CORE|Familial hypokalaemic periodic paralysis|Familial hypokalemic periodic paralysis
C0238358|T047|OAS|240093008|SNOMEDCT_CORE|Familial hypokalemic periodic paralysis|Familial hypokalemic periodic paralysis
C0238358|T047|PT|82732003|SNOMEDCT_CORE|Familial hypokalemic periodic paralysis|Familial hypokalemic periodic paralysis
C0238358|T047|FN|82732003|SNOMEDCT_CORE|Familial hypokalemic periodic paralysis|Familial hypokalemic periodic paralysis
C0238358|T047|OAP|240093008|SNOMEDCT_CORE|Hypokalaemic periodic paralysis|Familial hypokalemic periodic paralysis
C0238358|T047|SYGB|82732003|SNOMEDCT_CORE|Hypokalaemic periodic paralysis|Familial hypokalemic periodic paralysis
C0238358|T047|OAP|240093008|SNOMEDCT_CORE|Hypokalemic periodic paralysis|Familial hypokalemic periodic paralysis
C0238358|T047|SY|82732003|SNOMEDCT_CORE|Hypokalemic periodic paralysis|Familial hypokalemic periodic paralysis
C0238358|T047|OAF|240093008|SNOMEDCT_CORE|Hypokalemic periodic paralysis|Familial hypokalemic periodic paralysis
C0238358|T047|SY|82732003|SNOMEDCT_CORE|Periodic paralysis I|Familial hypokalemic periodic paralysis
C0238397|T190|PT|95441000|SNOMEDCT_CORE|Pulmonary artery stenosis|Pulmonary artery stenosis
C0238397|T190|FN|95441000|SNOMEDCT_CORE|Pulmonary artery stenosis|Pulmonary artery stenosis
C0238418|T047|PT|27717006|SNOMEDCT_CORE|Abscess of scrotum|Abscess of scrotum
C0238418|T047|FN|27717006|SNOMEDCT_CORE|Abscess of scrotum|Abscess of scrotum
C0238418|T047|SY|27717006|SNOMEDCT_CORE|Scrotal abscess|Abscess of scrotum
C0238425|T047|PTGB|417425009|SNOMEDCT_CORE|Haemoglobin SS disease with crisis|Hemoglobin SS disease with crisis
C0238425|T047|PT|417425009|SNOMEDCT_CORE|Hemoglobin SS disease with crisis|Hemoglobin SS disease with crisis
C0238425|T047|FN|417425009|SNOMEDCT_CORE|Hemoglobin SS disease with crisis|Hemoglobin SS disease with crisis
C0238425|T047|SYGB|417425009|SNOMEDCT_CORE|Sickle cell anaemia with crisis|Hemoglobin SS disease with crisis
C0238425|T047|IS|417425009|SNOMEDCT_CORE|SIckle cell anaemia with crisis|Hemoglobin SS disease with crisis
C0238425|T047|SY|417425009|SNOMEDCT_CORE|Sickle cell anemia with crisis|Hemoglobin SS disease with crisis
C0238425|T047|SY|417425009|SNOMEDCT_CORE|Sickle cell crisis|Hemoglobin SS disease with crisis
C0238441|T190|SY|22668006|SNOMEDCT_CORE|SGS - Subglottic stenosis|Subglottic stenosis
C0238441|T190|PT|22668006|SNOMEDCT_CORE|Subglottic stenosis|Subglottic stenosis
C0238441|T190|FN|22668006|SNOMEDCT_CORE|Subglottic stenosis|Subglottic stenosis
C0238460|T047|SY|4997005|SNOMEDCT_CORE|Factitious hyperthyroidism|Thyrotoxicosis factitia
C0238460|T047|SY|4997005|SNOMEDCT_CORE|Factitious hyperthyroidism from ingestion of excessive thyroid material|Thyrotoxicosis factitia
C0238460|T047|PT|4997005|SNOMEDCT_CORE|Thyrotoxicosis factitia|Thyrotoxicosis factitia
C0238460|T047|FN|4997005|SNOMEDCT_CORE|Thyrotoxicosis factitia|Thyrotoxicosis factitia
C0238462|T191|SY|255032005|SNOMEDCT_CORE|Medullary carcinoma of thyroid|Medullary thyroid carcinoma
C0238462|T191|PT|255032005|SNOMEDCT_CORE|Medullary thyroid carcinoma|Medullary thyroid carcinoma
C0238462|T191|FN|255032005|SNOMEDCT_CORE|Medullary thyroid carcinoma|Medullary thyroid carcinoma
C0238462|T191|SY|255032005|SNOMEDCT_CORE|MTC - Medullary thyroid carcinoma|Medullary thyroid carcinoma
C0238463|T191|PT|255029007|SNOMEDCT_CORE|Papillary thyroid carcinoma|Papillary thyroid carcinoma
C0238463|T191|FN|255029007|SNOMEDCT_CORE|Papillary thyroid carcinoma|Papillary thyroid carcinoma
C0238463|T191|SY|255029007|SNOMEDCT_CORE|PTC - papillary thyroid carcinoma|Papillary thyroid carcinoma
C0238463|T191|IS|255029007|SNOMEDCT_CORE|PTC - Papillary thyroid carcinoma|Papillary thyroid carcinoma
C0238469|T047|PT|33261009|SNOMEDCT_CORE|Abscess of tonsil|Abscess of tonsil
C0238469|T047|FN|33261009|SNOMEDCT_CORE|Abscess of tonsil|Abscess of tonsil
C0238522|T019|IS|30288003|SNOMEDCT_CORE|Roger's disease|Roger's disease
C0238551|T184|PT|301716002|SNOMEDCT_CORE|Left lower quadrant pain|Left lower quadrant pain
C0238551|T184|FN|301716002|SNOMEDCT_CORE|Left lower quadrant pain|Left lower quadrant pain
C0238552|T184|PT|301715003|SNOMEDCT_CORE|Left upper quadrant pain|Left upper quadrant pain
C0238552|T184|FN|301715003|SNOMEDCT_CORE|Left upper quadrant pain|Left upper quadrant pain
C0238634|T033|PT|301779004|SNOMEDCT_CORE|Anal inflammation|Anal inflammation
C0238634|T033|FN|301779004|SNOMEDCT_CORE|Anal inflammation|Anal inflammation
C0238634|T033|SY|301779004|SNOMEDCT_CORE|Inflammation of anus|Anal inflammation
C0238637|T184|PT|68653001|SNOMEDCT_CORE|Anal pain|Anal pain
C0238637|T184|OF|68653001|SNOMEDCT_CORE|Anal pain|Anal pain
C0238637|T184|FN|68653001|SNOMEDCT_CORE|Anal pain|Anal pain
C0238656|T184|PT|202490009|SNOMEDCT_CORE|Ankle joint pain|Ankle pain
C0238656|T184|FN|202490009|SNOMEDCT_CORE|Ankle joint pain|Ankle pain
C0238656|T184|PT|247373008|SNOMEDCT_CORE|Ankle pain|Ankle pain
C0238656|T184|FN|247373008|SNOMEDCT_CORE|Ankle pain|Ankle pain
C0238656|T184|SY|202490009|SNOMEDCT_CORE|Arthralgia of ankle|Ankle pain
C0238669|T190|PT|251036003|SNOMEDCT_CORE|Aortic root dilatation|Aortic root dilatation
C0238669|T190|FN|251036003|SNOMEDCT_CORE|Aortic root dilatation|Aortic root dilatation
C0238729|T033|SY|300863000|SNOMEDCT_CORE|Lump of axilla|Mass of axilla
C0238729|T033|PT|300863000|SNOMEDCT_CORE|Mass of axilla|Mass of axilla
C0238729|T033|FN|300863000|SNOMEDCT_CORE|Mass of axilla|Mass of axilla
C0238738|T047|PT|203095000|SNOMEDCT_CORE|Spasm of back muscles|Spasm of back muscles
C0238738|T047|FN|203095000|SNOMEDCT_CORE|Spasm of back muscles|Spasm of back muscles
C0238775|T033|SY|428090004|SNOMEDCT_CORE|Bladder mass|Mass of urinary bladder
C0238775|T033|SY|428090004|SNOMEDCT_CORE|Mass of bladder|Mass of urinary bladder
C0238775|T033|PT|428090004|SNOMEDCT_CORE|Mass of urinary bladder|Mass of urinary bladder
C0238775|T033|FN|428090004|SNOMEDCT_CORE|Mass of urinary bladder|Mass of urinary bladder
C0238902|T047|PT|230482003|SNOMEDCT_CORE|Carotidynia|Carotidynia
C0238902|T047|FN|230482003|SNOMEDCT_CORE|Carotidynia|Carotidynia
C0239134|T033|SY|28743005|SNOMEDCT_CORE|Bronchial cough|Productive cough
C0239134|T033|SY|28743005|SNOMEDCT_CORE|Chesty cough|Productive cough
C0239134|T033|SY|28743005|SNOMEDCT_CORE|Loose cough|Productive cough
C0239134|T033|SY|28743005|SNOMEDCT_CORE|Moist cough|Productive cough
C0239134|T033|SY|28743005|SNOMEDCT_CORE|Producing sputum|Productive cough
C0239134|T033|PT|28743005|SNOMEDCT_CORE|Productive cough|Productive cough
C0239134|T033|FN|28743005|SNOMEDCT_CORE|Productive cough|Productive cough
C0239233|T184|PT|442076002|SNOMEDCT_CORE|Early satiety|Early satiety
C0239233|T184|SY|442076002|SNOMEDCT_CORE|Early satiety|Early satiety
C0239233|T184|FN|442076002|SNOMEDCT_CORE|Early satiety|Early satiety
C0239266|T184|SY|74323005|SNOMEDCT_CORE|Elbow pain|Pain in elbow
C0239266|T184|PT|74323005|SNOMEDCT_CORE|Pain in elbow|Pain in elbow
C0239266|T184|FN|74323005|SNOMEDCT_CORE|Pain in elbow|Pain in elbow
C0239293|T046|PT|15238002|SNOMEDCT_CORE|Esophageal bleeding|Esophageal bleeding
C0239293|T046|FN|15238002|SNOMEDCT_CORE|Esophageal bleeding|Esophageal bleeding
C0239293|T046|SY|15238002|SNOMEDCT_CORE|Esophageal hemorrhage|Esophageal bleeding
C0239293|T046|SYGB|15238002|SNOMEDCT_CORE|Haemorrhage of oesophagus|Esophageal bleeding
C0239293|T046|SY|15238002|SNOMEDCT_CORE|Hemorrhage of esophagus|Esophageal bleeding
C0239293|T046|PTGB|15238002|SNOMEDCT_CORE|Oesophageal bleeding|Esophageal bleeding
C0239293|T046|SYGB|15238002|SNOMEDCT_CORE|Oesophageal haemorrhage|Esophageal bleeding
C0239295|T047|SY|20639004|SNOMEDCT_CORE|Candida of esophagus|Candidiasis of the esophagus
C0239295|T047|SY|20639004|SNOMEDCT_CORE|Candidiasis of esophagus|Candidiasis of the esophagus
C0239295|T047|SYGB|20639004|SNOMEDCT_CORE|Candidiasis of oesophagus|Candidiasis of the esophagus
C0239295|T047|PT|20639004|SNOMEDCT_CORE|Candidiasis of the esophagus|Candidiasis of the esophagus
C0239295|T047|FN|20639004|SNOMEDCT_CORE|Candidiasis of the esophagus|Candidiasis of the esophagus
C0239295|T047|PTGB|20639004|SNOMEDCT_CORE|Candidiasis of the oesophagus|Candidiasis of the esophagus
C0239295|T047|SY|20639004|SNOMEDCT_CORE|Candidosis of esophagus|Candidiasis of the esophagus
C0239295|T047|SYGB|20639004|SNOMEDCT_CORE|Candidosis of oesophagus|Candidiasis of the esophagus
C0239295|T047|SY|20639004|SNOMEDCT_CORE|Esophageal thrush|Candidiasis of the esophagus
C0239295|T047|SYGB|20639004|SNOMEDCT_CORE|Oesophageal thrush|Candidiasis of the esophagus
C0239340|T033|PT|102572006|SNOMEDCT_CORE|Edema of lower extremity|Edema of lower extremity
C0239340|T033|FN|102572006|SNOMEDCT_CORE|Edema of lower extremity|Edema of lower extremity
C0239340|T033|SY|102572006|SNOMEDCT_CORE|Edema of lower limb|Edema of lower extremity
C0239340|T033|PTGB|102572006|SNOMEDCT_CORE|Oedema of lower extremity|Edema of lower extremity
C0239340|T033|SYGB|102572006|SNOMEDCT_CORE|Oedema of lower limb|Edema of lower extremity
C0239377|T184|IS|102556003|SNOMEDCT_CORE|Arm pain|Pain in upper limb
C0239377|T184|IS|102556003|SNOMEDCT_CORE|Arm pain, NOS|Pain in upper limb
C0239377|T184|PT|102556003|SNOMEDCT_CORE|Pain in upper limb|Pain in upper limb
C0239377|T184|FN|102556003|SNOMEDCT_CORE|Pain in upper limb|Pain in upper limb
C0239377|T184|SY|102556003|SNOMEDCT_CORE|Pain of upper limb|Pain in upper limb
C0239505|T033|PT|299704007|SNOMEDCT_CORE|Lump on face|Lump on face
C0239505|T033|FN|299704007|SNOMEDCT_CORE|Lump on face|Lump on face
C0239505|T033|SY|299704007|SNOMEDCT_CORE|Mass of face|Lump on face
C0239511|T184|PT|309557009|SNOMEDCT_CORE|Numbness of face|Numbness of face
C0239511|T184|FN|309557009|SNOMEDCT_CORE|Numbness of face|Numbness of face
C0239589|T184|SY|18876004|SNOMEDCT_CORE|Finger pain|Pain in finger
C0239589|T184|PT|18876004|SNOMEDCT_CORE|Pain in finger|Pain in finger
C0239589|T184|FN|18876004|SNOMEDCT_CORE|Pain in finger|Pain in finger
C0239598|T033|PT|299060006|SNOMEDCT_CORE|Swelling of finger|Swelling of finger
C0239598|T033|FN|299060006|SNOMEDCT_CORE|Swelling of finger|Swelling of finger
C0239598|T033|SY|299060006|SNOMEDCT_CORE|Swollen finger|Swelling of finger
C0239649|T184|PT|309538000|SNOMEDCT_CORE|Numbness of foot|Numbness of foot
C0239649|T184|FN|309538000|SNOMEDCT_CORE|Numbness of foot|Numbness of foot
C0239652|T033|PTGB|309087008|SNOMEDCT_CORE|Paraesthesia of foot|Paresthesia of foot
C0239652|T033|PT|309087008|SNOMEDCT_CORE|Paresthesia of foot|Paresthesia of foot
C0239652|T033|FN|309087008|SNOMEDCT_CORE|Paresthesia of foot|Paresthesia of foot
C0239667|T184|PT|444899003|SNOMEDCT_CORE|Pain in forearm|Pain in forearm
C0239667|T184|FN|444899003|SNOMEDCT_CORE|Pain in forearm|Pain in forearm
C0239783|T184|SY|102570003|SNOMEDCT_CORE|Groin pain|Inguinal pain
C0239783|T184|PT|102570003|SNOMEDCT_CORE|Inguinal pain|Inguinal pain
C0239783|T184|FN|102570003|SNOMEDCT_CORE|Inguinal pain|Inguinal pain
C0239783|T184|IS|102570003|SNOMEDCT_CORE|Inguinodynia|Inguinal pain
C0239816|T047|SY|238539001|SNOMEDCT_CORE|Dermatitis of hand|Hand eczema
C0239816|T047|SY|238539001|SNOMEDCT_CORE|Hand dermatitis|Hand eczema
C0239816|T047|PT|238539001|SNOMEDCT_CORE|Hand eczema|Hand eczema
C0239816|T047|FN|238539001|SNOMEDCT_CORE|Hand eczema|Hand eczema
C0239832|T184|PT|309521004|SNOMEDCT_CORE|Numbness of hand|Numbness of hand
C0239832|T184|FN|309521004|SNOMEDCT_CORE|Numbness of hand|Numbness of hand
C0239833|T184|PT|53057004|SNOMEDCT_CORE|Hand pain|Hand pain
C0239833|T184|FN|53057004|SNOMEDCT_CORE|Hand pain|Hand pain
C0239833|T184|IS|53057004|SNOMEDCT_CORE|Pain in hand|Hand pain
C0239833|T184|SY|53057004|SNOMEDCT_CORE|Painful hand|Hand pain
C0239836|T184|PTGB|309086004|SNOMEDCT_CORE|Paraesthesia of hand|Paresthesia of hand
C0239836|T184|PT|309086004|SNOMEDCT_CORE|Paresthesia of hand|Paresthesia of hand
C0239836|T184|FN|309086004|SNOMEDCT_CORE|Paresthesia of hand|Paresthesia of hand
C0239886|T184|PT|267096005|SNOMEDCT_CORE|Frontal headache|Frontal headache
C0239886|T184|FN|267096005|SNOMEDCT_CORE|Frontal headache|Frontal headache
C0239937|T033|PTGB|197940006|SNOMEDCT_CORE|Microscopic haematuria|Microscopic hematuria
C0239937|T033|PT|197940006|SNOMEDCT_CORE|Microscopic hematuria|Microscopic hematuria
C0239937|T033|FN|197940006|SNOMEDCT_CORE|Microscopic hematuria|Microscopic hematuria
C0239954|T033|PT|299233007|SNOMEDCT_CORE|Deformity of hip joint|Deformity of hip joint
C0239954|T033|FN|299233007|SNOMEDCT_CORE|Deformity of hip joint|Deformity of hip joint
C0239957|T184|PT|249914008|SNOMEDCT_CORE|Hip stiff|Hip stiff
C0239957|T184|FN|249914008|SNOMEDCT_CORE|Hip stiff|Hip stiff
C0239981|T047|PTGB|119247004|SNOMEDCT_CORE|Hypoalbuminaemia|Hypoalbuminemia
C0239981|T047|PT|119247004|SNOMEDCT_CORE|Hypoalbuminemia|Hypoalbuminemia
C0239981|T047|OF|119247004|SNOMEDCT_CORE|Hypoalbuminemia|Hypoalbuminemia
C0239981|T047|FN|119247004|SNOMEDCT_CORE|Hypoalbuminemia|Hypoalbuminemia
C0239981|T047|SY|119247004|SNOMEDCT_CORE|Serum albumin low|Hypoalbuminemia
C0239997|T033|PT|288252009|SNOMEDCT_CORE|Maternal infection|Maternal infection
C0239997|T033|OF|288252009|SNOMEDCT_CORE|Maternal infection|Maternal infection
C0239997|T033|FN|288252009|SNOMEDCT_CORE|Maternal infection|Maternal infection
C0240007|T184|SY|281398003|SNOMEDCT_CORE|Groin lump|Groin mass
C0240007|T184|OF|281398003|SNOMEDCT_CORE|Groin lump|Groin mass
C0240007|T184|PT|281398003|SNOMEDCT_CORE|Groin mass|Groin mass
C0240007|T184|FN|281398003|SNOMEDCT_CORE|Groin mass|Groin mass
C0240007|T184|SY|281398003|SNOMEDCT_CORE|Mass of inguinal region|Groin mass
C0240066|T047|PT|35240004|SNOMEDCT_CORE|Iron deficiency|Iron deficiency
C0240066|T047|FN|35240004|SNOMEDCT_CORE|Iron deficiency|Iron deficiency
C0240066|T047|IS|35240004|SNOMEDCT_CORE|Iron deficiency, NOS|Iron deficiency
C0240111|T047|PT|371081002|SNOMEDCT_CORE|Arthritis of knee|Arthritis of knee
C0240111|T047|FN|371081002|SNOMEDCT_CORE|Arthritis of knee|Arthritis of knee
C0240129|T184|PT|249913002|SNOMEDCT_CORE|Knee stiff|Knee stiff
C0240129|T184|FN|249913002|SNOMEDCT_CORE|Knee stiff|Knee stiff
C0240140|T033|PT|248866005|SNOMEDCT_CORE|Labial adhesions|Labial adhesions
C0240140|T033|FN|248866005|SNOMEDCT_CORE|Labial adhesions|Labial adhesions
C0240225|T047|PT|300332007|SNOMEDCT_CORE|Liver mass|Liver mass
C0240225|T047|FN|300332007|SNOMEDCT_CORE|Liver mass|Liver mass
C0240318|T033|SY|94147001|SNOMEDCT_CORE|Mass of mediastinum|Mediastinal mass
C0240318|T033|FN|94147001|SNOMEDCT_CORE|Mass of mediastinum|Mediastinal mass
C0240318|T033|PT|94147001|SNOMEDCT_CORE|Mediastinal mass|Mediastinal mass
C0240318|T033|OF|94147001|SNOMEDCT_CORE|Mediastinal mass|Mediastinal mass
C0240318|T033|IS|94147001|SNOMEDCT_CORE|Mediastinal mass, NOS|Mediastinal mass
C0240557|T184|SY|70076002|SNOMEDCT_CORE|Irritation of nose|Irritation of nose
C0240596|T033|PT|247824007|SNOMEDCT_CORE|Fear of becoming fat|Fear of becoming fat
C0240596|T033|FN|247824007|SNOMEDCT_CORE|Fear of becoming fat|Fear of becoming fat
C0240596|T033|SY|247824007|SNOMEDCT_CORE|Fear of obesity|Fear of becoming fat
C0240611|T033|PT|289922002|SNOMEDCT_CORE|Mass of ovary|Mass of ovary
C0240611|T033|FN|289922002|SNOMEDCT_CORE|Mass of ovary|Mass of ovary
C0240611|T033|SY|289922002|SNOMEDCT_CORE|Ovarian mass|Mass of ovary
C0240671|T033|FN|409675001|SNOMEDCT_CORE|Partial thromboplastin time increased|Partial thromboplastin time increased
C0240671|T033|PT|409675001|SNOMEDCT_CORE|Partial thromboplastin time increased|Partial thromboplastin time increased
C0240717|T184|PT|225565007|SNOMEDCT_CORE|Perineal pain|Perineal pain
C0240717|T184|FN|225565007|SNOMEDCT_CORE|Perineal pain|Perineal pain
C0240735|T048|PT|192073007|SNOMEDCT_CORE|Change in personality|Change in personality
C0240735|T048|FN|192073007|SNOMEDCT_CORE|Change in personality|Change in personality
C0240873|T033|SY|248523006|SNOMEDCT_CORE|Rectal lump|Rectal mass
C0240873|T033|PT|248523006|SNOMEDCT_CORE|Rectal mass|Rectal mass
C0240873|T033|FN|248523006|SNOMEDCT_CORE|Rectal mass|Rectal mass
C0240937|T037|PT|274166008|SNOMEDCT_CORE|Scalp laceration|Scalp laceration
C0240937|T037|FN|274166008|SNOMEDCT_CORE|Scalp laceration|Scalp laceration
C0240941|T184|PT|277799005|SNOMEDCT_CORE|Pruritus of scalp|Pruritus of scalp
C0240941|T184|SY|277799005|SNOMEDCT_CORE|Scalp pruritus|Pruritus of scalp
C0240941|T184|FN|277799005|SNOMEDCT_CORE|Scalp pruritus|Pruritus of scalp
C0240941|T184|OF|277799005|SNOMEDCT_CORE|Scalp pruritus|Pruritus of scalp
C0240991|T184|PT|445458007|SNOMEDCT_CORE|Sensory ataxia|Sensory ataxia
C0240991|T184|FN|445458007|SNOMEDCT_CORE|Sensory ataxia|Sensory ataxia
C0241042|T184|PT|249918006|SNOMEDCT_CORE|Shoulder stiff|Shoulder stiff
C0241042|T184|FN|249918006|SNOMEDCT_CORE|Shoulder stiff|Shoulder stiff
C0241057|T184|IS|102604002|SNOMEDCT_CORE|Burning sensation of skin|Burning sensation of skin
C0241057|T184|OAP|102604002|SNOMEDCT_CORE|Sensation of burning of skin|Burning sensation of skin
C0241057|T184|OAF|102604002|SNOMEDCT_CORE|Sensation of burning of skin|Burning sensation of skin
C0241069|T047|FN|93448009|SNOMEDCT_CORE|Superficial ulcer of skin|Superficial ulcer of skin
C0241069|T047|PT|93448009|SNOMEDCT_CORE|Superficial ulcer of skin|Superficial ulcer of skin
C0241157|T033|SY|271760008|SNOMEDCT_CORE|Pussey spot|Pustule
C0241157|T033|PT|271760008|SNOMEDCT_CORE|Pustule|Pustule
C0241157|T033|FN|271760008|SNOMEDCT_CORE|Pustule|Pustule
C0241158|T033|SY|70582006|SNOMEDCT_CORE|Cicatrix of skin|Scar of skin
C0241158|T033|IS|70582006|SNOMEDCT_CORE|Cicatrix of skin, NOS|Scar of skin
C0241158|T033|PT|70582006|SNOMEDCT_CORE|Scar of skin|Scar of skin
C0241158|T033|FN|70582006|SNOMEDCT_CORE|Scar of skin|Scar of skin
C0241158|T033|IS|70582006|SNOMEDCT_CORE|Scar of skin, NOS|Scar of skin
C0241210|T048|SY|229721007|SNOMEDCT_CORE|Slow to talk|Speech delay
C0241210|T048|PT|229721007|SNOMEDCT_CORE|Speech delay|Speech delay
C0241210|T048|FN|229721007|SNOMEDCT_CORE|Speech delay|Speech delay
C0241310|T184|SY|162053006|SNOMEDCT_CORE|Hypogastric pain|Suprapubic pain
C0241310|T184|SY|162053006|SNOMEDCT_CORE|Pain of hypogastrium|Suprapubic pain
C0241310|T184|PT|162053006|SNOMEDCT_CORE|Suprapubic pain|Suprapubic pain
C0241310|T184|FN|162053006|SNOMEDCT_CORE|Suprapubic pain|Suprapubic pain
C0241353|T033|SY|87860000|SNOMEDCT_CORE|Lump in testis|Testicular mass
C0241353|T033|SY|87860000|SNOMEDCT_CORE|Mass of testicle|Testicular mass
C0241353|T033|FN|87860000|SNOMEDCT_CORE|Mass of testicle|Testicular mass
C0241353|T033|SY|87860000|SNOMEDCT_CORE|Mass of testis|Testicular mass
C0241353|T033|SY|87860000|SNOMEDCT_CORE|Testicular lump|Testicular mass
C0241353|T033|IS|87860000|SNOMEDCT_CORE|Testicular lump, NOS|Testicular mass
C0241353|T033|PT|87860000|SNOMEDCT_CORE|Testicular mass|Testicular mass
C0241353|T033|OF|87860000|SNOMEDCT_CORE|Testicular mass|Testicular mass
C0241353|T033|IS|87860000|SNOMEDCT_CORE|Testicular mass, NOS|Testicular mass
C0241374|T184|IS|78514002|SNOMEDCT_CORE|Meralgia|Thigh pain
C0241374|T184|FN|78514002|SNOMEDCT_CORE|Thigh pain|Thigh pain
C0241374|T184|PT|78514002|SNOMEDCT_CORE|Thigh pain|Thigh pain
C0241394|T184|PT|300955002|SNOMEDCT_CORE|Pain in thumb|Pain in thumb
C0241394|T184|FN|300955002|SNOMEDCT_CORE|Pain in thumb|Pain in thumb
C0241407|T037|FN|95898004|SNOMEDCT_CORE|Tick bite|Tick bite
C0241407|T037|PT|95898004|SNOMEDCT_CORE|Tick bite|Tick bite
C0241407|T037|IS|95898004|SNOMEDCT_CORE|Tick bite, NOS|Tick bite
C0241416|T184|PT|285365001|SNOMEDCT_CORE|Pain in toe|Pain in toe
C0241416|T184|FN|285365001|SNOMEDCT_CORE|Pain in toe|Pain in toe
C0241416|T184|SY|285365001|SNOMEDCT_CORE|Toe pain|Pain in toe
C0241426|T047|SY|399044006|SNOMEDCT_CORE|Burning tongue|Glossopyrosis
C0241426|T047|PT|399044006|SNOMEDCT_CORE|Glossopyrosis|Glossopyrosis
C0241426|T047|FN|399044006|SNOMEDCT_CORE|Glossopyrosis|Glossopyrosis
C0241436|T033|PT|441975003|SNOMEDCT_CORE|Mass of tongue|Mass of tongue
C0241436|T033|FN|441975003|SNOMEDCT_CORE|Mass of tongue|Mass of tongue
C0241558|T046|PTGB|405555006|SNOMEDCT_CORE|Haemorrhage of urethra|Hemorrhage of urethra
C0241558|T046|PT|405555006|SNOMEDCT_CORE|Hemorrhage of urethra|Hemorrhage of urethra
C0241558|T046|FN|405555006|SNOMEDCT_CORE|Hemorrhage of urethra|Hemorrhage of urethra
C0241616|T047|PT|297147009|SNOMEDCT_CORE|Atrophy of vagina|Atrophy of vagina
C0241616|T047|FN|297147009|SNOMEDCT_CORE|Atrophy of vagina|Atrophy of vagina
C0241619|T033|PT|24548005|SNOMEDCT_CORE|Cyst of vagina|Cyst of vagina
C0241619|T033|FN|24548005|SNOMEDCT_CORE|Cyst of vagina|Cyst of vagina
C0241619|T033|SY|24548005|SNOMEDCT_CORE|Vaginal cyst|Cyst of vagina
C0241633|T033|IS|31908003|SNOMEDCT_CORE|Dryness of vagina|Vaginal dryness
C0241633|T033|PT|31908003|SNOMEDCT_CORE|Vaginal dryness|Vaginal dryness
C0241633|T033|FN|31908003|SNOMEDCT_CORE|Vaginal dryness|Vaginal dryness
C0241716|T033|PT|289477004|SNOMEDCT_CORE|Mass of vulva|Mass of vulva
C0241716|T033|FN|289477004|SNOMEDCT_CORE|Mass of vulva|Mass of vulva
C0241745|T184|PT|298012000|SNOMEDCT_CORE|Wound pain|Wound pain
C0241745|T184|FN|298012000|SNOMEDCT_CORE|Wound pain|Wound pain
C0241880|T047|PT|26681001|SNOMEDCT_CORE|Endometriosis of pelvis|Endometriosis of pelvis
C0241880|T047|FN|26681001|SNOMEDCT_CORE|Endometriosis of pelvis|Endometriosis of pelvis
C0241880|T047|IS|26681001|SNOMEDCT_CORE|Endometriosis of pelvis, NOS|Endometriosis of pelvis
C0241880|T047|SY|26681001|SNOMEDCT_CORE|Pelvic endometriosis|Endometriosis of pelvis
C0241880|T047|IS|26681001|SNOMEDCT_CORE|Pelvic endometriosis, NOS|Endometriosis of pelvis
C0241910|T047|SY|197284004|SNOMEDCT_CORE|Autoimmune chronic active hepatitis|Autoimmune chronic active hepatitis
C0241910|T047|IS|197284004|SNOMEDCT_CORE|Autoimmune hepatitis|Autoimmune chronic active hepatitis
C0241961|T191|PT|254921004|SNOMEDCT_CORE|Angiomyolipoma of kidney|Angiomyolipoma of kidney
C0241961|T191|FN|254921004|SNOMEDCT_CORE|Angiomyolipoma of kidney|Angiomyolipoma of kidney
C0241961|T191|SY|254921004|SNOMEDCT_CORE|Hamartoma of kidney|Angiomyolipoma of kidney
C0241981|T033|SY|387603000|SNOMEDCT_CORE|Balance impairment|Impairment of balance
C0241981|T033|PT|387603000|SNOMEDCT_CORE|Impairment of balance|Impairment of balance
C0241981|T033|FN|387603000|SNOMEDCT_CORE|Impairment of balance|Impairment of balance
C0241981|T033|SY|282299006|SNOMEDCT_CORE|Loss of balance|Impairment of balance
C0241981|T033|SY|387603000|SNOMEDCT_CORE|Problem with balance|Impairment of balance
C0241981|T033|PT|282299006|SNOMEDCT_CORE|Unable to balance|Impairment of balance
C0241981|T033|FN|282299006|SNOMEDCT_CORE|Unable to balance|Impairment of balance
C0242073|T047|PT|67599009|SNOMEDCT_CORE|Pulmonary congestion|Pulmonary congestion
C0242073|T047|FN|67599009|SNOMEDCT_CORE|Pulmonary congestion|Pulmonary congestion
C0242073|T047|IS|67599009|SNOMEDCT_CORE|Pulmonary congestion, NOS|Pulmonary congestion
C0242084|T047|PT|233983001|SNOMEDCT_CORE|Ruptured cerebral aneurysm|Ruptured cerebral aneurysm
C0242084|T047|FN|233983001|SNOMEDCT_CORE|Ruptured cerebral aneurysm|Ruptured cerebral aneurysm
C0242129|T047|PT|371040005|SNOMEDCT_CORE|Thrombotic stroke|Thrombotic stroke
C0242129|T047|FN|371040005|SNOMEDCT_CORE|Thrombotic stroke|Thrombotic stroke
C0242147|T047|PT|431309003|SNOMEDCT_CORE|Acute urinary tract infection|Acute urinary tract infection
C0242147|T047|FN|431309003|SNOMEDCT_CORE|Acute urinary tract infection|Acute urinary tract infection
C0242147|T047|SY|431309003|SNOMEDCT_CORE|Acute UTI|Acute urinary tract infection
C0242147|T047|SY|431309003|SNOMEDCT_CORE|Urinary tract infection of sudden onset AND/OR short duration|Acute urinary tract infection
C0242172|T047|SY|198130006|SNOMEDCT_CORE|Female pelvic inflammation|Female pelvic inflammatory disease
C0242172|T047|PT|198130006|SNOMEDCT_CORE|Female pelvic inflammatory disease|Female pelvic inflammatory disease
C0242172|T047|FN|198130006|SNOMEDCT_CORE|Female pelvic inflammatory disease|Female pelvic inflammatory disease
C0242172|T047|IS|198130006|SNOMEDCT_CORE|Inflammatory disease of female pelvic organs AND/OR tissues|Female pelvic inflammatory disease
C0242172|T047|SY|198130006|SNOMEDCT_CORE|Pelvic inflammatory disease|Female pelvic inflammatory disease
C0242172|T047|IS|198130006|SNOMEDCT_CORE|PID|Female pelvic inflammatory disease
C0242172|T047|SY|198130006|SNOMEDCT_CORE|PID - pelvic inflammatory disease|Female pelvic inflammatory disease
C0242184|T046|SY|389086002|SNOMEDCT_CORE|Decreased oxygen supply|Hypoxia
C0242184|T046|PT|389086002|SNOMEDCT_CORE|Hypoxia|Hypoxia
C0242184|T046|FN|389086002|SNOMEDCT_CORE|Hypoxia|Hypoxia
C0242184|T046|SY|389086002|SNOMEDCT_CORE|Hypoxic|Hypoxia
C0242301|T047|SY|416675009|SNOMEDCT_CORE|Boil|Furuncle
C0242301|T047|PT|416675009|SNOMEDCT_CORE|Furuncle|Furuncle
C0242301|T047|FN|416675009|SNOMEDCT_CORE|Furuncle|Furuncle
C0242339|T047|PTGB|370992007|SNOMEDCT_CORE|Dyslipidaemia|Dyslipidemia
C0242339|T047|PT|370992007|SNOMEDCT_CORE|Dyslipidemia|Dyslipidemia
C0242339|T047|FN|370992007|SNOMEDCT_CORE|Dyslipidemia|Dyslipidemia
C0242339|T047|SY|370992007|SNOMEDCT_CORE|High blood cholesterol/triglycerides|Dyslipidemia
C0242342|T047|SY|32390006|SNOMEDCT_CORE|Simmond's disease|Simmonds' disease
C0242342|T047|IS|32390006|SNOMEDCT_CORE|Simmonds disease|Simmonds' disease
C0242342|T047|SY|32390006|SNOMEDCT_CORE|Simmonds' disease|Simmonds' disease
C0242343|T047|SY|32390006|SNOMEDCT_CORE|Deficient secretion of all pituitary hormones|Panhypopituitarism
C0242343|T047|PT|32390006|SNOMEDCT_CORE|Panhypopituitarism|Panhypopituitarism
C0242343|T047|FN|32390006|SNOMEDCT_CORE|Panhypopituitarism|Panhypopituitarism
C0242343|T047|IS|32390006|SNOMEDCT_CORE|Panhypopituitarism, NOS|Panhypopituitarism
C0242343|T047|SY|32390006|SNOMEDCT_CORE|Primary hypopituitarism|Panhypopituitarism
C0242350|T047|SY|397803000|SNOMEDCT_CORE|Erectile dysfunction|Impotence
C0242350|T047|OAS|398175007|SNOMEDCT_CORE|Erectile dysfunction|Impotence
C0242350|T047|SY|397803000|SNOMEDCT_CORE|Failure of erection|Impotence
C0242350|T047|PT|397803000|SNOMEDCT_CORE|Impotence|Impotence
C0242350|T047|FN|397803000|SNOMEDCT_CORE|Impotence|Impotence
C0242350|T047|OAP|398175007|SNOMEDCT_CORE|Male erectile disorder|Impotence
C0242350|T047|OAF|398175007|SNOMEDCT_CORE|Male erectile disorder|Impotence
C0242350|T047|SY|397803000|SNOMEDCT_CORE|Sexual impotence|Impotence
C0242362|T020|IS|73589001|SNOMEDCT_CORE|Herniation of anulus fibrosus|Intervertebral disc prolapse
C0242362|T020|IS|73589001|SNOMEDCT_CORE|Herniation of intervertebral disc|Intervertebral disc prolapse
C0242362|T020|SY|73589001|SNOMEDCT_CORE|Intervertebral disc extrusion|Intervertebral disc prolapse
C0242362|T020|PT|73589001|SNOMEDCT_CORE|Intervertebral disc prolapse|Intervertebral disc prolapse
C0242362|T020|FN|73589001|SNOMEDCT_CORE|Intervertebral disc prolapse|Intervertebral disc prolapse
C0242362|T020|SY|73589001|SNOMEDCT_CORE|Intervertebral disc protrusion|Intervertebral disc prolapse
C0242362|T020|SY|73589001|SNOMEDCT_CORE|IVDP - Intervertebral disc prolapse|Intervertebral disc prolapse
C0242362|T020|SY|73589001|SNOMEDCT_CORE|PID - Prolapsed intervertebral disc|Intervertebral disc prolapse
C0242362|T020|SY|73589001|SNOMEDCT_CORE|PIVD - Prolapsed intervertebral disc|Intervertebral disc prolapse
C0242362|T020|SY|73589001|SNOMEDCT_CORE|Prolapsed intervertebral disc|Intervertebral disc prolapse
C0242362|T020|SY|73589001|SNOMEDCT_CORE|Slipped disc|Intervertebral disc prolapse
C0242362|T020|SY|73589001|SNOMEDCT_CORE|Slipped intervertebral disc|Intervertebral disc prolapse
C0242379|T191|SY|363358000|SNOMEDCT_CORE|CA - Lung cancer|Malignant tumor of lung
C0242379|T191|IS|93880001|SNOMEDCT_CORE|Malignant neoplasm of lung|Malignant tumor of lung
C0242379|T191|IS|93880001|SNOMEDCT_CORE|Malignant neoplasm of lung, NOS|Malignant tumor of lung
C0242379|T191|PT|363358000|SNOMEDCT_CORE|Malignant tumor of lung|Malignant tumor of lung
C0242379|T191|FN|363358000|SNOMEDCT_CORE|Malignant tumor of lung|Malignant tumor of lung
C0242379|T191|PTGB|363358000|SNOMEDCT_CORE|Malignant tumour of lung|Malignant tumor of lung
C0242383|T047|SY|267718000|SNOMEDCT_CORE|AAMD - Age related macular degeneration|Age related macular degeneration
C0242383|T047|PT|267718000|SNOMEDCT_CORE|Age related macular degeneration|Age related macular degeneration
C0242383|T047|SY|267718000|SNOMEDCT_CORE|Age-related macular degeneration|Age related macular degeneration
C0242383|T047|FN|267718000|SNOMEDCT_CORE|Age-related macular degeneration|Age related macular degeneration
C0242383|T047|SY|267718000|SNOMEDCT_CORE|AMD - Age-related macular degeneration|Age related macular degeneration
C0242383|T047|SY|267718000|SNOMEDCT_CORE|ARMD - Age-related macular degeneration|Age related macular degeneration
C0242383|T047|SY|267718000|SNOMEDCT_CORE|Senile macular degeneration|Age related macular degeneration
C0242383|T047|SY|267718000|SNOMEDCT_CORE|Senile macular retinal degeneration|Age related macular degeneration
C0242383|T047|SY|267718000|SNOMEDCT_CORE|SMD - Senile macular degeneration|Age related macular degeneration
C0242420|T046|PT|6141006|SNOMEDCT_CORE|Retinal edema|Retinal edema
C0242420|T046|FN|6141006|SNOMEDCT_CORE|Retinal edema|Retinal edema
C0242420|T046|IS|6141006|SNOMEDCT_CORE|Retinal edema, NOS|Retinal edema
C0242420|T046|PTGB|6141006|SNOMEDCT_CORE|Retinal oedema|Retinal edema
C0242422|T047|PT|32798002|SNOMEDCT_CORE|Parkinsonism|Parkinsonism
C0242422|T047|FN|32798002|SNOMEDCT_CORE|Parkinsonism|Parkinsonism
C0242422|T047|IS|32798002|SNOMEDCT_CORE|Parkinsonism, NOS|Parkinsonism
C0242429|T184|PT|267102003|SNOMEDCT_CORE|Sore throat symptom|Sore throat symptom
C0242429|T184|FN|267102003|SNOMEDCT_CORE|Sore throat symptom|Sore throat symptom
C0242453|T184|PT|11441004|SNOMEDCT_CORE|Prostatism|Prostatism
C0242453|T184|FN|11441004|SNOMEDCT_CORE|Prostatism|Prostatism
C0242453|T184|IS|11441004|SNOMEDCT_CORE|Prostatism, NOS|Prostatism
C0242520|T047|IS|66944004|SNOMEDCT_CORE|Chronic thyroiditis, NOS|Chronic thyroiditis, NOS
C0242528|T047|PTGB|445009001|SNOMEDCT_CORE|Azotaemia|Azotemia
C0242528|T047|PT|445009001|SNOMEDCT_CORE|Azotemia|Azotemia
C0242528|T047|FN|445009001|SNOMEDCT_CORE|Azotemia|Azotemia
C0242584|T047|IS|2897005|SNOMEDCT_CORE|Auto-immune thrombocytopenia|Auto-immune thrombocytopenia
C0242647|T191|SY|277622004|SNOMEDCT_CORE|Maltoma|Mucosa-associated lymphoma
C0242647|T191|PT|277622004|SNOMEDCT_CORE|Mucosa-associated lymphoma|Mucosa-associated lymphoma
C0242647|T191|FN|277622004|SNOMEDCT_CORE|Mucosa-associated lymphoma|Mucosa-associated lymphoma
C0242666|T047|SY|1563006|SNOMEDCT_CORE|Protein S deficiency|Protein S deficiency disease
C0242666|T047|PT|1563006|SNOMEDCT_CORE|Protein S deficiency disease|Protein S deficiency disease
C0242666|T047|FN|1563006|SNOMEDCT_CORE|Protein S deficiency disease|Protein S deficiency disease
C0242669|T047|PT|109894007|SNOMEDCT_CORE|Retained placenta|Retained placenta
C0242669|T047|FN|109894007|SNOMEDCT_CORE|Retained placenta|Retained placenta
C0242770|T047|IS|129458007|SNOMEDCT_CORE|BOOP|Cryptogenic organizing pneumonia
C0242770|T047|IS|129458007|SNOMEDCT_CORE|BOOP - Bronchiolitis obliterans and organising pneumonitis|Cryptogenic organizing pneumonia
C0242770|T047|IS|129458007|SNOMEDCT_CORE|BOOP - Bronchiolitis obliterans and organizing pneumonitis|Cryptogenic organizing pneumonia
C0242770|T047|OAS|129458007|SNOMEDCT_CORE|BOOP - Bronchiolitis obliterans organising pneumonia|Cryptogenic organizing pneumonia
C0242770|T047|SYGB|719218000|SNOMEDCT_CORE|BOOP - Bronchiolitis obliterans organising pneumonia|Cryptogenic organizing pneumonia
C0242770|T047|OAS|129458007|SNOMEDCT_CORE|BOOP - Bronchiolitis obliterans organizing pneumonia|Cryptogenic organizing pneumonia
C0242770|T047|SY|719218000|SNOMEDCT_CORE|BOOP - Bronchiolitis obliterans organizing pneumonia|Cryptogenic organizing pneumonia
C0242770|T047|IS|129458007|SNOMEDCT_CORE|Bronchiolitis obliterans and organising pneumonitis|Cryptogenic organizing pneumonia
C0242770|T047|IS|129458007|SNOMEDCT_CORE|Bronchiolitis obliterans and organizing pneumonitis|Cryptogenic organizing pneumonia
C0242770|T047|OAP|129458007|SNOMEDCT_CORE|Bronchiolitis obliterans organising pneumonia|Cryptogenic organizing pneumonia
C0242770|T047|SYGB|719218000|SNOMEDCT_CORE|Bronchiolitis obliterans organising pneumonia|Cryptogenic organizing pneumonia
C0242770|T047|OAP|129458007|SNOMEDCT_CORE|Bronchiolitis obliterans organizing pneumonia|Cryptogenic organizing pneumonia
C0242770|T047|SY|719218000|SNOMEDCT_CORE|Bronchiolitis obliterans organizing pneumonia|Cryptogenic organizing pneumonia
C0242770|T047|OAF|129458007|SNOMEDCT_CORE|Bronchiolitis obliterans organizing pneumonia|Cryptogenic organizing pneumonia
C0242770|T047|OAS|129458007|SNOMEDCT_CORE|Bronchiolitis obliterans with organising pneumonia|Cryptogenic organizing pneumonia
C0242770|T047|OAS|129458007|SNOMEDCT_CORE|Bronchiolitis obliterans with organizing pneumonia|Cryptogenic organizing pneumonia
C0242770|T047|SY|719218000|SNOMEDCT_CORE|Bronchiolitis obliterans with usual interstitial pneumonitis|Cryptogenic organizing pneumonia
C0242770|T047|IS|129458007|SNOMEDCT_CORE|COP - Cryptogenic organising pneumonitis|Cryptogenic organizing pneumonia
C0242770|T047|SYGB|719218000|SNOMEDCT_CORE|COP - Cryptogenic organising pneumonitis|Cryptogenic organizing pneumonia
C0242770|T047|IS|129458007|SNOMEDCT_CORE|COP - Cryptogenic organizing pneumonitis|Cryptogenic organizing pneumonia
C0242770|T047|SY|719218000|SNOMEDCT_CORE|COP - Cryptogenic organizing pneumonitis|Cryptogenic organizing pneumonia
C0242770|T047|IS|129458007|SNOMEDCT_CORE|Cryptogenic organising pneumonia|Cryptogenic organizing pneumonia
C0242770|T047|PTGB|719218000|SNOMEDCT_CORE|Cryptogenic organising pneumonia|Cryptogenic organizing pneumonia
C0242770|T047|IS|129458007|SNOMEDCT_CORE|Cryptogenic organising pneumonitis|Cryptogenic organizing pneumonia
C0242770|T047|IS|129458007|SNOMEDCT_CORE|Cryptogenic organizing pneumonia|Cryptogenic organizing pneumonia
C0242770|T047|PT|719218000|SNOMEDCT_CORE|Cryptogenic organizing pneumonia|Cryptogenic organizing pneumonia
C0242770|T047|FN|719218000|SNOMEDCT_CORE|Cryptogenic organizing pneumonia|Cryptogenic organizing pneumonia
C0242770|T047|IS|129458007|SNOMEDCT_CORE|Cryptogenic organizing pneumonitis|Cryptogenic organizing pneumonia
C0242786|T046|PT|47200007|SNOMEDCT_CORE|High risk pregnancy|High risk pregnancy
C0242786|T046|FN|47200007|SNOMEDCT_CORE|High risk pregnancy|High risk pregnancy
C0242786|T046|SY|47200007|SNOMEDCT_CORE|HRP - High risk pregnancy|High risk pregnancy
C0242855|T047|PT|204342004|SNOMEDCT_CORE|Congenital atresia of pulmonary valve|Congenital atresia of pulmonary valve
C0242855|T047|SY|204342004|SNOMEDCT_CORE|Congenital atresia of the pulmonary valve|Congenital atresia of pulmonary valve
C0242855|T047|FN|204342004|SNOMEDCT_CORE|Congenital atresia of the pulmonary valve|Congenital atresia of pulmonary valve
C0243001|T047|PT|75100008|SNOMEDCT_CORE|Abdominal abscess|Abdominal abscess
C0243001|T047|FN|75100008|SNOMEDCT_CORE|Abdominal abscess|Abdominal abscess
C0243001|T047|IS|75100008|SNOMEDCT_CORE|Abdominal abscess, NOS|Abdominal abscess
C0243001|T047|SY|75100008|SNOMEDCT_CORE|Intra-abdominal abscess|Abdominal abscess
C0243026|T047|PT|91302008|SNOMEDCT_CORE|Sepsis|Sepsis
C0243026|T047|FN|91302008|SNOMEDCT_CORE|Sepsis|Sepsis
C0243026|T047|IS|91302008|SNOMEDCT_CORE|Sepsis, NOS|Sepsis
C0243026|T047|SY|91302008|SNOMEDCT_CORE|Systemic infection|Sepsis
C0243026|T047|OF|91302008|SNOMEDCT_CORE|Systemic infection|Sepsis
C0243026|T047|IS|91302008|SNOMEDCT_CORE|Systemic infection, NOS|Sepsis
C0259749|T047|PT|277879009|SNOMEDCT_CORE|Autonomic neuropathy|Autonomic neuropathy
C0259749|T047|FN|277879009|SNOMEDCT_CORE|Autonomic neuropathy|Autonomic neuropathy
C0259765|T047|SY|20425006|SNOMEDCT_CORE|Labyrinthine vertigo|Labyrinthine vertigo
C0259768|T046|SY|225553008|SNOMEDCT_CORE|Burst wound|Wound dehiscence
C0259768|T046|PT|225553008|SNOMEDCT_CORE|Wound dehiscence|Wound dehiscence
C0259768|T046|FN|225553008|SNOMEDCT_CORE|Wound dehiscence|Wound dehiscence
C0259768|T046|SY|225553008|SNOMEDCT_CORE|Wound opened up|Wound dehiscence
C0259768|T046|SY|225553008|SNOMEDCT_CORE|Wound reopened - observation|Wound dehiscence
C0259768|T046|SY|225553008|SNOMEDCT_CORE|Wound rupture|Wound dehiscence
C0259769|T033|SY|18070006|SNOMEDCT_CORE|Inspissated cerumen|Inspissated cerumen
C0259770|T190|SY|419893006|SNOMEDCT_CORE|EIC - Epidermal inclusion cyst|Epidermal inclusion cyst
C0259770|T190|SY|419893006|SNOMEDCT_CORE|Epidermal inclusion cyst|Epidermal inclusion cyst
C0259770|T190|SY|419893006|SNOMEDCT_CORE|Inclusion cyst|Epidermal inclusion cyst
C0259781|T191|PTGB|254805008|SNOMEDCT_CORE|Compound naevus of skin|Compound nevus of skin
C0259781|T191|PT|254805008|SNOMEDCT_CORE|Compound nevus of skin|Compound nevus of skin
C0259781|T191|FN|254805008|SNOMEDCT_CORE|Compound nevus of skin|Compound nevus of skin
C0259783|T191|PT|443937008|SNOMEDCT_CORE|Mixed glioma|Mixed glioma
C0259783|T191|PT|22217002|SNOMEDCT_CORE|Mixed glioma|Mixed glioma
C0259783|T191|FN|22217002|SNOMEDCT_CORE|Mixed glioma|Mixed glioma
C0259783|T191|FN|443937008|SNOMEDCT_CORE|Mixed glioma|Mixed glioma
C0259795|T037|FN|73817000|SNOMEDCT_CORE|Enteritis caused by radiation|Enteritis due to radiation
C0259795|T037|SY|73817000|SNOMEDCT_CORE|Enteritis caused by radiation|Enteritis due to radiation
C0259795|T037|PT|73817000|SNOMEDCT_CORE|Enteritis due to radiation|Enteritis due to radiation
C0259795|T037|OF|73817000|SNOMEDCT_CORE|Enteritis due to radiation|Enteritis due to radiation
C0259795|T037|SY|73817000|SNOMEDCT_CORE|Radiation enteritis|Enteritis due to radiation
C0259795|T037|SY|73817000|SNOMEDCT_CORE|Radiation induced enteritis|Enteritis due to radiation
C0259797|T037|PT|217697000|SNOMEDCT_CORE|Dog bite|Dog bite
C0259797|T037|OF|217697000|SNOMEDCT_CORE|Dog bite|Dog bite
C0259797|T037|FN|217697000|SNOMEDCT_CORE|Dog bite|Dog bite
C0259799|T047|SY|42513006|SNOMEDCT_CORE|PK - Punctate keratitis|Superficial punctate keratitis
C0259799|T047|SY|42513006|SNOMEDCT_CORE|Punctate epithelial keratitis|Superficial punctate keratitis
C0259799|T047|IS|42513006|SNOMEDCT_CORE|Punctate epithelial keratoconjunctivitis|Superficial punctate keratitis
C0259799|T047|SY|42513006|SNOMEDCT_CORE|Punctate keratitis|Superficial punctate keratitis
C0259799|T047|FN|42513006|SNOMEDCT_CORE|Punctate keratitis|Superficial punctate keratitis
C0259799|T047|PT|42513006|SNOMEDCT_CORE|Superficial punctate keratitis|Superficial punctate keratitis
C0260334|T047|OAP|196032009|SNOMEDCT_CORE|Pneumonitis due to inhalation of food or vomitus|Pneumonitis due to inhalation of food or vomitus
C0260334|T047|OAF|196032009|SNOMEDCT_CORE|Pneumonitis due to inhalation of food or vomitus|Pneumonitis due to inhalation of food or vomitus
C0260506|T033|PT|429006005|SNOMEDCT_CORE|Family history of malignant neoplasm of gastrointestinal tract|Family history of malignant neoplasm of gastrointestinal tract
C0260506|T033|FN|429006005|SNOMEDCT_CORE|Family history of malignant neoplasm of gastrointestinal tract|Family history of malignant neoplasm of gastrointestinal tract
C0260515|T033|PT|275937001|SNOMEDCT_CORE|Family history of cancer|Family history of cancer
C0260515|T033|OF|275937001|SNOMEDCT_CORE|Family history of cancer|Family history of cancer
C0260515|T033|FN|275937001|SNOMEDCT_CORE|Family history of cancer|Family history of cancer
C0260515|T033|IS|275937001|SNOMEDCT_CORE|FH: Cancer - *|Family history of cancer
C0260515|T033|SY|275937001|SNOMEDCT_CORE|FH: Malignant disease|Family history of cancer
C0260662|T033|SY|128540005|SNOMEDCT_CORE|Auditory alteration|Hearing problem
C0260662|T033|SY|128540005|SNOMEDCT_CORE|Disorder of hearing|Hearing problem
C0260662|T033|PT|128540005|SNOMEDCT_CORE|Hearing disorder|Hearing problem
C0260662|T033|OF|128540005|SNOMEDCT_CORE|Hearing disorder|Hearing problem
C0260662|T033|FN|128540005|SNOMEDCT_CORE|Hearing disorder|Hearing problem
C0260662|T033|PT|300228004|SNOMEDCT_CORE|Hearing problem|Hearing problem
C0260662|T033|FN|300228004|SNOMEDCT_CORE|Hearing problem|Hearing problem
C0261200|T037|PT|386662004|SNOMEDCT_CORE|Pedal cycle accident|Pedal cycle accident
C0261200|T037|OF|386662004|SNOMEDCT_CORE|Pedal cycle accident|Pedal cycle accident
C0261200|T037|FN|386662004|SNOMEDCT_CORE|Pedal cycle accident|Pedal cycle accident
C0261503|T037|PT|420057003|SNOMEDCT_CORE|Accidental poisoning by carbon monoxide|Accidental poisoning by carbon monoxide
C0261503|T037|OF|420057003|SNOMEDCT_CORE|Accidental poisoning by carbon monoxide|Accidental poisoning by carbon monoxide
C0261503|T037|FN|420057003|SNOMEDCT_CORE|Accidental poisoning caused by carbon monoxide|Accidental poisoning by carbon monoxide
C0261503|T037|SY|420057003|SNOMEDCT_CORE|Accidental poisoning caused by carbon monoxide|Accidental poisoning by carbon monoxide
C0261695|T037|PT|217839002|SNOMEDCT_CORE|Accidentally struck by falling object|Accidentally struck by falling object
C0261695|T037|OF|217839002|SNOMEDCT_CORE|Accidentally struck by falling object|Accidentally struck by falling object
C0261695|T037|FN|217839002|SNOMEDCT_CORE|Accidentally struck by falling object|Accidentally struck by falling object
C0261712|T037|FN|269716005|SNOMEDCT_CORE|Accident caused by machinery|Accident caused by machinery
C0261712|T037|PT|269716005|SNOMEDCT_CORE|Accident caused by machinery|Accident caused by machinery
C0261712|T037|OF|269716005|SNOMEDCT_CORE|Accident caused by machinery|Accident caused by machinery
C0261713|T037|PT|218016007|SNOMEDCT_CORE|Accidents caused by cutting and piercing instruments or objects|Accidents caused by cutting and piercing instruments or objects
C0261713|T037|OF|218016007|SNOMEDCT_CORE|Accidents caused by cutting and piercing instruments or objects|Accidents caused by cutting and piercing instruments or objects
C0261713|T037|FN|218016007|SNOMEDCT_CORE|Accidents caused by cutting and piercing instruments or objects|Accidents caused by cutting and piercing instruments or objects
C0261717|T037|PT|218034006|SNOMEDCT_CORE|Accidents caused by knives, swords and daggers|Accidents caused by knives, swords and daggers
C0261717|T037|OF|218034006|SNOMEDCT_CORE|Accidents caused by knives, swords and daggers|Accidents caused by knives, swords and daggers
C0261717|T037|FN|218034006|SNOMEDCT_CORE|Accidents caused by knives, swords and daggers|Accidents caused by knives, swords and daggers
C0261736|T037|PT|218129009|SNOMEDCT_CORE|Accidents caused by hot substance or object, caustic or corrosive material and steam|Accidents caused by hot substance or object, caustic or corrosive material and steam
C0261736|T037|OF|218129009|SNOMEDCT_CORE|Accidents caused by hot substance or object, caustic or corrosive material and steam|Accidents caused by hot substance or object, caustic or corrosive material and steam
C0261736|T037|FN|218129009|SNOMEDCT_CORE|Accidents caused by hot substance or object, caustic or corrosive material and steam|Accidents caused by hot substance or object, caustic or corrosive material and steam
C0261737|T037|PT|218130004|SNOMEDCT_CORE|Accident caused by hot liquid and vapor, including steam|Accident caused by hot liquid and vapor, including steam
C0261737|T037|FN|218130004|SNOMEDCT_CORE|Accident caused by hot liquid and vapor, including steam|Accident caused by hot liquid and vapor, including steam
C0261737|T037|PTGB|218130004|SNOMEDCT_CORE|Accident caused by hot liquid and vapour, including steam|Accident caused by hot liquid and vapor, including steam
C0261737|T037|IS|218130004|SNOMEDCT_CORE|Accidents caused by hot liquids and vapours,including steam|Accident caused by hot liquid and vapor, including steam
C0261737|T037|OF|218130004|SNOMEDCT_CORE|Accidents caused by hot liquids and vapours,including steam|Accident caused by hot liquid and vapor, including steam
C0261740|T037|FN|218164000|SNOMEDCT_CORE|Accident caused by electric current|Accident caused by electric current
C0261740|T037|PT|218164000|SNOMEDCT_CORE|Accident caused by electric current|Accident caused by electric current
C0261740|T037|SY|218164000|SNOMEDCT_CORE|Accidents caused by electric current|Accident caused by electric current
C0261740|T037|OF|218164000|SNOMEDCT_CORE|Accidents caused by electric current|Accident caused by electric current
C0261751|T037|FN|218218000|SNOMEDCT_CORE|Overexertion and strenuous movements|Overexertion and strenuous movements
C0261751|T037|PT|218218000|SNOMEDCT_CORE|Overexertion and strenuous movements|Overexertion and strenuous movements
C0261751|T037|OF|218218000|SNOMEDCT_CORE|Overexertion and strenuous movements|Overexertion and strenuous movements
C0262027|T037|PT|219235009|SNOMEDCT_CORE|Assault by striking by blunt or thrown object|Assault by striking by blunt or thrown object
C0262027|T037|OF|219235009|SNOMEDCT_CORE|Assault by striking by blunt or thrown object|Assault by striking by blunt or thrown object
C0262027|T037|FN|219235009|SNOMEDCT_CORE|Assault by striking by blunt or thrown object|Assault by striking by blunt or thrown object
C0262174|T033|PT|300197009|SNOMEDCT_CORE|Ear problem|Ear problem
C0262174|T033|FN|300197009|SNOMEDCT_CORE|Ear problem|Ear problem
C0262365|T033|SY|168750009|SNOMEDCT_CORE|Abnormal mammogram|Mammography abnormal
C0262365|T033|PT|168750009|SNOMEDCT_CORE|Mammography abnormal|Mammography abnormal
C0262365|T033|FN|168750009|SNOMEDCT_CORE|Mammography abnormal|Mammography abnormal
C0262374|T033|IS|69914001|SNOMEDCT_CORE|Anal stenosis|Stricture of anus
C0262374|T033|SY|69914001|SNOMEDCT_CORE|Anal stricture|Stricture of anus
C0262374|T033|IS|69914001|SNOMEDCT_CORE|Stenosis of anus|Stricture of anus
C0262374|T033|PT|69914001|SNOMEDCT_CORE|Stricture of anus|Stricture of anus
C0262374|T033|FN|69914001|SNOMEDCT_CORE|Stricture of anus|Stricture of anus
C0262384|T184|PT|102589003|SNOMEDCT_CORE|Atypical chest pain|Atypical chest pain
C0262384|T184|FN|102589003|SNOMEDCT_CORE|Atypical chest pain|Atypical chest pain
C0262399|T047|PT|239961006|SNOMEDCT_CORE|Bursitis of shoulder|Bursitis of shoulder
C0262399|T047|FN|239961006|SNOMEDCT_CORE|Bursitis of shoulder|Bursitis of shoulder
C0262399|T047|SY|239961006|SNOMEDCT_CORE|Bursitis of shoulder region|Bursitis of shoulder
C0262401|T191|SY|254609000|SNOMEDCT_CORE|Ampullary carcinoma|Carcinoma of ampulla of Vater
C0262401|T191|PT|254609000|SNOMEDCT_CORE|Carcinoma of ampulla of Vater|Carcinoma of ampulla of Vater
C0262401|T191|FN|254609000|SNOMEDCT_CORE|Carcinoma of ampulla of Vater|Carcinoma of ampulla of Vater
C0262404|T047|PT|95646004|SNOMEDCT_CORE|Cerebellar degeneration|Cerebellar degeneration
C0262404|T047|FN|95646004|SNOMEDCT_CORE|Cerebellar degeneration|Cerebellar degeneration
C0262404|T047|IS|95646004|SNOMEDCT_CORE|Cerebellar degeneration, NOS|Cerebellar degeneration
C0262414|T037|PT|125606003|SNOMEDCT_CORE|Fracture of cervical spine|Fracture of cervical spine
C0262414|T037|FN|125606003|SNOMEDCT_CORE|Fracture of cervical spine|Fracture of cervical spine
C0262414|T037|SY|125606003|SNOMEDCT_CORE|Fracture of cervical vertebra|Fracture of cervical spine
C0262414|T037|SY|125606003|SNOMEDCT_CORE|Fracture of neck|Fracture of cervical spine
C0262421|T047|PT|197928006|SNOMEDCT_CORE|Chronic urinary tract infection|Chronic urinary tract infection
C0262421|T047|FN|197928006|SNOMEDCT_CORE|Chronic urinary tract infection|Chronic urinary tract infection
C0262431|T046|SY|42942008|SNOMEDCT_CORE|Compression fracture of spine|Compression fracture of vertebral column
C0262431|T046|IS|42942008|SNOMEDCT_CORE|Compression fracture of spine, NOS|Compression fracture of vertebral column
C0262431|T046|PT|42942008|SNOMEDCT_CORE|Compression fracture of vertebral column|Compression fracture of vertebral column
C0262431|T046|FN|42942008|SNOMEDCT_CORE|Compression fracture of vertebral column|Compression fracture of vertebral column
C0262431|T046|IS|42942008|SNOMEDCT_CORE|Compression fracture of vertebral column, NOS|Compression fracture of vertebral column
C0262489|T037|PT|428257007|SNOMEDCT_CORE|Fracture of tibial plateau|Fracture of tibial plateau
C0262489|T037|FN|428257007|SNOMEDCT_CORE|Fracture of tibial plateau|Fracture of tibial plateau
C0262493|T191|SY|197433003|SNOMEDCT_CORE|Gallbladder polyp|Polyp of gallbladder
C0262493|T191|PT|197433003|SNOMEDCT_CORE|Polyp of gallbladder|Polyp of gallbladder
C0262493|T191|FN|197433003|SNOMEDCT_CORE|Polyp of gallbladder|Polyp of gallbladder
C0262505|T033|FN|235871004|SNOMEDCT_CORE|Hepatitis B carrier|Hepatitis B carrier
C0262505|T033|PT|235871004|SNOMEDCT_CORE|Hepatitis B carrier|Hepatitis B carrier
C0262537|T020|PT|236022004|SNOMEDCT_CORE|Left inguinal hernia|Left inguinal hernia
C0262537|T020|FN|236022004|SNOMEDCT_CORE|Left inguinal hernia|Left inguinal hernia
C0262537|T020|SY|236022004|SNOMEDCT_CORE|LIH - Left inguinal hernia|Left inguinal hernia
C0262538|T037|SY|263134008|SNOMEDCT_CORE|Complete tear of ligament|Ligament rupture
C0262538|T037|PT|263134008|SNOMEDCT_CORE|Ligament rupture|Ligament rupture
C0262538|T037|FN|263134008|SNOMEDCT_CORE|Ligament rupture|Ligament rupture
C0262538|T037|SY|263134008|SNOMEDCT_CORE|Ligament tear|Ligament rupture
C0262541|T037|PT|300956001|SNOMEDCT_CORE|Low back strain|Low back strain
C0262541|T037|FN|300956001|SNOMEDCT_CORE|Low back strain|Low back strain
C0262541|T037|SY|300956001|SNOMEDCT_CORE|Lumbar strain|Low back strain
C0262544|T037|PT|125608002|SNOMEDCT_CORE|Fracture of lumbar spine|Fracture of lumbar spine
C0262544|T037|FN|125608002|SNOMEDCT_CORE|Fracture of lumbar spine|Fracture of lumbar spine
C0262544|T037|SY|125608002|SNOMEDCT_CORE|Fracture of lumbar vertebra|Fracture of lumbar spine
C0262573|T037|SY|360450007|SNOMEDCT_CORE|Cervical strain|Strain of neck muscle
C0262573|T037|IS|360450007|SNOMEDCT_CORE|Neck strain|Strain of neck muscle
C0262573|T037|PT|360450007|SNOMEDCT_CORE|Strain of neck muscle|Strain of neck muscle
C0262573|T037|FN|360450007|SNOMEDCT_CORE|Strain of neck muscle|Strain of neck muscle
C0262578|T184|PT|102549009|SNOMEDCT_CORE|Cramp in lower leg associated with rest|Cramp in lower leg associated with rest
C0262578|T184|FN|102549009|SNOMEDCT_CORE|Cramp in lower leg associated with rest|Cramp in lower leg associated with rest
C0262578|T184|SY|102549009|SNOMEDCT_CORE|Night cramps|Cramp in lower leg associated with rest
C0262578|T184|OF|102549009|SNOMEDCT_CORE|Night cramps|Cramp in lower leg associated with rest
C0262578|T184|SY|102549009|SNOMEDCT_CORE|Nocturnal lower leg cramp|Cramp in lower leg associated with rest
C0262578|T184|SY|102549009|SNOMEDCT_CORE|Recumbency cramps|Cramp in lower leg associated with rest
C0262578|T184|SY|102549009|SNOMEDCT_CORE|Sleep related lower leg cramp|Cramp in lower leg associated with rest
C0262587|T191|PT|128474007|SNOMEDCT_CORE|Parathyroid adenoma|Parathyroid adenoma
C0262587|T191|FN|128474007|SNOMEDCT_CORE|Parathyroid adenoma|Parathyroid adenoma
C0262595|T047|PT|201340008|SNOMEDCT_CORE|Pigmented skin lesion|Pigmented skin lesion
C0262595|T047|FN|201340008|SNOMEDCT_CORE|Pigmented skin lesion|Pigmented skin lesion
C0262611|T047|PT|767678008|SNOMEDCT_CORE|Recurrent left inguinal hernia|Recurrent left inguinal hernia
C0262611|T047|FN|767678008|SNOMEDCT_CORE|Recurrent left inguinal hernia|Recurrent left inguinal hernia
C0262613|T033|SY|309088003|SNOMEDCT_CORE|Kidney mass|Renal mass
C0262613|T033|PT|309088003|SNOMEDCT_CORE|Renal mass|Renal mass
C0262613|T033|FN|309088003|SNOMEDCT_CORE|Renal mass|Renal mass
C0262617|T020|PT|236021006|SNOMEDCT_CORE|Right inguinal hernia|Right inguinal hernia
C0262617|T020|FN|236021006|SNOMEDCT_CORE|Right inguinal hernia|Right inguinal hernia
C0262617|T020|SY|236021006|SNOMEDCT_CORE|RIH - Right inguinal hernia|Right inguinal hernia
C0262627|T046|PT|56021002|SNOMEDCT_CORE|Seroma|Seroma
C0262627|T046|FN|56021002|SNOMEDCT_CORE|Seroma|Seroma
C0262633|T047|OAP|202852009|SNOMEDCT_CORE|Shoulder tendinitis|Shoulder tendinitis
C0262633|T047|OAF|202852009|SNOMEDCT_CORE|Shoulder tendinitis|Shoulder tendinitis
C0262633|T047|OAS|202852009|SNOMEDCT_CORE|Shoulder tendonitis|Shoulder tendonitis
C0262649|T037|SY|262520005|SNOMEDCT_CORE|Injury of thumb|Thumb injury
C0262649|T037|PT|262520005|SNOMEDCT_CORE|Thumb injury|Thumb injury
C0262649|T037|FN|262520005|SNOMEDCT_CORE|Thumb injury|Thumb injury
C0262655|T047|PT|197927001|SNOMEDCT_CORE|Recurrent urinary tract infection|Recurrent urinary tract infection
C0262655|T047|FN|197927001|SNOMEDCT_CORE|Recurrent urinary tract infection|Recurrent urinary tract infection
C0262655|T047|SY|197927001|SNOMEDCT_CORE|Recurrent UTI - urinary tract infection|Recurrent urinary tract infection
C0262666|T047|PT|69430001|SNOMEDCT_CORE|Abscess of vulva|Abscess of vulva
C0262666|T047|FN|69430001|SNOMEDCT_CORE|Abscess of vulva|Abscess of vulva
C0262666|T047|SY|69430001|SNOMEDCT_CORE|Vulval abscess|Abscess of vulva
C0262666|T047|SY|69430001|SNOMEDCT_CORE|Vulvar abscess|Abscess of vulva
C0262985|T047|PT|238564003|SNOMEDCT_CORE|Psoriasiform eczema|Psoriasiform eczema
C0262985|T047|FN|238564003|SNOMEDCT_CORE|Psoriasiform eczema|Psoriasiform eczema
C0263097|T047|PT|200751004|SNOMEDCT_CORE|Abscess of face|Abscess of face
C0263097|T047|FN|200751004|SNOMEDCT_CORE|Abscess of face|Abscess of face
C0263109|T047|PT|301802001|SNOMEDCT_CORE|Loin abscess|Loin abscess
C0263109|T047|FN|301802001|SNOMEDCT_CORE|Loin abscess|Loin abscess
C0263115|T047|PT|13802001|SNOMEDCT_CORE|Abscess of axilla|Abscess of axilla
C0263115|T047|FN|13802001|SNOMEDCT_CORE|Abscess of axilla|Abscess of axilla
C0263118|T047|PT|64576003|SNOMEDCT_CORE|Abscess of buttock|Abscess of buttock
C0263118|T047|FN|64576003|SNOMEDCT_CORE|Abscess of buttock|Abscess of buttock
C0263118|T047|SY|64576003|SNOMEDCT_CORE|Abscess of gluteal region|Abscess of buttock
C0263118|T047|SY|64576003|SNOMEDCT_CORE|Gluteal abscess|Abscess of buttock
C0263132|T047|PT|27561001|SNOMEDCT_CORE|Cellulitis of finger|Cellulitis of finger
C0263132|T047|FN|27561001|SNOMEDCT_CORE|Cellulitis of finger|Cellulitis of finger
C0263132|T047|IS|27561001|SNOMEDCT_CORE|Cellulitis of finger, NOS|Cellulitis of finger
C0263134|T047|PT|70637004|SNOMEDCT_CORE|Cellulitis of toe|Cellulitis of toe
C0263134|T047|FN|70637004|SNOMEDCT_CORE|Cellulitis of toe|Cellulitis of toe
C0263134|T047|IS|70637004|SNOMEDCT_CORE|Cellulitis of toe, NOS|Cellulitis of toe
C0263135|T047|PT|388982007|SNOMEDCT_CORE|Onychia of toe|Onychia of toe
C0263135|T047|FN|388982007|SNOMEDCT_CORE|Onychia of toe|Onychia of toe
C0263136|T047|PT|200652002|SNOMEDCT_CORE|Cellulitis of face|Cellulitis of face
C0263136|T047|FN|200652002|SNOMEDCT_CORE|Cellulitis of face|Cellulitis of face
C0263140|T047|PT|37098000|SNOMEDCT_CORE|Cellulitis of external nose|Cellulitis of external nose
C0263140|T047|FN|37098000|SNOMEDCT_CORE|Cellulitis of external nose|Cellulitis of external nose
C0263144|T047|PT|46876003|SNOMEDCT_CORE|Cellulitis of trunk|Cellulitis of trunk
C0263144|T047|FN|46876003|SNOMEDCT_CORE|Cellulitis of trunk|Cellulitis of trunk
C0263144|T047|IS|46876003|SNOMEDCT_CORE|Cellulitis of trunk, NOS|Cellulitis of trunk
C0263145|T047|PT|59883002|SNOMEDCT_CORE|Cellulitis of abdominal wall|Cellulitis of abdominal wall
C0263145|T047|FN|59883002|SNOMEDCT_CORE|Cellulitis of abdominal wall|Cellulitis of abdominal wall
C0263153|T047|PT|38217004|SNOMEDCT_CORE|Cellulitis of upper arm|Cellulitis of upper arm
C0263153|T047|FN|38217004|SNOMEDCT_CORE|Cellulitis of upper arm|Cellulitis of upper arm
C0263158|T047|PT|44428005|SNOMEDCT_CORE|Cellulitis of buttock|Cellulitis of buttock
C0263158|T047|FN|44428005|SNOMEDCT_CORE|Cellulitis of buttock|Cellulitis of buttock
C0263158|T047|SY|44428005|SNOMEDCT_CORE|Cellulitis of gluteal region|Cellulitis of buttock
C0263159|T047|SY|287001000|SNOMEDCT_CORE|Cellulitis of leg, except foot|Cellulitis of leg, excluding foot
C0263159|T047|PT|287001000|SNOMEDCT_CORE|Cellulitis of leg, excluding foot|Cellulitis of leg, excluding foot
C0263159|T047|FN|287001000|SNOMEDCT_CORE|Cellulitis of leg, excluding foot|Cellulitis of leg, excluding foot
C0263162|T047|PT|13301002|SNOMEDCT_CORE|Cellulitis of knee|Cellulitis of knee
C0263162|T047|FN|13301002|SNOMEDCT_CORE|Cellulitis of knee|Cellulitis of knee
C0263218|T191|SY|39629007|SNOMEDCT_CORE|Granuloma telangiectaticum of skin|Pyogenic granuloma of skin
C0263218|T191|PT|39629007|SNOMEDCT_CORE|Pyogenic granuloma of skin|Pyogenic granuloma of skin
C0263218|T191|FN|39629007|SNOMEDCT_CORE|Pyogenic granuloma of skin|Pyogenic granuloma of skin
C0263218|T191|IS|39629007|SNOMEDCT_CORE|Suppurative granuloma of skin|Pyogenic granuloma of skin
C0263233|T047|PT|62742006|SNOMEDCT_CORE|Cradle cap|Cradle cap
C0263233|T047|FN|62742006|SNOMEDCT_CORE|Cradle cap|Cradle cap
C0263240|T047|PT|51221005|SNOMEDCT_CORE|Chronic contact dermatitis|Chronic contact dermatitis
C0263240|T047|FN|51221005|SNOMEDCT_CORE|Chronic contact dermatitis|Chronic contact dermatitis
C0263240|T047|IS|51221005|SNOMEDCT_CORE|Chronic contact dermatitis, NOS|Chronic contact dermatitis
C0263324|T047|SY|240302002|SNOMEDCT_CORE|Erythema neonatorum|Erythroderma neonatorum
C0263324|T047|SY|240302002|SNOMEDCT_CORE|Erythema toxicum neonatorum|Erythroderma neonatorum
C0263324|T047|PT|240302002|SNOMEDCT_CORE|Erythroderma neonatorum|Erythroderma neonatorum
C0263324|T047|FN|240302002|SNOMEDCT_CORE|Erythroderma neonatorum|Erythroderma neonatorum
C0263324|T047|SY|240302002|SNOMEDCT_CORE|ETN - Erythema toxicum neonatorum|Erythroderma neonatorum
C0263324|T047|SY|240302002|SNOMEDCT_CORE|Neonatal erythema toxicum|Erythroderma neonatorum
C0263324|T047|SY|240302002|SNOMEDCT_CORE|Toxic erythema of newborn|Erythroderma neonatorum
C0263324|T047|SY|240302002|SNOMEDCT_CORE|Toxic erythema of the newborn|Erythroderma neonatorum
C0263338|T047|PT|51611005|SNOMEDCT_CORE|Chronic urticaria|Chronic urticaria
C0263338|T047|FN|51611005|SNOMEDCT_CORE|Chronic urticaria|Chronic urticaria
C0263338|T047|SY|51611005|SNOMEDCT_CORE|Recurrent periodic urticaria|Chronic urticaria
C0263352|T047|SY|55608001|SNOMEDCT_CORE|Lichen urticatus|Prurigo simplex
C0263352|T047|SY|55608001|SNOMEDCT_CORE|Papular urticaria|Prurigo simplex
C0263352|T047|PT|55608001|SNOMEDCT_CORE|Prurigo simplex|Prurigo simplex
C0263352|T047|FN|55608001|SNOMEDCT_CORE|Prurigo simplex|Prurigo simplex
C0263352|T047|SY|55608001|SNOMEDCT_CORE|Strophulus|Prurigo simplex
C0263353|T047|SY|63501000|SNOMEDCT_CORE|Hyde's disease|Prurigo nodularis
C0263353|T047|SY|63501000|SNOMEDCT_CORE|Nodular prurigo|Prurigo nodularis
C0263353|T047|SY|63501000|SNOMEDCT_CORE|Picker's nodules|Prurigo nodularis
C0263353|T047|PT|63501000|SNOMEDCT_CORE|Prurigo nodularis|Prurigo nodularis
C0263353|T047|FN|63501000|SNOMEDCT_CORE|Prurigo nodularis|Prurigo nodularis
C0263383|T020|PT|5132005|SNOMEDCT_CORE|Keratosis pilaris|Keratosis pilaris
C0263383|T020|FN|5132005|SNOMEDCT_CORE|Keratosis pilaris|Keratosis pilaris
C0263383|T020|SY|5132005|SNOMEDCT_CORE|KP - Keratosis pilaris|Keratosis pilaris
C0263415|T037|SYGB|43982006|SNOMEDCT_CORE|Actinic ageing|Solar degeneration
C0263415|T037|SY|43982006|SNOMEDCT_CORE|Actinic aging|Solar degeneration
C0263415|T037|SY|43982006|SNOMEDCT_CORE|Actinic degeneration|Solar degeneration
C0263415|T037|SY|43982006|SNOMEDCT_CORE|Actinic degeneration of skin|Solar degeneration
C0263415|T037|SY|43982006|SNOMEDCT_CORE|Actinic elastosis|Solar degeneration
C0263415|T037|SY|43982006|SNOMEDCT_CORE|Dermatoheliosis|Solar degeneration
C0263415|T037|SY|43982006|SNOMEDCT_CORE|Farmer's skin|Solar degeneration
C0263415|T037|SYGB|43982006|SNOMEDCT_CORE|Photoageing|Solar degeneration
C0263415|T037|SY|43982006|SNOMEDCT_CORE|Photoaging|Solar degeneration
C0263415|T037|SY|43982006|SNOMEDCT_CORE|Sailor's skin|Solar degeneration
C0263415|T037|PT|43982006|SNOMEDCT_CORE|Solar degeneration|Solar degeneration
C0263415|T037|FN|43982006|SNOMEDCT_CORE|Solar degeneration|Solar degeneration
C0263415|T037|SY|43982006|SNOMEDCT_CORE|Solar elastosis|Solar degeneration
C0263415|T037|SY|43982006|SNOMEDCT_CORE|Sun damaged skin|Solar degeneration
C0263437|T047|SY|49706007|SNOMEDCT_CORE|Acne neonatorum|Neonatal acne
C0263437|T047|IS|49706007|SNOMEDCT_CORE|Infantile acne|Neonatal acne
C0263437|T047|PT|49706007|SNOMEDCT_CORE|Neonatal acne|Neonatal acne
C0263437|T047|FN|49706007|SNOMEDCT_CORE|Neonatal acne|Neonatal acne
C0263449|T047|PT|238751002|SNOMEDCT_CORE|Perioral dermatitis|Perioral dermatitis
C0263449|T047|FN|238751002|SNOMEDCT_CORE|Perioral dermatitis|Perioral dermatitis
C0263449|T047|SY|238751002|SNOMEDCT_CORE|POD - Perioral dermatitis|Perioral dermatitis
C0263465|T047|PT|89105000|SNOMEDCT_CORE|Asteatosis cutis|Asteatosis cutis
C0263465|T047|FN|89105000|SNOMEDCT_CORE|Asteatosis cutis|Asteatosis cutis
C0263465|T047|SY|89105000|SNOMEDCT_CORE|Xerosis cutis|Asteatosis cutis
C0263518|T047|PT|39479004|SNOMEDCT_CORE|Telogen effluvium|Telogen effluvium
C0263518|T047|FN|39479004|SNOMEDCT_CORE|Telogen effluvium|Telogen effluvium
C0263525|T047|SY|773296007|SNOMEDCT_CORE|Infection of periungual skin due to ingrown nail|Paronychia due to ingrown nail
C0263525|T047|OAP|25055007|SNOMEDCT_CORE|Ingrowing nail with infection|Paronychia due to ingrown nail
C0263525|T047|SY|773296007|SNOMEDCT_CORE|Ingrowing nail with infection|Paronychia due to ingrown nail
C0263525|T047|OAF|25055007|SNOMEDCT_CORE|Ingrowing nail with infection|Paronychia due to ingrown nail
C0263525|T047|OAS|25055007|SNOMEDCT_CORE|Ingrowing toenail with infection|Paronychia due to ingrown nail
C0263525|T047|PT|773296007|SNOMEDCT_CORE|Paronychia due to ingrown nail|Paronychia due to ingrown nail
C0263525|T047|FN|773296007|SNOMEDCT_CORE|Paronychia due to ingrown nail|Paronychia due to ingrown nail
C0263536|T047|PT|30654002|SNOMEDCT_CORE|Hypertrophy of nail|Hypertrophy of nail
C0263536|T047|FN|30654002|SNOMEDCT_CORE|Hypertrophy of nail|Hypertrophy of nail
C0263536|T047|SY|30654002|SNOMEDCT_CORE|Nail hypertrophy|Hypertrophy of nail
C0263536|T047|SY|30654002|SNOMEDCT_CORE|Nail overgrowth|Hypertrophy of nail
C0263536|T047|SY|30654002|SNOMEDCT_CORE|Onychauxis|Hypertrophy of nail
C0263536|T047|SY|30654002|SNOMEDCT_CORE|OX - Onychauxic|Hypertrophy of nail
C0263537|T047|SY|52897009|SNOMEDCT_CORE|Hook nail|Onychogryposis
C0263537|T047|SY|52897009|SNOMEDCT_CORE|OG - Onychogryphosis|Onychogryposis
C0263537|T047|SY|52897009|SNOMEDCT_CORE|Onychogryphosis|Onychogryposis
C0263537|T047|PT|52897009|SNOMEDCT_CORE|Onychogryposis|Onychogryposis
C0263537|T047|FN|52897009|SNOMEDCT_CORE|Onychogryposis|Onychogryposis
C0263560|T047|IS|26649005|SNOMEDCT_CORE|Chronic ulcer of leg|Chronic ulcer of lower extremity
C0263560|T047|IS|26649005|SNOMEDCT_CORE|Chronic ulcer of leg, NOS|Chronic ulcer of lower extremity
C0263560|T047|PT|26649005|SNOMEDCT_CORE|Chronic ulcer of lower extremity|Chronic ulcer of lower extremity
C0263560|T047|FN|26649005|SNOMEDCT_CORE|Chronic ulcer of lower extremity|Chronic ulcer of lower extremity
C0263560|T047|IS|26649005|SNOMEDCT_CORE|Chronic ulcer of lower extremity, NOS|Chronic ulcer of lower extremity
C0263560|T047|IS|26649005|SNOMEDCT_CORE|Chronic ulcer of lower leg|Chronic ulcer of lower extremity
C0263560|T047|SY|26649005|SNOMEDCT_CORE|Chronic ulcer of lower limb|Chronic ulcer of lower extremity
C0263630|T047|PT|24782002|SNOMEDCT_CORE|Hypertrophic condition of skin|Hypertrophic condition of skin
C0263630|T047|FN|24782002|SNOMEDCT_CORE|Hypertrophic condition of skin|Hypertrophic condition of skin
C0263630|T047|IS|24782002|SNOMEDCT_CORE|Hypertrophic condition of skin, NOS|Hypertrophic condition of skin
C0263630|T047|SY|24782002|SNOMEDCT_CORE|Hypertrophic skin|Hypertrophic condition of skin
C0263637|T191|IS|195382003|SNOMEDCT_CORE|Angioma serpiginosum of skin|Angioma serpiginosum of skin
C0263661|T047|IS|88230002|SNOMEDCT_CORE|Disease of bone and joint, NOS|Disorder of skeletal system
C0263661|T047|SY|88230002|SNOMEDCT_CORE|Disease of bone AND/OR joint|Disorder of skeletal system
C0263661|T047|IS|88230002|SNOMEDCT_CORE|Disease of skeletal system|Disorder of skeletal system
C0263661|T047|OF|88230002|SNOMEDCT_CORE|Disease of skeletal system|Disorder of skeletal system
C0263661|T047|IS|88230002|SNOMEDCT_CORE|Disease of skeletal system, NOS|Disorder of skeletal system
C0263661|T047|PT|88230002|SNOMEDCT_CORE|Disorder of skeletal system|Disorder of skeletal system
C0263661|T047|FN|88230002|SNOMEDCT_CORE|Disorder of skeletal system|Disorder of skeletal system
C0263661|T047|IS|88230002|SNOMEDCT_CORE|Disorder of skeletal system, NOS|Disorder of skeletal system
C0263661|T047|SY|88230002|SNOMEDCT_CORE|Osteoarthropathy|Disorder of skeletal system
C0263661|T047|IS|88230002|SNOMEDCT_CORE|Osteoarthropathy, NOS|Disorder of skeletal system
C0263680|T047|PT|35908007|SNOMEDCT_CORE|Chronic arthritis|Chronic arthritis
C0263680|T047|FN|35908007|SNOMEDCT_CORE|Chronic arthritis|Chronic arthritis
C0263746|T047|PT|22193007|SNOMEDCT_CORE|Degenerative joint disease of hand|Degenerative joint disease of hand
C0263746|T047|FN|22193007|SNOMEDCT_CORE|Degenerative joint disease of hand|Degenerative joint disease of hand
C0263746|T047|SY|22193007|SNOMEDCT_CORE|Osteoarthritis - hand joint|Degenerative joint disease of hand
C0263746|T047|SY|22193007|SNOMEDCT_CORE|Osteoarthrosis of hand|Degenerative joint disease of hand
C0263750|T047|IS|82300000|SNOMEDCT_CORE|Degenerative joint disease of ankle and foot|Degenerative joint disease of ankle AND/OR foot
C0263750|T047|PT|82300000|SNOMEDCT_CORE|Degenerative joint disease of ankle AND/OR foot|Degenerative joint disease of ankle AND/OR foot
C0263750|T047|FN|82300000|SNOMEDCT_CORE|Degenerative joint disease of ankle AND/OR foot|Degenerative joint disease of ankle AND/OR foot
C0263750|T047|SY|82300000|SNOMEDCT_CORE|Osteoarthritis - ankle and/or foot|Degenerative joint disease of ankle AND/OR foot
C0263750|T047|SY|82300000|SNOMEDCT_CORE|Osteoarthritis - ankle/foot|Degenerative joint disease of ankle AND/OR foot
C0263750|T047|SY|82300000|SNOMEDCT_CORE|Osteoarthrosis of ankle and/or foot|Degenerative joint disease of ankle AND/OR foot
C0263752|T047|PTGB|201831003|SNOMEDCT_CORE|Localised, primary osteoarthritis of the shoulder region|Localized, primary osteoarthritis of the shoulder region
C0263752|T047|PT|201831003|SNOMEDCT_CORE|Localized, primary osteoarthritis of the shoulder region|Localized, primary osteoarthritis of the shoulder region
C0263752|T047|FN|201831003|SNOMEDCT_CORE|Localized, primary osteoarthritis of the shoulder region|Localized, primary osteoarthritis of the shoulder region
C0263752|T047|SYGB|201831003|SNOMEDCT_CORE|Primary localised osteoarthrosis of shoulder region|Localized, primary osteoarthritis of the shoulder region
C0263752|T047|SY|201831003|SNOMEDCT_CORE|Primary localized osteoarthrosis of shoulder region|Localized, primary osteoarthritis of the shoulder region
C0263755|T047|PTGB|201834006|SNOMEDCT_CORE|Localised, primary osteoarthritis of the hand|Localized, primary osteoarthritis of the hand
C0263755|T047|PT|201834006|SNOMEDCT_CORE|Localized, primary osteoarthritis of the hand|Localized, primary osteoarthritis of the hand
C0263755|T047|FN|201834006|SNOMEDCT_CORE|Localized, primary osteoarthritis of the hand|Localized, primary osteoarthritis of the hand
C0263755|T047|SYGB|201834006|SNOMEDCT_CORE|Primary localised osteoarthrosis of hand|Localized, primary osteoarthritis of the hand
C0263755|T047|SY|201834006|SNOMEDCT_CORE|Primary localized osteoarthrosis of hand|Localized, primary osteoarthritis of the hand
C0263756|T047|PTGB|77994009|SNOMEDCT_CORE|Primary localised osteoarthrosis of pelvic region|Primary localized osteoarthrosis of pelvic region
C0263756|T047|PT|77994009|SNOMEDCT_CORE|Primary localized osteoarthrosis of pelvic region|Primary localized osteoarthrosis of pelvic region
C0263756|T047|FN|77994009|SNOMEDCT_CORE|Primary localized osteoarthrosis of pelvic region|Primary localized osteoarthrosis of pelvic region
C0263758|T047|OAP|201836008|SNOMEDCT_CORE|Localised, primary osteoarthritis of the lower leg|Localised, primary osteoarthritis of the lower leg
C0263758|T047|OAP|201836008|SNOMEDCT_CORE|Localized, primary osteoarthritis of the lower leg|Localised, primary osteoarthritis of the lower leg
C0263758|T047|OAF|201836008|SNOMEDCT_CORE|Localized, primary osteoarthritis of the lower leg|Localised, primary osteoarthritis of the lower leg
C0263758|T047|OAS|201836008|SNOMEDCT_CORE|Primary localised osteoarthrosis of lower leg|Localised, primary osteoarthritis of the lower leg
C0263758|T047|OAS|201836008|SNOMEDCT_CORE|Primary localized osteoarthrosis of lower leg|Localised, primary osteoarthritis of the lower leg
C0263759|T047|SYGB|201837004|SNOMEDCT_CORE|Localised, primary osteoarthritis of the ankle and foot|Localized, primary osteoarthritis of the ankle and/or foot
C0263759|T047|PTGB|201837004|SNOMEDCT_CORE|Localised, primary osteoarthritis of the ankle and/or foot|Localized, primary osteoarthritis of the ankle and/or foot
C0263759|T047|SY|201837004|SNOMEDCT_CORE|Localized, primary osteoarthritis of the ankle and foot|Localized, primary osteoarthritis of the ankle and/or foot
C0263759|T047|OF|201837004|SNOMEDCT_CORE|Localized, primary osteoarthritis of the ankle and foot|Localized, primary osteoarthritis of the ankle and/or foot
C0263759|T047|PT|201837004|SNOMEDCT_CORE|Localized, primary osteoarthritis of the ankle and/or foot|Localized, primary osteoarthritis of the ankle and/or foot
C0263759|T047|FN|201837004|SNOMEDCT_CORE|Localized, primary osteoarthritis of the ankle and/or foot|Localized, primary osteoarthritis of the ankle and/or foot
C0263759|T047|SYGB|201837004|SNOMEDCT_CORE|Primary localised osteoarthrosis of ankle AND/OR foot|Localized, primary osteoarthritis of the ankle and/or foot
C0263759|T047|SY|201837004|SNOMEDCT_CORE|Primary localized osteoarthrosis of ankle AND/OR foot|Localized, primary osteoarthritis of the ankle and/or foot
C0263772|T047|SY|239872002|SNOMEDCT_CORE|Coxae malum senilis|Coxae malum senilis
C0263774|T047|PTGB|33262002|SNOMEDCT_CORE|Osteoarthrosis involving multiple sites but not designated as generalised|Osteoarthrosis involving multiple sites but not designated as generalized
C0263774|T047|PT|33262002|SNOMEDCT_CORE|Osteoarthrosis involving multiple sites but not designated as generalized|Osteoarthrosis involving multiple sites but not designated as generalized
C0263774|T047|FN|33262002|SNOMEDCT_CORE|Osteoarthrosis involving multiple sites but not designated as generalized|Osteoarthrosis involving multiple sites but not designated as generalized
C0263778|T047|SY|43829003|SNOMEDCT_CORE|Arthritis sicca|Chronic osteoarthritis
C0263778|T047|SY|43829003|SNOMEDCT_CORE|Arthroxerosis|Chronic osteoarthritis
C0263778|T047|PT|43829003|SNOMEDCT_CORE|Chronic osteoarthritis|Chronic osteoarthritis
C0263778|T047|FN|43829003|SNOMEDCT_CORE|Chronic osteoarthritis|Chronic osteoarthritis
C0263782|T047|PT|22591001|SNOMEDCT_CORE|Degeneration of cartilage AND/OR meniscus of knee|Degeneration of cartilage AND/OR meniscus of knee
C0263782|T047|FN|22591001|SNOMEDCT_CORE|Degeneration of cartilage AND/OR meniscus of knee|Degeneration of cartilage AND/OR meniscus of knee
C0263782|T047|SY|22591001|SNOMEDCT_CORE|Degeneration of cartilage or meniscus of knee|Degeneration of cartilage AND/OR meniscus of knee
C0263782|T047|IS|22591001|SNOMEDCT_CORE|Degeneration of cartilage or meniscus of knee, NOS|Degeneration of cartilage AND/OR meniscus of knee
C0263789|T047|PT|14949009|SNOMEDCT_CORE|Old disruption of ligament of knee|Old disruption of ligament of knee
C0263789|T047|FN|14949009|SNOMEDCT_CORE|Old disruption of ligament of knee|Old disruption of ligament of knee
C0263789|T047|IS|14949009|SNOMEDCT_CORE|Old disruption of ligament of knee, NOS|Old disruption of ligament of knee
C0263813|T037|PT|30556007|SNOMEDCT_CORE|Recurrent dislocation of shoulder region|Recurrent dislocation of shoulder region
C0263813|T037|FN|30556007|SNOMEDCT_CORE|Recurrent dislocation of shoulder region|Recurrent dislocation of shoulder region
C0263854|T047|PT|387801000|SNOMEDCT_CORE|Cervical arthritis|Cervical arthritis
C0263854|T047|FN|387801000|SNOMEDCT_CORE|Cervical arthritis|Cervical arthritis
C0263854|T047|SY|387800004|SNOMEDCT_CORE|Cervical osteoarthritis|Cervical arthritis
C0263854|T047|SY|387800004|SNOMEDCT_CORE|Cervical spondylarthritis|Cervical arthritis
C0263854|T047|SY|387801000|SNOMEDCT_CORE|Cervical spondylitis|Cervical arthritis
C0263854|T047|SY|387800004|SNOMEDCT_CORE|Osteoarthritis of cervical spine|Cervical arthritis
C0263856|T047|SY|34781003|SNOMEDCT_CORE|Vertebral artery compression syndrome|Vertebral artery compression syndrome
C0263872|T047|PT|68675004|SNOMEDCT_CORE|Degeneration of thoracic intervertebral disc|Degeneration of thoracic intervertebral disc
C0263872|T047|FN|68675004|SNOMEDCT_CORE|Degeneration of thoracic intervertebral disc|Degeneration of thoracic intervertebral disc
C0263874|T047|PT|26538006|SNOMEDCT_CORE|Degeneration of lumbar intervertebral disc|Degeneration of lumbar intervertebral disc
C0263874|T047|FN|26538006|SNOMEDCT_CORE|Degeneration of lumbar intervertebral disc|Degeneration of lumbar intervertebral disc
C0263875|T047|PT|60937000|SNOMEDCT_CORE|Degeneration of lumbosacral intervertebral disc|Degeneration of lumbosacral intervertebral disc
C0263875|T047|FN|60937000|SNOMEDCT_CORE|Degeneration of lumbosacral intervertebral disc|Degeneration of lumbosacral intervertebral disc
C0263884|T047|PT|11049006|SNOMEDCT_CORE|Cervical radiculitis|Cervical radiculitis
C0263884|T047|FN|11049006|SNOMEDCT_CORE|Cervical radiculitis|Cervical radiculitis
C0263898|T047|PT|46578006|SNOMEDCT_CORE|Lumbosacral radiculitis|Lumbosacral radiculitis
C0263898|T047|FN|46578006|SNOMEDCT_CORE|Lumbosacral radiculitis|Lumbosacral radiculitis
C0263898|T047|IS|46578006|SNOMEDCT_CORE|Lumbosacral radiculitis, NOS|Lumbosacral radiculitis
C0263904|T046|IS|29885006|SNOMEDCT_CORE|Instability of sacroiliac joint|Sacroiliac instability
C0263904|T046|PT|29885006|SNOMEDCT_CORE|Sacroiliac instability|Sacroiliac instability
C0263904|T046|FN|29885006|SNOMEDCT_CORE|Sacroiliac instability|Sacroiliac instability
C0263904|T046|OF|29885006|SNOMEDCT_CORE|Sacroiliac instability|Sacroiliac instability
C0263904|T046|SY|29885006|SNOMEDCT_CORE|Sacroiliac joint unstable|Sacroiliac instability
C0263907|T047|PT|6858004|SNOMEDCT_CORE|Capsulitis|Capsulitis
C0263907|T047|FN|6858004|SNOMEDCT_CORE|Capsulitis|Capsulitis
C0263907|T047|IS|6858004|SNOMEDCT_CORE|Capsulitis, NOS|Capsulitis
C0263910|T047|PT|55833001|SNOMEDCT_CORE|Disorder of bursa of shoulder region|Disorder of bursa of shoulder region
C0263910|T047|FN|55833001|SNOMEDCT_CORE|Disorder of bursa of shoulder region|Disorder of bursa of shoulder region
C0263910|T047|SY|55833001|SNOMEDCT_CORE|Disorder of bursae of shoulder region|Disorder of bursa of shoulder region
C0263910|T047|OF|55833001|SNOMEDCT_CORE|Disorder of bursae of shoulder region|Disorder of bursa of shoulder region
C0263910|T047|IS|55833001|SNOMEDCT_CORE|Disorder of bursae of shoulder region, NOS|Disorder of bursa of shoulder region
C0263910|T047|SY|55833001|SNOMEDCT_CORE|Disorder of shoulder bursa|Disorder of bursa of shoulder region
C0263910|T047|SY|55833001|SNOMEDCT_CORE|Shoulder bursa disorder|Disorder of bursa of shoulder region
C0263911|T047|PT|76318008|SNOMEDCT_CORE|Disorder of tendon of shoulder region|Disorder of tendon of shoulder region
C0263911|T047|FN|76318008|SNOMEDCT_CORE|Disorder of tendon of shoulder region|Disorder of tendon of shoulder region
C0263911|T047|IS|76318008|SNOMEDCT_CORE|Disorder of tendon of shoulder region, NOS|Disorder of tendon of shoulder region
C0263912|T047|IS|4106009|SNOMEDCT_CORE|Impingement syndrome|Rotator cuff syndrome
C0263912|T047|SY|4106009|SNOMEDCT_CORE|Rotator cuff rupture|Rotator cuff syndrome
C0263912|T047|PT|4106009|SNOMEDCT_CORE|Rotator cuff syndrome|Rotator cuff syndrome
C0263912|T047|FN|4106009|SNOMEDCT_CORE|Rotator cuff syndrome|Rotator cuff syndrome
C0263912|T047|IS|4106009|SNOMEDCT_CORE|Rotator cuff syndrome, NOS|Rotator cuff syndrome
C0263912|T047|SY|4106009|SNOMEDCT_CORE|Rotator cuff tear|Rotator cuff syndrome
C0263912|T047|SY|4106009|SNOMEDCT_CORE|Rupture of rotator cuff of shoulder|Rotator cuff syndrome
C0263922|T047|PT|81498004|SNOMEDCT_CORE|Bursitis of hip|Bursitis of hip
C0263922|T047|FN|81498004|SNOMEDCT_CORE|Bursitis of hip|Bursitis of hip
C0263929|T047|PT|73105000|SNOMEDCT_CORE|Pes anserinus bursitis|Pes anserinus bursitis
C0263929|T047|FN|73105000|SNOMEDCT_CORE|Pes anserinus bursitis|Pes anserinus bursitis
C0263933|T047|PT|11654001|SNOMEDCT_CORE|Achilles tendinitis|Achilles tendinitis
C0263933|T047|FN|11654001|SNOMEDCT_CORE|Achilles tendinitis|Achilles tendinitis
C0263933|T047|SY|11654001|SNOMEDCT_CORE|Achilles tendonitis|Achilles tendinitis
C0263936|T047|PT|53208009|SNOMEDCT_CORE|Peroneal tendinitis|Peroneal tendinitis
C0263936|T047|FN|53208009|SNOMEDCT_CORE|Peroneal tendinitis|Peroneal tendinitis
C0263936|T047|SY|53208009|SNOMEDCT_CORE|Peroneal tendonitis|Peroneal tendinitis
C0263957|T020|SY|7951001|SNOMEDCT_CORE|Bunionette|Tailor's bunion
C0263957|T020|PT|7951001|SNOMEDCT_CORE|Tailor's bunion|Tailor's bunion
C0263957|T020|FN|7951001|SNOMEDCT_CORE|Tailor's bunion|Tailor's bunion
C0263957|T020|SY|7951001|SNOMEDCT_CORE|Tailors bunion|Tailor's bunion
C0263962|T047|SY|425940002|SNOMEDCT_CORE|Capped elbow|Olecranon bursitis
C0263962|T047|SY|425940002|SNOMEDCT_CORE|Inflammation of bursa of olecranon|Olecranon bursitis
C0263962|T047|FN|425940002|SNOMEDCT_CORE|Inflammation of bursa of olecranon|Olecranon bursitis
C0263962|T047|SY|425940002|SNOMEDCT_CORE|Miner's elbow|Olecranon bursitis
C0263962|T047|IS|425940002|SNOMEDCT_CORE|Miners' elbow|Olecranon bursitis
C0263962|T047|PT|425940002|SNOMEDCT_CORE|Olecranon bursitis|Olecranon bursitis
C0263962|T047|SY|425940002|SNOMEDCT_CORE|Student's elbow|Olecranon bursitis
C0263970|T037|SY|429513001|SNOMEDCT_CORE|Rupture achilles tendon|Rupture of Achilles tendon
C0263970|T037|PT|429513001|SNOMEDCT_CORE|Rupture of Achilles tendon|Rupture of Achilles tendon
C0263970|T037|FN|429513001|SNOMEDCT_CORE|Rupture of Achilles tendon|Rupture of Achilles tendon
C0263978|T047|PT|19660004|SNOMEDCT_CORE|Disorder of soft tissue|Disorder of soft tissue
C0263978|T047|FN|19660004|SNOMEDCT_CORE|Disorder of soft tissue|Disorder of soft tissue
C0263978|T047|IS|19660004|SNOMEDCT_CORE|Disorder of soft tissue, NOS|Disorder of soft tissue
C0263978|T047|SY|19660004|SNOMEDCT_CORE|Soft tissue disorder|Disorder of soft tissue
C0264028|T047|PT|21120002|SNOMEDCT_CORE|Osteomyelitis of lower leg|Osteomyelitis of lower leg
C0264028|T047|FN|21120002|SNOMEDCT_CORE|Osteomyelitis of lower leg|Osteomyelitis of lower leg
C0264029|T047|IS|28769004|SNOMEDCT_CORE|Osteomyelitis of ankle and foot|Osteomyelitis of ankle AND/OR foot
C0264029|T047|PT|28769004|SNOMEDCT_CORE|Osteomyelitis of ankle AND/OR foot|Osteomyelitis of ankle AND/OR foot
C0264029|T047|FN|28769004|SNOMEDCT_CORE|Osteomyelitis of ankle AND/OR foot|Osteomyelitis of ankle AND/OR foot
C0264039|T047|PT|268017000|SNOMEDCT_CORE|Acute osteomyelitis of ankle and/or foot|Acute osteomyelitis of ankle and/or foot
C0264039|T047|FN|268017000|SNOMEDCT_CORE|Acute osteomyelitis of ankle and/or foot|Acute osteomyelitis of ankle and/or foot
C0264039|T047|SY|268017000|SNOMEDCT_CORE|Acute osteomyelitis of the ankle and foot|Acute osteomyelitis of ankle and/or foot
C0264039|T047|OF|268017000|SNOMEDCT_CORE|Acute osteomyelitis of the ankle and foot|Acute osteomyelitis of ankle and/or foot
C0264039|T047|OP|268017000|SNOMEDCT_CORE|Acute osteomyelitis of the ankle and/or foot|Acute osteomyelitis of ankle and/or foot
C0264039|T047|OF|268017000|SNOMEDCT_CORE|Acute osteomyelitis of the ankle and/or foot|Acute osteomyelitis of ankle and/or foot
C0264049|T047|PT|268019002|SNOMEDCT_CORE|Chronic osteomyelitis of ankle and/or foot|Chronic osteomyelitis of ankle and/or foot
C0264049|T047|FN|268019002|SNOMEDCT_CORE|Chronic osteomyelitis of ankle and/or foot|Chronic osteomyelitis of ankle and/or foot
C0264049|T047|IS|268019002|SNOMEDCT_CORE|Chronic osteomyelitis of the ankle and foot|Chronic osteomyelitis of ankle and/or foot
C0264049|T047|OF|268019002|SNOMEDCT_CORE|Chronic osteomyelitis of the ankle and foot|Chronic osteomyelitis of ankle and/or foot
C0264049|T047|OP|268019002|SNOMEDCT_CORE|Chronic osteomyelitis of the ankle and/or foot|Chronic osteomyelitis of ankle and/or foot
C0264049|T047|OF|268019002|SNOMEDCT_CORE|Chronic osteomyelitis of the ankle and/or foot|Chronic osteomyelitis of ankle and/or foot
C0264133|T020|IS|53226007|SNOMEDCT_CORE|Acquired flat foot|Talipes planus
C0264133|T020|IS|53226007|SNOMEDCT_CORE|Acquired pes planus|Talipes planus
C0264133|T020|IS|53226007|SNOMEDCT_CORE|Acquired talipes planus|Talipes planus
C0264133|T020|SY|53226007|SNOMEDCT_CORE|Fallen arch|Talipes planus
C0264133|T020|IS|53226007|SNOMEDCT_CORE|Fallen arches|Talipes planus
C0264133|T020|SY|53226007|SNOMEDCT_CORE|Flat foot|Talipes planus
C0264133|T020|SY|53226007|SNOMEDCT_CORE|Low medial arch of foot|Talipes planus
C0264133|T020|SY|53226007|SNOMEDCT_CORE|Pes planus|Talipes planus
C0264133|T020|OF|53226007|SNOMEDCT_CORE|Pes planus|Talipes planus
C0264133|T020|FN|53226007|SNOMEDCT_CORE|Talipes planus|Talipes planus
C0264133|T020|PT|53226007|SNOMEDCT_CORE|Talipes planus|Talipes planus
C0264134|T047|PT|6654000|SNOMEDCT_CORE|Acquired hallux rigidus|Acquired hallux rigidus
C0264134|T047|FN|6654000|SNOMEDCT_CORE|Acquired hallux rigidus|Acquired hallux rigidus
C0264134|T047|SY|6654000|SNOMEDCT_CORE|Hallux rigidus|Acquired hallux rigidus
C0264134|T047|SY|6654000|SNOMEDCT_CORE|Hallux rigidus - acquired|Acquired hallux rigidus
C0264134|T047|IS|6654000|SNOMEDCT_CORE|HL - Hallux limitus|Acquired hallux rigidus
C0264134|T047|SY|6654000|SNOMEDCT_CORE|HR - Hallux rigidus|Acquired hallux rigidus
C0264134|T047|SY|6654000|SNOMEDCT_CORE|Rigidity of 1st MTP joint|Acquired hallux rigidus
C0264150|T020|SY|88562000|SNOMEDCT_CORE|Acquired ankle and/or foot deformity|Acquired deformity of ankle AND/OR foot
C0264150|T020|IS|88562000|SNOMEDCT_CORE|Acquired deformity of ankle and foot, NOS|Acquired deformity of ankle AND/OR foot
C0264150|T020|PT|88562000|SNOMEDCT_CORE|Acquired deformity of ankle AND/OR foot|Acquired deformity of ankle AND/OR foot
C0264150|T020|FN|88562000|SNOMEDCT_CORE|Acquired deformity of ankle AND/OR foot|Acquired deformity of ankle AND/OR foot
C0264156|T020|OAS|68701004|SNOMEDCT_CORE|Acquired disparity of leg length|Acquired unequal leg length
C0264156|T020|PT|203601000|SNOMEDCT_CORE|Acquired unequal leg length|Acquired unequal leg length
C0264156|T020|OAP|68701004|SNOMEDCT_CORE|Acquired unequal leg length|Acquired unequal leg length
C0264156|T020|OF|203601000|SNOMEDCT_CORE|Acquired unequal leg length|Acquired unequal leg length
C0264156|T020|OF|68701004|SNOMEDCT_CORE|Acquired unequal leg length|Acquired unequal leg length
C0264156|T020|FN|203601000|SNOMEDCT_CORE|Acquired unequal leg length|Acquired unequal leg length
C0264156|T020|OAF|68701004|SNOMEDCT_CORE|Acquired unequal leg length|Acquired unequal leg length
C0264156|T020|SY|203601000|SNOMEDCT_CORE|Acquired unequal lower limb length|Acquired unequal leg length
C0264184|T047|PT|4046000|SNOMEDCT_CORE|Degenerative spondylolisthesis|Degenerative spondylolisthesis
C0264184|T047|FN|4046000|SNOMEDCT_CORE|Degenerative spondylolisthesis|Degenerative spondylolisthesis
C0264222|T047|PT|54398005|SNOMEDCT_CORE|Acute upper respiratory infection|Acute upper respiratory infection
C0264222|T047|FN|54398005|SNOMEDCT_CORE|Acute upper respiratory infection|Acute upper respiratory infection
C0264222|T047|SY|54398005|SNOMEDCT_CORE|Acute upper respiratory tract infection|Acute upper respiratory infection
C0264222|T047|SY|54398005|SNOMEDCT_CORE|Acute URI|Acute upper respiratory infection
C0264222|T047|SY|54398005|SNOMEDCT_CORE|AURTI - Acute upper respiratory tract infection|Acute upper respiratory infection
C0264222|T047|IS|54398005|SNOMEDCT_CORE|URTI - Acute upper respiratory infection|Acute upper respiratory infection
C0264230|T047|PT|80600003|SNOMEDCT_CORE|Acute suppuration of nasal sinus|Acute suppuration of nasal sinus
C0264230|T047|FN|80600003|SNOMEDCT_CORE|Acute suppuration of nasal sinus|Acute suppuration of nasal sinus
C0264230|T047|SY|80600003|SNOMEDCT_CORE|Acute suppurative inflammation of nasal sinus|Acute suppuration of nasal sinus
C0264230|T047|SY|80600003|SNOMEDCT_CORE|Acute suppurative sinusitis|Acute suppuration of nasal sinus
C0264231|T191|SY|32307003|SNOMEDCT_CORE|Nasal sinus polyp|Polyp of nasal sinus
C0264231|T191|SY|32307003|SNOMEDCT_CORE|Polyp of accessory sinus|Polyp of nasal sinus
C0264231|T191|IS|32307003|SNOMEDCT_CORE|Polyp of accessory sinus, NOS|Polyp of nasal sinus
C0264231|T191|PT|32307003|SNOMEDCT_CORE|Polyp of nasal sinus|Polyp of nasal sinus
C0264231|T191|FN|32307003|SNOMEDCT_CORE|Polyp of nasal sinus|Polyp of nasal sinus
C0264231|T191|IS|32307003|SNOMEDCT_CORE|Polyp of nasal sinus, NOS|Polyp of nasal sinus
C0264272|T184|PT|8442000|SNOMEDCT_CORE|Purulent rhinitis|Purulent rhinitis
C0264272|T184|FN|8442000|SNOMEDCT_CORE|Purulent rhinitis|Purulent rhinitis
C0264303|T019|PT|38086007|SNOMEDCT_CORE|Laryngomalacia|Laryngomalacia
C0264303|T019|FN|38086007|SNOMEDCT_CORE|Laryngomalacia|Laryngomalacia
C0264309|T047|IS|57781000|SNOMEDCT_CORE|Disease of vocal cords|Disorder of vocal cord
C0264309|T047|OF|57781000|SNOMEDCT_CORE|Disease of vocal cords|Disorder of vocal cord
C0264309|T047|IS|57781000|SNOMEDCT_CORE|Disease of vocal cords, NOS|Disorder of vocal cord
C0264309|T047|PT|57781000|SNOMEDCT_CORE|Disorder of vocal cord|Disorder of vocal cord
C0264309|T047|FN|57781000|SNOMEDCT_CORE|Disorder of vocal cord|Disorder of vocal cord
C0264314|T046|PT|57713008|SNOMEDCT_CORE|Chorditis|Chorditis
C0264314|T046|OF|57713008|SNOMEDCT_CORE|Chorditis|Chorditis
C0264314|T046|SY|57713008|SNOMEDCT_CORE|Inflammation of vocal cord|Chorditis
C0264314|T046|FN|57713008|SNOMEDCT_CORE|Inflammation of vocal cord|Chorditis
C0264314|T046|SY|57713008|SNOMEDCT_CORE|Singers' chorditis|Chorditis
C0264348|T047|PT|195949008|SNOMEDCT_CORE|Chronic asthmatic bronchitis|Chronic asthmatic bronchitis
C0264348|T047|FN|195949008|SNOMEDCT_CORE|Chronic asthmatic bronchitis|Chronic asthmatic bronchitis
C0264348|T047|SY|195949008|SNOMEDCT_CORE|Chronic wheezy bronchitis|Chronic asthmatic bronchitis
C0264390|T047|SY|196035006|SNOMEDCT_CORE|Aspiration pneumonia caused by vomit|Pneumonitis due to inhalation of vomitus
C0264390|T047|SY|196035006|SNOMEDCT_CORE|Aspiration pneumonia due to vomit|Pneumonitis due to inhalation of vomitus
C0264390|T047|SY|196035006|SNOMEDCT_CORE|Pneumonitis caused by inhalation of vomitus|Pneumonitis due to inhalation of vomitus
C0264390|T047|FN|196035006|SNOMEDCT_CORE|Pneumonitis caused by inhalation of vomitus|Pneumonitis due to inhalation of vomitus
C0264390|T047|PT|196035006|SNOMEDCT_CORE|Pneumonitis due to inhalation of vomitus|Pneumonitis due to inhalation of vomitus
C0264390|T047|OF|196035006|SNOMEDCT_CORE|Pneumonitis due to inhalation of vomitus|Pneumonitis due to inhalation of vomitus
C0264390|T047|SY|196035006|SNOMEDCT_CORE|Vomit inhalation pneumonitis|Pneumonitis due to inhalation of vomitus
C0264405|T047|PT|55570000|SNOMEDCT_CORE|Asthma without status asthmaticus|Asthma without status asthmaticus
C0264405|T047|FN|55570000|SNOMEDCT_CORE|Asthma without status asthmaticus|Asthma without status asthmaticus
C0264490|T047|PT|65710008|SNOMEDCT_CORE|Acute respiratory failure|Acute respiratory failure
C0264490|T047|FN|65710008|SNOMEDCT_CORE|Acute respiratory failure|Acute respiratory failure
C0264490|T047|SY|65710008|SNOMEDCT_CORE|ARF - Acute respiratory failure|Acute respiratory failure
C0264491|T047|SY|67905004|SNOMEDCT_CORE|Acute on chronic respiratory failure|Acute-on-chronic respiratory failure
C0264491|T047|PT|67905004|SNOMEDCT_CORE|Acute-on-chronic respiratory failure|Acute-on-chronic respiratory failure
C0264491|T047|FN|67905004|SNOMEDCT_CORE|Acute-on-chronic respiratory failure|Acute-on-chronic respiratory failure
C0264492|T047|PT|39871006|SNOMEDCT_CORE|Chronic respiratory failure|Chronic respiratory failure
C0264492|T047|FN|39871006|SNOMEDCT_CORE|Chronic respiratory failure|Chronic respiratory failure
C0264545|T047|SY|73725006|SNOMEDCT_CORE|Pleural cuirasse|Thickening of pleura
C0264545|T047|SY|73725006|SNOMEDCT_CORE|Pleural thickening|Thickening of pleura
C0264545|T047|PT|73725006|SNOMEDCT_CORE|Thickening of pleura|Thickening of pleura
C0264545|T047|FN|73725006|SNOMEDCT_CORE|Thickening of pleura|Thickening of pleura
C0264550|T047|SY|81075000|SNOMEDCT_CORE|Parapneumonic effusion|Pleural effusion associated with pulmonary infection
C0264550|T047|PT|81075000|SNOMEDCT_CORE|Pleural effusion associated with pulmonary infection|Pleural effusion associated with pulmonary infection
C0264550|T047|FN|81075000|SNOMEDCT_CORE|Pleural effusion associated with pulmonary infection|Pleural effusion associated with pulmonary infection
C0264588|T033|SY|29003001|SNOMEDCT_CORE|Spasmodic dysphonia|Spastic dysphonia
C0264588|T033|PT|29003001|SNOMEDCT_CORE|Spastic dysphonia|Spastic dysphonia
C0264588|T033|FN|29003001|SNOMEDCT_CORE|Spastic dysphonia|Spastic dysphonia
C0264588|T033|IS|29003001|SNOMEDCT_CORE|Spastic dysphonia, NOS|Spastic dysphonia
C0264611|T047|SY|74227009|SNOMEDCT_CORE|Apraxia of phonation|Apraxic aphonia
C0264611|T047|SY|74227009|SNOMEDCT_CORE|Apraxia of speech|Apraxic aphonia
C0264611|T047|PT|74227009|SNOMEDCT_CORE|Apraxic aphonia|Apraxic aphonia
C0264611|T047|FN|74227009|SNOMEDCT_CORE|Apraxic aphonia|Apraxic aphonia
C0264611|T047|SY|74227009|SNOMEDCT_CORE|Verbal apraxia|Apraxic aphonia
C0264637|T047|FN|10725009|SNOMEDCT_CORE|Benign hypertension|Benign hypertension
C0264637|T047|PT|10725009|SNOMEDCT_CORE|Benign hypertension|Benign hypertension
C0264642|T047|PT|73410007|SNOMEDCT_CORE|Benign secondary renovascular hypertension|Benign secondary renovascular hypertension
C0264642|T047|FN|73410007|SNOMEDCT_CORE|Benign secondary renovascular hypertension|Benign secondary renovascular hypertension
C0264642|T047|SY|73410007|SNOMEDCT_CORE|Secondary benign renovascular hypertension|Benign secondary renovascular hypertension
C0264650|T047|PT|5148006|SNOMEDCT_CORE|Hypertensive heart disease with congestive heart failure|Hypertensive heart disease with congestive heart failure
C0264650|T047|FN|5148006|SNOMEDCT_CORE|Hypertensive heart disease with congestive heart failure|Hypertensive heart disease with congestive heart failure
C0264652|T047|PT|46113002|SNOMEDCT_CORE|Hypertensive heart failure|Hypertensive heart failure
C0264652|T047|FN|46113002|SNOMEDCT_CORE|Hypertensive heart failure|Hypertensive heart failure
C0264652|T047|IS|46113002|SNOMEDCT_CORE|Hypertensive heart failure, NOS|Hypertensive heart failure
C0264653|T047|PT|49220004|SNOMEDCT_CORE|Hypertensive renal failure|Hypertensive renal failure
C0264653|T047|FN|49220004|SNOMEDCT_CORE|Hypertensive renal failure|Hypertensive renal failure
C0264694|T047|PTGB|413838009|SNOMEDCT_CORE|Chronic ischaemic heart disease|Chronic ischemic heart disease
C0264694|T047|PT|413838009|SNOMEDCT_CORE|Chronic ischemic heart disease|Chronic ischemic heart disease
C0264694|T047|FN|413838009|SNOMEDCT_CORE|Chronic ischemic heart disease|Chronic ischemic heart disease
C0264695|T047|PTGB|46109009|SNOMEDCT_CORE|Subendocardial ischaemia|Subendocardial ischemia
C0264695|T047|PT|46109009|SNOMEDCT_CORE|Subendocardial ischemia|Subendocardial ischemia
C0264695|T047|FN|46109009|SNOMEDCT_CORE|Subendocardial ischemia|Subendocardial ischemia
C0264699|T047|PT|62695002|SNOMEDCT_CORE|Acute anteroseptal myocardial infarction|Acute anteroseptal myocardial infarction
C0264699|T047|FN|62695002|SNOMEDCT_CORE|Acute anteroseptal myocardial infarction|Acute anteroseptal myocardial infarction
C0264700|T047|SY|73795002|SNOMEDCT_CORE|Acute inferior myocardial infarction|Acute myocardial infarction of inferior wall
C0264700|T047|SY|73795002|SNOMEDCT_CORE|Acute myocardial infarction of diaphragmatic wall|Acute myocardial infarction of inferior wall
C0264700|T047|PT|73795002|SNOMEDCT_CORE|Acute myocardial infarction of inferior wall|Acute myocardial infarction of inferior wall
C0264700|T047|FN|73795002|SNOMEDCT_CORE|Acute myocardial infarction of inferior wall|Acute myocardial infarction of inferior wall
C0264700|T047|IS|73795002|SNOMEDCT_CORE|Acute myocardial infarction of inferior wall, NOS|Acute myocardial infarction of inferior wall
C0264710|T047|IS|70422006|SNOMEDCT_CORE|Acute nontransmural infarction|Acute subendocardial infarction
C0264710|T047|PT|70422006|SNOMEDCT_CORE|Acute subendocardial infarction|Acute subendocardial infarction
C0264710|T047|FN|70422006|SNOMEDCT_CORE|Acute subendocardial infarction|Acute subendocardial infarction
C0264722|T047|PT|88805009|SNOMEDCT_CORE|Chronic congestive heart failure|Chronic congestive heart failure
C0264722|T047|FN|88805009|SNOMEDCT_CORE|Chronic congestive heart failure|Chronic congestive heart failure
C0264766|T047|PT|86466006|SNOMEDCT_CORE|Rheumatic mitral stenosis|Rheumatic mitral stenosis
C0264766|T047|FN|86466006|SNOMEDCT_CORE|Rheumatic mitral stenosis|Rheumatic mitral stenosis
C0264766|T047|IS|86466006|SNOMEDCT_CORE|Rheumatic mitral stenosis, NOS|Rheumatic mitral stenosis
C0264766|T047|SY|86466006|SNOMEDCT_CORE|Rheumatic mitral valve obstruction|Rheumatic mitral stenosis
C0264767|T047|SY|787001|SNOMEDCT_CORE|Rheumatic mitral stenosis with incompetence|Rheumatic mitral stenosis with regurgitation
C0264767|T047|SY|787001|SNOMEDCT_CORE|Rheumatic mitral stenosis with insufficiency|Rheumatic mitral stenosis with regurgitation
C0264767|T047|PT|787001|SNOMEDCT_CORE|Rheumatic mitral stenosis with regurgitation|Rheumatic mitral stenosis with regurgitation
C0264767|T047|FN|787001|SNOMEDCT_CORE|Rheumatic mitral stenosis with regurgitation|Rheumatic mitral stenosis with regurgitation
C0264774|T047|PT|194736003|SNOMEDCT_CORE|Mitral and aortic incompetence|Mitral and aortic incompetence
C0264774|T047|FN|194736003|SNOMEDCT_CORE|Mitral and aortic incompetence|Mitral and aortic incompetence
C0264774|T047|SY|194736003|SNOMEDCT_CORE|Mitral and aortic insufficiency|Mitral and aortic incompetence
C0264774|T047|SY|194736003|SNOMEDCT_CORE|Mitral and aortic regurgitation|Mitral and aortic incompetence
C0264776|T047|PT|49699002|SNOMEDCT_CORE|Rheumatic disease of tricuspid valve|Rheumatic disease of tricuspid valve
C0264776|T047|FN|49699002|SNOMEDCT_CORE|Rheumatic disease of tricuspid valve|Rheumatic disease of tricuspid valve
C0264776|T047|IS|49699002|SNOMEDCT_CORE|Rheumatic disease of tricuspid valve, NOS|Rheumatic disease of tricuspid valve
C0264776|T047|SY|49699002|SNOMEDCT_CORE|Rheumatic tricuspid valve disease|Rheumatic disease of tricuspid valve
C0264776|T047|IS|49699002|SNOMEDCT_CORE|Rheumatic tricuspid valve disease, NOS|Rheumatic disease of tricuspid valve
C0264778|T047|SY|67696008|SNOMEDCT_CORE|Rheumatic tricuspid insufficiency|Rheumatic tricuspid valve regurgitation
C0264778|T047|SY|67696008|SNOMEDCT_CORE|Rheumatic tricuspid regurgitation|Rheumatic tricuspid valve regurgitation
C0264778|T047|SY|67696008|SNOMEDCT_CORE|Rheumatic tricuspid valve incompetence|Rheumatic tricuspid valve regurgitation
C0264778|T047|SY|67696008|SNOMEDCT_CORE|Rheumatic tricuspid valve insufficiency|Rheumatic tricuspid valve regurgitation
C0264778|T047|PT|67696008|SNOMEDCT_CORE|Rheumatic tricuspid valve regurgitation|Rheumatic tricuspid valve regurgitation
C0264778|T047|FN|67696008|SNOMEDCT_CORE|Rheumatic tricuspid valve regurgitation|Rheumatic tricuspid valve regurgitation
C0264778|T047|SY|67696008|SNOMEDCT_CORE|Tricuspid incompetence - rheumatic|Rheumatic tricuspid valve regurgitation
C0264839|T047|PT|15544002|SNOMEDCT_CORE|Restrictive cardiomyopathy secondary to infiltrations|Restrictive cardiomyopathy secondary to infiltrations
C0264839|T047|FN|15544002|SNOMEDCT_CORE|Restrictive cardiomyopathy secondary to infiltrations|Restrictive cardiomyopathy secondary to infiltrations
C0264882|T047|SY|20721001|SNOMEDCT_CORE|Tricuspid valve disease|Tricuspid valve disorder
C0264882|T047|PT|20721001|SNOMEDCT_CORE|Tricuspid valve disorder|Tricuspid valve disorder
C0264882|T047|FN|20721001|SNOMEDCT_CORE|Tricuspid valve disorder|Tricuspid valve disorder
C0264882|T047|IS|20721001|SNOMEDCT_CORE|Tricuspid valve disorder, NOS|Tricuspid valve disorder
C0264886|T047|PT|44808001|SNOMEDCT_CORE|Conduction disorder of the heart|Conduction disorder of the heart
C0264886|T047|FN|44808001|SNOMEDCT_CORE|Conduction disorder of the heart|Conduction disorder of the heart
C0264886|T047|IS|44808001|SNOMEDCT_CORE|Conduction disorder of the heart, NOS|Conduction disorder of the heart
C0264886|T047|SY|44808001|SNOMEDCT_CORE|Disorder of heart conduction|Conduction disorder of the heart
C0264893|T047|SY|71792006|SNOMEDCT_CORE|Nodal arrhythmia|Nodal rhythm disorder
C0264893|T047|PT|71792006|SNOMEDCT_CORE|Nodal rhythm disorder|Nodal rhythm disorder
C0264893|T047|FN|71792006|SNOMEDCT_CORE|Nodal rhythm disorder|Nodal rhythm disorder
C0264907|T047|SY|54016002|SNOMEDCT_CORE|Mobitz type 1 second degree atrioventricular block|Mobitz type I incomplete atrioventricular block
C0264907|T047|PT|54016002|SNOMEDCT_CORE|Mobitz type I incomplete atrioventricular block|Mobitz type I incomplete atrioventricular block
C0264907|T047|FN|54016002|SNOMEDCT_CORE|Mobitz type I incomplete atrioventricular block|Mobitz type I incomplete atrioventricular block
C0264907|T047|SY|54016002|SNOMEDCT_CORE|Mobitz type I Wenckebach atrioventricular block|Mobitz type I incomplete atrioventricular block
C0264907|T047|SY|54016002|SNOMEDCT_CORE|Wenckebach's incomplete AV block|Mobitz type I incomplete atrioventricular block
C0264907|T047|SY|54016002|SNOMEDCT_CORE|Wenckebach's phenomenon|Mobitz type I incomplete atrioventricular block
C0264936|T047|PT|88223008|SNOMEDCT_CORE|Secondary pulmonary hypertension|Secondary pulmonary hypertension
C0264936|T047|FN|88223008|SNOMEDCT_CORE|Secondary pulmonary hypertension|Secondary pulmonary hypertension
C0264964|T047|PT|48273005|SNOMEDCT_CORE|Aneurysm of popliteal artery|Aneurysm of popliteal artery
C0264964|T047|FN|48273005|SNOMEDCT_CORE|Aneurysm of popliteal artery|Aneurysm of popliteal artery
C0264964|T047|SY|48273005|SNOMEDCT_CORE|Popliteal artery aneurysm|Aneurysm of popliteal artery
C0264993|T047|PT|399923009|SNOMEDCT_CORE|Rheumatoid arteritis|Rheumatoid arteritis
C0264993|T047|FN|399923009|SNOMEDCT_CORE|Rheumatoid arteritis|Rheumatoid arteritis
C0264995|T046|SY|2929001|SNOMEDCT_CORE|Arterial occlusion|Arterial occlusion
C0264995|T046|SY|2929001|SNOMEDCT_CORE|Blocked artery|Arterial occlusion
C0264995|T046|SY|2929001|SNOMEDCT_CORE|Obstruction of artery|Arterial occlusion
C0264995|T046|IS|2929001|SNOMEDCT_CORE|Obstruction of artery, NOS|Arterial occlusion
C0264995|T046|FN|2929001|SNOMEDCT_CORE|Occlusion of artery|Arterial occlusion
C0265000|T047|SY|13954005|SNOMEDCT_CORE|Arterial ulcer|Ischemic ulcer
C0265000|T047|PTGB|13954005|SNOMEDCT_CORE|Ischaemic ulcer|Ischemic ulcer
C0265000|T047|IS|13954005|SNOMEDCT_CORE|Ischaemic ulcer, NOS|Ischemic ulcer
C0265000|T047|PT|13954005|SNOMEDCT_CORE|Ischemic ulcer|Ischemic ulcer
C0265000|T047|FN|13954005|SNOMEDCT_CORE|Ischemic ulcer|Ischemic ulcer
C0265000|T047|IS|13954005|SNOMEDCT_CORE|Ischemic ulcer, NOS|Ischemic ulcer
C0265004|T047|PT|26660001|SNOMEDCT_CORE|Dilatation of aorta|Dilatation of aorta
C0265004|T047|FN|26660001|SNOMEDCT_CORE|Dilatation of aorta|Dilatation of aorta
C0265011|T020|PT|75878002|SNOMEDCT_CORE|Abdominal aortic aneurysm without rupture|Abdominal aortic aneurysm without rupture
C0265011|T020|FN|75878002|SNOMEDCT_CORE|Abdominal aortic aneurysm without rupture|Abdominal aortic aneurysm without rupture
C0265012|T047|SY|14336007|SNOMEDCT_CORE|Abdominal aortic aneurysm which has ruptured|Ruptured abdominal aortic aneurysm
C0265012|T047|PT|14336007|SNOMEDCT_CORE|Ruptured abdominal aortic aneurysm|Ruptured abdominal aortic aneurysm
C0265012|T047|FN|14336007|SNOMEDCT_CORE|Ruptured abdominal aortic aneurysm|Ruptured abdominal aortic aneurysm
C0265012|T047|SY|14336007|SNOMEDCT_CORE|Ruptured aneurysm of abdominal aorta|Ruptured abdominal aortic aneurysm
C0265027|T047|PTGB|195381005|SNOMEDCT_CORE|Non-neoplastic naevus|Non-neoplastic nevus
C0265027|T047|PT|195381005|SNOMEDCT_CORE|Non-neoplastic nevus|Non-neoplastic nevus
C0265027|T047|FN|195381005|SNOMEDCT_CORE|Non-neoplastic nevus|Non-neoplastic nevus
C0265034|T047|SYGB|90458007|SNOMEDCT_CORE|Internal haemorrhoid|Internal hemorrhoids
C0265034|T047|PTGB|90458007|SNOMEDCT_CORE|Internal haemorrhoids|Internal hemorrhoids
C0265034|T047|SY|90458007|SNOMEDCT_CORE|Internal hemorrhoid|Internal hemorrhoids
C0265034|T047|PT|90458007|SNOMEDCT_CORE|Internal hemorrhoids|Internal hemorrhoids
C0265034|T047|FN|90458007|SNOMEDCT_CORE|Internal hemorrhoids|Internal hemorrhoids
C0265034|T047|IS|90458007|SNOMEDCT_CORE|Internal hemorrhoids, NOS|Internal hemorrhoids
C0265035|T047|PTGB|38214006|SNOMEDCT_CORE|Internal haemorrhoids without complication|Internal hemorrhoids without complication
C0265035|T047|PT|38214006|SNOMEDCT_CORE|Internal hemorrhoids without complication|Internal hemorrhoids without complication
C0265035|T047|FN|38214006|SNOMEDCT_CORE|Internal hemorrhoids without complication|Internal hemorrhoids without complication
C0265037|T047|SYGB|80426004|SNOMEDCT_CORE|Internal prolapsed haemorrhoids|Prolapsed internal hemorrhoids
C0265037|T047|SY|80426004|SNOMEDCT_CORE|Internal prolapsed hemorrhoids|Prolapsed internal hemorrhoids
C0265037|T047|PTGB|80426004|SNOMEDCT_CORE|Prolapsed internal haemorrhoids|Prolapsed internal hemorrhoids
C0265037|T047|PT|80426004|SNOMEDCT_CORE|Prolapsed internal hemorrhoids|Prolapsed internal hemorrhoids
C0265037|T047|FN|80426004|SNOMEDCT_CORE|Prolapsed internal hemorrhoids|Prolapsed internal hemorrhoids
C0265040|T047|SYGB|23913003|SNOMEDCT_CORE|External haemorrhoid|External hemorrhoids
C0265040|T047|PTGB|23913003|SNOMEDCT_CORE|External haemorrhoids|External hemorrhoids
C0265040|T047|SY|23913003|SNOMEDCT_CORE|External hemorrhoid|External hemorrhoids
C0265040|T047|FN|23913003|SNOMEDCT_CORE|External hemorrhoids|External hemorrhoids
C0265040|T047|PT|23913003|SNOMEDCT_CORE|External hemorrhoids|External hemorrhoids
C0265040|T047|IS|23913003|SNOMEDCT_CORE|External hemorrhoids, NOS|External hemorrhoids
C0265041|T047|PTGB|38996000|SNOMEDCT_CORE|External haemorrhoids without complication|External hemorrhoids without complication
C0265041|T047|SYGB|38996000|SNOMEDCT_CORE|External haemorrhoids, simple|External hemorrhoids without complication
C0265041|T047|PT|38996000|SNOMEDCT_CORE|External hemorrhoids without complication|External hemorrhoids without complication
C0265041|T047|FN|38996000|SNOMEDCT_CORE|External hemorrhoids without complication|External hemorrhoids without complication
C0265041|T047|SY|38996000|SNOMEDCT_CORE|External hemorrhoids, simple|External hemorrhoids without complication
C0265057|T047|PT|40283005|SNOMEDCT_CORE|Thrombophlebitis of superficial veins of lower extremity|Thrombophlebitis of superficial veins of lower extremity
C0265057|T047|FN|40283005|SNOMEDCT_CORE|Thrombophlebitis of superficial veins of lower extremity|Thrombophlebitis of superficial veins of lower extremity
C0265072|T047|IS|79671001|SNOMEDCT_CORE|Inferior vena cava obstruction|Inferior vena cava syndrome
C0265072|T047|PT|79671001|SNOMEDCT_CORE|Inferior vena cava syndrome|Inferior vena cava syndrome
C0265072|T047|FN|79671001|SNOMEDCT_CORE|Inferior vena cava syndrome|Inferior vena cava syndrome
C0265072|T047|IS|79671001|SNOMEDCT_CORE|IVC - Inferior vena cava obstruction|Inferior vena cava syndrome
C0265080|T047|SYGB|195176009|SNOMEDCT_CORE|Non-traumatic intracranial subdural haemorrhage|Non-traumatic subdural hemorrhage
C0265080|T047|SY|195176009|SNOMEDCT_CORE|Non-traumatic intracranial subdural hemorrhage|Non-traumatic subdural hemorrhage
C0265080|T047|FN|195176009|SNOMEDCT_CORE|Non-traumatic intracranial subdural hemorrhage|Non-traumatic subdural hemorrhage
C0265080|T047|PTGB|195176009|SNOMEDCT_CORE|Non-traumatic subdural haemorrhage|Non-traumatic subdural hemorrhage
C0265080|T047|PT|195176009|SNOMEDCT_CORE|Non-traumatic subdural hemorrhage|Non-traumatic subdural hemorrhage
C0265080|T047|IS|195176009|SNOMEDCT_CORE|Subdural haemorrhage - nontraumatic|Non-traumatic subdural hemorrhage
C0265080|T047|OF|195176009|SNOMEDCT_CORE|Subdural hemorrhage - nontraumatic|Non-traumatic subdural hemorrhage
C0265080|T047|SY|195176009|SNOMEDCT_CORE|Subdural hemorrhage - nontraumatic|Non-traumatic subdural hemorrhage
C0265089|T047|SY|1055001|SNOMEDCT_CORE|Narrowing of precerebral artery|Stenosis of precerebral artery
C0265089|T047|IS|1055001|SNOMEDCT_CORE|Narrowing of precerebral artery, NOS|Stenosis of precerebral artery
C0265089|T047|PT|1055001|SNOMEDCT_CORE|Stenosis of precerebral artery|Stenosis of precerebral artery
C0265089|T047|FN|1055001|SNOMEDCT_CORE|Stenosis of precerebral artery|Stenosis of precerebral artery
C0265089|T047|IS|1055001|SNOMEDCT_CORE|Stenosis of precerebral artery, NOS|Stenosis of precerebral artery
C0265101|T047|PT|266254007|SNOMEDCT_CORE|Carotid artery occlusion|Carotid artery occlusion
C0265101|T047|OF|266254007|SNOMEDCT_CORE|Carotid artery occlusion|Carotid artery occlusion
C0265101|T047|SY|266254007|SNOMEDCT_CORE|Occlusion of carotid artery|Carotid artery occlusion
C0265101|T047|FN|266254007|SNOMEDCT_CORE|Occlusion of carotid artery|Carotid artery occlusion
C0265103|T047|SY|90520006|SNOMEDCT_CORE|Vertebral artery narrowing|Vertebral artery stenosis
C0265103|T047|PT|90520006|SNOMEDCT_CORE|Vertebral artery stenosis|Vertebral artery stenosis
C0265103|T047|FN|90520006|SNOMEDCT_CORE|Vertebral artery stenosis|Vertebral artery stenosis
C0265122|T047|IS|55855009|SNOMEDCT_CORE|Disease of pericardium|Disorder of pericardium
C0265122|T047|OF|55855009|SNOMEDCT_CORE|Disease of pericardium|Disorder of pericardium
C0265122|T047|IS|55855009|SNOMEDCT_CORE|Disease of pericardium, NOS|Disorder of pericardium
C0265122|T047|PT|55855009|SNOMEDCT_CORE|Disorder of pericardium|Disorder of pericardium
C0265122|T047|FN|55855009|SNOMEDCT_CORE|Disorder of pericardium|Disorder of pericardium
C0265122|T047|SY|55855009|SNOMEDCT_CORE|Pericardial disorder|Disorder of pericardium
C0265122|T047|IS|55855009|SNOMEDCT_CORE|Pericardial disorder, NOS|Disorder of pericardium
C0265143|T047|PT|23627006|SNOMEDCT_CORE|Chronic pericarditis|Chronic pericarditis
C0265143|T047|FN|23627006|SNOMEDCT_CORE|Chronic pericarditis|Chronic pericarditis
C0265191|T047|PT|28590005|SNOMEDCT_CORE|Chronic acquired lymphedema|Chronic acquired lymphedema
C0265191|T047|FN|28590005|SNOMEDCT_CORE|Chronic acquired lymphedema|Chronic acquired lymphedema
C0265191|T047|PTGB|28590005|SNOMEDCT_CORE|Chronic acquired lymphoedema|Chronic acquired lymphedema
C0265191|T047|SY|28590005|SNOMEDCT_CORE|Secondary lymphedema|Chronic acquired lymphedema
C0265191|T047|SYGB|28590005|SNOMEDCT_CORE|Secondary lymphoedema|Chronic acquired lymphedema
C0265527|T019|PT|51655004|SNOMEDCT_CORE|Congenital anomaly of skull|Congenital anomaly of skull
C0265527|T019|FN|51655004|SNOMEDCT_CORE|Congenital anomaly of skull|Congenital anomaly of skull
C0265527|T019|IS|51655004|SNOMEDCT_CORE|Congenital anomaly of skull, NOS|Congenital anomaly of skull
C0265527|T019|SY|51655004|SNOMEDCT_CORE|Congenital skull malformation|Congenital anomaly of skull
C0265527|T019|IS|51655004|SNOMEDCT_CORE|Congenital skull malformation, NOS|Congenital anomaly of skull
C0265529|T019|SY|21850008|SNOMEDCT_CORE|Asymmetric head|Plagiocephaly
C0265529|T019|SY|21850008|SNOMEDCT_CORE|Lateral curvatures of skull unequal|Plagiocephaly
C0265529|T019|PT|21850008|SNOMEDCT_CORE|Plagiocephaly|Plagiocephaly
C0265529|T019|FN|21850008|SNOMEDCT_CORE|Plagiocephaly|Plagiocephaly
C0265616|T019|SY|1239002|SNOMEDCT_CORE|Congenital anteversion of femoral neck|Congenital anteversion of femur
C0265616|T019|PT|1239002|SNOMEDCT_CORE|Congenital anteversion of femur|Congenital anteversion of femur
C0265616|T019|FN|1239002|SNOMEDCT_CORE|Congenital anteversion of femur|Congenital anteversion of femur
C0265647|T019|SY|23568008|SNOMEDCT_CORE|Congenital metatarsus adductus|Metatarsus adductus
C0265647|T019|SY|23568008|SNOMEDCT_CORE|Congenital metatarsus varus|Metatarsus adductus
C0265647|T019|PT|23568008|SNOMEDCT_CORE|Metatarsus adductus|Metatarsus adductus
C0265647|T019|FN|23568008|SNOMEDCT_CORE|Metatarsus adductus|Metatarsus adductus
C0265668|T019|PT|89689008|SNOMEDCT_CORE|Congenital genu valgum|Congenital genu valgum
C0265668|T019|FN|89689008|SNOMEDCT_CORE|Congenital genu valgum|Congenital genu valgum
C0265668|T019|SY|89689008|SNOMEDCT_CORE|Congenital knock-knee|Congenital genu valgum
C0265668|T019|SY|89689008|SNOMEDCT_CORE|Congenital valgus deformity of knee|Congenital genu valgum
C0265675|T019|PT|20944008|SNOMEDCT_CORE|Congenital postural scoliosis|Congenital postural scoliosis
C0265675|T019|FN|20944008|SNOMEDCT_CORE|Congenital postural scoliosis|Congenital postural scoliosis
C0265743|T019|PT|62667002|SNOMEDCT_CORE|Congenital deviation of nasal septum|Congenital deviation of nasal septum
C0265743|T019|FN|62667002|SNOMEDCT_CORE|Congenital deviation of nasal septum|Congenital deviation of nasal septum
C0265743|T019|SY|62667002|SNOMEDCT_CORE|Congenital nasal septum deviation|Congenital deviation of nasal septum
C0265743|T019|SY|62667002|SNOMEDCT_CORE|Deviated nasal septum - congenital|Congenital deviation of nasal septum
C0265808|T047|PT|12770006|SNOMEDCT_CORE|Cyanotic congenital heart disease|Cyanotic congenital heart disease
C0265808|T047|FN|12770006|SNOMEDCT_CORE|Cyanotic congenital heart disease|Cyanotic congenital heart disease
C0265808|T047|IS|12770006|SNOMEDCT_CORE|Cyanotic congenital heart disease, NOS|Cyanotic congenital heart disease
C0265840|T019|PT|83119008|SNOMEDCT_CORE|Congenital insufficiency of tricuspid valve|Congenital insufficiency of tricuspid valve
C0265840|T047|PT|83119008|SNOMEDCT_CORE|Congenital insufficiency of tricuspid valve|Congenital insufficiency of tricuspid valve
C0265840|T019|FN|83119008|SNOMEDCT_CORE|Congenital insufficiency of tricuspid valve|Congenital insufficiency of tricuspid valve
C0265840|T047|FN|83119008|SNOMEDCT_CORE|Congenital insufficiency of tricuspid valve|Congenital insufficiency of tricuspid valve
C0265840|T019|SY|83119008|SNOMEDCT_CORE|Congenital tricuspid regurgitation|Congenital insufficiency of tricuspid valve
C0265840|T047|SY|83119008|SNOMEDCT_CORE|Congenital tricuspid regurgitation|Congenital insufficiency of tricuspid valve
C0265840|T019|SY|83119008|SNOMEDCT_CORE|TR - Congenital tricuspid regurgitation|Congenital insufficiency of tricuspid valve
C0265840|T047|SY|83119008|SNOMEDCT_CORE|TR - Congenital tricuspid regurgitation|Congenital insufficiency of tricuspid valve
C0265890|T019|SY|18546004|SNOMEDCT_CORE|Congenital aortic stenosis|Congenital stenosis of aorta
C0265890|T019|SY|21234008|SNOMEDCT_CORE|Congenital narrowed aorta|Congenital stenosis of aorta
C0265890|T019|PT|21234008|SNOMEDCT_CORE|Congenital stenosis of aorta|Congenital stenosis of aorta
C0265890|T019|FN|21234008|SNOMEDCT_CORE|Congenital stenosis of aorta|Congenital stenosis of aorta
C0265890|T019|SY|21234008|SNOMEDCT_CORE|Congenital stricture of aorta|Congenital stenosis of aorta
C0265911|T019|IS|95441000|SNOMEDCT_CORE|Congenital narrowed pulmonary artery|Congenital stenosis of pulmonary artery
C0265911|T019|IS|95441000|SNOMEDCT_CORE|Congenital stenosis of pulmonary artery|Congenital stenosis of pulmonary artery
C0265911|T019|IS|95441000|SNOMEDCT_CORE|Congenital stricture of pulmonary artery|Congenital stenosis of pulmonary artery
C0266050|T047|SY|57650002|SNOMEDCT_CORE|Deciduous teeth retained|Failure of exfoliation of primary tooth
C0266050|T047|SY|57650002|SNOMEDCT_CORE|Delayed exfoliation of deciduous tooth|Failure of exfoliation of primary tooth
C0266050|T047|SY|57650002|SNOMEDCT_CORE|Delayed exfoliation of primary teeth|Failure of exfoliation of primary tooth
C0266050|T047|SY|57650002|SNOMEDCT_CORE|Delayed shedding of deciduous tooth|Failure of exfoliation of primary tooth
C0266050|T047|PT|57650002|SNOMEDCT_CORE|Failure of exfoliation of primary tooth|Failure of exfoliation of primary tooth
C0266050|T047|SY|57650002|SNOMEDCT_CORE|Failure of resorption of root of tooth|Failure of exfoliation of primary tooth
C0266050|T047|SY|57650002|SNOMEDCT_CORE|Persistent deciduous tooth|Failure of exfoliation of primary tooth
C0266050|T047|SY|57650002|SNOMEDCT_CORE|Persistent primary tooth|Failure of exfoliation of primary tooth
C0266050|T047|FN|57650002|SNOMEDCT_CORE|Persistent primary tooth|Failure of exfoliation of primary tooth
C0266050|T047|SY|57650002|SNOMEDCT_CORE|Primary teeth retained|Failure of exfoliation of primary tooth
C0266050|T047|SY|57650002|SNOMEDCT_CORE|Prolonged retention of deciduous tooth|Failure of exfoliation of primary tooth
C0266050|T047|SY|57650002|SNOMEDCT_CORE|Retained deciduous tooth|Failure of exfoliation of primary tooth
C0266126|T019|SY|69771008|SNOMEDCT_CORE|Congenital abnormality of esophagus|Congenital anomaly of esophagus
C0266126|T019|SYGB|69771008|SNOMEDCT_CORE|Congenital abnormality of oesophagus|Congenital anomaly of esophagus
C0266126|T019|PT|69771008|SNOMEDCT_CORE|Congenital anomaly of esophagus|Congenital anomaly of esophagus
C0266126|T019|FN|69771008|SNOMEDCT_CORE|Congenital anomaly of esophagus|Congenital anomaly of esophagus
C0266126|T019|IS|69771008|SNOMEDCT_CORE|Congenital anomaly of esophagus, NOS|Congenital anomaly of esophagus
C0266126|T019|PTGB|69771008|SNOMEDCT_CORE|Congenital anomaly of oesophagus|Congenital anomaly of esophagus
C0266126|T019|SY|69771008|SNOMEDCT_CORE|Congenital malformation of the esophagus|Congenital anomaly of esophagus
C0266126|T019|SYGB|69771008|SNOMEDCT_CORE|Congenital malformation of the oesophagus|Congenital anomaly of esophagus
C0266229|T019|IS|69914001|SNOMEDCT_CORE|Congenital stricture of anus|Congenital stricture of anus
C0266294|T019|OAS|55726006|SNOMEDCT_CORE|Congenital absence of one kidney|Unilateral agenesis of kidney
C0266294|T019|OAP|55726006|SNOMEDCT_CORE|Unilateral agenesis of kidney|Unilateral agenesis of kidney
C0266294|T019|OF|55726006|SNOMEDCT_CORE|Unilateral agenesis of kidney|Unilateral agenesis of kidney
C0266294|T019|OAF|55726006|SNOMEDCT_CORE|Unilateral agenesis of kidney|Unilateral agenesis of kidney
C0266294|T019|OAS|55726006|SNOMEDCT_CORE|Unilateral congenital absence of kidney|Unilateral agenesis of kidney
C0266503|T019|SY|77224008|SNOMEDCT_CORE|Lumbar spina bifida|Spina bifida of lumbar region
C0266503|T019|FN|77224008|SNOMEDCT_CORE|Spina bifida of lumbar region|Spina bifida of lumbar region
C0266503|T019|PT|77224008|SNOMEDCT_CORE|Spina bifida of lumbar region|Spina bifida of lumbar region
C0266534|T019|PT|28550007|SNOMEDCT_CORE|Congenital capsular cataract|Congenital capsular cataract
C0266534|T019|FN|28550007|SNOMEDCT_CORE|Congenital capsular cataract|Congenital capsular cataract
C0266573|T019|PT|268163008|SNOMEDCT_CORE|Congenital ptosis|Congenital ptosis
C0266573|T019|FN|268163008|SNOMEDCT_CORE|Congenital ptosis|Congenital ptosis
C0266573|T019|SY|268163008|SNOMEDCT_CORE|Congenital ptosis of upper eyelid|Congenital ptosis
C0266611|T019|SY|35547002|SNOMEDCT_CORE|Accessory auricle|Polyotia
C0266611|T019|SY|35547002|SNOMEDCT_CORE|Accessory auricle of ear|Polyotia
C0266611|T019|PT|35547002|SNOMEDCT_CORE|Polyotia|Polyotia
C0266611|T019|FN|35547002|SNOMEDCT_CORE|Polyotia|Polyotia
C0266611|T019|SY|35547002|SNOMEDCT_CORE|Supernumerary ear|Polyotia
C0266611|T019|SY|35547002|SNOMEDCT_CORE|Supernumerary external ear|Polyotia
C0266625|T019|OAS|204271000|SNOMEDCT_CORE|Congenital preauricular sinus|Preauricular sinus
C0266625|T019|OAP|204271000|SNOMEDCT_CORE|Preauricular sinus|Preauricular sinus
C0266625|T019|OAF|204271000|SNOMEDCT_CORE|Preauricular sinus|Preauricular sinus
C0266648|T046|SY|35999006|SNOMEDCT_CORE|Anembryonic pregnancy|Blighted ovum
C0266648|T046|PT|35999006|SNOMEDCT_CORE|Blighted ovum|Blighted ovum
C0266648|T046|FN|35999006|SNOMEDCT_CORE|Blighted ovum|Blighted ovum
C0266648|T046|SY|35999006|SNOMEDCT_CORE|Empty gestational sac with ongoing pregnancy|Blighted ovum
C0266648|T046|SY|35999006|SNOMEDCT_CORE|Pathologic ovum|Blighted ovum
C0266648|T046|SY|35999006|SNOMEDCT_CORE|Resorbed fetus|Blighted ovum
C0266648|T046|SY|35999006|SNOMEDCT_CORE|Resorbed foetus|Blighted ovum
C0266764|T046|SYGB|24095001|SNOMEDCT_CORE|Partial placenta praevia|Placenta previa partialis
C0266764|T046|SY|24095001|SNOMEDCT_CORE|Partial placenta previa|Placenta previa partialis
C0266764|T046|SY|24095001|SNOMEDCT_CORE|Partial previa|Placenta previa partialis
C0266764|T046|PTGB|24095001|SNOMEDCT_CORE|Placenta praevia partialis|Placenta previa partialis
C0266764|T046|PT|24095001|SNOMEDCT_CORE|Placenta previa partialis|Placenta previa partialis
C0266764|T046|FN|24095001|SNOMEDCT_CORE|Placenta previa partialis|Placenta previa partialis
C0266771|T190|SY|91153002|SNOMEDCT_CORE|Marginal placenta|Placenta marginalis
C0266771|T190|SY|91153002|SNOMEDCT_CORE|Placenta circummarginata|Placenta marginalis
C0266771|T190|PT|91153002|SNOMEDCT_CORE|Placenta marginalis|Placenta marginalis
C0266771|T190|FN|91153002|SNOMEDCT_CORE|Placenta marginalis|Placenta marginalis
C0266771|T190|SY|91153002|SNOMEDCT_CORE|Placenta marginata|Placenta marginalis
C0266813|T033|SYGB|59614000|SNOMEDCT_CORE|Faecal occult blood positive|Occult blood in stools
C0266813|T033|OAP|167669009|SNOMEDCT_CORE|Faecal occult blood: positive|Occult blood in stools
C0266813|T033|SY|59614000|SNOMEDCT_CORE|Fecal occult blood positive|Occult blood in stools
C0266813|T033|OAP|167669009|SNOMEDCT_CORE|Fecal occult blood: positive|Occult blood in stools
C0266813|T033|OAF|167669009|SNOMEDCT_CORE|Fecal occult blood: positive|Occult blood in stools
C0266813|T033|IS|59614000|SNOMEDCT_CORE|Guaiac-positive stools|Occult blood in stools
C0266813|T033|SY|59614000|SNOMEDCT_CORE|Occult blood in stool|Occult blood in stools
C0266813|T033|PT|59614000|SNOMEDCT_CORE|Occult blood in stools|Occult blood in stools
C0266813|T033|OF|59614000|SNOMEDCT_CORE|Occult blood in stools|Occult blood in stools
C0266813|T033|FN|59614000|SNOMEDCT_CORE|Occult blood in stools|Occult blood in stools
C0266816|T047|OAP|25868003|SNOMEDCT_CORE|Soy protein sensitivity|Soy protein sensitivity
C0266816|T047|OAF|25868003|SNOMEDCT_CORE|Soy protein sensitivity|Soy protein sensitivity
C0266816|T047|OAP|25868003|SNOMEDCT_CORE|Soya protein sensitivity|Soy protein sensitivity
C0266836|T184|PT|35363006|SNOMEDCT_CORE|Infantile colic|Infantile colic
C0266836|T184|FN|35363006|SNOMEDCT_CORE|Infantile colic|Infantile colic
C0266836|T184|SY|35363006|SNOMEDCT_CORE|Infantile colic - symptom|Infantile colic
C0266836|T184|SY|35363006|SNOMEDCT_CORE|Three month colic|Infantile colic
C0266846|T047|OAP|50047001|SNOMEDCT_CORE|Compound dental caries|Dental caries extending into dentin
C0266846|T047|OAF|50047001|SNOMEDCT_CORE|Compound dental caries|Dental caries extending into dentin
C0266846|T047|OAS|50047001|SNOMEDCT_CORE|Compound dental cavity|Dental caries extending into dentin
C0266846|T047|OAS|50047001|SNOMEDCT_CORE|Dental caries confined to enamel and dentine|Dental caries extending into dentin
C0266846|T047|PT|442551007|SNOMEDCT_CORE|Dental caries extending into dentin|Dental caries extending into dentin
C0266846|T047|FN|442551007|SNOMEDCT_CORE|Dental caries extending into dentin|Dental caries extending into dentin
C0266846|T047|OAS|50047001|SNOMEDCT_CORE|Dental caries extending into dentine|Dental caries extending into dentin
C0266846|T047|SY|442551007|SNOMEDCT_CORE|Dental caries extending into dentine|Dental caries extending into dentin
C0266846|T047|OF|442551007|SNOMEDCT_CORE|Dental caries extending into dentine|Dental caries extending into dentin
C0266846|T047|OAS|50047001|SNOMEDCT_CORE|Dentin caries|Dental caries extending into dentin
C0266846|T047|SY|442551007|SNOMEDCT_CORE|Dentin caries|Dental caries extending into dentin
C0266846|T047|SY|442551007|SNOMEDCT_CORE|Dentine caries|Dental caries extending into dentin
C0266924|T047|PT|4264000|SNOMEDCT_CORE|Chronic pericoronitis|Chronic pericoronitis
C0266924|T047|FN|4264000|SNOMEDCT_CORE|Chronic pericoronitis|Chronic pericoronitis
C0266929|T047|SY|5689008|SNOMEDCT_CORE|Chronic pericementitis|Chronic periodontitis
C0266929|T047|SY|5689008|SNOMEDCT_CORE|Chronic periodontal disease|Chronic periodontitis
C0266929|T047|PT|5689008|SNOMEDCT_CORE|Chronic periodontitis|Chronic periodontitis
C0266929|T047|FN|5689008|SNOMEDCT_CORE|Chronic periodontitis|Chronic periodontitis
C0266941|T047|PT|75630004|SNOMEDCT_CORE|Derangement of temporomandibular joint|Derangement of temporomandibular joint
C0266941|T190|PT|75630004|SNOMEDCT_CORE|Derangement of temporomandibular joint|Derangement of temporomandibular joint
C0266941|T047|FN|75630004|SNOMEDCT_CORE|Derangement of temporomandibular joint|Derangement of temporomandibular joint
C0266941|T190|FN|75630004|SNOMEDCT_CORE|Derangement of temporomandibular joint|Derangement of temporomandibular joint
C0266941|T047|SY|75630004|SNOMEDCT_CORE|Temporomandibular joint derangement|Derangement of temporomandibular joint
C0266941|T190|SY|75630004|SNOMEDCT_CORE|Temporomandibular joint derangement|Derangement of temporomandibular joint
C0266941|T047|SY|75630004|SNOMEDCT_CORE|Temporomandibular joint internal derangement|Derangement of temporomandibular joint
C0266941|T190|SY|75630004|SNOMEDCT_CORE|Temporomandibular joint internal derangement|Derangement of temporomandibular joint
C0266950|T047|PT|44402007|SNOMEDCT_CORE|Loss of teeth due to extraction|Loss of teeth due to extraction
C0266950|T047|FN|44402007|SNOMEDCT_CORE|Loss of teeth due to extraction|Loss of teeth due to extraction
C0266950|T047|SY|44402007|SNOMEDCT_CORE|Surgical edentia|Loss of teeth due to extraction
C0266980|T047|SY|11625007|SNOMEDCT_CORE|Lingual torus|Torus mandibularis
C0266980|T047|FN|11625007|SNOMEDCT_CORE|Torus mandibularis|Torus mandibularis
C0266980|T047|PT|11625007|SNOMEDCT_CORE|Torus mandibularis|Torus mandibularis
C0266989|T047|IS|42982001|SNOMEDCT_CORE|Sialoangitis, NOS|Sialoangitis, NOS
C0266998|T047|IS|41188003|SNOMEDCT_CORE|Disease of oral soft tissues|Disorder of oral soft tissues
C0266998|T047|OF|41188003|SNOMEDCT_CORE|Disease of oral soft tissues|Disorder of oral soft tissues
C0266998|T047|SY|41188003|SNOMEDCT_CORE|Disease of the oral soft tissues|Disorder of oral soft tissues
C0266998|T047|IS|41188003|SNOMEDCT_CORE|Disease of the oral soft tissues, NOS|Disorder of oral soft tissues
C0266998|T047|PT|41188003|SNOMEDCT_CORE|Disorder of oral soft tissues|Disorder of oral soft tissues
C0266998|T047|FN|41188003|SNOMEDCT_CORE|Disorder of oral soft tissues|Disorder of oral soft tissues
C0266998|T047|SY|41188003|SNOMEDCT_CORE|Oral soft tissue disease|Disorder of oral soft tissues
C0267026|T047|PT|46795000|SNOMEDCT_CORE|Actinic cheilitis|Actinic cheilitis
C0267026|T047|FN|46795000|SNOMEDCT_CORE|Actinic cheilitis|Actinic cheilitis
C0267026|T047|SY|46795000|SNOMEDCT_CORE|Solar keratosis of lip|Actinic cheilitis
C0267071|T047|PT|71457002|SNOMEDCT_CORE|Oropharyngeal dysphagia|Oropharyngeal dysphagia
C0267071|T047|FN|71457002|SNOMEDCT_CORE|Oropharyngeal dysphagia|Oropharyngeal dysphagia
C0267071|T047|IS|71457002|SNOMEDCT_CORE|Pharyngeal dysphagia|Oropharyngeal dysphagia
C0267071|T047|SY|71457002|SNOMEDCT_CORE|Transfer dysphagia|Oropharyngeal dysphagia
C0267072|T047|PT|40890009|SNOMEDCT_CORE|Esophageal dysphagia|Esophageal dysphagia
C0267072|T047|FN|40890009|SNOMEDCT_CORE|Esophageal dysphagia|Esophageal dysphagia
C0267072|T047|PTGB|40890009|SNOMEDCT_CORE|Oesophageal dysphagia|Esophageal dysphagia
C0267081|T047|SY|66889002|SNOMEDCT_CORE|Acquired Schatzki's ring|Terminal esophageal web
C0267081|T047|SY|66889002|SNOMEDCT_CORE|Esophageal ring|Terminal esophageal web
C0267081|T047|SY|66889002|SNOMEDCT_CORE|LOMR - Lower esophageal mucosal ring|Terminal esophageal web
C0267081|T047|SYGB|66889002|SNOMEDCT_CORE|LOMR - Lower oesophageal mucosal ring|Terminal esophageal web
C0267081|T047|SY|66889002|SNOMEDCT_CORE|Lower esophageal mucosal ring|Terminal esophageal web
C0267081|T047|SYGB|66889002|SNOMEDCT_CORE|Lower oesophageal mucosal ring|Terminal esophageal web
C0267081|T047|SYGB|66889002|SNOMEDCT_CORE|Oesophageal ring|Terminal esophageal web
C0267081|T047|SY|66889002|SNOMEDCT_CORE|Schatzki ring|Terminal esophageal web
C0267081|T047|SY|66889002|SNOMEDCT_CORE|Schatzki's ring|Terminal esophageal web
C0267081|T047|SY|66889002|SNOMEDCT_CORE|SR - Schatzki ring|Terminal esophageal web
C0267081|T047|SY|66889002|SNOMEDCT_CORE|Terminal esophageal ring|Terminal esophageal web
C0267081|T047|PT|66889002|SNOMEDCT_CORE|Terminal esophageal web|Terminal esophageal web
C0267081|T047|FN|66889002|SNOMEDCT_CORE|Terminal esophageal web|Terminal esophageal web
C0267081|T047|SYGB|66889002|SNOMEDCT_CORE|Terminal oesophageal ring|Terminal esophageal web
C0267081|T047|PTGB|66889002|SNOMEDCT_CORE|Terminal oesophageal web|Terminal esophageal web
C0267092|T047|PT|14223005|SNOMEDCT_CORE|Esophageal varices without bleeding|Esophageal varices without bleeding
C0267092|T047|FN|14223005|SNOMEDCT_CORE|Esophageal varices without bleeding|Esophageal varices without bleeding
C0267092|T047|PTGB|14223005|SNOMEDCT_CORE|Oesophageal varices without bleeding|Esophageal varices without bleeding
C0267112|T047|SY|18665000|SNOMEDCT_CORE|Acute erosion of stomach|Acute gastric mucosal erosion
C0267112|T047|IS|18665000|SNOMEDCT_CORE|Acute erosive gastritis|Acute gastric mucosal erosion
C0267112|T047|PT|18665000|SNOMEDCT_CORE|Acute gastric mucosal erosion|Acute gastric mucosal erosion
C0267112|T047|FN|18665000|SNOMEDCT_CORE|Acute gastric mucosal erosion|Acute gastric mucosal erosion
C0267112|T047|IS|18665000|SNOMEDCT_CORE|Acute gastric mucosal erosion, NOS|Acute gastric mucosal erosion
C0267127|T047|SY|57246001|SNOMEDCT_CORE|Bleeding chronic gastric ulcer|Chronic gastric ulcer with hemorrhage
C0267127|T047|PTGB|57246001|SNOMEDCT_CORE|Chronic gastric ulcer with haemorrhage|Chronic gastric ulcer with hemorrhage
C0267127|T047|PT|57246001|SNOMEDCT_CORE|Chronic gastric ulcer with hemorrhage|Chronic gastric ulcer with hemorrhage
C0267127|T047|FN|57246001|SNOMEDCT_CORE|Chronic gastric ulcer with hemorrhage|Chronic gastric ulcer with hemorrhage
C0267130|T047|PT|31301004|SNOMEDCT_CORE|Chronic gastric ulcer with perforation|Chronic gastric ulcer with perforation
C0267130|T047|FN|31301004|SNOMEDCT_CORE|Chronic gastric ulcer with perforation|Chronic gastric ulcer with perforation
C0267130|T047|SY|31301004|SNOMEDCT_CORE|Perforated chronic gastric ulcer|Chronic gastric ulcer with perforation
C0267142|T047|PTGB|59913009|SNOMEDCT_CORE|Gastric ulcer without haemorrhage, without perforation AND without obstruction|Gastric ulcer without hemorrhage, without perforation AND without obstruction
C0267142|T047|PT|59913009|SNOMEDCT_CORE|Gastric ulcer without hemorrhage, without perforation AND without obstruction|Gastric ulcer without hemorrhage, without perforation AND without obstruction
C0267142|T047|FN|59913009|SNOMEDCT_CORE|Gastric ulcer without hemorrhage, without perforation AND without obstruction|Gastric ulcer without hemorrhage, without perforation AND without obstruction
C0267142|T047|IS|59913009|SNOMEDCT_CORE|Gastric ulcer, NOS without hemorrhage or perforation and without obstruction|Gastric ulcer without hemorrhage, without perforation AND without obstruction
C0267166|T047|SY|196731005|SNOMEDCT_CORE|Gastritis and duodenitis|Gastroduodenitis
C0267166|T047|OF|196731005|SNOMEDCT_CORE|Gastritis and duodenitis|Gastroduodenitis
C0267166|T047|PT|196731005|SNOMEDCT_CORE|Gastroduodenitis|Gastroduodenitis
C0267166|T047|FN|196731005|SNOMEDCT_CORE|Gastroduodenitis|Gastroduodenitis
C0267167|T033|SY|3696007|SNOMEDCT_CORE|Functional dyspepsia|Nonulcer dyspepsia
C0267167|T033|SY|3696007|SNOMEDCT_CORE|Non ulcer dyspepsia|Nonulcer dyspepsia
C0267167|T033|SY|3696007|SNOMEDCT_CORE|Non-ulcer dyspepsia|Nonulcer dyspepsia
C0267167|T033|PT|3696007|SNOMEDCT_CORE|Nonulcer dyspepsia|Nonulcer dyspepsia
C0267167|T033|FN|3696007|SNOMEDCT_CORE|Nonulcer dyspepsia|Nonulcer dyspepsia
C0267174|T047|SY|13267003|SNOMEDCT_CORE|Gastric motor dysfunction|Gastric motor function disorder
C0267174|T047|IS|13267003|SNOMEDCT_CORE|Gastric motor dysfunction, NOS|Gastric motor function disorder
C0267174|T047|PT|13267003|SNOMEDCT_CORE|Gastric motor function disorder|Gastric motor function disorder
C0267174|T047|FN|13267003|SNOMEDCT_CORE|Gastric motor function disorder|Gastric motor function disorder
C0267174|T047|IS|13267003|SNOMEDCT_CORE|Gastric motor function disorder, NOS|Gastric motor function disorder
C0267174|T047|SY|13267003|SNOMEDCT_CORE|Idiopathic gastric motility disorder|Gastric motor function disorder
C0267176|T047|OAP|34140002|SNOMEDCT_CORE|Diabetic gastroparesis|Gastroparesis due to diabetes mellitus
C0267176|T047|OAF|34140002|SNOMEDCT_CORE|Diabetic gastroparesis|Gastroparesis due to diabetes mellitus
C0267176|T047|OF|713704004|SNOMEDCT_CORE|Gastroparesis co-occurrent and due to diabetes mellitus|Gastroparesis due to diabetes mellitus
C0267176|T047|IS|713704004|SNOMEDCT_CORE|Gastroparesis co-occurrent and due to diabetes mellitus|Gastroparesis due to diabetes mellitus
C0267176|T047|PT|713704004|SNOMEDCT_CORE|Gastroparesis due to diabetes mellitus|Gastroparesis due to diabetes mellitus
C0267176|T047|FN|713704004|SNOMEDCT_CORE|Gastroparesis due to diabetes mellitus|Gastroparesis due to diabetes mellitus
C0267176|T047|SY|713704004|SNOMEDCT_CORE|Gastroparesis with diabetes mellitus|Gastroparesis due to diabetes mellitus
C0267209|T047|PT|24807004|SNOMEDCT_CORE|Bleeding gastric varices|Bleeding gastric varices
C0267209|T047|FN|24807004|SNOMEDCT_CORE|Bleeding gastric varices|Bleeding gastric varices
C0267211|T020|SY|43935004|SNOMEDCT_CORE|GAVE - Gastric antral vascular ectasia|Vascular ectasia of gastric antrum
C0267211|T020|PT|43935004|SNOMEDCT_CORE|Vascular ectasia of gastric antrum|Vascular ectasia of gastric antrum
C0267211|T020|FN|43935004|SNOMEDCT_CORE|Vascular ectasia of gastric antrum|Vascular ectasia of gastric antrum
C0267211|T020|SY|43935004|SNOMEDCT_CORE|Watermelon stomach|Vascular ectasia of gastric antrum
C0267211|T020|OF|43935004|SNOMEDCT_CORE|Watermelon stomach|Vascular ectasia of gastric antrum
C0267267|T046|SY|89469000|SNOMEDCT_CORE|Bleeding chronic duodenal ulcer|Chronic duodenal ulcer with hemorrhage
C0267267|T046|PTGB|89469000|SNOMEDCT_CORE|Chronic duodenal ulcer with haemorrhage|Chronic duodenal ulcer with hemorrhage
C0267267|T046|PT|89469000|SNOMEDCT_CORE|Chronic duodenal ulcer with hemorrhage|Chronic duodenal ulcer with hemorrhage
C0267267|T046|FN|89469000|SNOMEDCT_CORE|Chronic duodenal ulcer with hemorrhage|Chronic duodenal ulcer with hemorrhage
C0267272|T047|PT|49916007|SNOMEDCT_CORE|Chronic duodenal ulcer with perforation|Chronic duodenal ulcer with perforation
C0267272|T047|FN|49916007|SNOMEDCT_CORE|Chronic duodenal ulcer with perforation|Chronic duodenal ulcer with perforation
C0267272|T047|SY|49916007|SNOMEDCT_CORE|Perforated chronic duodenal ulcer|Chronic duodenal ulcer with perforation
C0267288|T047|PTGB|12274003|SNOMEDCT_CORE|Acute peptic ulcer with haemorrhage|Acute peptic ulcer with hemorrhage
C0267288|T047|PT|12274003|SNOMEDCT_CORE|Acute peptic ulcer with hemorrhage|Acute peptic ulcer with hemorrhage
C0267288|T047|FN|12274003|SNOMEDCT_CORE|Acute peptic ulcer with hemorrhage|Acute peptic ulcer with hemorrhage
C0267300|T047|PTGB|49232000|SNOMEDCT_CORE|Chronic peptic ulcer with haemorrhage|Chronic peptic ulcer with hemorrhage
C0267300|T047|PT|49232000|SNOMEDCT_CORE|Chronic peptic ulcer with hemorrhage|Chronic peptic ulcer with hemorrhage
C0267300|T047|FN|49232000|SNOMEDCT_CORE|Chronic peptic ulcer with hemorrhage|Chronic peptic ulcer with hemorrhage
C0267319|T047|PTGB|38365000|SNOMEDCT_CORE|Peptic ulcer without haemorrhage, without perforation AND without obstruction|Peptic ulcer without hemorrhage, without perforation AND without obstruction
C0267319|T047|PT|38365000|SNOMEDCT_CORE|Peptic ulcer without hemorrhage, without perforation AND without obstruction|Peptic ulcer without hemorrhage, without perforation AND without obstruction
C0267319|T047|FN|38365000|SNOMEDCT_CORE|Peptic ulcer without hemorrhage, without perforation AND without obstruction|Peptic ulcer without hemorrhage, without perforation AND without obstruction
C0267319|T047|IS|38365000|SNOMEDCT_CORE|Peptic ulcer, NOS without hemorrhage or perforation and without obstruction|Peptic ulcer without hemorrhage, without perforation AND without obstruction
C0267364|T191|PT|89452002|SNOMEDCT_CORE|Hyperplastic polyp of intestine|Hyperplastic polyp of intestine
C0267364|T191|FN|89452002|SNOMEDCT_CORE|Hyperplastic polyp of intestine|Hyperplastic polyp of intestine
C0267364|T191|IS|89452002|SNOMEDCT_CORE|Hyperplastic polyp of intestine, NOS|Hyperplastic polyp of intestine
C0267364|T191|SY|89452002|SNOMEDCT_CORE|Metaplastic polyp of intestine|Hyperplastic polyp of intestine
C0267364|T191|IS|89452002|SNOMEDCT_CORE|Metaplastic polyp of intestine, NOS|Hyperplastic polyp of intestine
C0267367|T047|PT|235853006|SNOMEDCT_CORE|Angiodysplasia of intestine|Angiodysplasia of intestine
C0267367|T047|FN|235853006|SNOMEDCT_CORE|Angiodysplasia of intestine|Angiodysplasia of intestine
C0267367|T047|SY|235853006|SNOMEDCT_CORE|Intestinal vascular dysplasia|Angiodysplasia of intestine
C0267380|T047|SY|38106008|SNOMEDCT_CORE|Crohn disease of ileum|Crohn's disease of ileum
C0267380|T047|PT|38106008|SNOMEDCT_CORE|Crohn's disease of ileum|Crohn's disease of ileum
C0267380|T047|FN|38106008|SNOMEDCT_CORE|Crohn's disease of ileum|Crohn's disease of ileum
C0267380|T047|SY|38106008|SNOMEDCT_CORE|Crohn's ileitis|Crohn's disease of ileum
C0267383|T047|SY|71833008|SNOMEDCT_CORE|Crohn disease of small AND large intestines|Regional ileocolitis
C0267383|T047|IS|71833008|SNOMEDCT_CORE|Crohn's disease of small and large intestines|Regional ileocolitis
C0267383|T047|FN|71833008|SNOMEDCT_CORE|Crohn's disease of small AND large intestines|Regional ileocolitis
C0267383|T047|PT|71833008|SNOMEDCT_CORE|Crohn's disease of small AND large intestines|Regional ileocolitis
C0267383|T047|SY|71833008|SNOMEDCT_CORE|Crohn's disease of small intestine and colon|Regional ileocolitis
C0267383|T047|FN|196983007|SNOMEDCT_CORE|Regional ileocolitis|Regional ileocolitis
C0267383|T047|IS|71833008|SNOMEDCT_CORE|Regional ileocolitis|Regional ileocolitis
C0267383|T047|PT|196983007|SNOMEDCT_CORE|Regional ileocolitis|Regional ileocolitis
C0267390|T047|SY|52506002|SNOMEDCT_CORE|Chronic ulcerative proctosigmoiditis|Chronic ulcerative rectosigmoiditis
C0267390|T047|PT|52506002|SNOMEDCT_CORE|Chronic ulcerative rectosigmoiditis|Chronic ulcerative rectosigmoiditis
C0267390|T047|FN|52506002|SNOMEDCT_CORE|Chronic ulcerative rectosigmoiditis|Chronic ulcerative rectosigmoiditis
C0267390|T047|SY|52506002|SNOMEDCT_CORE|Ulcerative colitis confined to rectum and sigmoid colon|Chronic ulcerative rectosigmoiditis
C0267390|T047|SY|52506002|SNOMEDCT_CORE|Ulcerative proctosigmoiditis|Chronic ulcerative rectosigmoiditis
C0267390|T047|SY|52506002|SNOMEDCT_CORE|Ulcerative rectosigmoiditis|Chronic ulcerative rectosigmoiditis
C0267412|T046|PT|95446005|SNOMEDCT_CORE|Thrombosis of mesenteric vein|Thrombosis of mesenteric vein
C0267412|T046|FN|95446005|SNOMEDCT_CORE|Thrombosis of mesenteric vein|Thrombosis of mesenteric vein
C0267418|T047|PT|12574004|SNOMEDCT_CORE|Noninfectious gastroenteritis|Noninfectious gastroenteritis
C0267418|T047|FN|12574004|SNOMEDCT_CORE|Noninfectious gastroenteritis|Noninfectious gastroenteritis
C0267418|T047|IS|12574004|SNOMEDCT_CORE|Noninfectious gastroenteritis, NOS|Noninfectious gastroenteritis
C0267465|T047|PT|56226004|SNOMEDCT_CORE|Stricture of intestine|Stricture of intestine
C0267465|T047|FN|56226004|SNOMEDCT_CORE|Stricture of intestine|Stricture of intestine
C0267478|T047|PT|67766009|SNOMEDCT_CORE|Intestinal adhesions with obstruction|Intestinal adhesions with obstruction
C0267478|T047|FN|67766009|SNOMEDCT_CORE|Intestinal adhesions with obstruction|Intestinal adhesions with obstruction
C0267510|T047|PT|85920003|SNOMEDCT_CORE|Constipation by outlet obstruction|Constipation by outlet obstruction
C0267510|T047|OF|85920003|SNOMEDCT_CORE|Constipation by outlet obstruction|Constipation by outlet obstruction
C0267510|T047|SY|85920003|SNOMEDCT_CORE|Constipation due to outlet obstruction|Constipation by outlet obstruction
C0267510|T047|FN|85920003|SNOMEDCT_CORE|Constipation due to outlet obstruction|Constipation by outlet obstruction
C0267561|T190|SY|58103005|SNOMEDCT_CORE|Fistula of perianal skin|Perianal fistula
C0267561|T190|PT|58103005|SNOMEDCT_CORE|Perianal fistula|Perianal fistula
C0267561|T190|FN|58103005|SNOMEDCT_CORE|Perianal fistula|Perianal fistula
C0267566|T046|PT|91669008|SNOMEDCT_CORE|Perirectal abscess|Perirectal abscess
C0267566|T046|FN|91669008|SNOMEDCT_CORE|Perirectal abscess|Perirectal abscess
C0267572|T047|PT|67038005|SNOMEDCT_CORE|Nonspecific ulcerative proctitis|Nonspecific ulcerative proctitis
C0267572|T047|FN|67038005|SNOMEDCT_CORE|Nonspecific ulcerative proctitis|Nonspecific ulcerative proctitis
C0267573|T191|PT|88580009|SNOMEDCT_CORE|Anal polyp|Anal polyp
C0267573|T191|FN|88580009|SNOMEDCT_CORE|Anal polyp|Anal polyp
C0267596|T046|SY|12063002|SNOMEDCT_CORE|Bleeding per rectum|Rectal hemorrhage
C0267596|T046|SY|12063002|SNOMEDCT_CORE|Blood per rectum|Rectal hemorrhage
C0267596|T046|IS|12063002|SNOMEDCT_CORE|Hemorrhage of rectum|Rectal hemorrhage
C0267596|T046|SY|12063002|SNOMEDCT_CORE|PR - Bleeding per rectum|Rectal hemorrhage
C0267596|T046|SY|12063002|SNOMEDCT_CORE|PR - Blood per rectum|Rectal hemorrhage
C0267596|T046|SY|12063002|SNOMEDCT_CORE|PRB - Rectal bleeding|Rectal hemorrhage
C0267596|T046|SY|12063002|SNOMEDCT_CORE|Proctorrhagia|Rectal hemorrhage
C0267596|T046|SY|12063002|SNOMEDCT_CORE|RB - Rectal bleeding|Rectal hemorrhage
C0267596|T046|SY|12063002|SNOMEDCT_CORE|Rectal bleeding|Rectal hemorrhage
C0267596|T046|PTGB|12063002|SNOMEDCT_CORE|Rectal haemorrhage|Rectal hemorrhage
C0267596|T046|PT|12063002|SNOMEDCT_CORE|Rectal hemorrhage|Rectal hemorrhage
C0267596|T046|FN|12063002|SNOMEDCT_CORE|Rectal hemorrhage|Rectal hemorrhage
C0267596|T046|SY|12063002|SNOMEDCT_CORE|Rectorrhagia|Rectal hemorrhage
C0267613|T047|IS|18526009|SNOMEDCT_CORE|Disease of appendix|Disorder of appendix
C0267613|T047|OF|18526009|SNOMEDCT_CORE|Disease of appendix|Disorder of appendix
C0267613|T047|IS|18526009|SNOMEDCT_CORE|Disease of appendix, NOS|Disorder of appendix
C0267613|T047|PT|18526009|SNOMEDCT_CORE|Disorder of appendix|Disorder of appendix
C0267613|T047|FN|18526009|SNOMEDCT_CORE|Disorder of appendix|Disorder of appendix
C0267664|T046|PT|17551007|SNOMEDCT_CORE|Chronic diarrhea of unknown origin|Chronic diarrhea of unknown origin
C0267664|T046|FN|17551007|SNOMEDCT_CORE|Chronic diarrhea of unknown origin|Chronic diarrhea of unknown origin
C0267664|T046|PTGB|17551007|SNOMEDCT_CORE|Chronic diarrhoea of unknown origin|Chronic diarrhea of unknown origin
C0267672|T047|PT|85502002|SNOMEDCT_CORE|Bilateral inguinal hernia|Bilateral inguinal hernia
C0267672|T047|FN|85502002|SNOMEDCT_CORE|Bilateral inguinal hernia|Bilateral inguinal hernia
C0267704|T020|OAF|7544003|SNOMEDCT_CORE|Umbilical hernia without obstruction AND without gangrene|Umbilical hernia without obstruction AND without gangrene
C0267704|T020|OAP|7544003|SNOMEDCT_CORE|Umbilical hernia without obstruction AND without gangrene|Umbilical hernia without obstruction AND without gangrene
C0267704|T020|IS|7544003|SNOMEDCT_CORE|Umbilical hernia without obstruction or gangrene|Umbilical hernia without obstruction AND without gangrene
C0267716|T046|PT|236037000|SNOMEDCT_CORE|Incisional hernia|Incisional hernia
C0267716|T046|FN|236037000|SNOMEDCT_CORE|Incisional hernia|Incisional hernia
C0267771|T047|SY|69559004|SNOMEDCT_CORE|Mass of retroperitoneal structure|Retroperitoneal mass
C0267771|T047|FN|69559004|SNOMEDCT_CORE|Mass of retroperitoneal structure|Retroperitoneal mass
C0267771|T047|PT|69559004|SNOMEDCT_CORE|Retroperitoneal mass|Retroperitoneal mass
C0267771|T047|OF|69559004|SNOMEDCT_CORE|Retroperitoneal mass|Retroperitoneal mass
C0267797|T047|PT|37871000|SNOMEDCT_CORE|Acute hepatitis|Acute hepatitis
C0267797|T047|FN|37871000|SNOMEDCT_CORE|Acute hepatitis|Acute hepatitis
C0267797|T047|IS|37871000|SNOMEDCT_CORE|Acute hepatitis, NOS|Acute hepatitis
C0267809|T047|PT|89580002|SNOMEDCT_CORE|Cryptogenic cirrhosis|Cryptogenic cirrhosis
C0267809|T047|FN|89580002|SNOMEDCT_CORE|Cryptogenic cirrhosis|Cryptogenic cirrhosis
C0267834|T047|SY|85057007|SNOMEDCT_CORE|Cyst of liver|Liver cyst
C0267834|T047|FN|85057007|SNOMEDCT_CORE|Cyst of liver|Liver cyst
C0267834|T047|SY|85057007|SNOMEDCT_CORE|Hepatic cyst|Liver cyst
C0267834|T047|PT|85057007|SNOMEDCT_CORE|Liver cyst|Liver cyst
C0267834|T047|OF|85057007|SNOMEDCT_CORE|Liver cyst|Liver cyst
C0267853|T047|PT|25924004|SNOMEDCT_CORE|Calculus of gallbladder with cholecystitis|Calculus of gallbladder with cholecystitis
C0267853|T047|FN|25924004|SNOMEDCT_CORE|Calculus of gallbladder with cholecystitis|Calculus of gallbladder with cholecystitis
C0267853|T047|IS|25924004|SNOMEDCT_CORE|Calculus of gallbladder with cholecystitis, NOS|Calculus of gallbladder with cholecystitis
C0267853|T047|SY|25924004|SNOMEDCT_CORE|Cholelithiasis with cholecystitis|Calculus of gallbladder with cholecystitis
C0267853|T047|IS|25924004|SNOMEDCT_CORE|Cholelithiasis with cholecystitis, NOS|Calculus of gallbladder with cholecystitis
C0267861|T047|PT|70342003|SNOMEDCT_CORE|Cholelithiasis without obstruction|Cholelithiasis without obstruction
C0267861|T047|FN|70342003|SNOMEDCT_CORE|Cholelithiasis without obstruction|Cholelithiasis without obstruction
C0267861|T047|SY|70342003|SNOMEDCT_CORE|Cholelithiasis, non obstructive|Cholelithiasis without obstruction
C0267871|T047|PT|4661003|SNOMEDCT_CORE|Calculus of bile duct with obstruction|Calculus of bile duct with obstruction
C0267871|T047|FN|4661003|SNOMEDCT_CORE|Calculus of bile duct with obstruction|Calculus of bile duct with obstruction
C0267917|T047|PT|6215006|SNOMEDCT_CORE|Acute cholangitis|Acute cholangitis
C0267917|T047|FN|6215006|SNOMEDCT_CORE|Acute cholangitis|Acute cholangitis
C0267920|T047|PT|65001009|SNOMEDCT_CORE|Recurrent pyogenic cholangitis|Recurrent pyogenic cholangitis
C0267920|T047|FN|65001009|SNOMEDCT_CORE|Recurrent pyogenic cholangitis|Recurrent pyogenic cholangitis
C0267922|T047|PT|10184002|SNOMEDCT_CORE|Recurrent cholangitis|Recurrent cholangitis
C0267922|T047|FN|10184002|SNOMEDCT_CORE|Recurrent cholangitis|Recurrent cholangitis
C0267937|T047|PT|197458008|SNOMEDCT_CORE|Acute recurrent pancreatitis|Acute recurrent pancreatitis
C0267937|T047|FN|197458008|SNOMEDCT_CORE|Acute recurrent pancreatitis|Acute recurrent pancreatitis
C0267988|T047|PTGB|37064009|SNOMEDCT_CORE|Hyperproteinaemia|Hyperproteinemia
C0267988|T047|PT|37064009|SNOMEDCT_CORE|Hyperproteinemia|Hyperproteinemia
C0267988|T047|FN|37064009|SNOMEDCT_CORE|Hyperproteinemia|Hyperproteinemia
C0267988|T047|IS|37064009|SNOMEDCT_CORE|Hyperproteinemia, NOS|Hyperproteinemia
C0268000|T046|PT|43498006|SNOMEDCT_CORE|Body fluid retention|Body fluid retention
C0268000|T046|FN|43498006|SNOMEDCT_CORE|Body fluid retention|Body fluid retention
C0268000|T046|IS|43498006|SNOMEDCT_CORE|Fluid retention|Body fluid retention
C0268108|T047|FN|68451005|SNOMEDCT_CORE|Chronic arthritis due to gout|Chronic gouty arthritis
C0268108|T047|SY|68451005|SNOMEDCT_CORE|Chronic arthritis due to gout|Chronic gouty arthritis
C0268108|T047|PT|68451005|SNOMEDCT_CORE|Chronic gouty arthritis|Chronic gouty arthritis
C0268108|T047|OF|68451005|SNOMEDCT_CORE|Chronic gouty arthritis|Chronic gouty arthritis
C0268109|T047|PT|73877009|SNOMEDCT_CORE|Chronic tophaceous gout|Chronic tophaceous gout
C0268109|T047|FN|73877009|SNOMEDCT_CORE|Chronic tophaceous gout|Chronic tophaceous gout
C0268366|T047|SYGB|58588007|SNOMEDCT_CORE|Generalised elastorrhexis|Systematized elastorrhexis
C0268366|T047|SY|58588007|SNOMEDCT_CORE|Generalized elastorrhexis|Systematized elastorrhexis
C0268366|T047|SYGB|58588007|SNOMEDCT_CORE|Systematised elastorrhexis|Systematized elastorrhexis
C0268366|T047|SY|58588007|SNOMEDCT_CORE|Systematized elastorrhexis|Systematized elastorrhexis
C0268366|T047|SY|58588007|SNOMEDCT_CORE|Systemic elastorrhexis|Systematized elastorrhexis
C0268392|T047|PTGB|56871000|SNOMEDCT_CORE|Localised amyloidosis|Localized amyloidosis
C0268392|T047|PT|56871000|SNOMEDCT_CORE|Localized amyloidosis|Localized amyloidosis
C0268392|T047|FN|56871000|SNOMEDCT_CORE|Localized amyloidosis|Localized amyloidosis
C0268392|T047|IS|56871000|SNOMEDCT_CORE|Localized amyloidosis, NOS|Localized amyloidosis
C0268617|T047|PTGB|52311001|SNOMEDCT_CORE|Homocystinaemia|Homocystinemia
C0268617|T047|PT|52311001|SNOMEDCT_CORE|Homocystinemia|Homocystinemia
C0268617|T047|FN|52311001|SNOMEDCT_CORE|Homocystinemia|Homocystinemia
C0268617|T047|IS|52311001|SNOMEDCT_CORE|Homocystinemia, NOS|Homocystinemia
C0268679|T047|SY|64117007|SNOMEDCT_CORE|Cyanocobalamine deficiency|Vitamin B12 deficiency
C0268679|T047|SYGB|64117007|SNOMEDCT_CORE|Cyanocobalamine deficiency|Vitamin B12 deficiency
C0268679|T047|PT|64117007|SNOMEDCT_CORE|Vitamin B12 deficiency|Vitamin B12 deficiency
C0268679|T047|PTGB|64117007|SNOMEDCT_CORE|Vitamin B12 deficiency|Vitamin B12 deficiency
C0268679|T047|FN|64117007|SNOMEDCT_CORE|Vitamin B12 deficiency|Vitamin B12 deficiency
C0268769|T047|PT|190829000|SNOMEDCT_CORE|Chronic gouty nephropathy|Chronic gouty nephropathy
C0268769|T047|SY|190829000|SNOMEDCT_CORE|Chronic urate nephropathy|Chronic gouty nephropathy
C0268769|T047|FN|190829000|SNOMEDCT_CORE|Chronic urate nephropathy|Chronic gouty nephropathy
C0268781|T047|PT|11480007|SNOMEDCT_CORE|Idiopathic granulomatous interstitial nephropathy|Idiopathic granulomatous interstitial nephropathy
C0268781|T047|FN|11480007|SNOMEDCT_CORE|Idiopathic granulomatous interstitial nephropathy|Idiopathic granulomatous interstitial nephropathy
C0268781|T047|IS|11480007|SNOMEDCT_CORE|Idiopathic granulomatous interstitial nephropathy, NOS|Idiopathic granulomatous interstitial nephropathy
C0268800|T047|IS|77945009|SNOMEDCT_CORE|Cyst of kidney|Simple renal cyst
C0268800|T047|IS|77945009|SNOMEDCT_CORE|Renal cyst|Simple renal cyst
C0268800|T047|SY|77945009|SNOMEDCT_CORE|Simple cyst of kidney|Simple renal cyst
C0268800|T047|PT|77945009|SNOMEDCT_CORE|Simple renal cyst|Simple renal cyst
C0268800|T047|FN|77945009|SNOMEDCT_CORE|Simple renal cyst|Simple renal cyst
C0268800|T047|SY|77945009|SNOMEDCT_CORE|Single renal cyst|Simple renal cyst
C0268804|T047|PT|40068008|SNOMEDCT_CORE|Hydroureteronephrosis|Hydroureteronephrosis
C0268804|T047|FN|40068008|SNOMEDCT_CORE|Hydroureteronephrosis|Hydroureteronephrosis
C0268821|T047|SY|4009004|SNOMEDCT_CORE|Lower urinary tract infection|Lower urinary tract infectious disease
C0268821|T047|PT|4009004|SNOMEDCT_CORE|Lower urinary tract infectious disease|Lower urinary tract infectious disease
C0268821|T047|FN|4009004|SNOMEDCT_CORE|Lower urinary tract infectious disease|Lower urinary tract infectious disease
C0268821|T047|IS|4009004|SNOMEDCT_CORE|Lower urinary tract infectious disease, NOS|Lower urinary tract infectious disease
C0268821|T047|SY|4009004|SNOMEDCT_CORE|UTI - Lower urinary tract infection|Lower urinary tract infectious disease
C0268842|T047|SY|28626004|SNOMEDCT_CORE|Colovesical fistula|Vesicocolic fistula
C0268842|T047|SY|28626004|SNOMEDCT_CORE|CVF - Colovesical fistula|Vesicocolic fistula
C0268842|T047|PT|28626004|SNOMEDCT_CORE|Vesicocolic fistula|Vesicocolic fistula
C0268842|T047|FN|28626004|SNOMEDCT_CORE|Vesicocolic fistula|Vesicocolic fistula
C0268848|T047|IS|79184009|SNOMEDCT_CORE|Increased trabeculation of bladder|Increased trabeculation of bladder
C0268849|T047|PT|786460007|SNOMEDCT_CORE|Detrusor overactivity|Detrusor overactivity
C0268849|T047|FN|786460007|SNOMEDCT_CORE|Detrusor overactivity|Detrusor overactivity
C0268849|T047|OAS|236633002|SNOMEDCT_CORE|Overactive detrusor|Detrusor overactivity
C0268849|T047|SY|786460007|SNOMEDCT_CORE|Overactive detrusor|Detrusor overactivity
C0268936|T046|PTGB|89966002|SNOMEDCT_CORE|Haematoma of scrotum|Hematoma of scrotum
C0268936|T046|PT|89966002|SNOMEDCT_CORE|Hematoma of scrotum|Hematoma of scrotum
C0268936|T046|FN|89966002|SNOMEDCT_CORE|Hematoma of scrotum|Hematoma of scrotum
C0268936|T046|SYGB|89966002|SNOMEDCT_CORE|Scrotal haematoma|Hematoma of scrotum
C0268936|T046|SY|89966002|SNOMEDCT_CORE|Scrotal hematoma|Hematoma of scrotum
C0269084|T047|SY|30833006|SNOMEDCT_CORE|Vestibulodynia|Vulvar vestibulitis
C0269084|T047|SY|30833006|SNOMEDCT_CORE|Vulval vestibulitis|Vulvar vestibulitis
C0269084|T047|PT|30833006|SNOMEDCT_CORE|Vulvar vestibulitis|Vulvar vestibulitis
C0269084|T047|FN|30833006|SNOMEDCT_CORE|Vulvar vestibulitis|Vulvar vestibulitis
C0269125|T020|PT|48230001|SNOMEDCT_CORE|First degree uterine prolapse|First degree uterine prolapse
C0269125|T020|FN|48230001|SNOMEDCT_CORE|First degree uterine prolapse|First degree uterine prolapse
C0269126|T020|PT|9283009|SNOMEDCT_CORE|Second degree uterine prolapse|Second degree uterine prolapse
C0269126|T020|FN|9283009|SNOMEDCT_CORE|Second degree uterine prolapse|Second degree uterine prolapse
C0269130|T033|OAP|11374003|SNOMEDCT_CORE|Relaxation of vaginal outlet AND/OR pelvis|Relaxation of vaginal outlet AND/OR pelvis
C0269130|T033|OAF|11374003|SNOMEDCT_CORE|Relaxation of vaginal outlet AND/OR pelvis|Relaxation of vaginal outlet AND/OR pelvis
C0269130|T033|IS|11374003|SNOMEDCT_CORE|Relaxation of vaginal outlet or pelvis|Relaxation of vaginal outlet AND/OR pelvis
C0269151|T047|PT|79734007|SNOMEDCT_CORE|Noninflammatory disorder of ovary|Noninflammatory disorder of ovary
C0269151|T047|FN|79734007|SNOMEDCT_CORE|Noninflammatory disorder of ovary|Noninflammatory disorder of ovary
C0269151|T047|IS|79734007|SNOMEDCT_CORE|Noninflammatory disorder of ovary, NOS|Noninflammatory disorder of ovary
C0269165|T047|PT|64552006|SNOMEDCT_CORE|Noninflammatory disorder of fallopian tube|Noninflammatory disorder of fallopian tube
C0269165|T047|FN|64552006|SNOMEDCT_CORE|Noninflammatory disorder of fallopian tube|Noninflammatory disorder of fallopian tube
C0269165|T047|IS|64552006|SNOMEDCT_CORE|Noninflammatory disorder of fallopian tube, NOS|Noninflammatory disorder of fallopian tube
C0269175|T047|PT|15848008|SNOMEDCT_CORE|Noninflammatory disorder of broad ligament|Noninflammatory disorder of broad ligament
C0269175|T047|FN|15848008|SNOMEDCT_CORE|Noninflammatory disorder of broad ligament|Noninflammatory disorder of broad ligament
C0269175|T047|IS|15848008|SNOMEDCT_CORE|Noninflammatory disorder of broad ligament, NOS|Noninflammatory disorder of broad ligament
C0269199|T190|PT|83536006|SNOMEDCT_CORE|Stenosis of cervix|Stenosis of cervix
C0269199|T190|FN|83536006|SNOMEDCT_CORE|Stenosis of cervix|Stenosis of cervix
C0269199|T190|SY|83536006|SNOMEDCT_CORE|Stricture of cervix|Stenosis of cervix
C0269216|T047|PT|28271003|SNOMEDCT_CORE|Noninflammatory disorder of vulva|Noninflammatory disorder of vulva
C0269216|T047|FN|28271003|SNOMEDCT_CORE|Noninflammatory disorder of vulva|Noninflammatory disorder of vulva
C0269216|T047|IS|28271003|SNOMEDCT_CORE|Noninflammatory disorder of vulva, NOS|Noninflammatory disorder of vulva
C0269226|T046|PT|23186000|SNOMEDCT_CORE|Menstrual migraine|Menstrual migraine
C0269226|T046|FN|23186000|SNOMEDCT_CORE|Menstrual migraine|Menstrual migraine
C0269229|T047|PT|5084002|SNOMEDCT_CORE|Primary female infertility|Primary female infertility
C0269229|T047|FN|5084002|SNOMEDCT_CORE|Primary female infertility|Primary female infertility
C0269230|T047|PT|30238006|SNOMEDCT_CORE|Secondary female infertility|Secondary female infertility
C0269230|T047|FN|30238006|SNOMEDCT_CORE|Secondary female infertility|Secondary female infertility
C0269596|T046|SYGB|106004004|SNOMEDCT_CORE|Haemorrhage of pregnancy|Hemorrhagic complication of pregnancy
C0269596|T046|PTGB|106004004|SNOMEDCT_CORE|Haemorrhagic complication of pregnancy|Hemorrhagic complication of pregnancy
C0269596|T046|SY|106004004|SNOMEDCT_CORE|Hemorrhage of pregnancy|Hemorrhagic complication of pregnancy
C0269596|T046|PT|106004004|SNOMEDCT_CORE|Hemorrhagic complication of pregnancy|Hemorrhagic complication of pregnancy
C0269596|T046|FN|106004004|SNOMEDCT_CORE|Hemorrhagic complication of pregnancy|Hemorrhagic complication of pregnancy
C0269608|T046|PTGB|34842007|SNOMEDCT_CORE|Antepartum haemorrhage|Antepartum hemorrhage
C0269608|T046|FN|34842007|SNOMEDCT_CORE|Antepartum hemorrhage|Antepartum hemorrhage
C0269608|T046|PT|34842007|SNOMEDCT_CORE|Antepartum hemorrhage|Antepartum hemorrhage
C0269608|T046|IS|34842007|SNOMEDCT_CORE|Antepartum hemorrhage, NOS|Antepartum hemorrhage
C0269608|T046|SYGB|34842007|SNOMEDCT_CORE|APH - Antepartum haemorrhage|Antepartum hemorrhage
C0269608|T046|SY|34842007|SNOMEDCT_CORE|APH - Antepartum hemorrhage|Antepartum hemorrhage
C0269622|T047|PT|23717007|SNOMEDCT_CORE|Benign essential hypertension complicating AND/OR reason for care during pregnancy|Benign essential hypertension complicating AND/OR reason for care during pregnancy
C0269622|T047|FN|23717007|SNOMEDCT_CORE|Benign essential hypertension complicating AND/OR reason for care during pregnancy|Benign essential hypertension complicating AND/OR reason for care during pregnancy
C0269622|T047|IS|23717007|SNOMEDCT_CORE|Benign essential hypertension complicating or reason for care during pregnancy|Benign essential hypertension complicating AND/OR reason for care during pregnancy
C0269658|T046|PT|41114007|SNOMEDCT_CORE|Mild pre-eclampsia|Mild pre-eclampsia
C0269658|T046|FN|41114007|SNOMEDCT_CORE|Mild pre-eclampsia|Mild pre-eclampsia
C0269658|T046|SYGB|41114007|SNOMEDCT_CORE|Mild pre-eclamptic toxaemia|Mild pre-eclampsia
C0269658|T046|SY|41114007|SNOMEDCT_CORE|Mild pre-eclamptic toxemia|Mild pre-eclampsia
C0269658|T046|SY|41114007|SNOMEDCT_CORE|Mild proteinuric hypertension of pregnancy|Mild pre-eclampsia
C0269658|T046|SYGB|41114007|SNOMEDCT_CORE|PET - Mild pre-eclamptic toxaemia|Mild pre-eclampsia
C0269658|T046|SY|41114007|SNOMEDCT_CORE|PET - Mild pre-eclamptic toxemia|Mild pre-eclampsia
C0269661|T046|SY|90325002|SNOMEDCT_CORE|Vomiting as reason for care in pregnancy|Vomiting of pregnancy
C0269661|T046|IS|90325002|SNOMEDCT_CORE|Vomiting as reason for care in pregnancy, NOS|Vomiting of pregnancy
C0269661|T046|PT|90325002|SNOMEDCT_CORE|Vomiting of pregnancy|Vomiting of pregnancy
C0269661|T046|FN|90325002|SNOMEDCT_CORE|Vomiting of pregnancy|Vomiting of pregnancy
C0269661|T046|IS|90325002|SNOMEDCT_CORE|Vomiting of pregnancy, NOS|Vomiting of pregnancy
C0269672|T046|SY|44772007|SNOMEDCT_CORE|Excessive weight gain in pregnancy|Maternal obesity syndrome
C0269672|T046|PT|44772007|SNOMEDCT_CORE|Maternal obesity syndrome|Maternal obesity syndrome
C0269672|T046|FN|44772007|SNOMEDCT_CORE|Maternal obesity syndrome|Maternal obesity syndrome
C0269672|T046|SY|44772007|SNOMEDCT_CORE|Maternal obesity without hypertension|Maternal obesity syndrome
C0269673|T047|SY|75150001|SNOMEDCT_CORE|Nephropathy in pregnancy AND/OR puerperium without hypertension|Renal disease in pregnancy AND/OR puerperium without hypertension
C0269673|T047|IS|75150001|SNOMEDCT_CORE|Nephropathy, NOS, in pregnancy or puerperium without hypertension|Renal disease in pregnancy AND/OR puerperium without hypertension
C0269673|T047|PT|75150001|SNOMEDCT_CORE|Renal disease in pregnancy AND/OR puerperium without hypertension|Renal disease in pregnancy AND/OR puerperium without hypertension
C0269673|T047|FN|75150001|SNOMEDCT_CORE|Renal disease in pregnancy AND/OR puerperium without hypertension|Renal disease in pregnancy AND/OR puerperium without hypertension
C0269673|T047|IS|75150001|SNOMEDCT_CORE|Renal disease, NOS, in pregnancy or puerperium without hypertension|Renal disease in pregnancy AND/OR puerperium without hypertension
C0269674|T046|PT|34165000|SNOMEDCT_CORE|Gestational proteinuria|Gestational proteinuria
C0269674|T046|FN|34165000|SNOMEDCT_CORE|Gestational proteinuria|Gestational proteinuria
C0269684|T047|PTGB|45828008|SNOMEDCT_CORE|Anaemia in mother complicating pregnancy, childbirth AND/OR puerperium|Anemia in mother complicating pregnancy, childbirth AND/OR puerperium
C0269684|T047|PT|45828008|SNOMEDCT_CORE|Anemia in mother complicating pregnancy, childbirth AND/OR puerperium|Anemia in mother complicating pregnancy, childbirth AND/OR puerperium
C0269684|T047|FN|45828008|SNOMEDCT_CORE|Anemia in mother complicating pregnancy, childbirth AND/OR puerperium|Anemia in mother complicating pregnancy, childbirth AND/OR puerperium
C0269684|T047|IS|45828008|SNOMEDCT_CORE|Anemia in mother complicating pregnancy, childbirth or puerperium|Anemia in mother complicating pregnancy, childbirth AND/OR puerperium
C0269702|T046|PT|17532001|SNOMEDCT_CORE|Breech malpresentation successfully converted to cephalic presentation|Breech malpresentation successfully converted to cephalic presentation
C0269702|T046|FN|17532001|SNOMEDCT_CORE|Breech malpresentation successfully converted to cephalic presentation|Breech malpresentation successfully converted to cephalic presentation
C0269733|T033|OAS|64756007|SNOMEDCT_CORE|Pregnancy with history of previous caesarean section|Previous caesarean section
C0269733|T033|OAS|64756007|SNOMEDCT_CORE|Pregnancy with history of previous cesarean section|Previous caesarean section
C0269733|T033|OAP|64756007|SNOMEDCT_CORE|Previous caesarean section|Previous caesarean section
C0269733|T033|OAP|64756007|SNOMEDCT_CORE|Previous cesarean section|Previous caesarean section
C0269733|T033|OAF|64756007|SNOMEDCT_CORE|Previous cesarean section|Previous caesarean section
C0269733|T033|IS|64756007|SNOMEDCT_CORE|Previous cesarean section, NOS|Previous caesarean section
C0269764|T047|PT|106009009|SNOMEDCT_CORE|Fetal condition affecting obstetrical care of mother|Fetal condition affecting obstetrical care of mother
C0269764|T047|FN|106009009|SNOMEDCT_CORE|Fetal condition affecting obstetrical care of mother|Fetal condition affecting obstetrical care of mother
C0269764|T047|PTGB|106009009|SNOMEDCT_CORE|Foetal condition affecting obstetrical care of mother|Fetal condition affecting obstetrical care of mother
C0269791|T047|PT|20845005|SNOMEDCT_CORE|Meconium in amniotic fluid affecting management of mother|Meconium in amniotic fluid affecting management of mother
C0269791|T047|FN|20845005|SNOMEDCT_CORE|Meconium in amniotic fluid affecting management of mother|Meconium in amniotic fluid affecting management of mother
C0269806|T046|PT|42571002|SNOMEDCT_CORE|Failed induction of labor|Failed induction of labor
C0269806|T046|FN|42571002|SNOMEDCT_CORE|Failed induction of labor|Failed induction of labor
C0269806|T046|IS|42571002|SNOMEDCT_CORE|Failed induction of labor, NOS|Failed induction of labor
C0269806|T046|PTGB|42571002|SNOMEDCT_CORE|Failed induction of labour|Failed induction of labor
C0269806|T046|SY|42571002|SNOMEDCT_CORE|Unsuccessful attempt to induce labor|Failed induction of labor
C0269806|T046|SYGB|42571002|SNOMEDCT_CORE|Unsuccessful attempt to induce labour|Failed induction of labor
C0269806|T046|SY|42571002|SNOMEDCT_CORE|Unsuccessfully induced labor|Failed induction of labor
C0269806|T046|SYGB|42571002|SNOMEDCT_CORE|Unsuccessfully induced labour|Failed induction of labor
C0269808|T046|PT|77854008|SNOMEDCT_CORE|Failed medical induction of labor|Failed medical induction of labor
C0269808|T046|FN|77854008|SNOMEDCT_CORE|Failed medical induction of labor|Failed medical induction of labor
C0269808|T046|PTGB|77854008|SNOMEDCT_CORE|Failed medical induction of labour|Failed medical induction of labor
C0269824|T033|PT|70068004|SNOMEDCT_CORE|Persistent occipitoposterior position|Persistent occipitoposterior position
C0269824|T033|FN|70068004|SNOMEDCT_CORE|Persistent occipitoposterior position|Persistent occipitoposterior position
C0269824|T033|SY|70068004|SNOMEDCT_CORE|POP - Persistent occipitoposterior position|Persistent occipitoposterior position
C0269825|T046|SY|89700002|SNOMEDCT_CORE|Impacted shoulders|Shoulder girdle dystocia
C0269825|T046|SY|89700002|SNOMEDCT_CORE|Shoulder dystocia|Shoulder girdle dystocia
C0269825|T046|PT|89700002|SNOMEDCT_CORE|Shoulder girdle dystocia|Shoulder girdle dystocia
C0269825|T046|FN|89700002|SNOMEDCT_CORE|Shoulder girdle dystocia|Shoulder girdle dystocia
C0269827|T047|OAF|14331002|SNOMEDCT_CORE|Failed vacuum extraction delivery|Failed vacuum extractor
C0269827|T047|OAS|14331002|SNOMEDCT_CORE|Failed vacuum extraction delivery|Failed vacuum extractor
C0269827|T047|OAP|14331002|SNOMEDCT_CORE|Failed vacuum extractor|Failed vacuum extractor
C0269827|T047|OF|14331002|SNOMEDCT_CORE|Failed vacuum extractor|Failed vacuum extractor
C0269859|T037|PT|398019008|SNOMEDCT_CORE|Perineal laceration during delivery|Perineal laceration during delivery
C0269859|T037|FN|398019008|SNOMEDCT_CORE|Perineal laceration during delivery|Perineal laceration during delivery
C0269859|T037|SY|398019008|SNOMEDCT_CORE|Perineal tear resulting from childbirth|Perineal laceration during delivery
C0269863|T037|PT|57759005|SNOMEDCT_CORE|First degree perineal laceration|First degree perineal laceration
C0269863|T037|FN|57759005|SNOMEDCT_CORE|First degree perineal laceration|First degree perineal laceration
C0269863|T037|IS|57759005|SNOMEDCT_CORE|First degree perineal laceration, NOS|First degree perineal laceration
C0269863|T037|SY|57759005|SNOMEDCT_CORE|Laceration of superficial layers of perineal structures|First degree perineal laceration
C0269863|T037|SY|57759005|SNOMEDCT_CORE|Obstetrical laceration, first degree|First degree perineal laceration
C0269870|T037|IS|6234006|SNOMEDCT_CORE|Laceration of inner and muscular layers of perineal structures|Second degree perineal laceration
C0269870|T037|SY|6234006|SNOMEDCT_CORE|Laceration of inner AND/OR muscular layers of perineal structures|Second degree perineal laceration
C0269870|T037|SY|6234006|SNOMEDCT_CORE|Obstetrical laceration, second degree|Second degree perineal laceration
C0269870|T037|PT|6234006|SNOMEDCT_CORE|Second degree perineal laceration|Second degree perineal laceration
C0269870|T037|FN|6234006|SNOMEDCT_CORE|Second degree perineal laceration|Second degree perineal laceration
C0269870|T037|IS|6234006|SNOMEDCT_CORE|Second degree perineal laceration, NOS|Second degree perineal laceration
C0269874|T037|IS|10217006|SNOMEDCT_CORE|Laceration of tissues between vaginal and perineal muscular layers and rectal mucosa|Third degree perineal laceration
C0269874|T037|SY|10217006|SNOMEDCT_CORE|Laceration of tissues between vaginal AND/OR perineal muscular layers and rectal mucosa|Third degree perineal laceration
C0269874|T037|SY|10217006|SNOMEDCT_CORE|Obstetrical laceration, third degree|Third degree perineal laceration
C0269874|T037|PT|10217006|SNOMEDCT_CORE|Third degree perineal laceration|Third degree perineal laceration
C0269874|T037|FN|10217006|SNOMEDCT_CORE|Third degree perineal laceration|Third degree perineal laceration
C0269874|T037|IS|10217006|SNOMEDCT_CORE|Third degree perineal laceration, NOS|Third degree perineal laceration
C0269899|T046|PTGB|27214003|SNOMEDCT_CORE|Atonic postpartum haemorrhage|Atonic postpartum hemorrhage
C0269899|T046|PT|27214003|SNOMEDCT_CORE|Atonic postpartum hemorrhage|Atonic postpartum hemorrhage
C0269899|T046|FN|27214003|SNOMEDCT_CORE|Atonic postpartum hemorrhage|Atonic postpartum hemorrhage
C0269899|T046|IS|27214003|SNOMEDCT_CORE|Atonic postpartum hemorrhage, NOS|Atonic postpartum hemorrhage
C0269899|T046|SYGB|27214003|SNOMEDCT_CORE|Haemorrhage within 24 hours following delivery of placenta|Atonic postpartum hemorrhage
C0269899|T046|SY|27214003|SNOMEDCT_CORE|Hemorrhage within 24 hours following delivery of placenta|Atonic postpartum hemorrhage
C0269899|T046|SYGB|27214003|SNOMEDCT_CORE|Immediate postpartum haemorrhage|Atonic postpartum hemorrhage
C0269899|T046|SY|27214003|SNOMEDCT_CORE|Immediate postpartum hemorrhage|Atonic postpartum hemorrhage
C0269901|T046|SYGB|44216000|SNOMEDCT_CORE|Haemorrhage from retained portion of placenta AND/OR membranes|Retained products of conception, following delivery with hemorrhage
C0269901|T046|SY|44216000|SNOMEDCT_CORE|Hemorrhage from retained portion of placenta AND/OR membranes|Retained products of conception, following delivery with hemorrhage
C0269901|T046|IS|44216000|SNOMEDCT_CORE|Hemorrhage from retained portion of placenta or membranes|Retained products of conception, following delivery with hemorrhage
C0269901|T046|SYGB|44216000|SNOMEDCT_CORE|Postpartum haemorrhage with retained placenta|Retained products of conception, following delivery with hemorrhage
C0269901|T046|SY|44216000|SNOMEDCT_CORE|Postpartum hemorrhage with retained placenta|Retained products of conception, following delivery with hemorrhage
C0269901|T046|PTGB|44216000|SNOMEDCT_CORE|Retained products of conception, following delivery with haemorrhage|Retained products of conception, following delivery with hemorrhage
C0269901|T046|PT|44216000|SNOMEDCT_CORE|Retained products of conception, following delivery with hemorrhage|Retained products of conception, following delivery with hemorrhage
C0269901|T046|FN|44216000|SNOMEDCT_CORE|Retained products of conception, following delivery with hemorrhage|Retained products of conception, following delivery with hemorrhage
C0269901|T046|IS|44216000|SNOMEDCT_CORE|Retained products of conception, NOS, following delivery with hemorrhage|Retained products of conception, following delivery with hemorrhage
C0269966|T033|SY|398262004|SNOMEDCT_CORE|Breakdown of perineum|Disruption of episiotomy wound in the puerperium
C0269966|T033|PT|398262004|SNOMEDCT_CORE|Disruption of episiotomy wound in the puerperium|Disruption of episiotomy wound in the puerperium
C0269966|T033|FN|398262004|SNOMEDCT_CORE|Disruption of episiotomy wound in the puerperium|Disruption of episiotomy wound in the puerperium
C0269966|T033|SY|398262004|SNOMEDCT_CORE|Episiotomy breakdown|Disruption of episiotomy wound in the puerperium
C0269985|T047|OAS|86216003|SNOMEDCT_CORE|Mastitis associated with breastfeeding|Mastitis associated with lactation
C0269985|T047|SY|700038005|SNOMEDCT_CORE|Mastitis associated with breastfeeding|Mastitis associated with lactation
C0269985|T047|OAP|86216003|SNOMEDCT_CORE|Mastitis associated with lactation|Mastitis associated with lactation
C0269985|T047|PT|700038005|SNOMEDCT_CORE|Mastitis associated with lactation|Mastitis associated with lactation
C0269985|T047|OAF|86216003|SNOMEDCT_CORE|Mastitis associated with lactation|Mastitis associated with lactation
C0269985|T047|FN|700038005|SNOMEDCT_CORE|Mastitis associated with lactation|Mastitis associated with lactation
C0269985|T047|OAS|86216003|SNOMEDCT_CORE|Mastitis, associated with childbirth|Mastitis associated with lactation
C0269985|T047|OF|86216003|SNOMEDCT_CORE|Mastitis, associated with childbirth|Mastitis associated with lactation
C0269985|T047|IS|86216003|SNOMEDCT_CORE|Mastitis, NOS, associated with childbirth|Mastitis associated with lactation
C0269985|T047|OAS|86216003|SNOMEDCT_CORE|Postpartum mastitis|Mastitis associated with lactation
C0269985|T047|SY|700038005|SNOMEDCT_CORE|Postpartum mastitis|Mastitis associated with lactation
C0269985|T047|IS|86216003|SNOMEDCT_CORE|Postpartum mastitis, NOS|Mastitis associated with lactation
C0269985|T047|OAS|86216003|SNOMEDCT_CORE|Puerperal mastitis|Mastitis associated with lactation
C0269985|T047|SY|700038005|SNOMEDCT_CORE|Puerperal mastitis|Mastitis associated with lactation
C0269985|T047|IS|86216003|SNOMEDCT_CORE|Puerperal mastitis, NOS|Mastitis associated with lactation
C0270057|T046|IS|5984000|SNOMEDCT_CORE|Fetus or newborn affected by malpresentation, malposition or disproportion during labor and delivery|Fetus or newborn affected by malpresentation, malposition or disproportion during labor and delivery
C0270063|T046|PTGB|82719008|SNOMEDCT_CORE|Fetal or neonatal effect of maternal anaesthesia and/or analgesia|Fetal or neonatal effect of maternal anesthesia and/or analgesia
C0270063|T046|PT|82719008|SNOMEDCT_CORE|Fetal or neonatal effect of maternal anesthesia and/or analgesia|Fetal or neonatal effect of maternal anesthesia and/or analgesia
C0270063|T046|FN|82719008|SNOMEDCT_CORE|Fetal or neonatal effect of maternal anesthesia and/or analgesia|Fetal or neonatal effect of maternal anesthesia and/or analgesia
C0270063|T046|IS|82719008|SNOMEDCT_CORE|Fetus OR newborn affected by maternal anaesthesia AND/OR analgesia|Fetal or neonatal effect of maternal anesthesia and/or analgesia
C0270063|T046|OP|82719008|SNOMEDCT_CORE|Fetus OR newborn affected by maternal anesthesia AND/OR analgesia|Fetal or neonatal effect of maternal anesthesia and/or analgesia
C0270063|T046|OF|82719008|SNOMEDCT_CORE|Fetus OR newborn affected by maternal anesthesia AND/OR analgesia|Fetal or neonatal effect of maternal anesthesia and/or analgesia
C0270063|T046|IS|82719008|SNOMEDCT_CORE|Fetus or newborn affected by maternal anesthesia or analgesia|Fetal or neonatal effect of maternal anesthesia and/or analgesia
C0270063|T046|SYGB|82719008|SNOMEDCT_CORE|Foetal or neonatal effect of maternal anaesthesia and/or analgesia|Fetal or neonatal effect of maternal anesthesia and/or analgesia
C0270063|T046|OP|82719008|SNOMEDCT_CORE|Foetus OR newborn affected by maternal anaesthesia AND/OR analgesia|Fetal or neonatal effect of maternal anesthesia and/or analgesia
C0270078|T047|SY|276658003|SNOMEDCT_CORE|Extreme immaturity|Extreme prematurity of infant
C0270078|T047|FN|276658003|SNOMEDCT_CORE|Extreme immaturity|Extreme prematurity of infant
C0270078|T047|PT|276658003|SNOMEDCT_CORE|Extreme prematurity of infant|Extreme prematurity of infant
C0270078|T047|IS|276658003|SNOMEDCT_CORE|Very premature baby|Extreme prematurity of infant
C0270094|T037|PT|206209004|SNOMEDCT_CORE|Fracture of clavicle due to birth trauma|Fracture of clavicle due to birth trauma
C0270094|T037|FN|206209004|SNOMEDCT_CORE|Fracture of clavicle due to birth trauma|Fracture of clavicle due to birth trauma
C0270105|T037|PT|53785005|SNOMEDCT_CORE|Injury to brachial plexus as birth trauma|Injury to brachial plexus as birth trauma
C0270105|T037|FN|53785005|SNOMEDCT_CORE|Injury to brachial plexus as birth trauma|Injury to brachial plexus as birth trauma
C0270124|T047|PT|90562004|SNOMEDCT_CORE|Fetal distress, in liveborn infant|Fetal distress, in liveborn infant
C0270124|T047|OF|90562004|SNOMEDCT_CORE|Fetal distress, in liveborn infant|Fetal distress, in liveborn infant
C0270124|T047|FN|90562004|SNOMEDCT_CORE|Fetal distress, in liveborn infant|Fetal distress, in liveborn infant
C0270124|T047|IS|90562004|SNOMEDCT_CORE|Fetal distress, NOS, in liveborn infant|Fetal distress, in liveborn infant
C0270124|T047|SY|90562004|SNOMEDCT_CORE|Fetal intrauterine distress, not clear if noted before OR after onset of labor in liveborn infant|Fetal distress, in liveborn infant
C0270124|T047|IS|90562004|SNOMEDCT_CORE|Fetal intrauterine distress, not clear if noted before or after onset of labor in liveborn infant|Fetal distress, in liveborn infant
C0270124|T047|SYGB|90562004|SNOMEDCT_CORE|Fetal intrauterine distress, not clear if noted before OR after onset of labour in liveborn infant|Fetal distress, in liveborn infant
C0270124|T047|PTGB|90562004|SNOMEDCT_CORE|Foetal distress, in liveborn infant|Fetal distress, in liveborn infant
C0270124|T047|IS|90562004|SNOMEDCT_CORE|Foetal distress, NOS, in liveborn infant|Fetal distress, in liveborn infant
C0270124|T047|SYGB|90562004|SNOMEDCT_CORE|Foetal intrauterine distress, not clear if noted before OR after onset of labour in liveborn infant|Fetal distress, in liveborn infant
C0270139|T046|PT|7996008|SNOMEDCT_CORE|Fetal intrauterine distress first noted during labor AND/OR delivery in liveborn infant|Fetal intrauterine distress first noted during labor AND/OR delivery in liveborn infant
C0270139|T046|OF|7996008|SNOMEDCT_CORE|Fetal intrauterine distress first noted during labor AND/OR delivery in liveborn infant|Fetal intrauterine distress first noted during labor AND/OR delivery in liveborn infant
C0270139|T046|FN|7996008|SNOMEDCT_CORE|Fetal intrauterine distress first noted during labor AND/OR delivery in liveborn infant|Fetal intrauterine distress first noted during labor AND/OR delivery in liveborn infant
C0270139|T046|IS|7996008|SNOMEDCT_CORE|Fetal intrauterine distress first noted during labor or delivery in liveborn infant|Fetal intrauterine distress first noted during labor AND/OR delivery in liveborn infant
C0270139|T046|PTGB|7996008|SNOMEDCT_CORE|Fetal intrauterine distress first noted during labour AND/OR delivery in liveborn infant|Fetal intrauterine distress first noted during labor AND/OR delivery in liveborn infant
C0270139|T046|SYGB|7996008|SNOMEDCT_CORE|Foetal intrauterine distress first noted during labour AND/OR delivery in liveborn infant|Fetal intrauterine distress first noted during labor AND/OR delivery in liveborn infant
C0270146|T047|SY|17849001|SNOMEDCT_CORE|Fetus and newborn respiratory conditions|Respiratory condition of fetus OR newborn
C0270146|T047|SY|17849001|SNOMEDCT_CORE|Foetus and newborn respiratory conditions|Respiratory condition of fetus OR newborn
C0270146|T047|SY|17849001|SNOMEDCT_CORE|Perinatal respiratory disorders|Respiratory condition of fetus OR newborn
C0270146|T047|PT|17849001|SNOMEDCT_CORE|Respiratory condition of fetus OR newborn|Respiratory condition of fetus OR newborn
C0270146|T047|FN|17849001|SNOMEDCT_CORE|Respiratory condition of fetus OR newborn|Respiratory condition of fetus OR newborn
C0270146|T047|IS|17849001|SNOMEDCT_CORE|Respiratory condition of fetus or newborn, NOS|Respiratory condition of fetus OR newborn
C0270146|T047|SY|17849001|SNOMEDCT_CORE|Respiratory condition of foetus OR newborn|Respiratory condition of fetus OR newborn
C0270191|T046|SYGB|70611002|SNOMEDCT_CORE|Intraventricular haemorrhage from any perinatal cause|Perinatal intraventricular hemorrhage
C0270191|T046|SY|70611002|SNOMEDCT_CORE|Intraventricular hemorrhage from any perinatal cause|Perinatal intraventricular hemorrhage
C0270191|T046|SYGB|70611002|SNOMEDCT_CORE|Neonatal intraventricular haemorrhage|Perinatal intraventricular hemorrhage
C0270191|T046|SY|70611002|SNOMEDCT_CORE|Neonatal intraventricular hemorrhage|Perinatal intraventricular hemorrhage
C0270191|T046|PTGB|70611002|SNOMEDCT_CORE|Perinatal intraventricular haemorrhage|Perinatal intraventricular hemorrhage
C0270191|T046|PT|70611002|SNOMEDCT_CORE|Perinatal intraventricular hemorrhage|Perinatal intraventricular hemorrhage
C0270191|T046|FN|70611002|SNOMEDCT_CORE|Perinatal intraventricular hemorrhage|Perinatal intraventricular hemorrhage
C0270202|T047|SYGB|32858009|SNOMEDCT_CORE|ABO haemolytic disease of the newborn|Hemolytic disease of fetus OR newborn due to ABO immunization
C0270202|T047|SYGB|32858009|SNOMEDCT_CORE|ABO HDN - ABO haemolytic disease of the newborn|Hemolytic disease of fetus OR newborn due to ABO immunization
C0270202|T047|SY|32858009|SNOMEDCT_CORE|ABO HDN - ABO hemolytic disease of the newborn|Hemolytic disease of fetus OR newborn due to ABO immunization
C0270202|T047|SY|32858009|SNOMEDCT_CORE|ABO hemolytic disease of the newborn|Hemolytic disease of fetus OR newborn due to ABO immunization
C0270202|T047|SYGB|32858009|SNOMEDCT_CORE|ABO isoimmunisation of the newborn|Hemolytic disease of fetus OR newborn due to ABO immunization
C0270202|T047|SY|32858009|SNOMEDCT_CORE|ABO isoimmunization of the newborn|Hemolytic disease of fetus OR newborn due to ABO immunization
C0270202|T047|SYGB|32858009|SNOMEDCT_CORE|Anaemia due to ABO incompatibility in the newborn|Hemolytic disease of fetus OR newborn due to ABO immunization
C0270202|T047|SY|32858009|SNOMEDCT_CORE|Anemia due to ABO incompatibility in the newborn|Hemolytic disease of fetus OR newborn due to ABO immunization
C0270202|T047|SYGB|32858009|SNOMEDCT_CORE|Erythroblastosis fetalis due to ABO isoimmunisation|Hemolytic disease of fetus OR newborn due to ABO immunization
C0270202|T047|SY|32858009|SNOMEDCT_CORE|Erythroblastosis fetalis due to ABO isoimmunization|Hemolytic disease of fetus OR newborn due to ABO immunization
C0270202|T047|SYGB|32858009|SNOMEDCT_CORE|Erythroblastosis foetalis due to ABO isoimmunisation|Hemolytic disease of fetus OR newborn due to ABO immunization
C0270202|T047|IS|32858009|SNOMEDCT_CORE|Erythroblastosis foetalis due to ABO isoimmunization|Hemolytic disease of fetus OR newborn due to ABO immunization
C0270202|T047|SYGB|32858009|SNOMEDCT_CORE|Haemolytic disease due to ABO isoimmunisation|Hemolytic disease of fetus OR newborn due to ABO immunization
C0270202|T047|SYGB|32858009|SNOMEDCT_CORE|Haemolytic disease of fetus OR newborn due to ABO immunisation|Hemolytic disease of fetus OR newborn due to ABO immunization
C0270202|T047|PTGB|32858009|SNOMEDCT_CORE|Haemolytic disease of foetus OR newborn due to ABO immunisation|Hemolytic disease of fetus OR newborn due to ABO immunization
C0270202|T047|SY|32858009|SNOMEDCT_CORE|Hemolytic disease due to ABO isoimmunization|Hemolytic disease of fetus OR newborn due to ABO immunization
C0270202|T047|PT|32858009|SNOMEDCT_CORE|Hemolytic disease of fetus OR newborn due to ABO immunization|Hemolytic disease of fetus OR newborn due to ABO immunization
C0270202|T047|IS|32858009|SNOMEDCT_CORE|Hemolytic disease of fetus or newborn due to ABO immunization|Hemolytic disease of fetus OR newborn due to ABO immunization
C0270202|T047|FN|32858009|SNOMEDCT_CORE|Hemolytic disease of fetus OR newborn due to ABO immunization|Hemolytic disease of fetus OR newborn due to ABO immunization
C0270202|T047|SYGB|32858009|SNOMEDCT_CORE|Jaundice due to ABO isoimmunisation of the newborn|Hemolytic disease of fetus OR newborn due to ABO immunization
C0270202|T047|SY|32858009|SNOMEDCT_CORE|Jaundice due to ABO isoimmunization of the newborn|Hemolytic disease of fetus OR newborn due to ABO immunization
C0270207|T046|SYGB|24911006|SNOMEDCT_CORE|Perinatal haemolytic jaundice|Perinatal jaundice from excessive hemolysis
C0270207|T046|PTGB|24911006|SNOMEDCT_CORE|Perinatal jaundice from excessive haemolysis|Perinatal jaundice from excessive hemolysis
C0270207|T046|PT|24911006|SNOMEDCT_CORE|Perinatal jaundice from excessive hemolysis|Perinatal jaundice from excessive hemolysis
C0270207|T046|FN|24911006|SNOMEDCT_CORE|Perinatal jaundice from excessive hemolysis|Perinatal jaundice from excessive hemolysis
C0270207|T046|IS|24911006|SNOMEDCT_CORE|Perinatal jaundice from excessive hemolysis, NOS|Perinatal jaundice from excessive hemolysis
C0270215|T046|SY|82696006|SNOMEDCT_CORE|Breast milk inhibitor jaundice|Neonatal jaundice due to delayed conjugation from breast milk inhibitor
C0270215|T046|SY|82696006|SNOMEDCT_CORE|Breast milk jaundice|Neonatal jaundice due to delayed conjugation from breast milk inhibitor
C0270215|T046|SY|82696006|SNOMEDCT_CORE|Breast-feeding inhibitor causing neonatal jaundice|Neonatal jaundice due to delayed conjugation from breast milk inhibitor
C0270215|T046|IS|82696006|SNOMEDCT_CORE|Breast-feeding inhibitors causing neonatal jaundice|Neonatal jaundice due to delayed conjugation from breast milk inhibitor
C0270215|T046|PT|82696006|SNOMEDCT_CORE|Neonatal jaundice due to delayed conjugation from breast milk inhibitor|Neonatal jaundice due to delayed conjugation from breast milk inhibitor
C0270215|T046|FN|82696006|SNOMEDCT_CORE|Neonatal jaundice due to delayed conjugation from breast milk inhibitor|Neonatal jaundice due to delayed conjugation from breast milk inhibitor
C0270215|T046|OP|82696006|SNOMEDCT_CORE|Neonatal jaundice due to delayed conjugation from breast milk inhibitors|Neonatal jaundice due to delayed conjugation from breast milk inhibitor
C0270215|T046|OF|82696006|SNOMEDCT_CORE|Neonatal jaundice due to delayed conjugation from breast milk inhibitors|Neonatal jaundice due to delayed conjugation from breast milk inhibitor
C0270221|T047|SY|21584002|SNOMEDCT_CORE|Infant of a diabetic mother syndrome|Syndrome of infant of diabetic mother
C0270221|T047|SY|21584002|SNOMEDCT_CORE|Maternal diabetes syndrome|Syndrome of infant of diabetic mother
C0270221|T047|PT|21584002|SNOMEDCT_CORE|Syndrome of infant of diabetic mother|Syndrome of infant of diabetic mother
C0270221|T047|FN|21584002|SNOMEDCT_CORE|Syndrome of infant of diabetic mother|Syndrome of infant of diabetic mother
C0270256|T046|PT|13629008|SNOMEDCT_CORE|Hypothermia of newborn|Hypothermia of newborn
C0270256|T046|FN|13629008|SNOMEDCT_CORE|Hypothermia of newborn|Hypothermia of newborn
C0270256|T046|IS|13629008|SNOMEDCT_CORE|Hypothermia of newborn, NOS|Hypothermia of newborn
C0270302|T048|PT|53467004|SNOMEDCT_CORE|Anxiety disorder of childhood|Anxiety disorder of childhood
C0270302|T048|FN|53467004|SNOMEDCT_CORE|Anxiety disorder of childhood|Anxiety disorder of childhood
C0270302|T048|IS|53467004|SNOMEDCT_CORE|Anxiety disorder of childhood, NOS|Anxiety disorder of childhood
C0270307|T048|PT|13438001|SNOMEDCT_CORE|Overanxious disorder of childhood|Overanxious disorder of childhood
C0270307|T048|FN|13438001|SNOMEDCT_CORE|Overanxious disorder of childhood|Overanxious disorder of childhood
C0270312|T048|PT|18003009|SNOMEDCT_CORE|Gender identity disorder of adulthood|Gender identity disorder of adulthood
C0270312|T048|FN|18003009|SNOMEDCT_CORE|Gender identity disorder of adulthood|Gender identity disorder of adulthood
C0270312|T048|IS|18003009|SNOMEDCT_CORE|Gender identity disorder of adulthood, NOS|Gender identity disorder of adulthood
C0270327|T048|SY|8009008|SNOMEDCT_CORE|Bed wetting|Nocturnal enuresis
C0270327|T048|IS|8009008|SNOMEDCT_CORE|Bed-wetting|Nocturnal enuresis
C0270327|T048|SY|8009008|SNOMEDCT_CORE|Bedwetting|Nocturnal enuresis
C0270327|T048|PT|8009008|SNOMEDCT_CORE|Nocturnal enuresis|Nocturnal enuresis
C0270327|T048|OF|8009008|SNOMEDCT_CORE|Nocturnal enuresis|Nocturnal enuresis
C0270327|T048|FN|8009008|SNOMEDCT_CORE|Nocturnal enuresis|Nocturnal enuresis
C0270327|T048|SY|8009008|SNOMEDCT_CORE|Nocturnal incontinence of urine|Nocturnal enuresis
C0270327|T048|IS|8009008|SNOMEDCT_CORE|Nocturnal only enuresis|Nocturnal enuresis
C0270327|T048|SY|8009008|SNOMEDCT_CORE|Wets bed|Nocturnal enuresis
C0270330|T048|PT|1145003|SNOMEDCT_CORE|Developmental speech disorder|Developmental speech disorder
C0270330|T048|FN|1145003|SNOMEDCT_CORE|Developmental speech disorder|Developmental speech disorder
C0270330|T048|IS|1145003|SNOMEDCT_CORE|Developmental speech disorder, NOS|Developmental speech disorder
C0270330|T048|SY|1145003|SNOMEDCT_CORE|DSD - Developmental speech disorder|Developmental speech disorder
C0270380|T048|PT|427327003|SNOMEDCT_CORE|Sedative dependence|Sedative dependence
C0270380|T048|FN|427327003|SNOMEDCT_CORE|Sedative dependence|Sedative dependence
C0270398|T048|PT|31658008|SNOMEDCT_CORE|Chronic paranoid schizophrenia|Chronic paranoid schizophrenia
C0270398|T048|FN|31658008|SNOMEDCT_CORE|Chronic paranoid schizophrenia|Chronic paranoid schizophrenia
C0270400|T048|PT|63181006|SNOMEDCT_CORE|Paranoid schizophrenia in remission|Paranoid schizophrenia in remission
C0270400|T048|FN|63181006|SNOMEDCT_CORE|Paranoid schizophrenia in remission|Paranoid schizophrenia in remission
C0270400|T048|SY|63181006|SNOMEDCT_CORE|Paranoid schizophrenia, in remission|Paranoid schizophrenia in remission
C0270403|T048|PT|29599000|SNOMEDCT_CORE|Chronic undifferentiated schizophrenia|Chronic undifferentiated schizophrenia
C0270403|T048|FN|29599000|SNOMEDCT_CORE|Chronic undifferentiated schizophrenia|Chronic undifferentiated schizophrenia
C0270425|T048|PT|85248005|SNOMEDCT_CORE|Bipolar disorder in remission|Bipolar disorder in remission
C0270425|T048|FN|85248005|SNOMEDCT_CORE|Bipolar disorder in remission|Bipolar disorder in remission
C0270425|T048|SY|85248005|SNOMEDCT_CORE|Bipolar disorder, in remission|Bipolar disorder in remission
C0270456|T048|PT|832007|SNOMEDCT_CORE|Moderate major depression|Moderate major depression
C0270456|T048|FN|832007|SNOMEDCT_CORE|Moderate major depression|Moderate major depression
C0270457|T048|PT|75084000|SNOMEDCT_CORE|Severe major depression without psychotic features|Severe major depression without psychotic features
C0270457|T048|FN|75084000|SNOMEDCT_CORE|Severe major depression without psychotic features|Severe major depression without psychotic features
C0270458|T048|SY|73867007|SNOMEDCT_CORE|Psychotic depression|Severe major depression with psychotic features
C0270458|T048|IS|73867007|SNOMEDCT_CORE|Psychotic depression, NOS|Severe major depression with psychotic features
C0270458|T048|PT|73867007|SNOMEDCT_CORE|Severe major depression with psychotic features|Severe major depression with psychotic features
C0270458|T048|FN|73867007|SNOMEDCT_CORE|Severe major depression with psychotic features|Severe major depression with psychotic features
C0270458|T048|IS|73867007|SNOMEDCT_CORE|Severe major depression with psychotic features, NOS|Severe major depression with psychotic features
C0270461|T048|PT|42810003|SNOMEDCT_CORE|Major depression in remission|Major depression in remission
C0270461|T048|FN|42810003|SNOMEDCT_CORE|Major depression in remission|Major depression in remission
C0270461|T048|IS|42810003|SNOMEDCT_CORE|Major depression in remission, NOS|Major depression in remission
C0270461|T048|SY|42810003|SNOMEDCT_CORE|Major depression, in remission|Major depression in remission
C0270470|T048|SY|19527009|SNOMEDCT_CORE|Major depression, single episode, in complete remission|Single episode of major depression in full remission
C0270470|T048|OF|19527009|SNOMEDCT_CORE|Major depression, single episode, in complete remission|Single episode of major depression in full remission
C0270470|T048|SY|19527009|SNOMEDCT_CORE|Major depression, single episode, in full remission|Single episode of major depression in full remission
C0270470|T048|PT|19527009|SNOMEDCT_CORE|Single episode of major depression in full remission|Single episode of major depression in full remission
C0270470|T048|FN|19527009|SNOMEDCT_CORE|Single episode of major depression in full remission|Single episode of major depression in full remission
C0270477|T048|PT|68019004|SNOMEDCT_CORE|Recurrent major depression in remission|Recurrent major depression in remission
C0270477|T048|FN|68019004|SNOMEDCT_CORE|Recurrent major depression in remission|Recurrent major depression in remission
C0270480|T048|PT|2506003|SNOMEDCT_CORE|Early onset dysthymia|Early onset dysthymia
C0270480|T048|FN|2506003|SNOMEDCT_CORE|Early onset dysthymia|Early onset dysthymia
C0270497|T048|PT|84760002|SNOMEDCT_CORE|Schizoaffective disorder, depressive type|Schizoaffective disorder, depressive type
C0270497|T048|FN|84760002|SNOMEDCT_CORE|Schizoaffective disorder, depressive type|Schizoaffective disorder, depressive type
C0270497|T048|SY|84760002|SNOMEDCT_CORE|Schizophreniform psychosis, depressive type|Schizoaffective disorder, depressive type
C0270543|T047|PT|44455001|SNOMEDCT_CORE|Hypersomnia disorder related to a known organic factor|Hypersomnia disorder related to a known organic factor
C0270543|T047|FN|44455001|SNOMEDCT_CORE|Hypersomnia disorder related to a known organic factor|Hypersomnia disorder related to a known organic factor
C0270549|T048|SYGB|21897009|SNOMEDCT_CORE|GAD - Generalised anxiety disorder|Generalized anxiety disorder
C0270549|T048|SY|21897009|SNOMEDCT_CORE|GAD - Generalized anxiety disorder|Generalized anxiety disorder
C0270549|T048|PTGB|21897009|SNOMEDCT_CORE|Generalised anxiety disorder|Generalized anxiety disorder
C0270549|T048|PT|21897009|SNOMEDCT_CORE|Generalized anxiety disorder|Generalized anxiety disorder
C0270549|T048|FN|21897009|SNOMEDCT_CORE|Generalized anxiety disorder|Generalized anxiety disorder
C0270611|T037|IS|81308009|SNOMEDCT_CORE|Brain damage, NOS|Brain tissue injury
C0270611|T037|IS|127294003|SNOMEDCT_CORE|Brain injury|Brain tissue injury
C0270611|T037|SY|127294003|SNOMEDCT_CORE|Brain tissue injury|Brain tissue injury
C0270611|T037|SY|127294003|SNOMEDCT_CORE|Intracerebral injury|Brain tissue injury
C0270697|T184|PT|398987004|SNOMEDCT_CORE|Headache following lumbar puncture|Headache following lumbar puncture
C0270697|T184|FN|398987004|SNOMEDCT_CORE|Headache following lumbar puncture|Headache following lumbar puncture
C0270697|T184|SY|398987004|SNOMEDCT_CORE|Lumbar puncture headache|Headache following lumbar puncture
C0270697|T184|SY|398987004|SNOMEDCT_CORE|Post-lumbar puncture headache|Headache following lumbar puncture
C0270697|T184|SY|398987004|SNOMEDCT_CORE|Postspinal headache|Headache following lumbar puncture
C0270697|T184|SY|398987004|SNOMEDCT_CORE|Spinal headache|Headache following lumbar puncture
C0270736|T047|OAS|192839001|SNOMEDCT_CORE|Benign essential tremor|Essential tremor
C0270736|T047|OAP|192839001|SNOMEDCT_CORE|Essential tremor|Essential tremor
C0270736|T047|PT|609558009|SNOMEDCT_CORE|Essential tremor|Essential tremor
C0270736|T047|FN|609558009|SNOMEDCT_CORE|Essential tremor|Essential tremor
C0270736|T047|OAF|192839001|SNOMEDCT_CORE|Essential tremor|Essential tremor
C0270790|T184|SY|91327001|SNOMEDCT_CORE|Quadriparesis|Tetraparesis
C0270790|T184|FN|91327001|SNOMEDCT_CORE|Quadriparesis|Tetraparesis
C0270790|T184|PT|91327001|SNOMEDCT_CORE|Tetraparesis|Tetraparesis
C0270804|T047|SY|58193001|SNOMEDCT_CORE|Congenital diplegia|Diplegic cerebral palsy
C0270804|T047|OAF|275469001|SNOMEDCT_CORE|Congenital diplegia|Diplegic cerebral palsy
C0270804|T047|PT|58193001|SNOMEDCT_CORE|Diplegic cerebral palsy|Diplegic cerebral palsy
C0270804|T047|FN|58193001|SNOMEDCT_CORE|Diplegic cerebral palsy|Diplegic cerebral palsy
C0270804|T047|SY|58193001|SNOMEDCT_CORE|Spastic diplegic cerebral palsy|Diplegic cerebral palsy
C0270805|T019|SY|43486001|SNOMEDCT_CORE|Congenital hemiplegia|Hemiplegic cerebral palsy
C0270805|T047|SY|43486001|SNOMEDCT_CORE|Congenital hemiplegia|Hemiplegic cerebral palsy
C0270805|T019|PT|43486001|SNOMEDCT_CORE|Hemiplegic cerebral palsy|Hemiplegic cerebral palsy
C0270805|T047|PT|43486001|SNOMEDCT_CORE|Hemiplegic cerebral palsy|Hemiplegic cerebral palsy
C0270805|T019|FN|43486001|SNOMEDCT_CORE|Hemiplegic cerebral palsy|Hemiplegic cerebral palsy
C0270805|T047|FN|43486001|SNOMEDCT_CORE|Hemiplegic cerebral palsy|Hemiplegic cerebral palsy
C0270805|T019|SY|43486001|SNOMEDCT_CORE|Spastic hemiplegic cerebral palsy|Hemiplegic cerebral palsy
C0270805|T047|SY|43486001|SNOMEDCT_CORE|Spastic hemiplegic cerebral palsy|Hemiplegic cerebral palsy
C0270805|T019|IS|43486001|SNOMEDCT_CORE|Unilateral spastic cerebral palsy|Hemiplegic cerebral palsy
C0270805|T047|IS|43486001|SNOMEDCT_CORE|Unilateral spastic cerebral palsy|Hemiplegic cerebral palsy
C0270834|T047|PT|4103001|SNOMEDCT_CORE|Complex partial seizure with impairment of consciousness|Complex partial seizure with impairment of consciousness
C0270834|T047|OF|4103001|SNOMEDCT_CORE|Complex partial seizure with impairment of consciousness|Complex partial seizure with impairment of consciousness
C0270834|T047|FN|4103001|SNOMEDCT_CORE|Complex partial seizure with impairment of consciousness|Complex partial seizure with impairment of consciousness
C0270834|T047|SY|4103001|SNOMEDCT_CORE|Complex partial seizures with consciousness impaired|Complex partial seizure with impairment of consciousness
C0270864|T047|OAP|11060002|SNOMEDCT_CORE|Disease related peripheral neuropathy|Disease related peripheral neuropathy
C0270864|T047|OAF|11060002|SNOMEDCT_CORE|Disease related peripheral neuropathy|Disease related peripheral neuropathy
C0270864|T047|IS|11060002|SNOMEDCT_CORE|Disease related peripheral neuropathy, NOS|Disease related peripheral neuropathy
C0270897|T037|SY|78141002|SNOMEDCT_CORE|Erb-Duchenne brachial plexus injury|Erb-Duchenne paralysis
C0270897|T037|PT|78141002|SNOMEDCT_CORE|Erb-Duchenne paralysis|Erb-Duchenne paralysis
C0270897|T037|FN|78141002|SNOMEDCT_CORE|Erb-Duchenne paralysis|Erb-Duchenne paralysis
C0270897|T037|SY|78141002|SNOMEDCT_CORE|Erb's palsy|Erb-Duchenne paralysis
C0270897|T037|SY|78141002|SNOMEDCT_CORE|Erb's paralysis|Erb-Duchenne paralysis
C0270906|T047|PT|58497009|SNOMEDCT_CORE|Tardy ulnar nerve palsy|Tardy ulnar nerve palsy
C0270906|T047|OF|58497009|SNOMEDCT_CORE|Tardy ulnar nerve palsy|Tardy ulnar nerve palsy
C0270906|T047|FN|58497009|SNOMEDCT_CORE|Tardy ulnar nerve palsy|Tardy ulnar nerve palsy
C0270910|T047|PT|22722001|SNOMEDCT_CORE|Idiopathic peripheral neuropathy|Idiopathic peripheral neuropathy
C0270910|T047|FN|22722001|SNOMEDCT_CORE|Idiopathic peripheral neuropathy|Idiopathic peripheral neuropathy
C0270910|T047|IS|22722001|SNOMEDCT_CORE|Idiopathic peripheral neuropathy, NOS|Idiopathic peripheral neuropathy
C0270923|T047|PT|385006|SNOMEDCT_CORE|Secondary peripheral neuropathy|Secondary peripheral neuropathy
C0270923|T047|FN|385006|SNOMEDCT_CORE|Secondary peripheral neuropathy|Secondary peripheral neuropathy
C0270923|T047|IS|385006|SNOMEDCT_CORE|Secondary peripheral neuropathy, NOS|Secondary peripheral neuropathy
C0270933|T047|PT|21018002|SNOMEDCT_CORE|Inflammatory neuropathy|Inflammatory neuropathy
C0270933|T047|FN|21018002|SNOMEDCT_CORE|Inflammatory neuropathy|Inflammatory neuropathy
C0270933|T047|IS|21018002|SNOMEDCT_CORE|Inflammatory neuropathy, NOS|Inflammatory neuropathy
C0270971|T047|SY|33010005|SNOMEDCT_CORE|Congenital hypotonia|Floppy infant syndrome
C0270971|T047|PT|33010005|SNOMEDCT_CORE|Floppy infant syndrome|Floppy infant syndrome
C0270971|T047|FN|33010005|SNOMEDCT_CORE|Floppy infant syndrome|Floppy infant syndrome
C0270994|T047|SY|26715006|SNOMEDCT_CORE|Steroid myopathy|Steroid-induced myopathy
C0270994|T047|PT|26715006|SNOMEDCT_CORE|Steroid-induced myopathy|Steroid-induced myopathy
C0270994|T047|FN|26715006|SNOMEDCT_CORE|Steroid-induced myopathy|Steroid-induced myopathy
C0270997|T047|PT|62619007|SNOMEDCT_CORE|Ill-defined disorder of eye|Ill-defined disorder of eye
C0270997|T047|FN|62619007|SNOMEDCT_CORE|Ill-defined disorder of eye|Ill-defined disorder of eye
C0270997|T047|IS|62619007|SNOMEDCT_CORE|Ill-defined disorder of eye, NOS|Ill-defined disorder of eye
C0271036|T020|PT|66485003|SNOMEDCT_CORE|Retinal scar|Retinal scar
C0271036|T020|FN|66485003|SNOMEDCT_CORE|Retinal scar|Retinal scar
C0271036|T020|IS|66485003|SNOMEDCT_CORE|Retinal scar, NOS|Retinal scar
C0271050|T184|PTGB|28391008|SNOMEDCT_CORE|Localised retinal oedema|Localized retinal edema
C0271050|T184|PT|28391008|SNOMEDCT_CORE|Localized retinal edema|Localized retinal edema
C0271050|T184|FN|28391008|SNOMEDCT_CORE|Localized retinal edema|Localized retinal edema
C0271051|T047|SY|37231002|SNOMEDCT_CORE|Macular edema|Macular retinal edema
C0271051|T047|SYGB|37231002|SNOMEDCT_CORE|Macular oedema|Macular retinal edema
C0271051|T047|PT|37231002|SNOMEDCT_CORE|Macular retinal edema|Macular retinal edema
C0271051|T047|FN|37231002|SNOMEDCT_CORE|Macular retinal edema|Macular retinal edema
C0271051|T047|PTGB|37231002|SNOMEDCT_CORE|Macular retinal oedema|Macular retinal edema
C0271055|T047|SY|19620000|SNOMEDCT_CORE|Retinal detachment due to full thickness retinal tear|Rhegmatogenous retinal detachment
C0271055|T047|SY|19620000|SNOMEDCT_CORE|Retinal detachment with break|Rhegmatogenous retinal detachment
C0271055|T047|PT|19620000|SNOMEDCT_CORE|Rhegmatogenous retinal detachment|Rhegmatogenous retinal detachment
C0271055|T047|FN|19620000|SNOMEDCT_CORE|Rhegmatogenous retinal detachment|Rhegmatogenous retinal detachment
C0271066|T047|SY|75971007|SNOMEDCT_CORE|Choroidal neovascular membrane|Choroidal retinal neovascularization
C0271066|T047|PTGB|75971007|SNOMEDCT_CORE|Choroidal retinal neovascularisation|Choroidal retinal neovascularization
C0271066|T047|PT|75971007|SNOMEDCT_CORE|Choroidal retinal neovascularization|Choroidal retinal neovascularization
C0271066|T047|FN|75971007|SNOMEDCT_CORE|Choroidal retinal neovascularization|Choroidal retinal neovascularization
C0271066|T047|SYGB|75971007|SNOMEDCT_CORE|CNV - Choroidal neovascularisation|Choroidal retinal neovascularization
C0271066|T047|SY|75971007|SNOMEDCT_CORE|CNV - Choroidal neovascularization|Choroidal retinal neovascularization
C0271066|T047|SY|75971007|SNOMEDCT_CORE|CNVM - Choroidal neovascular membrane|Choroidal retinal neovascularization
C0271066|T047|SYGB|75971007|SNOMEDCT_CORE|SRNV-Subretinal neovascularisation|Choroidal retinal neovascularization
C0271066|T047|SY|75971007|SNOMEDCT_CORE|SRNV-Subretinal neovascularization|Choroidal retinal neovascularization
C0271066|T047|SYGB|75971007|SNOMEDCT_CORE|Subretinal neovascularisation|Choroidal retinal neovascularization
C0271066|T047|SY|75971007|SNOMEDCT_CORE|Subretinal neovascularization|Choroidal retinal neovascularization
C0271074|T047|PT|46674002|SNOMEDCT_CORE|Nondiabetic proliferative retinopathy|Nondiabetic proliferative retinopathy
C0271074|T047|FN|46674002|SNOMEDCT_CORE|Nondiabetic proliferative retinopathy|Nondiabetic proliferative retinopathy
C0271074|T047|IS|46674002|SNOMEDCT_CORE|Nondiabetic proliferative retinopathy, NOS|Nondiabetic proliferative retinopathy
C0271083|T020|SY|414875008|SNOMEDCT_CORE|Atrophic age-related macular degeneration|Nonexudative age-related macular degeneration
C0271083|T020|SY|414875008|SNOMEDCT_CORE|Atrophic senile macular retinal degeneration|Nonexudative age-related macular degeneration
C0271083|T020|SY|414875008|SNOMEDCT_CORE|Dry senile macular degeneration|Nonexudative age-related macular degeneration
C0271083|T020|SY|414875008|SNOMEDCT_CORE|Dry senile macular retinal degeneration|Nonexudative age-related macular degeneration
C0271083|T020|SY|414875008|SNOMEDCT_CORE|Geographic atrophy of the macula|Nonexudative age-related macular degeneration
C0271083|T020|PT|414875008|SNOMEDCT_CORE|Nonexudative age-related macular degeneration|Nonexudative age-related macular degeneration
C0271083|T020|FN|414875008|SNOMEDCT_CORE|Nonexudative age-related macular degeneration|Nonexudative age-related macular degeneration
C0271083|T020|SY|414875008|SNOMEDCT_CORE|Nonexudative senile macular degeneration|Nonexudative age-related macular degeneration
C0271083|T020|SY|414875008|SNOMEDCT_CORE|Nonexudative senile macular retinal degeneration|Nonexudative age-related macular degeneration
C0271083|T020|SY|414875008|SNOMEDCT_CORE|Nonneovascular age-related macular degeneration|Nonexudative age-related macular degeneration
C0271084|T047|SY|414173003|SNOMEDCT_CORE|Disciform macular degeneration|Exudative age-related macular degeneration
C0271084|T047|SY|414173003|SNOMEDCT_CORE|Disciform senile macular retinal degeneration|Exudative age-related macular degeneration
C0271084|T047|SY|414173003|SNOMEDCT_CORE|EMD - Exudative macular degeneration|Exudative age-related macular degeneration
C0271084|T047|FN|414173003|SNOMEDCT_CORE|Exudative age-related macular degeneration|Exudative age-related macular degeneration
C0271084|T047|PT|414173003|SNOMEDCT_CORE|Exudative age-related macular degeneration|Exudative age-related macular degeneration
C0271084|T047|SY|414173003|SNOMEDCT_CORE|Exudative senile macular retinal degeneration|Exudative age-related macular degeneration
C0271084|T047|SY|414173003|SNOMEDCT_CORE|Junius-Kuhnt degeneration|Exudative age-related macular degeneration
C0271084|T047|SY|414173003|SNOMEDCT_CORE|Kuhnt Junius degeneration|Exudative age-related macular degeneration
C0271084|T047|SY|414173003|SNOMEDCT_CORE|Neovascular age-related macular degeneration|Exudative age-related macular degeneration
C0271084|T047|SYGB|414173003|SNOMEDCT_CORE|Subretinal neovascularisation of macula|Exudative age-related macular degeneration
C0271084|T047|SY|414173003|SNOMEDCT_CORE|Subretinal neovascularization of macula|Exudative age-related macular degeneration
C0271084|T047|SY|414173003|SNOMEDCT_CORE|Wet senile macular degeneration|Exudative age-related macular degeneration
C0271088|T047|OAP|30523006|SNOMEDCT_CORE|Degenerative drusen|Degenerative drusen
C0271088|T047|OAF|30523006|SNOMEDCT_CORE|Degenerative drusen|Degenerative drusen
C0271143|T047|OAP|81416004|SNOMEDCT_CORE|Open angle with borderline findings|Open angle with borderline findings
C0271143|T047|OAF|81416004|SNOMEDCT_CORE|Open angle with borderline findings|Open angle with borderline findings
C0271143|T047|IS|81416004|SNOMEDCT_CORE|Open angle with borderline findings, NOS|Open angle with borderline findings
C0271163|T047|IS|52421005|SNOMEDCT_CORE|Immature cataract|Incipient cataract
C0271163|T047|PT|52421005|SNOMEDCT_CORE|Incipient cataract|Incipient cataract
C0271163|T047|FN|52421005|SNOMEDCT_CORE|Incipient cataract|Incipient cataract
C0271163|T047|SY|52421005|SNOMEDCT_CORE|Water clefts|Incipient cataract
C0271166|T020|PT|193589009|SNOMEDCT_CORE|Nuclear senile cataract|Nuclear senile cataract
C0271166|T020|FN|193589009|SNOMEDCT_CORE|Nuclear senile cataract|Nuclear senile cataract
C0271168|T047|PT|11422002|SNOMEDCT_CORE|Combined form of senile cataract|Combined form of senile cataract
C0271168|T047|FN|11422002|SNOMEDCT_CORE|Combined form of senile cataract|Combined form of senile cataract
C0271176|T047|IS|51044000|SNOMEDCT_CORE|After cataract not obscuring vision|After-cataract not obscuring vision following extraction of cataract
C0271176|T047|OP|51044000|SNOMEDCT_CORE|After-cataract not obscuring vision|After-cataract not obscuring vision following extraction of cataract
C0271176|T047|OF|51044000|SNOMEDCT_CORE|After-cataract not obscuring vision|After-cataract not obscuring vision following extraction of cataract
C0271176|T047|PT|51044000|SNOMEDCT_CORE|After-cataract not obscuring vision following extraction of cataract|After-cataract not obscuring vision following extraction of cataract
C0271176|T047|FN|51044000|SNOMEDCT_CORE|After-cataract not obscuring vision following extraction of cataract|After-cataract not obscuring vision following extraction of cataract
C0271193|T047|PT|33048000|SNOMEDCT_CORE|Peripheral visual field defect|Peripheral visual field defect
C0271193|T047|FN|33048000|SNOMEDCT_CORE|Peripheral visual field defect|Peripheral visual field defect
C0271202|T047|SY|34063005|SNOMEDCT_CORE|HH - Homonymous hemianopia|Homonymous hemianopia
C0271202|T047|SY|34063005|SNOMEDCT_CORE|Homonymous bilateral visual field defects|Homonymous hemianopia
C0271202|T047|PT|34063005|SNOMEDCT_CORE|Homonymous hemianopia|Homonymous hemianopia
C0271202|T047|FN|34063005|SNOMEDCT_CORE|Homonymous hemianopia|Homonymous hemianopia
C0271202|T047|IS|34063005|SNOMEDCT_CORE|Homonymous hemianopsia|Homonymous hemianopia
C0271215|T047|PT|65956007|SNOMEDCT_CORE|Legal blindness|Legal blindness
C0271215|T047|FN|65956007|SNOMEDCT_CORE|Legal blindness|Legal blindness
C0271225|T047|PT|91408006|SNOMEDCT_CORE|Impairment level: blindness, one eye - low vision other eye|Impairment level: blindness, one eye - low vision other eye
C0271225|T047|FN|91408006|SNOMEDCT_CORE|Impairment level: blindness, one eye - low vision other eye|Impairment level: blindness, one eye - low vision other eye
C0271234|T047|PT|193722001|SNOMEDCT_CORE|Low vision, both eyes|Low vision, both eyes
C0271234|T047|FN|193722001|SNOMEDCT_CORE|Low vision, both eyes|Low vision, both eyes
C0271240|T047|SY|22950006|SNOMEDCT_CORE|Blind eye|Blindness of one eye
C0271240|T047|FN|22950006|SNOMEDCT_CORE|Blindness of one eye|Blindness of one eye
C0271240|T047|PT|22950006|SNOMEDCT_CORE|Blindness of one eye|Blindness of one eye
C0271240|T047|IS|22950006|SNOMEDCT_CORE|Blindness of one eye, NOS|Blindness of one eye
C0271240|T047|SY|22950006|SNOMEDCT_CORE|Blindness, unilateral|Blindness of one eye
C0271285|T047|SY|373426005|SNOMEDCT_CORE|Anterior basement membrane dystrophy|Epithelial basement membrane dystrophy
C0271285|T047|OAS|32935005|SNOMEDCT_CORE|Cogan microcystic dystrophy|Epithelial basement membrane dystrophy
C0271285|T047|SY|373426005|SNOMEDCT_CORE|Cogan microcystic epithelial dystrophy|Epithelial basement membrane dystrophy
C0271285|T047|OAS|32935005|SNOMEDCT_CORE|Cogan-Guerry syndrome|Epithelial basement membrane dystrophy
C0271285|T047|OAS|32935005|SNOMEDCT_CORE|Cogan's corneal dystrophy|Epithelial basement membrane dystrophy
C0271285|T047|OAS|32935005|SNOMEDCT_CORE|Corneal epithelial basement membrane dystrophy|Epithelial basement membrane dystrophy
C0271285|T047|OAS|32935005|SNOMEDCT_CORE|EBMD - Corneal epithelial basement membrane dystrophy|Epithelial basement membrane dystrophy
C0271285|T047|PT|373426005|SNOMEDCT_CORE|Epithelial basement membrane dystrophy|Epithelial basement membrane dystrophy
C0271285|T047|FN|373426005|SNOMEDCT_CORE|Epithelial basement membrane dystrophy|Epithelial basement membrane dystrophy
C0271285|T047|OAS|32935005|SNOMEDCT_CORE|Map-dot-fingerprint corneal dystrophy|Epithelial basement membrane dystrophy
C0271285|T047|SY|373426005|SNOMEDCT_CORE|Map-dot-fingerprint dystrophy|Epithelial basement membrane dystrophy
C0271285|T047|OAS|32935005|SNOMEDCT_CORE|MDF - Map dot fingerprint corneal dystrophy|Epithelial basement membrane dystrophy
C0271285|T047|SY|373426005|SNOMEDCT_CORE|MDF - Map dot fingerprint dystrophy|Epithelial basement membrane dystrophy
C0271285|T047|OAS|32935005|SNOMEDCT_CORE|MDF - Map-dot-fingerprint corneal dystrophy|Epithelial basement membrane dystrophy
C0271285|T047|OAS|32935005|SNOMEDCT_CORE|Microcystoid epithelial dystrophy|Epithelial basement membrane dystrophy
C0271285|T047|OAP|32935005|SNOMEDCT_CORE|Microscopic cystic corneal dystrophy|Epithelial basement membrane dystrophy
C0271285|T047|SY|373426005|SNOMEDCT_CORE|Microscopic cystic corneal dystrophy|Epithelial basement membrane dystrophy
C0271285|T047|OAF|32935005|SNOMEDCT_CORE|Microscopic cystic corneal dystrophy|Epithelial basement membrane dystrophy
C0271294|T047|PT|26045000|SNOMEDCT_CORE|Chronic allergic conjunctivitis|Chronic allergic conjunctivitis
C0271294|T047|FN|26045000|SNOMEDCT_CORE|Chronic allergic conjunctivitis|Chronic allergic conjunctivitis
C0271294|T047|IS|26045000|SNOMEDCT_CORE|Chronic allergic conjunctivitis, NOS|Chronic allergic conjunctivitis
C0271308|T047|IS|68670009|SNOMEDCT_CORE|Allergic blepharitis|Contact dermatitis of eyelid
C0271308|T047|IS|68670009|SNOMEDCT_CORE|Allergic dermatitis of eyelid|Contact dermatitis of eyelid
C0271308|T047|IS|68670009|SNOMEDCT_CORE|Contact allergy eyelid|Contact dermatitis of eyelid
C0271308|T047|PT|68670009|SNOMEDCT_CORE|Contact dermatitis of eyelid|Contact dermatitis of eyelid
C0271308|T047|FN|68670009|SNOMEDCT_CORE|Contact dermatitis of eyelid|Contact dermatitis of eyelid
C0271308|T047|SY|68670009|SNOMEDCT_CORE|Contact eczema eyelid|Contact dermatitis of eyelid
C0271311|T047|IS|60332004|SNOMEDCT_CORE|Trichiasis without entropion|Trichiasis without entropion
C0271355|T047|SY|398925009|SNOMEDCT_CORE|Abducens nerve disease|Abducens nerve disorder
C0271355|T047|PT|398925009|SNOMEDCT_CORE|Abducens nerve disorder|Abducens nerve disorder
C0271355|T047|FN|398925009|SNOMEDCT_CORE|Abducens nerve disorder|Abducens nerve disorder
C0271355|T047|SY|398925009|SNOMEDCT_CORE|Lateral rectus muscle innervation disorder|Abducens nerve disorder
C0271355|T047|SY|398925009|SNOMEDCT_CORE|Sixth cranial nerve disease|Abducens nerve disorder
C0271355|T047|SY|398925009|SNOMEDCT_CORE|Sixth cranial nerve disorder|Abducens nerve disorder
C0271370|T047|OAS|3171005|SNOMEDCT_CORE|Partial oculomotor nerve palsy|Partial oculomotor nerve palsy
C0271370|T047|PT|194118007|SNOMEDCT_CORE|Partial oculomotor nerve palsy|Partial oculomotor nerve palsy
C0271370|T047|FN|194118007|SNOMEDCT_CORE|Partial oculomotor nerve palsy|Partial oculomotor nerve palsy
C0271370|T047|OAS|3171005|SNOMEDCT_CORE|Partial third cranial nerve paralysis|Partial oculomotor nerve palsy
C0271370|T047|OAP|3171005|SNOMEDCT_CORE|Partial third nerve palsy|Partial oculomotor nerve palsy
C0271370|T047|OAF|3171005|SNOMEDCT_CORE|Partial third nerve palsy|Partial oculomotor nerve palsy
C0271370|T047|IS|194118007|SNOMEDCT_CORE|Pupil-sparing third nerve palsy|Partial oculomotor nerve palsy
C0271370|T047|SY|194118007|SNOMEDCT_CORE|Third nerve palsy - partial|Partial oculomotor nerve palsy
C0271370|T047|IS|194118007|SNOMEDCT_CORE|Third nerve palsy with pupil sparing|Partial oculomotor nerve palsy
C0271375|T047|SY|20610004|SNOMEDCT_CORE|4th nerve palsy|Fourth nerve palsy
C0271375|T047|IS|20610004|SNOMEDCT_CORE|Disorder of trochlear nerve|Fourth nerve palsy
C0271375|T047|IS|20610004|SNOMEDCT_CORE|Fourth cranial nerve disease|Fourth nerve palsy
C0271375|T047|IS|20610004|SNOMEDCT_CORE|Fourth cranial nerve disorder|Fourth nerve palsy
C0271375|T047|SY|20610004|SNOMEDCT_CORE|Fourth cranial nerve palsy|Fourth nerve palsy
C0271375|T047|SY|20610004|SNOMEDCT_CORE|Fourth cranial nerve paralysis|Fourth nerve palsy
C0271375|T047|SY|20610004|SNOMEDCT_CORE|Fourth cranial nerve paresis|Fourth nerve palsy
C0271375|T047|PT|20610004|SNOMEDCT_CORE|Fourth nerve palsy|Fourth nerve palsy
C0271375|T047|FN|20610004|SNOMEDCT_CORE|Fourth nerve palsy|Fourth nerve palsy
C0271375|T047|SY|20610004|SNOMEDCT_CORE|IV nerve palsy|Fourth nerve palsy
C0271375|T047|IS|20610004|SNOMEDCT_CORE|Superior oblique muscle innervation disorder|Fourth nerve palsy
C0271375|T047|SY|20610004|SNOMEDCT_CORE|Superior oblique palsy|Fourth nerve palsy
C0271375|T047|IS|20610004|SNOMEDCT_CORE|Trochlear nerve disease|Fourth nerve palsy
C0271375|T047|IS|20610004|SNOMEDCT_CORE|Trochlear nerve disorder|Fourth nerve palsy
C0271375|T047|SY|20610004|SNOMEDCT_CORE|Trochlear nerve palsy|Fourth nerve palsy
C0271375|T047|SY|20610004|SNOMEDCT_CORE|Trochlear nerve paralysis|Fourth nerve palsy
C0271375|T047|SY|20610004|SNOMEDCT_CORE|Trochlear nerve weakness|Fourth nerve palsy
C0271379|T047|SY|194131002|SNOMEDCT_CORE|CI - Convergence insufficiency|Convergence insufficiency
C0271379|T047|PT|194131002|SNOMEDCT_CORE|Convergence insufficiency|Convergence insufficiency
C0271379|T047|FN|194131002|SNOMEDCT_CORE|Convergence insufficiency|Convergence insufficiency
C0271381|T033|PT|40631009|SNOMEDCT_CORE|Skew deviation|Skew deviation
C0271381|T033|FN|40631009|SNOMEDCT_CORE|Skew deviation|Skew deviation
C0271413|T046|SYGB|88050005|SNOMEDCT_CORE|Haematoma of auricle|Hematoma of pinna
C0271413|T046|PTGB|88050005|SNOMEDCT_CORE|Haematoma of pinna|Hematoma of pinna
C0271413|T046|SY|88050005|SNOMEDCT_CORE|Hematoma of auricle|Hematoma of pinna
C0271413|T046|PT|88050005|SNOMEDCT_CORE|Hematoma of pinna|Hematoma of pinna
C0271413|T046|FN|88050005|SNOMEDCT_CORE|Hematoma of pinna|Hematoma of pinna
C0271420|T047|IS|18070006|SNOMEDCT_CORE|Excess wax in ear|Excess wax in ear
C0271429|T047|PT|3110003|SNOMEDCT_CORE|Acute otitis media|Acute otitis media
C0271429|T047|FN|3110003|SNOMEDCT_CORE|Acute otitis media|Acute otitis media
C0271429|T047|IS|3110003|SNOMEDCT_CORE|Acute otitis media, NOS|Acute otitis media
C0271429|T047|SY|3110003|SNOMEDCT_CORE|AOM - Acute otitis media|Acute otitis media
C0271432|T047|SY|35183001|SNOMEDCT_CORE|Acute MEE - Acute middle ear effusion|Acute transudative otitis media
C0271432|T047|SY|35183001|SNOMEDCT_CORE|Acute middle ear effusion|Acute transudative otitis media
C0271432|T047|IS|35183001|SNOMEDCT_CORE|Acute otitis media with effusion|Acute transudative otitis media
C0271432|T047|PT|35183001|SNOMEDCT_CORE|Acute transudative otitis media|Acute transudative otitis media
C0271432|T047|FN|35183001|SNOMEDCT_CORE|Acute transudative otitis media|Acute transudative otitis media
C0271441|T047|PT|21186006|SNOMEDCT_CORE|Chronic otitis media|Chronic otitis media
C0271441|T047|FN|21186006|SNOMEDCT_CORE|Chronic otitis media|Chronic otitis media
C0271441|T047|IS|21186006|SNOMEDCT_CORE|Chronic otitis media, NOS|Chronic otitis media
C0271446|T047|PT|275481002|SNOMEDCT_CORE|Non-suppurative otitis media|Non-suppurative otitis media
C0271446|T047|FN|275481002|SNOMEDCT_CORE|Non-suppurative otitis media|Non-suppurative otitis media
C0271453|T047|PT|80327007|SNOMEDCT_CORE|Serous otitis media|Serous otitis media
C0271453|T047|FN|80327007|SNOMEDCT_CORE|Serous otitis media|Serous otitis media
C0271454|T047|IS|38394007|SNOMEDCT_CORE|Chronic non-suppurative otitis media with effusion - purulent|Chronic purulent otitis media
C0271454|T047|SY|38394007|SNOMEDCT_CORE|Chronic otitis media with effusion, purulent|Chronic purulent otitis media
C0271454|T047|PT|38394007|SNOMEDCT_CORE|Chronic purulent otitis media|Chronic purulent otitis media
C0271454|T047|FN|38394007|SNOMEDCT_CORE|Chronic purulent otitis media|Chronic purulent otitis media
C0271454|T047|SY|38394007|SNOMEDCT_CORE|Chronic secretory otitis media, purulent|Chronic purulent otitis media
C0271454|T047|SY|38394007|SNOMEDCT_CORE|Chronic suppurative otitis media|Chronic purulent otitis media
C0271454|T047|SY|38394007|SNOMEDCT_CORE|CSOM - Chronic suppurative otitis media|Chronic purulent otitis media
C0271468|T047|SY|69494008|SNOMEDCT_CORE|Auditory tube disorder|Eustachian tube disorder
C0271468|T047|SY|69494008|SNOMEDCT_CORE|Disease of Eustachian tube|Eustachian tube disorder
C0271468|T047|SY|69494008|SNOMEDCT_CORE|Disorder of Eustachian tube|Eustachian tube disorder
C0271468|T047|PT|56713002|SNOMEDCT_CORE|Dysfunction of eustachian tube|Eustachian tube disorder
C0271468|T047|FN|56713002|SNOMEDCT_CORE|Dysfunction of eustachian tube|Eustachian tube disorder
C0271468|T047|SY|69494008|SNOMEDCT_CORE|ET - Eustachian tube disorder|Eustachian tube disorder
C0271468|T047|SY|56713002|SNOMEDCT_CORE|ETD - Eustachian tube dysfunction|Eustachian tube disorder
C0271468|T047|IS|56713002|SNOMEDCT_CORE|Eustachian tube dis.|Eustachian tube disorder
C0271468|T047|IS|69494008|SNOMEDCT_CORE|Eustachian tube dis.|Eustachian tube disorder
C0271468|T047|PT|69494008|SNOMEDCT_CORE|Eustachian tube disorder|Eustachian tube disorder
C0271468|T047|FN|69494008|SNOMEDCT_CORE|Eustachian tube disorder|Eustachian tube disorder
C0271468|T047|IS|69494008|SNOMEDCT_CORE|Eustachian tube disorder, NOS|Eustachian tube disorder
C0271468|T047|SY|56713002|SNOMEDCT_CORE|Eustachian tube dysfunction|Eustachian tube disorder
C0271476|T047|SY|52404001|SNOMEDCT_CORE|Mastoid empyema|Mastoid empyemia
C0271476|T047|IS|52404001|SNOMEDCT_CORE|Mastoid empyemia|Mastoid empyemia
C0271503|T047|PT|65680009|SNOMEDCT_CORE|Sensorineural hearing loss of combined sites|Sensorineural hearing loss of combined sites
C0271503|T047|OF|65680009|SNOMEDCT_CORE|Sensorineural hearing loss of combined sites|Sensorineural hearing loss of combined sites
C0271503|T047|FN|65680009|SNOMEDCT_CORE|Sensorineural hearing loss of combined sites|Sensorineural hearing loss of combined sites
C0271561|T047|OAS|44008002|SNOMEDCT_CORE|GHD|Growth hormone deficiency
C0271561|T047|SY|397827003|SNOMEDCT_CORE|GHD - Growth hormone deficiency|Growth hormone deficiency
C0271561|T047|OAS|44008002|SNOMEDCT_CORE|Growth hormone deficiency|Growth hormone deficiency
C0271561|T047|PT|397827003|SNOMEDCT_CORE|Growth hormone deficiency|Growth hormone deficiency
C0271561|T047|FN|397827003|SNOMEDCT_CORE|Growth hormone deficiency|Growth hormone deficiency
C0271561|T047|IS|44008002|SNOMEDCT_CORE|Growth hormone deficiency, NOS|Growth hormone deficiency
C0271561|T047|SY|397827003|SNOMEDCT_CORE|Growth hormone insufficiency|Growth hormone deficiency
C0271561|T047|OAP|44008002|SNOMEDCT_CORE|Somatotropin deficiency|Growth hormone deficiency
C0271561|T047|OAF|44008002|SNOMEDCT_CORE|Somatotropin deficiency|Growth hormone deficiency
C0271561|T047|IS|44008002|SNOMEDCT_CORE|Somatotropin deficiency, NOS|Growth hormone deficiency
C0271561|T047|OAS|44008002|SNOMEDCT_CORE|STH deficiency|Growth hormone deficiency
C0271578|T047|SY|16041008|SNOMEDCT_CORE|Female hypogonadism|Female hypogonadism syndrome
C0271578|T047|PT|16041008|SNOMEDCT_CORE|Female hypogonadism syndrome|Female hypogonadism syndrome
C0271578|T047|FN|16041008|SNOMEDCT_CORE|Female hypogonadism syndrome|Female hypogonadism syndrome
C0271578|T047|IS|16041008|SNOMEDCT_CORE|Female hypogonadism syndrome, NOS|Female hypogonadism syndrome
C0271622|T047|PT|111551000|SNOMEDCT_CORE|Testicular hypofunction|Testicular hypofunction
C0271622|T047|FN|111551000|SNOMEDCT_CORE|Testicular hypofunction|Testicular hypofunction
C0271623|T047|SY|33927004|SNOMEDCT_CORE|Gonadotrophin deficiency|Hypogonadotropic hypogonadism
C0271623|T047|PT|33927004|SNOMEDCT_CORE|Hypogonadotropic hypogonadism|Hypogonadotropic hypogonadism
C0271623|T047|FN|33927004|SNOMEDCT_CORE|Hypogonadotropic hypogonadism|Hypogonadotropic hypogonadism
C0271623|T047|SY|33927004|SNOMEDCT_CORE|Secondary hypogonadism|Hypogonadotropic hypogonadism
C0271623|T047|IS|33927004|SNOMEDCT_CORE|Secondary hypogonadism, NOS|Hypogonadotropic hypogonadism
C0271638|T047|SY|81531005|SNOMEDCT_CORE|Diabetes mellitus type 2 in obese|Type 2 diabetes mellitus in obese
C0271638|T047|FN|81531005|SNOMEDCT_CORE|Diabetes mellitus type 2 in obese|Type 2 diabetes mellitus in obese
C0271638|T047|IS|81531005|SNOMEDCT_CORE|NIDDM in obese|Type 2 diabetes mellitus in obese
C0271638|T047|PT|81531005|SNOMEDCT_CORE|Type 2 diabetes mellitus in obese|Type 2 diabetes mellitus in obese
C0271650|T047|SY|9414007|SNOMEDCT_CORE|Chemical diabetes|Impaired glucose tolerance
C0271650|T047|SY|9414007|SNOMEDCT_CORE|IGT - Impaired glucose tolerance|Impaired glucose tolerance
C0271650|T047|PT|9414007|SNOMEDCT_CORE|Impaired glucose tolerance|Impaired glucose tolerance
C0271650|T047|FN|9414007|SNOMEDCT_CORE|Impaired glucose tolerance|Impaired glucose tolerance
C0271650|T047|IS|9414007|SNOMEDCT_CORE|Impaired glucose tolerance, NOS|Impaired glucose tolerance
C0271650|T047|SY|9414007|SNOMEDCT_CORE|Latent diabetes|Impaired glucose tolerance
C0271650|T047|SY|9414007|SNOMEDCT_CORE|Prediabetic nonclinical diabetes|Impaired glucose tolerance
C0271663|T047|MTH_SY|46894009|SNOMEDCT_CORE|GDM, class A<sub>2</sub>|Gestational diabetes mellitus, class A>2<
C0271663|T047|SY|46894009|SNOMEDCT_CORE|GDM, class A>2<|Gestational diabetes mellitus, class A>2<
C0271663|T047|MTH_SY|46894009|SNOMEDCT_CORE|GDM, class A2|Gestational diabetes mellitus, class A>2<
C0271663|T047|MTH_FN|46894009|SNOMEDCT_CORE|Gestational diabetes mellitus, class A<sub>2</sub>|Gestational diabetes mellitus, class A>2<
C0271663|T047|MTH_PT|46894009|SNOMEDCT_CORE|Gestational diabetes mellitus, class A<sub>2</sub>|Gestational diabetes mellitus, class A>2<
C0271663|T047|PT|46894009|SNOMEDCT_CORE|Gestational diabetes mellitus, class A>2<|Gestational diabetes mellitus, class A>2<
C0271663|T047|FN|46894009|SNOMEDCT_CORE|Gestational diabetes mellitus, class A>2<|Gestational diabetes mellitus, class A>2<
C0271663|T047|MTH_PT|46894009|SNOMEDCT_CORE|Gestational diabetes mellitus, class A2|Gestational diabetes mellitus, class A>2<
C0271663|T047|MTH_FN|46894009|SNOMEDCT_CORE|Gestational diabetes mellitus, class A2|Gestational diabetes mellitus, class A>2<
C0271678|T047|PT|230577008|SNOMEDCT_CORE|Diabetic mononeuropathy|Diabetic mononeuropathy
C0271678|T047|OF|230577008|SNOMEDCT_CORE|Diabetic mononeuropathy|Diabetic mononeuropathy
C0271678|T047|IS|230577008|SNOMEDCT_CORE|Mononeuropathy co-occurrent and due to diabetes mellitus|Diabetic mononeuropathy
C0271678|T047|OF|230577008|SNOMEDCT_CORE|Mononeuropathy co-occurrent and due to diabetes mellitus|Diabetic mononeuropathy
C0271678|T047|SY|230577008|SNOMEDCT_CORE|Mononeuropathy due to diabetes mellitus|Diabetic mononeuropathy
C0271678|T047|FN|230577008|SNOMEDCT_CORE|Mononeuropathy due to diabetes mellitus|Diabetic mononeuropathy
C0271680|T047|SY|49455004|SNOMEDCT_CORE|Diabetic polyneuropathy|Polyneuropathy due to diabetes mellitus
C0271680|T047|OF|49455004|SNOMEDCT_CORE|Diabetic polyneuropathy|Polyneuropathy due to diabetes mellitus
C0271680|T047|IS|49455004|SNOMEDCT_CORE|Diabetic polyneuropathy, NOS|Polyneuropathy due to diabetes mellitus
C0271680|T047|IS|49455004|SNOMEDCT_CORE|Polyneuropathy co-occurrent and due to diabetes mellitus|Polyneuropathy due to diabetes mellitus
C0271680|T047|OF|49455004|SNOMEDCT_CORE|Polyneuropathy co-occurrent and due to diabetes mellitus|Polyneuropathy due to diabetes mellitus
C0271680|T047|PT|49455004|SNOMEDCT_CORE|Polyneuropathy due to diabetes mellitus|Polyneuropathy due to diabetes mellitus
C0271680|T047|FN|49455004|SNOMEDCT_CORE|Polyneuropathy due to diabetes mellitus|Polyneuropathy due to diabetes mellitus
C0271686|T047|IS|50620007|SNOMEDCT_CORE|Autonomic neuropathy co-occurrent and due to diabetes mellitus|Autonomic neuropathy due to diabetes mellitus
C0271686|T047|OF|50620007|SNOMEDCT_CORE|Autonomic neuropathy co-occurrent and due to diabetes mellitus|Autonomic neuropathy due to diabetes mellitus
C0271686|T047|SY|50620007|SNOMEDCT_CORE|Autonomic neuropathy due to diabetes|Autonomic neuropathy due to diabetes mellitus
C0271686|T047|PT|50620007|SNOMEDCT_CORE|Autonomic neuropathy due to diabetes mellitus|Autonomic neuropathy due to diabetes mellitus
C0271686|T047|FN|50620007|SNOMEDCT_CORE|Autonomic neuropathy due to diabetes mellitus|Autonomic neuropathy due to diabetes mellitus
C0271686|T047|SY|50620007|SNOMEDCT_CORE|Autonomic neuropathy with diabetes mellitus|Autonomic neuropathy due to diabetes mellitus
C0271686|T047|SY|50620007|SNOMEDCT_CORE|Diabetic autonomic neuropathy|Autonomic neuropathy due to diabetes mellitus
C0271686|T047|OF|50620007|SNOMEDCT_CORE|Diabetic autonomic neuropathy|Autonomic neuropathy due to diabetes mellitus
C0271710|T047|SYGB|317006|SNOMEDCT_CORE|Hypoglycaemic reaction|Reactive hypoglycemia
C0271710|T047|SY|317006|SNOMEDCT_CORE|Hypoglycemic reaction|Reactive hypoglycemia
C0271710|T047|PTGB|317006|SNOMEDCT_CORE|Reactive hypoglycaemia|Reactive hypoglycemia
C0271710|T047|PT|317006|SNOMEDCT_CORE|Reactive hypoglycemia|Reactive hypoglycemia
C0271710|T047|FN|317006|SNOMEDCT_CORE|Reactive hypoglycemia|Reactive hypoglycemia
C0271725|T047|SY|41299009|SNOMEDCT_CORE|Drug-induced Cushing's syndrome|Iatrogenic Cushing's disease
C0271725|T047|SY|41299009|SNOMEDCT_CORE|Iatrogenic Cushing disease|Iatrogenic Cushing's disease
C0271725|T047|PT|41299009|SNOMEDCT_CORE|Iatrogenic Cushing's disease|Iatrogenic Cushing's disease
C0271725|T047|FN|41299009|SNOMEDCT_CORE|Iatrogenic Cushing's disease|Iatrogenic Cushing's disease
C0271725|T047|SY|41299009|SNOMEDCT_CORE|Iatrogenic Cushing's syndrome|Iatrogenic Cushing's disease
C0271725|T047|SY|41299009|SNOMEDCT_CORE|Iatrogenic syndrome of excess cortisol|Iatrogenic Cushing's disease
C0271761|T047|SY|36241006|SNOMEDCT_CORE|Multinodular non-toxic goiter|Non-toxic multinodular goiter
C0271761|T047|SYGB|36241006|SNOMEDCT_CORE|Multinodular non-toxic goitre|Non-toxic multinodular goiter
C0271761|T047|PT|36241006|SNOMEDCT_CORE|Non-toxic multinodular goiter|Non-toxic multinodular goiter
C0271761|T047|FN|36241006|SNOMEDCT_CORE|Non-toxic multinodular goiter|Non-toxic multinodular goiter
C0271761|T047|PTGB|36241006|SNOMEDCT_CORE|Non-toxic multinodular goitre|Non-toxic multinodular goiter
C0271790|T047|SY|54823002|SNOMEDCT_CORE|Borderline hypothyroidism|Subclinical hypothyroidism
C0271790|T047|SY|54823002|SNOMEDCT_CORE|Compensated euthyroidism|Subclinical hypothyroidism
C0271790|T047|PT|54823002|SNOMEDCT_CORE|Subclinical hypothyroidism|Subclinical hypothyroidism
C0271790|T047|FN|54823002|SNOMEDCT_CORE|Subclinical hypothyroidism|Subclinical hypothyroidism
C0271803|T047|PT|88273006|SNOMEDCT_CORE|Iatrogenic hypothyroidism|Iatrogenic hypothyroidism
C0271803|T047|FN|88273006|SNOMEDCT_CORE|Iatrogenic hypothyroidism|Iatrogenic hypothyroidism
C0271847|T047|PT|19034001|SNOMEDCT_CORE|Hyperparathyroidism due to renal insufficiency|Hyperparathyroidism due to renal insufficiency
C0271847|T047|FN|19034001|SNOMEDCT_CORE|Hyperparathyroidism due to renal insufficiency|Hyperparathyroidism due to renal insufficiency
C0271847|T047|SY|19034001|SNOMEDCT_CORE|Secondary hyperparathyroidism of renal origin|Hyperparathyroidism due to renal insufficiency
C0271864|T047|SY|37605006|SNOMEDCT_CORE|Osteopenia of the elderly|Senile osteopenia
C0271864|T047|PT|37605006|SNOMEDCT_CORE|Senile osteopenia|Senile osteopenia
C0271864|T047|FN|37605006|SNOMEDCT_CORE|Senile osteopenia|Senile osteopenia
C0271892|T047|PT|5876000|SNOMEDCT_CORE|Acquired pancytopenia|Acquired pancytopenia
C0271892|T047|FN|5876000|SNOMEDCT_CORE|Acquired pancytopenia|Acquired pancytopenia
C0271892|T047|SY|5876000|SNOMEDCT_CORE|Pancytopenia - acquired|Acquired pancytopenia
C0271901|T047|SYGB|44666001|SNOMEDCT_CORE|Hypochromic microcytic anaemia|Microcytic hypochromic anemia
C0271901|T047|SY|44666001|SNOMEDCT_CORE|Hypochromic microcytic anemia|Microcytic hypochromic anemia
C0271901|T047|PTGB|44666001|SNOMEDCT_CORE|Microcytic hypochromic anaemia|Microcytic hypochromic anemia
C0271901|T047|FN|44666001|SNOMEDCT_CORE|Microcytic hypochromic anemia|Microcytic hypochromic anemia
C0271901|T047|PT|44666001|SNOMEDCT_CORE|Microcytic hypochromic anemia|Microcytic hypochromic anemia
C0271930|T047|PTGB|27342004|SNOMEDCT_CORE|Anaemia of pregnancy|Anemia of pregnancy
C0271930|T047|PT|27342004|SNOMEDCT_CORE|Anemia of pregnancy|Anemia of pregnancy
C0271930|T047|FN|27342004|SNOMEDCT_CORE|Anemia of pregnancy|Anemia of pregnancy
C0271932|T047|PTGB|49708008|SNOMEDCT_CORE|Anaemia of chronic renal failure|Anemia of chronic renal failure
C0271932|T047|SYGB|49708008|SNOMEDCT_CORE|Anaemia of chronic renal insufficiency|Anemia of chronic renal failure
C0271932|T047|PT|49708008|SNOMEDCT_CORE|Anemia of chronic renal failure|Anemia of chronic renal failure
C0271932|T047|FN|49708008|SNOMEDCT_CORE|Anemia of chronic renal failure|Anemia of chronic renal failure
C0271932|T047|SY|49708008|SNOMEDCT_CORE|Anemia of chronic renal insufficiency|Anemia of chronic renal failure
C0272009|T047|PTGB|79035003|SNOMEDCT_CORE|Anaemia due to unknown mechanism|Anemia due to unknown mechanism
C0272009|T047|IS|79035003|SNOMEDCT_CORE|Anaemia due to unknown mechanism, NOS|Anemia due to unknown mechanism
C0272009|T047|PT|79035003|SNOMEDCT_CORE|Anemia due to unknown mechanism|Anemia due to unknown mechanism
C0272009|T047|FN|79035003|SNOMEDCT_CORE|Anemia due to unknown mechanism|Anemia due to unknown mechanism
C0272009|T047|IS|79035003|SNOMEDCT_CORE|Anemia due to unknown mechanism, NOS|Anemia due to unknown mechanism
C0272153|T047|PTGB|32984002|SNOMEDCT_CORE|Neonatal polycythaemia|Neonatal polycythemia
C0272153|T047|PT|32984002|SNOMEDCT_CORE|Neonatal polycythemia|Neonatal polycythemia
C0272153|T047|FN|32984002|SNOMEDCT_CORE|Neonatal polycythemia|Neonatal polycythemia
C0272153|T047|SY|32984002|SNOMEDCT_CORE|Plethora of newborn|Neonatal polycythemia
C0272153|T047|SYGB|32984002|SNOMEDCT_CORE|Polycythaemia neonatorum|Neonatal polycythemia
C0272153|T047|SY|32984002|SNOMEDCT_CORE|Polycythemia neonatorum|Neonatal polycythemia
C0272210|T047|OAP|16944002|SNOMEDCT_CORE|Mononucleosis syndrome|Mononucleosis syndrome
C0272210|T047|OAF|16944002|SNOMEDCT_CORE|Mononucleosis syndrome|Mononucleosis syndrome
C0272210|T047|IS|16944002|SNOMEDCT_CORE|Mononucleosis syndrome, NOS|Mononucleosis syndrome
C0272286|T047|FN|2897005|SNOMEDCT_CORE|Immune thrombocytopenia|Immune thrombocytopenia
C0272286|T047|PT|2897005|SNOMEDCT_CORE|Immune thrombocytopenia|Immune thrombocytopenia
C0272286|T047|SY|2897005|SNOMEDCT_CORE|Thrombocytopenia due to immune destruction|Immune thrombocytopenia
C0272286|T047|IS|2897005|SNOMEDCT_CORE|Thrombocytopenia due to immune destruction, NOS|Immune thrombocytopenia
C0272286|T047|IS|2897005|SNOMEDCT_CORE|Thrombocytopenia due to platelet alloimmunization|Immune thrombocytopenia
C0272290|T047|PT|19307009|SNOMEDCT_CORE|Drug-induced immune thrombocytopenia|Drug-induced immune thrombocytopenia
C0272290|T047|FN|19307009|SNOMEDCT_CORE|Drug-induced immune thrombocytopenia|Drug-induced immune thrombocytopenia
C0272290|T047|SY|19307009|SNOMEDCT_CORE|Drug-induced ITP|Drug-induced immune thrombocytopenia
C0272290|T047|SY|19307009|SNOMEDCT_CORE|Drug-induced thrombocytopenic purpura|Drug-induced immune thrombocytopenia
C0272316|T047|PT|16922007|SNOMEDCT_CORE|Hereditary coagulation factor deficiency|Hereditary coagulation factor deficiency
C0272316|T047|FN|16922007|SNOMEDCT_CORE|Hereditary coagulation factor deficiency|Hereditary coagulation factor deficiency
C0272316|T047|IS|16922007|SNOMEDCT_CORE|Hereditary coagulation factor deficiency, NOS|Hereditary coagulation factor deficiency
C0272386|T047|SY|46689006|SNOMEDCT_CORE|Enlargement of tonsils|Hypertrophy of tonsils
C0272386|T047|PT|46689006|SNOMEDCT_CORE|Hypertrophy of tonsils|Hypertrophy of tonsils
C0272386|T047|FN|46689006|SNOMEDCT_CORE|Hypertrophy of tonsils|Hypertrophy of tonsils
C0272386|T047|SY|46689006|SNOMEDCT_CORE|Tonsillar enlargement|Hypertrophy of tonsils
C0272386|T047|SY|46689006|SNOMEDCT_CORE|Tonsillar hypertrophy|Hypertrophy of tonsils
C0272388|T047|PT|6461009|SNOMEDCT_CORE|Amygdalolith|Amygdalolith
C0272388|T047|FN|6461009|SNOMEDCT_CORE|Amygdalolith|Amygdalolith
C0272388|T047|SY|6461009|SNOMEDCT_CORE|Calculus of tonsil|Amygdalolith
C0272388|T047|SY|6461009|SNOMEDCT_CORE|Tonsil stone|Amygdalolith
C0272388|T047|SY|6461009|SNOMEDCT_CORE|Tonsillar calculus|Amygdalolith
C0272388|T047|SY|6461009|SNOMEDCT_CORE|Tonsillith|Amygdalolith
C0272388|T047|SY|6461009|SNOMEDCT_CORE|Tonsillolith|Amygdalolith
C0272388|T047|SY|6461009|SNOMEDCT_CORE|Tonsillolithiasis|Amygdalolith
C0272452|T037|PT|69866009|SNOMEDCT_CORE|Closed fracture of vault of skull without intracranial injury|Closed fracture of vault of skull without intracranial injury
C0272452|T037|FN|69866009|SNOMEDCT_CORE|Closed fracture of vault of skull without intracranial injury|Closed fracture of vault of skull without intracranial injury
C0272504|T037|PT|42157000|SNOMEDCT_CORE|Closed fracture of vertebral column|Closed fracture of vertebral column
C0272504|T037|FN|42157000|SNOMEDCT_CORE|Closed fracture of vertebral column|Closed fracture of vertebral column
C0272504|T037|IS|42157000|SNOMEDCT_CORE|Closed fracture of vertebral column, NOS|Closed fracture of vertebral column
C0272530|T037|SY|89825003|SNOMEDCT_CORE|Closed fracture of dorsal vertebra without spinal cord injury|Closed fracture of thoracic vertebra without spinal cord injury
C0272530|T037|PT|89825003|SNOMEDCT_CORE|Closed fracture of thoracic vertebra without spinal cord injury|Closed fracture of thoracic vertebra without spinal cord injury
C0272530|T037|FN|89825003|SNOMEDCT_CORE|Closed fracture of thoracic vertebra without spinal cord injury|Closed fracture of thoracic vertebra without spinal cord injury
C0272532|T037|PT|17463000|SNOMEDCT_CORE|Closed fracture of lumbar vertebra without spinal cord injury|Closed fracture of lumbar vertebra without spinal cord injury
C0272532|T037|FN|17463000|SNOMEDCT_CORE|Closed fracture of lumbar vertebra without spinal cord injury|Closed fracture of lumbar vertebra without spinal cord injury
C0272567|T037|PT|1261007|SNOMEDCT_CORE|Fracture of multiple ribs|Fracture of multiple ribs
C0272567|T037|FN|1261007|SNOMEDCT_CORE|Fracture of multiple ribs|Fracture of multiple ribs
C0272567|T037|IS|1261007|SNOMEDCT_CORE|Fracture of multiple ribs, NOS|Fracture of multiple ribs
C0272567|T037|SY|1261007|SNOMEDCT_CORE|Multiple fractures of ribs|Fracture of multiple ribs
C0272576|T037|PT|91037003|SNOMEDCT_CORE|Closed fracture of pelvis|Closed fracture of pelvis
C0272576|T037|FN|91037003|SNOMEDCT_CORE|Closed fracture of pelvis|Closed fracture of pelvis
C0272576|T037|IS|91037003|SNOMEDCT_CORE|Closed fracture of pelvis, NOS|Closed fracture of pelvis
C0272609|T037|PT|43295006|SNOMEDCT_CORE|Closed fracture of humerus|Closed fracture of humerus
C0272609|T037|FN|43295006|SNOMEDCT_CORE|Closed fracture of humerus|Closed fracture of humerus
C0272609|T037|IS|43295006|SNOMEDCT_CORE|Closed fracture of humerus, NOS|Closed fracture of humerus
C0272609|T037|SY|43295006|SNOMEDCT_CORE|Closed fracture of upper arm|Closed fracture of humerus
C0272609|T037|IS|43295006|SNOMEDCT_CORE|Closed fracture of upper arm, NOS|Closed fracture of humerus
C0272622|T037|PT|111640008|SNOMEDCT_CORE|Closed fracture of radius|Closed fracture of radius
C0272622|T037|FN|111640008|SNOMEDCT_CORE|Closed fracture of radius|Closed fracture of radius
C0272624|T037|PT|53627009|SNOMEDCT_CORE|Closed fracture of radius AND ulna|Closed fracture of radius AND ulna
C0272624|T037|IS|53627009|SNOMEDCT_CORE|Closed fracture of radius and ulna|Closed fracture of radius AND ulna
C0272624|T037|FN|53627009|SNOMEDCT_CORE|Closed fracture of radius AND ulna|Closed fracture of radius AND ulna
C0272624|T037|SY|53627009|SNOMEDCT_CORE|Closed fracture of the radius and ulna|Closed fracture of radius AND ulna
C0272637|T037|PT|28078000|SNOMEDCT_CORE|Closed fracture of shaft of bone of forearm|Closed fracture of shaft of bone of forearm
C0272637|T037|FN|28078000|SNOMEDCT_CORE|Closed fracture of shaft of bone of forearm|Closed fracture of shaft of bone of forearm
C0272637|T037|IS|28078000|SNOMEDCT_CORE|Closed fracture of shaft of bone of forearm, NOS|Closed fracture of shaft of bone of forearm
C0272637|T037|SY|28078000|SNOMEDCT_CORE|Closed fracture of shaft of radius and/or ulna|Closed fracture of shaft of bone of forearm
C0272638|T037|PT|3228009|SNOMEDCT_CORE|Closed fracture of shaft of radius|Closed fracture of shaft of radius
C0272638|T037|FN|3228009|SNOMEDCT_CORE|Closed fracture of shaft of radius|Closed fracture of shaft of radius
C0272638|T037|SY|3228009|SNOMEDCT_CORE|Closed fracture of the radial shaft|Closed fracture of shaft of radius
C0272644|T037|PT|17222009|SNOMEDCT_CORE|Closed fracture of distal end of radius|Closed fracture of distal end of radius
C0272644|T037|FN|17222009|SNOMEDCT_CORE|Closed fracture of distal end of radius|Closed fracture of distal end of radius
C0272644|T037|IS|17222009|SNOMEDCT_CORE|Closed fracture of distal end of radius, NOS|Closed fracture of distal end of radius
C0272644|T037|SY|17222009|SNOMEDCT_CORE|Closed fracture of lower end of radius|Closed fracture of distal end of radius
C0272644|T037|IS|17222009|SNOMEDCT_CORE|Closed fracture of lower end of radius, NOS|Closed fracture of distal end of radius
C0272647|T037|PT|50397009|SNOMEDCT_CORE|Closed fracture of distal end of ulna|Closed fracture of distal end of ulna
C0272647|T037|FN|50397009|SNOMEDCT_CORE|Closed fracture of distal end of ulna|Closed fracture of distal end of ulna
C0272647|T037|SY|50397009|SNOMEDCT_CORE|Closed fracture of lower end of ulna|Closed fracture of distal end of ulna
C0272647|T037|SY|50397009|SNOMEDCT_CORE|Closed fracture of lower epiphysis|Closed fracture of distal end of ulna
C0272654|T037|SY|31975004|SNOMEDCT_CORE|Fracture of navicular bone of wrist|Fracture of scaphoid bone of wrist
C0272654|T037|FN|31975004|SNOMEDCT_CORE|Fracture of navicular bone of wrist|Fracture of scaphoid bone of wrist
C0272654|T037|SY|31975004|SNOMEDCT_CORE|Fracture of scaphoid bone|Fracture of scaphoid bone of wrist
C0272654|T037|PT|31975004|SNOMEDCT_CORE|Fracture of scaphoid bone of wrist|Fracture of scaphoid bone of wrist
C0272677|T037|PT|208393000|SNOMEDCT_CORE|Fracture of metacarpal bone|Fracture of metacarpal bone
C0272677|T037|FN|208393000|SNOMEDCT_CORE|Fracture of metacarpal bone|Fracture of metacarpal bone
C0272677|T037|SY|208393000|SNOMEDCT_CORE|Fracture of metacarpus|Fracture of metacarpal bone
C0272677|T037|SY|208393000|SNOMEDCT_CORE|Hand fracture - metacarpal bone|Fracture of metacarpal bone
C0272686|T037|PT|54641008|SNOMEDCT_CORE|Closed fracture of base of metacarpal bone other than first metacarpal|Closed fracture of base of metacarpal bone other than first metacarpal
C0272686|T037|FN|54641008|SNOMEDCT_CORE|Closed fracture of base of metacarpal bone other than first metacarpal|Closed fracture of base of metacarpal bone other than first metacarpal
C0272686|T037|IS|54641008|SNOMEDCT_CORE|Closed fracture of base of other metacarpal bone|Closed fracture of base of metacarpal bone other than first metacarpal
C0272687|T037|PT|46422008|SNOMEDCT_CORE|Closed fracture of shaft of metacarpal bone|Closed fracture of shaft of metacarpal bone
C0272687|T037|FN|46422008|SNOMEDCT_CORE|Closed fracture of shaft of metacarpal bone|Closed fracture of shaft of metacarpal bone
C0272688|T037|PT|7551007|SNOMEDCT_CORE|Closed fracture of neck of metacarpal bone|Closed fracture of neck of metacarpal bone
C0272688|T037|FN|7551007|SNOMEDCT_CORE|Closed fracture of neck of metacarpal bone|Closed fracture of neck of metacarpal bone
C0272694|T037|PT|405817008|SNOMEDCT_CORE|Fracture of phalanx of hand|Fracture of phalanx of hand
C0272694|T037|FN|405817008|SNOMEDCT_CORE|Fracture of phalanx of hand|Fracture of phalanx of hand
C0272696|T037|PT|36778005|SNOMEDCT_CORE|Fracture of distal phalanx of finger|Fracture of distal phalanx of finger
C0272696|T037|FN|36778005|SNOMEDCT_CORE|Fracture of distal phalanx of finger|Fracture of distal phalanx of finger
C0272698|T037|SY|24424003|SNOMEDCT_CORE|Closed fracture of finger|Closed fracture of phalanx of finger
C0272698|T037|IS|24424003|SNOMEDCT_CORE|Closed fracture of finger, NOS|Closed fracture of phalanx of finger
C0272698|T037|PT|24424003|SNOMEDCT_CORE|Closed fracture of phalanx of finger|Closed fracture of phalanx of finger
C0272698|T037|FN|24424003|SNOMEDCT_CORE|Closed fracture of phalanx of finger|Closed fracture of phalanx of finger
C0272698|T037|IS|24424003|SNOMEDCT_CORE|Closed fracture of phalanx of finger, NOS|Closed fracture of phalanx of finger
C0272699|T037|OAP|22713002|SNOMEDCT_CORE|Closed fracture of middle AND/OR proximal phalanx of finger|Closed fracture of middle AND/OR proximal phalanx of finger
C0272699|T037|OAF|22713002|SNOMEDCT_CORE|Closed fracture of middle AND/OR proximal phalanx of finger|Closed fracture of middle AND/OR proximal phalanx of finger
C0272699|T037|IS|22713002|SNOMEDCT_CORE|Closed fracture of middle or proximal phalanx of finger|Closed fracture of middle AND/OR proximal phalanx of finger
C0272700|T037|SY|76865005|SNOMEDCT_CORE|Closed fracture finger distal phalanx|Closed fracture of distal phalanx of finger
C0272700|T037|PT|76865005|SNOMEDCT_CORE|Closed fracture of distal phalanx of finger|Closed fracture of distal phalanx of finger
C0272700|T037|FN|76865005|SNOMEDCT_CORE|Closed fracture of distal phalanx of finger|Closed fracture of distal phalanx of finger
C0272701|T037|PT|68360003|SNOMEDCT_CORE|Closed fracture of multiple sites of phalanges of hand|Closed fracture of multiple sites of phalanges of hand
C0272701|T037|FN|68360003|SNOMEDCT_CORE|Closed fracture of multiple sites of phalanges of hand|Closed fracture of multiple sites of phalanges of hand
C0272702|T037|SY|21698002|SNOMEDCT_CORE|Open fracture of finger|Open fracture of phalanx of finger
C0272702|T037|IS|21698002|SNOMEDCT_CORE|Open fracture of finger, NOS|Open fracture of phalanx of finger
C0272702|T037|PT|21698002|SNOMEDCT_CORE|Open fracture of phalanx of finger|Open fracture of phalanx of finger
C0272702|T037|FN|21698002|SNOMEDCT_CORE|Open fracture of phalanx of finger|Open fracture of phalanx of finger
C0272702|T037|IS|21698002|SNOMEDCT_CORE|Open fracture of phalanx of finger, NOS|Open fracture of phalanx of finger
C0272709|T037|PT|32805004|SNOMEDCT_CORE|Fractures of multiple bones of lower limb|Fractures of multiple bones of lower limb
C0272709|T037|FN|32805004|SNOMEDCT_CORE|Fractures of multiple bones of lower limb|Fractures of multiple bones of lower limb
C0272709|T037|IS|32805004|SNOMEDCT_CORE|Fractures of multiple bones of lower limb, NOS|Fractures of multiple bones of lower limb
C0272729|T037|PT|25415003|SNOMEDCT_CORE|Closed fracture of femur|Closed fracture of femur
C0272729|T037|FN|25415003|SNOMEDCT_CORE|Closed fracture of femur|Closed fracture of femur
C0272729|T037|IS|25415003|SNOMEDCT_CORE|Closed fracture of femur, NOS|Closed fracture of femur
C0272729|T037|SY|25415003|SNOMEDCT_CORE|Closed fracture of thigh|Closed fracture of femur
C0272729|T037|SY|25415003|SNOMEDCT_CORE|Closed fracture of upper leg|Closed fracture of femur
C0272731|T037|PT|79484004|SNOMEDCT_CORE|Closed transcervical fracture of femur|Closed transcervical fracture of femur
C0272731|T037|FN|79484004|SNOMEDCT_CORE|Closed transcervical fracture of femur|Closed transcervical fracture of femur
C0272731|T037|IS|79484004|SNOMEDCT_CORE|Closed transcervical fracture of femur, NOS|Closed transcervical fracture of femur
C0272732|T037|PT|20100009|SNOMEDCT_CORE|Closed fracture of intracapsular section of femur|Closed fracture of intracapsular section of femur
C0272732|T037|FN|20100009|SNOMEDCT_CORE|Closed fracture of intracapsular section of femur|Closed fracture of intracapsular section of femur
C0272732|T037|IS|20100009|SNOMEDCT_CORE|Closed fracture of intracapsular section of femur, NOS|Closed fracture of intracapsular section of femur
C0272744|T037|PT|89820008|SNOMEDCT_CORE|Closed intertrochanteric fracture|Closed intertrochanteric fracture
C0272744|T037|FN|89820008|SNOMEDCT_CORE|Closed intertrochanteric fracture|Closed intertrochanteric fracture
C0272751|T037|PT|359820003|SNOMEDCT_CORE|Closed fracture of neck of femur|Closed fracture of neck of femur
C0272751|T037|FN|359820003|SNOMEDCT_CORE|Closed fracture of neck of femur|Closed fracture of neck of femur
C0272753|T037|PT|54441004|SNOMEDCT_CORE|Fracture of shaft of femur|Fracture of shaft of femur
C0272753|T037|FN|54441004|SNOMEDCT_CORE|Fracture of shaft of femur|Fracture of shaft of femur
C0272754|T037|PT|66926007|SNOMEDCT_CORE|Closed fracture of femoral condyle of femur|Closed fracture of femoral condyle of femur
C0272754|T037|FN|66926007|SNOMEDCT_CORE|Closed fracture of femoral condyle of femur|Closed fracture of femoral condyle of femur
C0272759|T037|PT|413877007|SNOMEDCT_CORE|Closed fracture of tibia AND fibula|Closed fracture of tibia AND fibula
C0272759|T037|FN|413877007|SNOMEDCT_CORE|Closed fracture of tibia AND fibula|Closed fracture of tibia AND fibula
C0272760|T037|PT|414943006|SNOMEDCT_CORE|Open fracture of tibia AND fibula|Open fracture of tibia AND fibula
C0272760|T037|FN|414943006|SNOMEDCT_CORE|Open fracture of tibia AND fibula|Open fracture of tibia AND fibula
C0272767|T037|PT|6990005|SNOMEDCT_CORE|Fracture of shaft of tibia|Fracture of shaft of tibia
C0272767|T037|FN|6990005|SNOMEDCT_CORE|Fracture of shaft of tibia|Fracture of shaft of tibia
C0272769|T037|PT|42188001|SNOMEDCT_CORE|Closed fracture of ankle|Closed fracture of ankle
C0272769|T037|FN|42188001|SNOMEDCT_CORE|Closed fracture of ankle|Closed fracture of ankle
C0272773|T037|SY|263244000|SNOMEDCT_CORE|Pott's fracture of ankle|Pott's fracture of ankle
C0272774|T037|PT|15574005|SNOMEDCT_CORE|Fracture of foot|Fracture of foot
C0272774|T037|FN|15574005|SNOMEDCT_CORE|Fracture of foot|Fracture of foot
C0272774|T037|IS|15574005|SNOMEDCT_CORE|Fracture of foot, NOS|Fracture of foot
C0272775|T037|PT|342070009|SNOMEDCT_CORE|Closed fracture of foot|Closed fracture of foot
C0272775|T037|FN|342070009|SNOMEDCT_CORE|Closed fracture of foot|Closed fracture of foot
C0272790|T037|PT|70204006|SNOMEDCT_CORE|Closed fracture of fifth metatarsal bone|Closed fracture of fifth metatarsal bone
C0272790|T037|FN|70204006|SNOMEDCT_CORE|Closed fracture of fifth metatarsal bone|Closed fracture of fifth metatarsal bone
C0272839|T037|SY|19494006|SNOMEDCT_CORE|Current tear of meniscus of knee|Current tear of semilunar cartilage
C0272839|T037|IS|19494006|SNOMEDCT_CORE|Current tear of meniscus of knee, NOS|Current tear of semilunar cartilage
C0272839|T037|PT|19494006|SNOMEDCT_CORE|Current tear of semilunar cartilage|Current tear of semilunar cartilage
C0272839|T037|FN|19494006|SNOMEDCT_CORE|Current tear of semilunar cartilage|Current tear of semilunar cartilage
C0272839|T037|IS|19494006|SNOMEDCT_CORE|Current tear of semilunar cartilage, NOS|Current tear of semilunar cartilage
C0272839|T037|SY|19494006|SNOMEDCT_CORE|Tear of meniscus of knee joint|Current tear of semilunar cartilage
C0272839|T037|IS|19494006|SNOMEDCT_CORE|Tear of meniscus of knee joint, NOS|Current tear of semilunar cartilage
C0272869|T037|PT|3199001|SNOMEDCT_CORE|Sprain of shoulder|Sprain of shoulder
C0272869|T037|FN|3199001|SNOMEDCT_CORE|Sprain of shoulder|Sprain of shoulder
C0272869|T037|SY|3199001|SNOMEDCT_CORE|Sprain of shoulder joint|Sprain of shoulder
C0272869|T037|IS|3199001|SNOMEDCT_CORE|Sprain of shoulder, NOS|Sprain of shoulder
C0272876|T037|OAP|47874006|SNOMEDCT_CORE|Sprain of arm|Sprain of arm
C0272876|T037|OAF|47874006|SNOMEDCT_CORE|Sprain of arm|Sprain of arm
C0272876|T037|IS|47874006|SNOMEDCT_CORE|Sprain of arm, NOS|Sprain of arm, NOS
C0272889|T037|SY|17883008|SNOMEDCT_CORE|Hip sprain|Sprain of hip
C0272889|T037|PT|17883008|SNOMEDCT_CORE|Sprain of hip|Sprain of hip
C0272889|T037|FN|17883008|SNOMEDCT_CORE|Sprain of hip|Sprain of hip
C0272889|T037|SY|17883008|SNOMEDCT_CORE|Sprain of hip joint|Sprain of hip
C0272889|T037|IS|17883008|SNOMEDCT_CORE|Sprain of hip, NOS|Sprain of hip
C0272890|T037|SY|17883008|SNOMEDCT_CORE|Thigh sprain|Thigh sprain
C0272891|T037|SY|54888009|SNOMEDCT_CORE|Knee sprain|Sprain of knee
C0272891|T037|PT|54888009|SNOMEDCT_CORE|Sprain of knee|Sprain of knee
C0272891|T037|FN|54888009|SNOMEDCT_CORE|Sprain of knee|Sprain of knee
C0272891|T037|SY|54888009|SNOMEDCT_CORE|Sprain of knee joint|Sprain of knee
C0272891|T037|IS|54888009|SNOMEDCT_CORE|Sprain of knee, NOS|Sprain of knee
C0272891|T037|SY|54888009|SNOMEDCT_CORE|Sprain of ligament of knee joint|Sprain of knee
C0272893|T037|PT|262994004|SNOMEDCT_CORE|Leg sprain|Leg sprain
C0272893|T037|FN|262994004|SNOMEDCT_CORE|Leg sprain|Leg sprain
C0272910|T037|FN|66540002|SNOMEDCT_CORE|Back strain of thoracic region|Strain of thoracic region
C0272910|T037|SY|66540002|SNOMEDCT_CORE|Back strain of thoracic region|Strain of thoracic region
C0272910|T037|PT|66540002|SNOMEDCT_CORE|Strain of thoracic region|Strain of thoracic region
C0272910|T037|IS|66540002|SNOMEDCT_CORE|Strain of thoracic region, NOS|Strain of thoracic region
C0272914|T037|SY|209548004|SNOMEDCT_CORE|Lumbosacral sprain|Sprain of ligament of lumbosacral joint
C0272914|T037|OAP|40129004|SNOMEDCT_CORE|Sprain of ligament of lumbosacral joint|Sprain of ligament of lumbosacral joint
C0272914|T037|PT|209548004|SNOMEDCT_CORE|Sprain of ligament of lumbosacral joint|Sprain of ligament of lumbosacral joint
C0272914|T037|OAF|40129004|SNOMEDCT_CORE|Sprain of ligament of lumbosacral joint|Sprain of ligament of lumbosacral joint
C0272914|T037|FN|209548004|SNOMEDCT_CORE|Sprain of ligament of lumbosacral joint|Sprain of ligament of lumbosacral joint
C0272914|T037|OAS|40129004|SNOMEDCT_CORE|Sprain of lumbosacral joint AND/OR ligament|Sprain of ligament of lumbosacral joint
C0272914|T037|IS|40129004|SNOMEDCT_CORE|Sprain of lumbosacral joint or ligament|Sprain of ligament of lumbosacral joint
C0272914|T037|SY|209548004|SNOMEDCT_CORE|Sprain, lumbosacral ligament|Sprain of ligament of lumbosacral joint
C0272914|T037|OF|209548004|SNOMEDCT_CORE|Sprain, lumbosacral ligament|Sprain of ligament of lumbosacral joint
C0272925|T037|IS|54355006|SNOMEDCT_CORE|Head injury, NOS, without skull fracture|Intracranial injury, without skull fracture
C0272925|T037|SY|54355006|SNOMEDCT_CORE|Head injury, without skull fracture|Intracranial injury, without skull fracture
C0272925|T037|IS|54355006|SNOMEDCT_CORE|Intracranial injury, NOS, without skull fracture|Intracranial injury, without skull fracture
C0272925|T037|PT|54355006|SNOMEDCT_CORE|Intracranial injury, without skull fracture|Intracranial injury, without skull fracture
C0272925|T037|FN|54355006|SNOMEDCT_CORE|Intracranial injury, without skull fracture|Intracranial injury, without skull fracture
C0272927|T037|PT|9015001|SNOMEDCT_CORE|Brain injury without open intracranial wound|Brain injury without open intracranial wound
C0272927|T037|FN|9015001|SNOMEDCT_CORE|Brain injury without open intracranial wound|Brain injury without open intracranial wound
C0272927|T037|IS|9015001|SNOMEDCT_CORE|Brain injury without open intracranial wound, NOS|Brain injury without open intracranial wound
C0272927|T037|SY|9015001|SNOMEDCT_CORE|Closed traumatic brain injury|Brain injury without open intracranial wound
C0272936|T037|PT|28188001|SNOMEDCT_CORE|Brain injury with open intracranial wound|Brain injury with open intracranial wound
C0272936|T037|FN|28188001|SNOMEDCT_CORE|Brain injury with open intracranial wound|Brain injury with open intracranial wound
C0272936|T037|IS|28188001|SNOMEDCT_CORE|Brain injury with open intracranial wound, NOS|Brain injury with open intracranial wound
C0272950|T037|PT|23713006|SNOMEDCT_CORE|Contusion of cerebral cortex|Contusion of cerebral cortex
C0272950|T037|FN|23713006|SNOMEDCT_CORE|Contusion of cerebral cortex|Contusion of cerebral cortex
C0272950|T037|IS|23713006|SNOMEDCT_CORE|Contusion of cerebral cortex, NOS|Contusion of cerebral cortex
C0272950|T037|SY|23713006|SNOMEDCT_CORE|Cortex contusion|Contusion of cerebral cortex
C0273287|T037|PT|58411009|SNOMEDCT_CORE|Broken tooth with complication|Broken tooth with complication
C0273287|T037|FN|58411009|SNOMEDCT_CORE|Broken tooth with complication|Broken tooth with complication
C0273333|T037|PT|16809003|SNOMEDCT_CORE|Open wound of abdominal wall with complication|Open wound of abdominal wall with complication
C0273333|T037|FN|16809003|SNOMEDCT_CORE|Open wound of abdominal wall with complication|Open wound of abdominal wall with complication
C0273333|T037|IS|16809003|SNOMEDCT_CORE|Open wound of abdominal wall with complication, NOS|Open wound of abdominal wall with complication
C0273402|T037|PT|32976001|SNOMEDCT_CORE|Open wound of leg with complication|Open wound of leg with complication
C0273402|T037|FN|32976001|SNOMEDCT_CORE|Open wound of leg with complication|Open wound of leg with complication
C0273444|T037|SY|50793006|SNOMEDCT_CORE|Crush injury of hand|Crushing injury of hand
C0273444|T037|SY|50793006|SNOMEDCT_CORE|Crush injury to hand|Crushing injury of hand
C0273444|T037|PT|50793006|SNOMEDCT_CORE|Crushing injury of hand|Crushing injury of hand
C0273444|T037|FN|50793006|SNOMEDCT_CORE|Crushing injury of hand|Crushing injury of hand
C0273445|T037|SY|10380004|SNOMEDCT_CORE|Crush injury of finger|Crushing injury of finger
C0273445|T037|SY|10380004|SNOMEDCT_CORE|Crush injury to finger|Crushing injury of finger
C0273445|T037|PT|10380004|SNOMEDCT_CORE|Crushing injury of finger|Crushing injury of finger
C0273445|T037|FN|10380004|SNOMEDCT_CORE|Crushing injury of finger|Crushing injury of finger
C0273448|T037|SY|74682007|SNOMEDCT_CORE|Crush injury of toe|Crushing injury of toe
C0273448|T037|OAP|211609000|SNOMEDCT_CORE|Crush injury, toe|Crushing injury of toe
C0273448|T037|OAF|211609000|SNOMEDCT_CORE|Crush injury, toe|Crushing injury of toe
C0273448|T037|PT|74682007|SNOMEDCT_CORE|Crushing injury of toe|Crushing injury of toe
C0273448|T037|FN|74682007|SNOMEDCT_CORE|Crushing injury of toe|Crushing injury of toe
C0273529|T037|OAP|212361009|SNOMEDCT_CORE|Injury of nerves at shoulder and upper arm level|Injury of nerves at shoulder and upper arm level
C0273529|T037|OAF|212361009|SNOMEDCT_CORE|Injury of nerves at shoulder and upper arm level|Injury of nerves at shoulder and upper arm level
C0273530|T037|SY|4412009|SNOMEDCT_CORE|Digital nerve injury|Injury of digital nerve
C0273530|T037|PT|4412009|SNOMEDCT_CORE|Injury of digital nerve|Injury of digital nerve
C0273530|T037|FN|4412009|SNOMEDCT_CORE|Injury of digital nerve|Injury of digital nerve
C0273940|T037|IS|17771000|SNOMEDCT_CORE|Burn of face and head, NOS|Burn of face AND/OR head
C0273940|T037|OAF|17771000|SNOMEDCT_CORE|Burn of face AND/OR head|Burn of face AND/OR head
C0273940|T037|OAP|17771000|SNOMEDCT_CORE|Burn of face AND/OR head|Burn of face AND/OR head
C0273982|T037|PT|60713008|SNOMEDCT_CORE|Burn of neck|Burn of neck
C0273982|T037|FN|60713008|SNOMEDCT_CORE|Burn of neck|Burn of neck
C0273982|T037|IS|60713008|SNOMEDCT_CORE|Burn of neck, NOS|Burn of neck
C0274035|T037|PT|6055000|SNOMEDCT_CORE|Burn of upper limb|Burn of upper limb
C0274035|T037|FN|6055000|SNOMEDCT_CORE|Burn of upper limb|Burn of upper limb
C0274035|T037|IS|6055000|SNOMEDCT_CORE|Burn of upper limb, NOS|Burn of upper limb
C0274089|T037|PT|14893008|SNOMEDCT_CORE|Burn of hand|Burn of hand
C0274089|T037|FN|14893008|SNOMEDCT_CORE|Burn of hand|Burn of hand
C0274089|T037|IS|14893008|SNOMEDCT_CORE|Burn of hand, NOS|Burn of hand
C0274091|T037|PT|54296007|SNOMEDCT_CORE|Partial thickness burn of hand|Partial thickness burn of hand
C0274091|T037|FN|54296007|SNOMEDCT_CORE|Partial thickness burn of hand|Partial thickness burn of hand
C0274091|T037|SY|54296007|SNOMEDCT_CORE|Second degree burn of hand|Partial thickness burn of hand
C0274091|T037|OF|54296007|SNOMEDCT_CORE|Second degree burn of hand|Partial thickness burn of hand
C0274137|T037|PT|84677008|SNOMEDCT_CORE|Burn of lower limb|Burn of lower limb
C0274137|T037|FN|84677008|SNOMEDCT_CORE|Burn of lower limb|Burn of lower limb
C0274137|T037|IS|84677008|SNOMEDCT_CORE|Burn of lower limb, NOS|Burn of lower limb
C0274137|T037|SY|84677008|SNOMEDCT_CORE|Leg - burn|Burn of lower limb
C0274137|T037|SY|84677008|SNOMEDCT_CORE|Leg burns|Burn of lower limb
C0274167|T037|PT|11980003|SNOMEDCT_CORE|Burn of foot|Burn of foot
C0274167|T037|FN|11980003|SNOMEDCT_CORE|Burn of foot|Burn of foot
C0274167|T037|IS|11980003|SNOMEDCT_CORE|Burn of foot, NOS|Burn of foot
C0274210|T037|PT|60897004|SNOMEDCT_CORE|Contusion of nose|Contusion of nose
C0274210|T037|FN|60897004|SNOMEDCT_CORE|Contusion of nose|Contusion of nose
C0274210|T037|SY|60897004|SNOMEDCT_CORE|Contusion, nose|Contusion of nose
C0274210|T037|SY|60897004|SNOMEDCT_CORE|Nose - bruise|Contusion of nose
C0274220|T037|PT|68893001|SNOMEDCT_CORE|Contusion of buttock|Contusion of buttock
C0274220|T037|FN|68893001|SNOMEDCT_CORE|Contusion of buttock|Contusion of buttock
C0274236|T037|SY|91603007|SNOMEDCT_CORE|Contusion of leg|Contusion of lower limb
C0274236|T037|IS|91603007|SNOMEDCT_CORE|Contusion of leg, NOS|Contusion of lower limb
C0274236|T037|PT|91603007|SNOMEDCT_CORE|Contusion of lower limb|Contusion of lower limb
C0274236|T037|FN|91603007|SNOMEDCT_CORE|Contusion of lower limb|Contusion of lower limb
C0274236|T037|IS|91603007|SNOMEDCT_CORE|Contusion of lower limb, NOS|Contusion of lower limb
C0274278|T037|PT|74472004|SNOMEDCT_CORE|Late effect of intracranial injury without skull fracture|Late effect of intracranial injury without skull fracture
C0274278|T037|FN|74472004|SNOMEDCT_CORE|Late effect of intracranial injury without skull fracture|Late effect of intracranial injury without skull fracture
C0274278|T037|IS|74472004|SNOMEDCT_CORE|Sequelae of intracranial injury|Late effect of intracranial injury without skull fracture
C0274301|T047|SY|45376003|SNOMEDCT_CORE|Adverse effect, caused by correct medicinal substance properly administered|Adverse effect, due to correct medicinal substance properly administered
C0274301|T047|FN|45376003|SNOMEDCT_CORE|Adverse effect, caused by correct medicinal substance properly administered|Adverse effect, due to correct medicinal substance properly administered
C0274301|T047|PT|45376003|SNOMEDCT_CORE|Adverse effect, due to correct medicinal substance properly administered|Adverse effect, due to correct medicinal substance properly administered
C0274301|T047|OF|45376003|SNOMEDCT_CORE|Adverse effect, due to correct medicinal substance properly administered|Adverse effect, due to correct medicinal substance properly administered
C0274301|T047|IS|45376003|SNOMEDCT_CORE|Adverse effect, NOS, due to correct medicinal substance properly administered|Adverse effect, due to correct medicinal substance properly administered
C0274311|T046|PT|88797001|SNOMEDCT_CORE|Complication of surgical procedure|Complication of surgical procedure
C0274311|T046|FN|88797001|SNOMEDCT_CORE|Complication of surgical procedure|Complication of surgical procedure
C0274311|T046|IS|88797001|SNOMEDCT_CORE|Complication of surgical procedure, NOS|Complication of surgical procedure
C0274311|T046|SY|88797001|SNOMEDCT_CORE|Misadventure of surgical procedure|Complication of surgical procedure
C0274311|T046|IS|88797001|SNOMEDCT_CORE|Misadventure of surgical procedure, NOS|Complication of surgical procedure
C0274348|T033|PTGB|111744007|SNOMEDCT_CORE|Mechanical complication of internal orthopaedic device|Mechanical complication of internal orthopedic device
C0274348|T033|PT|111744007|SNOMEDCT_CORE|Mechanical complication of internal orthopedic device|Mechanical complication of internal orthopedic device
C0274348|T033|FN|111744007|SNOMEDCT_CORE|Mechanical complication of internal orthopedic device|Mechanical complication of internal orthopedic device
C0274357|T046|SY|45945004|SNOMEDCT_CORE|Mechanical complication due to breast implant|Mechanical complication due to breast prosthesis
C0274357|T046|PT|45945004|SNOMEDCT_CORE|Mechanical complication due to breast prosthesis|Mechanical complication due to breast prosthesis
C0274357|T046|FN|45945004|SNOMEDCT_CORE|Mechanical complication due to breast prosthesis|Mechanical complication due to breast prosthesis
C0274357|T046|IS|45945004|SNOMEDCT_CORE|Mechanical complication due to breast prosthesis, NOS|Mechanical complication due to breast prosthesis
C0274363|T046|SY|31871009|SNOMEDCT_CORE|Infection and inflammation reaction due to internal prosthetic device, implant or graft|Infection AND/OR inflammatory reaction due to internal prosthetic device, implant AND/OR graft
C0274363|T046|PT|31871009|SNOMEDCT_CORE|Infection AND/OR inflammatory reaction due to internal prosthetic device, implant AND/OR graft|Infection AND/OR inflammatory reaction due to internal prosthetic device, implant AND/OR graft
C0274363|T046|FN|31871009|SNOMEDCT_CORE|Infection AND/OR inflammatory reaction due to internal prosthetic device, implant AND/OR graft|Infection AND/OR inflammatory reaction due to internal prosthetic device, implant AND/OR graft
C0274363|T046|IS|31871009|SNOMEDCT_CORE|Infection or inflammatory reaction due to internal prosthetic device, implant or graft, NOS|Infection AND/OR inflammatory reaction due to internal prosthetic device, implant AND/OR graft
C0274369|T184|OAP|79608006|SNOMEDCT_CORE|Pain due to any device, implant AND/OR graft|Pain due to any device, implant AND/OR graft
C0274369|T184|OAF|79608006|SNOMEDCT_CORE|Pain due to any device, implant AND/OR graft|Pain due to any device, implant AND/OR graft
C0274369|T184|IS|79608006|SNOMEDCT_CORE|Pain due to any device, implant or graft|Pain due to any device, implant AND/OR graft
C0274419|T046|PT|33603003|SNOMEDCT_CORE|Complication of renal dialysis|Complication of renal dialysis
C0274419|T046|FN|33603003|SNOMEDCT_CORE|Complication of renal dialysis|Complication of renal dialysis
C0274610|T037|PT|11196001|SNOMEDCT_CORE|Poisoning by opiate AND/OR related narcotic|Poisoning by opiate AND/OR related narcotic
C0274610|T037|OF|11196001|SNOMEDCT_CORE|Poisoning by opiate AND/OR related narcotic|Poisoning by opiate AND/OR related narcotic
C0274610|T037|FN|11196001|SNOMEDCT_CORE|Poisoning caused by opiate AND/OR related narcotic|Poisoning by opiate AND/OR related narcotic
C0274610|T037|SY|11196001|SNOMEDCT_CORE|Poisoning caused by opiate AND/OR related narcotic|Poisoning by opiate AND/OR related narcotic
C0274638|T037|PT|85337000|SNOMEDCT_CORE|Poisoning by sedative AND/OR hypnotic|Poisoning by sedative AND/OR hypnotic
C0274638|T037|OF|85337000|SNOMEDCT_CORE|Poisoning by sedative AND/OR hypnotic|Poisoning by sedative AND/OR hypnotic
C0274638|T037|IS|85337000|SNOMEDCT_CORE|Poisoning by sedative or hypnotic, NOS|Poisoning by sedative AND/OR hypnotic
C0274638|T037|SY|85337000|SNOMEDCT_CORE|Poisoning by sleeping drug|Poisoning by sedative AND/OR hypnotic
C0274638|T037|IS|85337000|SNOMEDCT_CORE|Poisoning by sleeping drug, NOS|Poisoning by sedative AND/OR hypnotic
C0274638|T037|SY|85337000|SNOMEDCT_CORE|Poisoning by sleeping pill|Poisoning by sedative AND/OR hypnotic
C0274638|T037|IS|85337000|SNOMEDCT_CORE|Poisoning by sleeping pill, NOS|Poisoning by sedative AND/OR hypnotic
C0274638|T037|SY|85337000|SNOMEDCT_CORE|Poisoning by sleeping tablet|Poisoning by sedative AND/OR hypnotic
C0274638|T037|IS|85337000|SNOMEDCT_CORE|Poisoning by sleeping tablet, NOS|Poisoning by sedative AND/OR hypnotic
C0274638|T037|FN|85337000|SNOMEDCT_CORE|Poisoning caused by sedative AND/OR hypnotic|Poisoning by sedative AND/OR hypnotic
C0274638|T037|SY|85337000|SNOMEDCT_CORE|Poisoning caused by sedative AND/OR hypnotic|Poisoning by sedative AND/OR hypnotic
C0274638|T037|SY|85337000|SNOMEDCT_CORE|Poisoning caused by sleeping drug|Poisoning by sedative AND/OR hypnotic
C0274638|T037|SY|85337000|SNOMEDCT_CORE|Poisoning caused by sleeping pill|Poisoning by sedative AND/OR hypnotic
C0274638|T037|SY|85337000|SNOMEDCT_CORE|Poisoning caused by sleeping tablet|Poisoning by sedative AND/OR hypnotic
C0274797|T037|PT|36265009|SNOMEDCT_CORE|Poisoning by local anti-inflammatory drug|Poisoning by local anti-inflammatory drug
C0274797|T037|OF|36265009|SNOMEDCT_CORE|Poisoning by local anti-inflammatory drug|Poisoning by local anti-inflammatory drug
C0274797|T037|IS|36265009|SNOMEDCT_CORE|Poisoning by local anti-inflammatory drug, NOS|Poisoning by local anti-inflammatory drug
C0274797|T037|FN|36265009|SNOMEDCT_CORE|Poisoning caused by local anti-inflammatory drug|Poisoning by local anti-inflammatory drug
C0274797|T037|SY|36265009|SNOMEDCT_CORE|Poisoning caused by local anti-inflammatory drug|Poisoning by local anti-inflammatory drug
C0274817|T037|IS|7895008|SNOMEDCT_CORE|Poisoning by drug or medicinal substance, NEC|Poisoning by drug or medicinal substance, NEC
C0274979|T037|SY|25440005|SNOMEDCT_CORE|Dioxin poisoning|Tetrachlorodibenzodioxin poisoning
C0274979|T037|SY|25440005|SNOMEDCT_CORE|TCDD poisoning|Tetrachlorodibenzodioxin poisoning
C0274979|T037|PT|25440005|SNOMEDCT_CORE|Tetrachlorodibenzodioxin poisoning|Tetrachlorodibenzodioxin poisoning
C0274979|T037|FN|25440005|SNOMEDCT_CORE|Tetrachlorodibenzodioxin poisoning|Tetrachlorodibenzodioxin poisoning
C0275120|T037|PT|7456000|SNOMEDCT_CORE|Poisoning by wasp sting|Poisoning by wasp sting
C0275120|T037|OF|7456000|SNOMEDCT_CORE|Poisoning by wasp sting|Poisoning by wasp sting
C0275120|T037|IS|7456000|SNOMEDCT_CORE|Poisoning by wasp sting, NOS|Poisoning by wasp sting
C0275120|T037|SY|7456000|SNOMEDCT_CORE|Poisoning caused by wasp sting|Poisoning by wasp sting
C0275120|T037|FN|7456000|SNOMEDCT_CORE|Poisoning caused by wasp sting|Poisoning by wasp sting
C0275120|T037|SY|7456000|SNOMEDCT_CORE|Toxic reaction caused by wasp sting|Poisoning by wasp sting
C0275551|T047|PT|11836002|SNOMEDCT_CORE|Primary bacterial peritonitis|Primary bacterial peritonitis
C0275551|T047|FN|11836002|SNOMEDCT_CORE|Primary bacterial peritonitis|Primary bacterial peritonitis
C0275551|T047|SY|11836002|SNOMEDCT_CORE|SBP - Spontaneous bacterial peritonitis|Primary bacterial peritonitis
C0275551|T047|SY|11836002|SNOMEDCT_CORE|Spontaneous bacterial peritonitis|Primary bacterial peritonitis
C0275804|T047|PT|41582007|SNOMEDCT_CORE|Streptococcal tonsillitis|Streptococcal tonsillitis
C0275804|T047|FN|41582007|SNOMEDCT_CORE|Streptococcal tonsillitis|Streptococcal tonsillitis
C0275858|T047|PT|67125004|SNOMEDCT_CORE|Latent syphilis with positive serology|Latent syphilis with positive serology
C0275858|T047|FN|67125004|SNOMEDCT_CORE|Latent syphilis with positive serology|Latent syphilis with positive serology
C0275982|T047|SY|18081009|SNOMEDCT_CORE|Campylobacter diarrhea|Enteric campylobacteriosis
C0275982|T047|SYGB|18081009|SNOMEDCT_CORE|Campylobacter diarrhoea|Enteric campylobacteriosis
C0275982|T047|SY|18081009|SNOMEDCT_CORE|Campylobacter intestinal infection|Enteric campylobacteriosis
C0275982|T047|PT|18081009|SNOMEDCT_CORE|Enteric campylobacteriosis|Enteric campylobacteriosis
C0275982|T047|FN|18081009|SNOMEDCT_CORE|Enteric campylobacteriosis|Enteric campylobacteriosis
C0276026|T047|PT|70036007|SNOMEDCT_CORE|Haemophilus influenzae pneumonia|Haemophilus influenzae pneumonia
C0276026|T047|FN|70036007|SNOMEDCT_CORE|Haemophilus influenzae pneumonia|Haemophilus influenzae pneumonia
C0276026|T047|IS|70036007|SNOMEDCT_CORE|Hemophilus influenzae pneumonia|Haemophilus influenzae pneumonia
C0276088|T047|OAS|9323009|SNOMEDCT_CORE|E. coli septicaemia|Escherichia coli septicemia
C0276088|T047|OAS|9323009|SNOMEDCT_CORE|E. coli septicemia|Escherichia coli septicemia
C0276088|T047|OAS|9323009|SNOMEDCT_CORE|Escherichia coli septicaemia|Escherichia coli septicemia
C0276088|T047|OAS|9323009|SNOMEDCT_CORE|Escherichia coli septicemia|Escherichia coli septicemia
C0276088|T047|OAP|9323009|SNOMEDCT_CORE|Septicaemia due to E. Coli|Escherichia coli septicemia
C0276088|T047|OAS|9323009|SNOMEDCT_CORE|Septicaemia due to Escherichia coli|Escherichia coli septicemia
C0276088|T047|OAS|9323009|SNOMEDCT_CORE|Septicaemic colibacillosis|Escherichia coli septicemia
C0276088|T047|OAP|9323009|SNOMEDCT_CORE|Septicemia due to E. Coli|Escherichia coli septicemia
C0276088|T047|OF|9323009|SNOMEDCT_CORE|Septicemia due to E. Coli|Escherichia coli septicemia
C0276088|T047|OAS|9323009|SNOMEDCT_CORE|Septicemia due to Escherichia coli|Escherichia coli septicemia
C0276088|T047|OAF|9323009|SNOMEDCT_CORE|Septicemia due to Escherichia coli|Escherichia coli septicemia
C0276088|T047|OAS|9323009|SNOMEDCT_CORE|Septicemic colibacillosis|Escherichia coli septicemia
C0276089|T047|SY|51530003|SNOMEDCT_CORE|Escherichia coli pneumonia|Pneumonia due to Escherichia coli
C0276089|T047|SY|51530003|SNOMEDCT_CORE|Pneumonia caused by E. coli|Pneumonia due to Escherichia coli
C0276089|T047|FN|51530003|SNOMEDCT_CORE|Pneumonia caused by Escherichia coli|Pneumonia due to Escherichia coli
C0276089|T047|SY|51530003|SNOMEDCT_CORE|Pneumonia caused by Escherichia coli|Pneumonia due to Escherichia coli
C0276089|T047|SY|51530003|SNOMEDCT_CORE|Pneumonia due to E. coli|Pneumonia due to Escherichia coli
C0276089|T047|PT|51530003|SNOMEDCT_CORE|Pneumonia due to Escherichia coli|Pneumonia due to Escherichia coli
C0276089|T047|OF|51530003|SNOMEDCT_CORE|Pneumonia due to Escherichia coli|Pneumonia due to Escherichia coli
C0276141|T047|PT|16146001|SNOMEDCT_CORE|Viral bronchitis|Viral bronchitis
C0276141|T047|FN|16146001|SNOMEDCT_CORE|Viral bronchitis|Viral bronchitis
C0276141|T047|IS|16146001|SNOMEDCT_CORE|Viral bronchitis, NOS|Viral bronchitis
C0276143|T047|PT|1532007|SNOMEDCT_CORE|Viral pharyngitis|Viral pharyngitis
C0276143|T047|FN|1532007|SNOMEDCT_CORE|Viral pharyngitis|Viral pharyngitis
C0276143|T047|IS|1532007|SNOMEDCT_CORE|Viral pharyngitis, NOS|Viral pharyngitis
C0276156|T047|PT|41207000|SNOMEDCT_CORE|Adenoviral pneumonia|Adenoviral pneumonia
C0276156|T047|FN|41207000|SNOMEDCT_CORE|Adenoviral pneumonia|Adenoviral pneumonia
C0276223|T047|PT|37323009|SNOMEDCT_CORE|Recurrent herpes simplex|Recurrent herpes simplex
C0276223|T047|FN|37323009|SNOMEDCT_CORE|Recurrent herpes simplex|Recurrent herpes simplex
C0276262|T020|SY|240539000|SNOMEDCT_CORE|Flat wart|Plane wart
C0276262|T020|PT|240539000|SNOMEDCT_CORE|Plane wart|Plane wart
C0276262|T020|FN|240539000|SNOMEDCT_CORE|Plane wart|Plane wart
C0276262|T020|SY|240539000|SNOMEDCT_CORE|Verruca plana|Plane wart
C0276333|T047|SY|64917006|SNOMEDCT_CORE|Parainfluenza pneumonia|Parainfluenza virus pneumonia
C0276333|T047|PT|64917006|SNOMEDCT_CORE|Parainfluenza virus pneumonia|Parainfluenza virus pneumonia
C0276333|T047|FN|64917006|SNOMEDCT_CORE|Parainfluenza virus pneumonia|Parainfluenza virus pneumonia
C0276333|T047|SY|64917006|SNOMEDCT_CORE|Parainfluenzal pneumonia|Parainfluenza virus pneumonia
C0276333|T047|SY|64917006|SNOMEDCT_CORE|Pneumonia due to parainfluenza virus|Parainfluenza virus pneumonia
C0276351|T047|OAP|78431007|SNOMEDCT_CORE|Influenza due to Influenza virus, type A, human|Influenza due to Influenza virus, type A, human
C0276351|T047|OAF|78431007|SNOMEDCT_CORE|Influenza due to Influenza virus, type A, human|Influenza due to Influenza virus, type A, human
C0276353|T047|FN|24662006|SNOMEDCT_CORE|Influenza caused by Influenza B virus|Influenza due to Influenza B virus
C0276353|T047|SY|24662006|SNOMEDCT_CORE|Influenza caused by Influenza B virus|Influenza due to Influenza B virus
C0276353|T047|OF|24662006|SNOMEDCT_CORE|Influenza caused by Influenza virus, type B|Influenza due to Influenza B virus
C0276353|T047|IS|24662006|SNOMEDCT_CORE|Influenza caused by Influenza virus, type B|Influenza due to Influenza B virus
C0276353|T047|PT|24662006|SNOMEDCT_CORE|Influenza due to Influenza B virus|Influenza due to Influenza B virus
C0276353|T047|OP|24662006|SNOMEDCT_CORE|Influenza due to Influenza virus, type B|Influenza due to Influenza B virus
C0276353|T047|OF|24662006|SNOMEDCT_CORE|Influenza due to Influenza virus, type B|Influenza due to Influenza B virus
C0276535|T191|SY|109385007|SNOMEDCT_CORE|Epidemic Kaposi's sarcoma|Epidemic Kaposi's sarcoma
C0276609|T047|SY|76795007|SNOMEDCT_CORE|Acute hepatitis B|Acute type B viral hepatitis
C0276609|T047|PT|76795007|SNOMEDCT_CORE|Acute type B viral hepatitis|Acute type B viral hepatitis
C0276609|T047|FN|76795007|SNOMEDCT_CORE|Acute type B viral hepatitis|Acute type B viral hepatitis
C0276610|T047|PT|186639003|SNOMEDCT_CORE|Chronic viral hepatitis B without delta-agent|Chronic viral hepatitis B without delta-agent
C0276610|T047|FN|186639003|SNOMEDCT_CORE|Chronic viral hepatitis B without delta-agent|Chronic viral hepatitis B without delta-agent
C0276619|T047|SY|24789006|SNOMEDCT_CORE|Norwalk virus food poisoning|Viral gastroenteritis due to Norwalk-like agent
C0276619|T047|SY|24789006|SNOMEDCT_CORE|Norwalk virus gastroenteritis|Viral gastroenteritis due to Norwalk-like agent
C0276619|T047|SY|24789006|SNOMEDCT_CORE|Norwalk-like virus gastroenteritis|Viral gastroenteritis due to Norwalk-like agent
C0276619|T047|SY|24789006|SNOMEDCT_CORE|Small round structured virus gastroenteritis|Viral gastroenteritis due to Norwalk-like agent
C0276619|T047|FN|24789006|SNOMEDCT_CORE|Viral gastroenteritis caused by Norwalk-like agent|Viral gastroenteritis due to Norwalk-like agent
C0276619|T047|SY|24789006|SNOMEDCT_CORE|Viral gastroenteritis caused by Norwalk-like agent|Viral gastroenteritis due to Norwalk-like agent
C0276619|T047|PT|24789006|SNOMEDCT_CORE|Viral gastroenteritis due to Norwalk-like agent|Viral gastroenteritis due to Norwalk-like agent
C0276619|T047|OP|24789006|SNOMEDCT_CORE|Viral gastroenteritis due to Norwalk-like agents|Viral gastroenteritis due to Norwalk-like agent
C0276619|T047|OF|24789006|SNOMEDCT_CORE|Viral gastroenteritis due to Norwalk-like agents|Viral gastroenteritis due to Norwalk-like agent
C0276682|T047|SY|414821002|SNOMEDCT_CORE|Neonatal candida infection|Neonatal candidiasis
C0276682|T047|PT|414821002|SNOMEDCT_CORE|Neonatal candidiasis|Neonatal candidiasis
C0276682|T047|FN|414821002|SNOMEDCT_CORE|Neonatal candidiasis|Neonatal candidiasis
C0276682|T047|SY|414821002|SNOMEDCT_CORE|Neonatal candidosis|Neonatal candidiasis
C0276682|T047|SY|414821002|SNOMEDCT_CORE|Neonatal thrush|Neonatal candidiasis
C0276683|T047|PT|1085006|SNOMEDCT_CORE|Candidiasis of vulva|Candidiasis of vulva
C0276683|T047|FN|1085006|SNOMEDCT_CORE|Candidiasis of vulva|Candidiasis of vulva
C0276683|T047|SY|1085006|SNOMEDCT_CORE|Vulval candidiasis|Candidiasis of vulva
C0276683|T047|SY|1085006|SNOMEDCT_CORE|Vulval candidosis|Candidiasis of vulva
C0276683|T047|SY|1085006|SNOMEDCT_CORE|Vulval thrush|Candidiasis of vulva
C0277348|T047|SY|74949007|SNOMEDCT_CORE|Anoplurosis|Infestation by Anoplura
C0277348|T047|PT|74949007|SNOMEDCT_CORE|Infestation by Anoplura|Infestation by Anoplura
C0277348|T047|OF|74949007|SNOMEDCT_CORE|Infestation by Anoplura|Infestation by Anoplura
C0277348|T047|IS|74949007|SNOMEDCT_CORE|Infestation by Anoplura, NOS|Infestation by Anoplura
C0277348|T047|SY|74949007|SNOMEDCT_CORE|Infestation by sucking lice|Infestation by Anoplura
C0277348|T047|IS|74949007|SNOMEDCT_CORE|Infestation by sucking lice, NOS|Infestation by Anoplura
C0277348|T047|FN|74949007|SNOMEDCT_CORE|Infestation caused by Anoplura|Infestation by Anoplura
C0277348|T047|SY|74949007|SNOMEDCT_CORE|Infestation caused by Anoplura|Infestation by Anoplura
C0277348|T047|SY|74949007|SNOMEDCT_CORE|Infestation caused by sucking lice|Infestation by Anoplura
C0277525|T047|SY|12463005|SNOMEDCT_CORE|Gastric flu|Infectious gastroenteritis
C0277525|T047|PT|12463005|SNOMEDCT_CORE|Infectious gastroenteritis|Infectious gastroenteritis
C0277525|T047|FN|12463005|SNOMEDCT_CORE|Infectious gastroenteritis|Infectious gastroenteritis
C0277525|T047|IS|12463005|SNOMEDCT_CORE|Infectious gastroenteritis, NOS|Infectious gastroenteritis
C0277525|T047|SY|12463005|SNOMEDCT_CORE|Septic gastroenteritis|Infectious gastroenteritis
C0277525|T047|IS|12463005|SNOMEDCT_CORE|Septic gastroenteritis, NOS|Infectious gastroenteritis
C0277526|T047|PT|46799006|SNOMEDCT_CORE|Dysenteric diarrhea|Dysenteric diarrhea
C0277526|T047|FN|46799006|SNOMEDCT_CORE|Dysenteric diarrhea|Dysenteric diarrhea
C0277526|T047|PTGB|46799006|SNOMEDCT_CORE|Dysenteric diarrhoea|Dysenteric diarrhea
C0277526|T047|SY|46799006|SNOMEDCT_CORE|Dysentery|Dysenteric diarrhea
C0277534|T047|SY|57419008|SNOMEDCT_CORE|Gastroenteritis - presumed infectious origin|Gastroenteritis presumed infectious
C0277534|T047|PT|57419008|SNOMEDCT_CORE|Gastroenteritis presumed infectious|Gastroenteritis presumed infectious
C0277534|T047|FN|57419008|SNOMEDCT_CORE|Gastroenteritis presumed infectious|Gastroenteritis presumed infectious
C0277663|T037|PT|891003|SNOMEDCT_CORE|Suicide by self-administered drug|Suicide by self-administered drug
C0277663|T037|OF|891003|SNOMEDCT_CORE|Suicide by self-administered drug|Suicide by self-administered drug
C0277663|T037|FN|891003|SNOMEDCT_CORE|Suicide by self-administered drug|Suicide by self-administered drug
C0277725|T033|PT|90774003|SNOMEDCT_CORE|Victim of physical assault|Victim of physical assault
C0277725|T033|FN|90774003|SNOMEDCT_CORE|Victim of physical assault|Victim of physical assault
C0277725|T033|IS|90774003|SNOMEDCT_CORE|Victim of physical assault, NOS|Victim of physical assault
C0277730|T033|SY|56890008|SNOMEDCT_CORE|Sexual assault victim|Victim of sexual aggression
C0277730|T033|PT|56890008|SNOMEDCT_CORE|Victim of sexual aggression|Victim of sexual aggression
C0277730|T033|FN|56890008|SNOMEDCT_CORE|Victim of sexual aggression|Victim of sexual aggression
C0277851|T033|OAS|271772002|SNOMEDCT_CORE|Ankle gives way|Ankle instability
C0277851|T033|PT|813001|SNOMEDCT_CORE|Ankle instability|Ankle instability
C0277851|T033|FN|813001|SNOMEDCT_CORE|Ankle instability|Ankle instability
C0277851|T033|OAS|271772002|SNOMEDCT_CORE|Ankle joint instability|Ankle instability
C0277851|T033|OAP|271772002|SNOMEDCT_CORE|Unstable ankle|Ankle instability
C0277851|T033|OAF|271772002|SNOMEDCT_CORE|Unstable ankle|Ankle instability
C0277877|T033|SY|409609008|SNOMEDCT_CORE|Pulmonary infiltrate|Radiologic infiltrate of lung
C0277877|T033|PT|409609008|SNOMEDCT_CORE|Radiologic infiltrate of lung|Radiologic infiltrate of lung
C0277877|T033|FN|409609008|SNOMEDCT_CORE|Radiologic infiltrate of lung|Radiologic infiltrate of lung
C0277919|T047|PT|238788004|SNOMEDCT_CORE|Venous stasis syndrome|Venous stasis syndrome
C0277919|T047|FN|238788004|SNOMEDCT_CORE|Venous stasis syndrome|Venous stasis syndrome
C0278008|T184|IS|88111009|SNOMEDCT_CORE|Abnormal bowel habits|Altered bowel function
C0278008|T184|PT|88111009|SNOMEDCT_CORE|Altered bowel function|Altered bowel function
C0278008|T184|FN|88111009|SNOMEDCT_CORE|Altered bowel function|Altered bowel function
C0278008|T184|SY|88111009|SNOMEDCT_CORE|Altered bowel habit|Altered bowel function
C0278008|T184|SY|88111009|SNOMEDCT_CORE|Altered bowel habits|Altered bowel function
C0278008|T184|SY|88111009|SNOMEDCT_CORE|Change in bowel habit|Altered bowel function
C0278008|T184|SY|88111009|SNOMEDCT_CORE|Change in bowel pattern|Altered bowel function
C0278061|T048|IS|1855002|SNOMEDCT_CORE|Abnormal mental state|Altered mental status
C0278061|T048|IS|1855002|SNOMEDCT_CORE|Altered mental status|Altered mental status
C0278061|T048|PT|419284004|SNOMEDCT_CORE|Altered mental status|Altered mental status
C0278061|T048|FN|419284004|SNOMEDCT_CORE|Altered mental status|Altered mental status
C0278076|T048|SY|568005|SNOMEDCT_CORE|Habit disorder|Habit disorder
C0278097|T048|PT|5413009|SNOMEDCT_CORE|Abnormal male sexual function|Abnormal male sexual function
C0278097|T048|FN|5413009|SNOMEDCT_CORE|Abnormal male sexual function|Abnormal male sexual function
C0278097|T048|SY|5413009|SNOMEDCT_CORE|Male sexual dysfunction|Abnormal male sexual function
C0278100|T048|PT|28154007|SNOMEDCT_CORE|Abnormal female sexual function|Abnormal female sexual function
C0278100|T048|FN|28154007|SNOMEDCT_CORE|Abnormal female sexual function|Abnormal female sexual function
C0278151|T033|PT|32402008|SNOMEDCT_CORE|Facial spasm|Facial spasm
C0278151|T033|FN|32402008|SNOMEDCT_CORE|Facial spasm|Facial spasm
C0278151|T033|IS|32402008|SNOMEDCT_CORE|Facial spasm, NOS|Facial spasm
C0278152|T047|SY|13753008|SNOMEDCT_CORE|Facial hemispasm|Hemifacial spasm
C0278152|T047|PT|13753008|SNOMEDCT_CORE|Hemifacial spasm|Hemifacial spasm
C0278152|T047|FN|13753008|SNOMEDCT_CORE|Hemifacial spasm|Hemifacial spasm
C0278701|T191|PT|408647009|SNOMEDCT_CORE|Adenocarcinoma of stomach|Adenocarcinoma of stomach
C0278701|T191|FN|408647009|SNOMEDCT_CORE|Adenocarcinoma of stomach|Adenocarcinoma of stomach
C0278701|T191|SY|408647009|SNOMEDCT_CORE|Cancer of stomach, adenocarcinoma|Adenocarcinoma of stomach
C0278996|T191|PT|255056009|SNOMEDCT_CORE|Malignant tumor of head and neck|Malignant tumor of head and neck
C0278996|T191|OF|255056009|SNOMEDCT_CORE|Malignant tumor of head and neck|Malignant tumor of head and neck
C0278996|T191|FN|255056009|SNOMEDCT_CORE|Malignant tumor of head and/or neck|Malignant tumor of head and neck
C0278996|T191|SY|255056009|SNOMEDCT_CORE|Malignant tumor of head and/or neck|Malignant tumor of head and neck
C0278996|T191|PTGB|255056009|SNOMEDCT_CORE|Malignant tumour of head and neck|Malignant tumor of head and neck
C0278996|T191|SYGB|255056009|SNOMEDCT_CORE|Malignant tumour of head and/or neck|Malignant tumor of head and neck
C0279530|T191|PT|428281000|SNOMEDCT_CORE|Malignant neoplasm of bone|Malignant neoplasm of bone
C0279530|T191|FN|428281000|SNOMEDCT_CORE|Malignant neoplasm of bone|Malignant neoplasm of bone
C0279563|T191|PT|109888004|SNOMEDCT_CORE|Lobular carcinoma in situ of breast|Lobular carcinoma in situ of breast
C0279563|T191|FN|109888004|SNOMEDCT_CORE|Lobular carcinoma in situ of breast|Lobular carcinoma in situ of breast
C0279680|T191|SY|255109008|SNOMEDCT_CORE|TCC - Transitional cell carcinoma of bladder|Transitional cell carcinoma of bladder
C0279680|T191|PT|255109008|SNOMEDCT_CORE|Transitional cell carcinoma of bladder|Transitional cell carcinoma of bladder
C0279680|T191|FN|255109008|SNOMEDCT_CORE|Transitional cell carcinoma of bladder|Transitional cell carcinoma of bladder
C0279702|T191|PT|254915003|SNOMEDCT_CORE|Clear cell carcinoma of kidney|Clear cell carcinoma of kidney
C0279702|T191|FN|254915003|SNOMEDCT_CORE|Clear cell carcinoma of kidney|Clear cell carcinoma of kidney
C0279702|T191|SY|254915003|SNOMEDCT_CORE|Clear cell renal cell carcinoma|Clear cell carcinoma of kidney
C0279702|T191|IS|254915003|SNOMEDCT_CORE|Grawitz tumor|Clear cell carcinoma of kidney
C0279702|T191|IS|254915003|SNOMEDCT_CORE|Grawitz tumour|Clear cell carcinoma of kidney
C0280300|T191|SY|276954004|SNOMEDCT_CORE|SCC - Squamous cell carcinoma of floor of mouth|Squamous cell carcinoma of floor of mouth
C0280300|T191|PT|276954004|SNOMEDCT_CORE|Squamous cell carcinoma of floor of mouth|Squamous cell carcinoma of floor of mouth
C0280300|T191|FN|276954004|SNOMEDCT_CORE|Squamous cell carcinoma of floor of mouth|Squamous cell carcinoma of floor of mouth
C0280302|T191|SY|255071008|SNOMEDCT_CORE|SCC - Squamous cell carcinoma of lip|Squamous cell carcinoma of lip
C0280302|T191|PT|255071008|SNOMEDCT_CORE|Squamous cell carcinoma of lip|Squamous cell carcinoma of lip
C0280302|T191|FN|255071008|SNOMEDCT_CORE|Squamous cell carcinoma of lip|Squamous cell carcinoma of lip
C0280324|T191|SY|405822008|SNOMEDCT_CORE|Cancer of the larynx, squamous cell|Squamous cell carcinoma of larynx
C0280324|T191|PT|405822008|SNOMEDCT_CORE|Squamous cell carcinoma of larynx|Squamous cell carcinoma of larynx
C0280324|T191|FN|405822008|SNOMEDCT_CORE|Squamous cell carcinoma of larynx|Squamous cell carcinoma of larynx
C0280793|T191|SY|22217002|SNOMEDCT_CORE|Oligoastrocytoma|Oligoastrocytoma
C0280803|T191|SY|307649006|SNOMEDCT_CORE|Microglioma|Primary central nervous system lymphoma
C0280803|T191|FN|307649006|SNOMEDCT_CORE|Microglioma|Primary central nervous system lymphoma
C0280803|T191|SY|307649006|SNOMEDCT_CORE|PCNSL - Primary CNS lymphoma|Primary central nervous system lymphoma
C0280803|T191|PT|307649006|SNOMEDCT_CORE|Primary central nervous system lymphoma|Primary central nervous system lymphoma
C0280803|T191|SY|307649006|SNOMEDCT_CORE|Primary CNS lymphoma|Primary central nervous system lymphoma
C0281797|T047|PT|202776005|SNOMEDCT_CORE|Cervical root syndrome|Cervical root syndrome
C0281797|T047|FN|202776005|SNOMEDCT_CORE|Cervical root syndrome|Cervical root syndrome
C0281856|T184|PTGB|82991003|SNOMEDCT_CORE|Generalised aches and pains|Generalized aches and pains
C0281856|T184|SYGB|82991003|SNOMEDCT_CORE|Generalised body aches|Generalized aches and pains
C0281856|T184|SYGB|82991003|SNOMEDCT_CORE|Generalised pain|Generalized aches and pains
C0281856|T184|PT|82991003|SNOMEDCT_CORE|Generalized aches and pains|Generalized aches and pains
C0281856|T184|FN|82991003|SNOMEDCT_CORE|Generalized aches and pains|Generalized aches and pains
C0281856|T184|SY|82991003|SNOMEDCT_CORE|Generalized body aches|Generalized aches and pains
C0281856|T184|IS|82991003|SNOMEDCT_CORE|Generalized body pains|Generalized aches and pains
C0281856|T184|SY|82991003|SNOMEDCT_CORE|Generalized pain|Generalized aches and pains
C0281860|T046|PTGB|239160006|SNOMEDCT_CORE|Wound haematoma|Wound hematoma
C0281860|T046|PT|239160006|SNOMEDCT_CORE|Wound hematoma|Wound hematoma
C0281860|T046|FN|239160006|SNOMEDCT_CORE|Wound hematoma|Wound hematoma
C0281883|T037|SY|127287001|SNOMEDCT_CORE|Pertrochanteric fracture of neck of femur|Pertrochanteric fracture of neck of femur
C0281899|T020|PT|202708005|SNOMEDCT_CORE|Prolapsed lumbar intervertebral disc|Prolapsed lumbar intervertebral disc
C0281899|T020|FN|202708005|SNOMEDCT_CORE|Prolapsed lumbar intervertebral disc|Prolapsed lumbar intervertebral disc
C0281926|T037|PT|263247007|SNOMEDCT_CORE|Fracture of calcaneus|Fracture of calcaneus
C0281926|T037|FN|263247007|SNOMEDCT_CORE|Fracture of calcaneus|Fracture of calcaneus
C0281926|T037|SY|263247007|SNOMEDCT_CORE|Fracture of os calcis|Fracture of calcaneus
C0281926|T037|SY|263247007|SNOMEDCT_CORE|Heel bone fracture|Fracture of calcaneus
C0281936|T047|PT|429196001|SNOMEDCT_CORE|Partial obstruction of small bowel|Partial obstruction of small bowel
C0281936|T047|FN|429196001|SNOMEDCT_CORE|Partial obstruction of small bowel|Partial obstruction of small bowel
C0281936|T047|SY|429196001|SNOMEDCT_CORE|Partial obstruction of small intestine|Partial obstruction of small bowel
C0281936|T047|SY|429196001|SNOMEDCT_CORE|Partial small bowel obstruction|Partial obstruction of small bowel
C0281981|T033|SY|297960002|SNOMEDCT_CORE|Lump of skin|Mass of skin
C0281981|T033|PT|297960002|SNOMEDCT_CORE|Mass of skin|Mass of skin
C0281981|T033|FN|297960002|SNOMEDCT_CORE|Mass of skin|Mass of skin
C0282005|T184|PT|271687003|SNOMEDCT_CORE|Swelling of scrotum|Swelling of scrotum
C0282005|T184|FN|271687003|SNOMEDCT_CORE|Swelling of scrotum|Swelling of scrotum
C0282005|T184|SY|271687003|SNOMEDCT_CORE|Swollen scrotum|Swelling of scrotum
C0282015|T037|SY|90070003|SNOMEDCT_CORE|Pneumothorax due to trauma|Traumatic pneumothorax
C0282015|T037|FN|90070003|SNOMEDCT_CORE|Pneumothorax due to trauma|Traumatic pneumothorax
C0282015|T037|PT|90070003|SNOMEDCT_CORE|Traumatic pneumothorax|Traumatic pneumothorax
C0282015|T037|OF|90070003|SNOMEDCT_CORE|Traumatic pneumothorax|Traumatic pneumothorax
C0282015|T037|IS|90070003|SNOMEDCT_CORE|Traumatic pneumothorax, NOS|Traumatic pneumothorax
C0282126|T048|IS|78667006|SNOMEDCT_CORE|Neurotic depression|Neurotic depression
C0282350|T037|SY|213017001|SNOMEDCT_CORE|SA - Sexual abuse|Sexual abuse
C0282350|T037|PT|213017001|SNOMEDCT_CORE|Sexual abuse|Sexual abuse
C0282350|T037|OF|213017001|SNOMEDCT_CORE|Sexual abuse|Sexual abuse
C0282350|T037|FN|213017001|SNOMEDCT_CORE|Sexual abuse|Sexual abuse
C0282488|T047|SY|197834003|SNOMEDCT_CORE|IC - Interstitial cystitis|IC - Interstitial cystitis
C0282488|T047|SY|197834003|SNOMEDCT_CORE|Interstitial cystitis|IC - Interstitial cystitis
C0282504|T047|PT|426232007|SNOMEDCT_CORE|Environmental allergy|Environmental allergy
C0282504|T047|FN|426232007|SNOMEDCT_CORE|Environmental allergy|Environmental allergy
C0282504|T047|OF|426232007|SNOMEDCT_CORE|Environmental allergy|Environmental allergy
C0282612|T191|SY|254901000|SNOMEDCT_CORE|PIN - Prostatic intraepithelial neoplasia|Prostatic intraepithelial neoplasia
C0282612|T191|PT|254901000|SNOMEDCT_CORE|Prostatic intraepithelial neoplasia|Prostatic intraepithelial neoplasia
C0282612|T191|FN|254901000|SNOMEDCT_CORE|Prostatic intraepithelial neoplasia|Prostatic intraepithelial neoplasia
C0300946|T047|SY|48813009|SNOMEDCT_CORE|Alymphocytosis|Alymphocytosis
C0302142|T190|PT|417893002|SNOMEDCT_CORE|Deformity|Deformity
C0302142|T190|FN|417893002|SNOMEDCT_CORE|Deformity|Deformity
C0302180|T047|PT|19672005|SNOMEDCT_CORE|Condyloma|Condyloma
C0302180|T047|FN|19672005|SNOMEDCT_CORE|Condyloma|Condyloma
C0302180|T047|IS|19672005|SNOMEDCT_CORE|Condyloma, NOS|Condyloma
C0302313|T033|SY|203522001|SNOMEDCT_CORE|Osteolytic lesion|Osteolytic lesion
C0302472|T047|PT|396335001|SNOMEDCT_CORE|Acute and chronic cholecystitis|Acute and chronic cholecystitis
C0302472|T047|FN|396335001|SNOMEDCT_CORE|Acute and chronic cholecystitis|Acute and chronic cholecystitis
C0302472|T047|SY|396335001|SNOMEDCT_CORE|Acute on chronic cholecystitis|Acute and chronic cholecystitis
C0302491|T046|PT|274146004|SNOMEDCT_CORE|Pathological fracture of vertebra|Pathological fracture of vertebra
C0302491|T046|FN|274146004|SNOMEDCT_CORE|Pathological fracture of vertebra|Pathological fracture of vertebra
C0302592|T191|PT|285432005|SNOMEDCT_CORE|Carcinoma of cervix|Carcinoma of cervix
C0302592|T191|FN|285432005|SNOMEDCT_CORE|Carcinoma of cervix|Carcinoma of cervix
C0302832|T048|IS|37746008|SNOMEDCT_CORE|Obsessional neurosis|Obsessional neurosis
C0302885|T019|IS|38804009|SNOMEDCT_CORE|Testicular dysgenesis|Testicular dysgenesis
C0302885|T019|IS|38804009|SNOMEDCT_CORE|Testicular dysplasia|Testicular dysgenesis
C0311210|T047|PT|36857002|SNOMEDCT_CORE|Onychia of finger|Onychia of finger
C0311210|T047|FN|36857002|SNOMEDCT_CORE|Onychia of finger|Onychia of finger
C0311210|T047|IS|36857002|SNOMEDCT_CORE|Panaritium of finger|Onychia of finger
C0311210|T047|IS|36857002|SNOMEDCT_CORE|Paronychia of finger|Onychia of finger
C0311210|T047|IS|36857002|SNOMEDCT_CORE|Perionychia of finger|Onychia of finger
C0311211|T047|PT|388983002|SNOMEDCT_CORE|Paronychia of toe|Paronychia of toe
C0311211|T047|FN|388983002|SNOMEDCT_CORE|Paronychia of toe|Paronychia of toe
C0311211|T047|SY|388983002|SNOMEDCT_CORE|Perionychia of toe|Paronychia of toe
C0311223|T047|PT|399114005|SNOMEDCT_CORE|Adhesive capsulitis of shoulder|Adhesive capsulitis of shoulder
C0311223|T047|FN|399114005|SNOMEDCT_CORE|Adhesive capsulitis of shoulder|Adhesive capsulitis of shoulder
C0311223|T047|SY|399114005|SNOMEDCT_CORE|Frozen shoulder|Adhesive capsulitis of shoulder
C0311223|T047|SY|399114005|SNOMEDCT_CORE|Pericapsulitis of shoulder|Adhesive capsulitis of shoulder
C0311245|T019|SY|82525005|SNOMEDCT_CORE|Congenital cyst of kidney|Multiple congenital cysts of kidney
C0311245|T047|SY|82525005|SNOMEDCT_CORE|Congenital cyst of kidney|Multiple congenital cysts of kidney
C0311245|T019|SY|82525005|SNOMEDCT_CORE|Congenital cystic disease of kidney|Multiple congenital cysts of kidney
C0311245|T047|SY|82525005|SNOMEDCT_CORE|Congenital cystic disease of kidney|Multiple congenital cysts of kidney
C0311245|T019|SY|82525005|SNOMEDCT_CORE|Congenital cystic kidney disease|Multiple congenital cysts of kidney
C0311245|T047|SY|82525005|SNOMEDCT_CORE|Congenital cystic kidney disease|Multiple congenital cysts of kidney
C0311245|T019|FN|82525005|SNOMEDCT_CORE|Congenital cystic kidney disease|Multiple congenital cysts of kidney
C0311245|T047|FN|82525005|SNOMEDCT_CORE|Congenital cystic kidney disease|Multiple congenital cysts of kidney
C0311245|T019|SY|82525005|SNOMEDCT_CORE|Congenital polycystic kidney disease|Multiple congenital cysts of kidney
C0311245|T047|SY|82525005|SNOMEDCT_CORE|Congenital polycystic kidney disease|Multiple congenital cysts of kidney
C0311245|T019|PT|82525005|SNOMEDCT_CORE|Multiple congenital cysts of kidney|Multiple congenital cysts of kidney
C0311245|T047|PT|82525005|SNOMEDCT_CORE|Multiple congenital cysts of kidney|Multiple congenital cysts of kidney
C0311245|T019|SY|82525005|SNOMEDCT_CORE|Sponge kidney|Multiple congenital cysts of kidney
C0311245|T047|SY|82525005|SNOMEDCT_CORE|Sponge kidney|Multiple congenital cysts of kidney
C0311310|T047|IS|237044002|SNOMEDCT_CORE|Chronic female pelvic cellulitis|Chronic female pelvic cellulitis
C0311334|T047|PTGB|65120008|SNOMEDCT_CORE|Generalised convulsive epilepsy|Generalized convulsive epilepsy
C0311334|T047|PTGB|4619009|SNOMEDCT_CORE|Generalised-onset seizures|Generalized convulsive epilepsy
C0311334|T047|PT|65120008|SNOMEDCT_CORE|Generalized convulsive epilepsy|Generalized convulsive epilepsy
C0311334|T047|FN|65120008|SNOMEDCT_CORE|Generalized convulsive epilepsy|Generalized convulsive epilepsy
C0311334|T047|IS|65120008|SNOMEDCT_CORE|Generalized convulsive epilepsy, NOS|Generalized convulsive epilepsy
C0311334|T047|PT|4619009|SNOMEDCT_CORE|Generalized-onset seizures|Generalized convulsive epilepsy
C0311334|T047|FN|4619009|SNOMEDCT_CORE|Generalized-onset seizures|Generalized convulsive epilepsy
C0311334|T047|IS|4619009|SNOMEDCT_CORE|Generalized-onset seizures, NOS|Generalized convulsive epilepsy
C0311335|T047|SY|13973009|SNOMEDCT_CORE|Convulsive status epilepticus|Grand mal status
C0311335|T047|PT|13973009|SNOMEDCT_CORE|Grand mal status|Grand mal status
C0311335|T047|FN|13973009|SNOMEDCT_CORE|Grand mal status|Grand mal status
C0311337|T047|SY|30085007|SNOMEDCT_CORE|Interdigital neuralgia|Morton's metatarsalgia
C0311337|T047|SY|30085007|SNOMEDCT_CORE|Interdigital neuroma|Morton's metatarsalgia
C0311337|T047|SY|30085007|SNOMEDCT_CORE|Morton metatarsalgia|Morton's metatarsalgia
C0311337|T047|SY|30085007|SNOMEDCT_CORE|Morton neuroma|Morton's metatarsalgia
C0311337|T047|SY|30085007|SNOMEDCT_CORE|Morton's disease|Morton's metatarsalgia
C0311337|T047|PT|30085007|SNOMEDCT_CORE|Morton's metatarsalgia|Morton's metatarsalgia
C0311337|T047|FN|30085007|SNOMEDCT_CORE|Morton's metatarsalgia|Morton's metatarsalgia
C0311337|T047|SY|30085007|SNOMEDCT_CORE|Morton's neuralgia|Morton's metatarsalgia
C0311337|T047|SY|30085007|SNOMEDCT_CORE|Morton's neuroma|Morton's metatarsalgia
C0311337|T047|SY|30085007|SNOMEDCT_CORE|Morton's toe|Morton's metatarsalgia
C0311337|T047|SY|30085007|SNOMEDCT_CORE|Mortons neuroma|Morton's metatarsalgia
C0311341|T047|SY|44219007|SNOMEDCT_CORE|PEX - Pseudoexfoliation|Pseudoexfoliation of lens capsule
C0311341|T047|SY|44219007|SNOMEDCT_CORE|Pseudoexfoliation lens capsule|Pseudoexfoliation of lens capsule
C0311341|T047|PT|44219007|SNOMEDCT_CORE|Pseudoexfoliation of lens capsule|Pseudoexfoliation of lens capsule
C0311341|T047|FN|44219007|SNOMEDCT_CORE|Pseudoexfoliation of lens capsule|Pseudoexfoliation of lens capsule
C0311341|T047|SY|44219007|SNOMEDCT_CORE|PXF - Pseudoexfoliation of lens capsule|Pseudoexfoliation of lens capsule
C0311349|T047|IS|40608009|SNOMEDCT_CORE|Constant vertical heterotropia|Constant vertical heterotropia
C0311370|T047|SY|19267009|SNOMEDCT_CORE|Lupus anticoagulant|Lupus anticoagulant disorder
C0311370|T047|PT|19267009|SNOMEDCT_CORE|Lupus anticoagulant disorder|Lupus anticoagulant disorder
C0311370|T047|FN|19267009|SNOMEDCT_CORE|Lupus anticoagulant disorder|Lupus anticoagulant disorder
C0311370|T047|SY|19267009|SNOMEDCT_CORE|Lupus anticoagulant inhibitor syndrome|Lupus anticoagulant disorder
C0311370|T047|SY|19267009|SNOMEDCT_CORE|SLE inhibitor syndrome|Lupus anticoagulant disorder
C0311389|T047|IS|31822004|SNOMEDCT_CORE|Urethritis, NOS|Urethritis, NOS
C0311394|T033|IS|228158008|SNOMEDCT_CORE|Difficulty walking|Walking disability
C0311394|T033|SY|228158008|SNOMEDCT_CORE|Impaired walking|Walking disability
C0311394|T033|PT|228158008|SNOMEDCT_CORE|Walking disability|Walking disability
C0311394|T033|FN|228158008|SNOMEDCT_CORE|Walking disability|Walking disability
C0314719|T184|OAP|1249004|SNOMEDCT_CORE|Dry eye|Dryness of eye
C0314719|T184|OAF|1249004|SNOMEDCT_CORE|Dry eye|Dryness of eye
C0314719|T184|IS|1249004|SNOMEDCT_CORE|Dryness of eye|Dryness of eye
C0332544|T184|SY|161833006|SNOMEDCT_CORE|Abnormal increase in weight|Abnormal weight gain
C0332544|T184|PT|161833006|SNOMEDCT_CORE|Abnormal weight gain|Abnormal weight gain
C0332544|T184|FN|161833006|SNOMEDCT_CORE|Abnormal weight gain|Abnormal weight gain
C0332563|T033|SY|25694009|SNOMEDCT_CORE|Papula|Papule
C0332563|T033|SY|25694009|SNOMEDCT_CORE|Papulae|Papule
C0332563|T033|OAP|443871003|SNOMEDCT_CORE|Papule|Papule
C0332563|T033|PT|25694009|SNOMEDCT_CORE|Papule|Papule
C0332563|T033|FN|25694009|SNOMEDCT_CORE|Papule|Papule
C0332563|T033|OAF|443871003|SNOMEDCT_CORE|Papule|Papule
C0332563|T033|IS|25694009|SNOMEDCT_CORE|Papule, NOS|Papule
C0332679|T037|PT|125665001|SNOMEDCT_CORE|Crushing injury|Crushing injury
C0332679|T037|FN|125665001|SNOMEDCT_CORE|Crushing injury|Crushing injury
C0332679|T037|SY|125665001|SNOMEDCT_CORE|Crushing injury - disorder|Crushing injury
C0332687|T037|PT|403191005|SNOMEDCT_CORE|Partial thickness burn|Partial thickness burn
C0332687|T037|FN|403191005|SNOMEDCT_CORE|Partial thickness burn|Partial thickness burn
C0332687|T037|SY|403191005|SNOMEDCT_CORE|Second degree burn|Partial thickness burn
C0332687|T037|OF|403191005|SNOMEDCT_CORE|Second degree burn|Partial thickness burn
C0332743|T046|PT|134194006|SNOMEDCT_CORE|Delayed union of fracture|Delayed union of fracture
C0332743|T046|OF|134194006|SNOMEDCT_CORE|Delayed union of fracture|Delayed union of fracture
C0332743|T046|PT|28087009|SNOMEDCT_CORE|Delayed union of fracture|Delayed union of fracture
C0332743|T046|FN|28087009|SNOMEDCT_CORE|Delayed union of fracture|Delayed union of fracture
C0332743|T046|FN|134194006|SNOMEDCT_CORE|Delayed union of fracture|Delayed union of fracture
C0332743|T046|SY|28087009|SNOMEDCT_CORE|Fracture, delayed union|Delayed union of fracture
C0332743|T046|OF|28087009|SNOMEDCT_CORE|Fracture, delayed union|Delayed union of fracture
C0332743|T046|IS|28087009|SNOMEDCT_CORE|Fracture, delayed union, NOS|Delayed union of fracture
C0332798|T037|PT|125643001|SNOMEDCT_CORE|Open wound|Open wound
C0332798|T037|FN|125643001|SNOMEDCT_CORE|Open wound|Open wound
C0332798|T037|SY|125643001|SNOMEDCT_CORE|Open wound of body region|Open wound
C0332815|T037|PT|429305003|SNOMEDCT_CORE|Nonvenomous insect bite|Nonvenomous insect bite
C0332815|T037|FN|429305003|SNOMEDCT_CORE|Nonvenomous insect bite|Nonvenomous insect bite
C0333014|T047|PT|197794008|SNOMEDCT_CORE|Staghorn calculus|Staghorn calculus
C0333014|T047|FN|197794008|SNOMEDCT_CORE|Staghorn calculus|Staghorn calculus
C0333128|T047|SY|247467008|SNOMEDCT_CORE|Blackhead|Blackhead
C0333355|T046|PT|95361005|SNOMEDCT_CORE|Inflammatory disease of mucous membrane|Inflammatory disease of mucous membrane
C0333355|T046|FN|95361005|SNOMEDCT_CORE|Inflammatory disease of mucous membrane|Inflammatory disease of mucous membrane
C0333355|T046|SY|95361005|SNOMEDCT_CORE|Mucitis|Inflammatory disease of mucous membrane
C0333355|T046|IS|95361005|SNOMEDCT_CORE|Mucitis, NOS|Inflammatory disease of mucous membrane
C0333355|T046|SY|95361005|SNOMEDCT_CORE|Mucosal inflammation|Inflammatory disease of mucous membrane
C0333355|T046|IS|95361005|SNOMEDCT_CORE|Mucosal inflammation, NOS|Inflammatory disease of mucous membrane
C0333355|T046|SY|95361005|SNOMEDCT_CORE|Mucositis|Inflammatory disease of mucous membrane
C0333355|T046|IS|95361005|SNOMEDCT_CORE|Mucositis, NOS|Inflammatory disease of mucous membrane
C0333355|T046|SY|95361005|SNOMEDCT_CORE|Mucous membrane inflammation|Inflammatory disease of mucous membrane
C0333355|T046|IS|95361005|SNOMEDCT_CORE|Mucous membrane inflammation disorder|Inflammatory disease of mucous membrane
C0333355|T046|IS|95361005|SNOMEDCT_CORE|Mucous membrane inflammation, NOS|Inflammatory disease of mucous membrane
C0333559|T047|SY|230698000|SNOMEDCT_CORE|LACI - Lacunar infarction|Lacunar infarction
C0333559|T047|PT|230698000|SNOMEDCT_CORE|Lacunar infarction|Lacunar infarction
C0333559|T047|FN|230698000|SNOMEDCT_CORE|Lacunar infarction|Lacunar infarction
C0333559|T047|SY|230698000|SNOMEDCT_CORE|LI - Lacunar infarction|Lacunar infarction
C0333616|T046|SY|238699007|SNOMEDCT_CORE|Post-inflammatory hypermelanosis|Post-inflammatory hyperpigmentation
C0333616|T046|PT|238699007|SNOMEDCT_CORE|Post-inflammatory hyperpigmentation|Post-inflammatory hyperpigmentation
C0333616|T046|FN|238699007|SNOMEDCT_CORE|Post-inflammatory hyperpigmentation|Post-inflammatory hyperpigmentation
C0333616|T046|SY|238699007|SNOMEDCT_CORE|Postinflammatory hyperpigmentation|Post-inflammatory hyperpigmentation
C0334082|T047|OF|239107007|SNOMEDCT_CORE|Epidermal naevus|Epidermal nevus
C0334082|T047|PTGB|239107007|SNOMEDCT_CORE|Epidermal naevus|Epidermal nevus
C0334082|T047|FN|239107007|SNOMEDCT_CORE|Epidermal nevus|Epidermal nevus
C0334082|T047|PT|239107007|SNOMEDCT_CORE|Epidermal nevus|Epidermal nevus
C0334245|T191|PT|400066006|SNOMEDCT_CORE|Intraepithelial squamous cell carcinoma|Intraepithelial squamous cell carcinoma
C0334245|T191|FN|400066006|SNOMEDCT_CORE|Intraepithelial squamous cell carcinoma|Intraepithelial squamous cell carcinoma
C0334246|T191|PT|403906006|SNOMEDCT_CORE|Metastatic squamous cell carcinoma|Metastatic squamous cell carcinoma
C0334246|T191|FN|403906006|SNOMEDCT_CORE|Metastatic squamous cell carcinoma|Metastatic squamous cell carcinoma
C0334292|T191|SY|19665009|SNOMEDCT_CORE|Tubular adenoma|Tubular adenoma
C0334292|T191|PT|444408007|SNOMEDCT_CORE|Tubular adenoma|Tubular adenoma
C0334292|T191|OF|19665009|SNOMEDCT_CORE|Tubular adenoma|Tubular adenoma
C0334292|T191|FN|444408007|SNOMEDCT_CORE|Tubular adenoma|Tubular adenoma
C0334292|T191|OF|19665009|SNOMEDCT_CORE|Tubular adenoma, no ICD-O subtype|Tubular adenoma
C0334292|T191|PT|19665009|SNOMEDCT_CORE|Tubular adenoma, no ICD-O subtype|Tubular adenoma
C0334292|T191|SY|19665009|SNOMEDCT_CORE|Tubular adenoma, no International Classification of Diseases for Oncology subtype|Tubular adenoma
C0334292|T191|FN|19665009|SNOMEDCT_CORE|Tubular adenoma, no International Classification of Diseases for Oncology subtype|Tubular adenoma
C0334292|T191|IS|19665009|SNOMEDCT_CORE|Tubular adenoma, NOS|Tubular adenoma
C0334463|T191|PT|34360000|SNOMEDCT_CORE|Fibrous histiocytoma, malignant|Malignant fibrous histiocytoma
C0334463|T191|FN|34360000|SNOMEDCT_CORE|Fibrous histiocytoma, malignant|Malignant fibrous histiocytoma
C0334463|T191|SY|34360000|SNOMEDCT_CORE|Fibroxanthoma, malignant|Malignant fibrous histiocytoma
C0334463|T191|SY|34360000|SNOMEDCT_CORE|Malignant fibrous histiocytoma|Malignant fibrous histiocytoma
C0334463|T191|PT|443439001|SNOMEDCT_CORE|Malignant fibrous histiocytoma|Malignant fibrous histiocytoma
C0334463|T191|FN|443439001|SNOMEDCT_CORE|Malignant fibrous histiocytoma|Malignant fibrous histiocytoma
C0334463|T191|SY|34360000|SNOMEDCT_CORE|Malignant fibroxanthoma|Malignant fibrous histiocytoma
C0334463|T191|SY|34360000|SNOMEDCT_CORE|Undifferentiated high grade pleomorphic sarcoma|Malignant fibrous histiocytoma
C0334634|T191|IS|74654000|SNOMEDCT_CORE|Malignant lymphoma, centrocytic|Mantle cell lymphoma
C0334634|T191|IS|74654000|SNOMEDCT_CORE|Malignant lymphoma, lymphocytic, intermediate differentiation, diffuse|Mantle cell lymphoma
C0334634|T191|PT|74654000|SNOMEDCT_CORE|Mantle cell lymphoma|Mantle cell lymphoma
C0334634|T191|FN|74654000|SNOMEDCT_CORE|Mantle cell lymphoma|Mantle cell lymphoma
C0334634|T191|IS|74654000|SNOMEDCT_CORE|Mantle zone lymphoma|Mantle cell lymphoma
C0334638|T191|SY|74654000|SNOMEDCT_CORE|Malignant lymphomatous polyposis|Malignant lymphomatous polyposis
C0334678|T191|SYGB|128845005|SNOMEDCT_CORE|Refractory anaemia without sideroblasts|Refractory anemia without sideroblasts
C0334678|T191|SY|128845005|SNOMEDCT_CORE|Refractory anemia without sideroblasts|Refractory anemia without sideroblasts
C0337212|T033|PT|86591008|SNOMEDCT_CORE|Fall from ladder|Fall from ladder
C0337212|T033|OF|86591008|SNOMEDCT_CORE|Fall from ladder|Fall from ladder
C0337212|T033|FN|86591008|SNOMEDCT_CORE|Fall from ladder|Fall from ladder
C0337212|T033|SY|86591008|SNOMEDCT_CORE|Fall off ladder|Fall from ladder
C0337212|T033|IS|86591008|SNOMEDCT_CORE|Fall on and from ladder|Fall from ladder
C0337234|T033|PT|41411008|SNOMEDCT_CORE|Fall from playground equipment|Fall from playground equipment
C0337234|T033|OF|41411008|SNOMEDCT_CORE|Fall from playground equipment|Fall from playground equipment
C0337234|T033|FN|41411008|SNOMEDCT_CORE|Fall from playground equipment|Fall from playground equipment
C0337234|T033|IS|41411008|SNOMEDCT_CORE|Fall from playground equipment, NOS|Fall from playground equipment
C0337234|T033|IS|41411008|SNOMEDCT_CORE|Fall involving playground equipment|Fall from playground equipment
C0337234|T033|SY|41411008|SNOMEDCT_CORE|Fall involving playground equipment|Fall from playground equipment
C0337253|T037|PT|71893005|SNOMEDCT_CORE|Struck by falling object|Struck by falling object
C0337253|T037|OF|71893005|SNOMEDCT_CORE|Struck by falling object|Struck by falling object
C0337253|T037|FN|71893005|SNOMEDCT_CORE|Struck by falling object|Struck by falling object
C0337253|T037|IS|71893005|SNOMEDCT_CORE|Struck by falling object, NOS|Struck by falling object
C0337616|T033|PT|4506002|SNOMEDCT_CORE|Educational problem|Educational problem
C0337616|T033|FN|4506002|SNOMEDCT_CORE|Educational problem|Educational problem
C0337629|T033|OAP|5015009|SNOMEDCT_CORE|Economic problem|Economic problem
C0337629|T033|OAF|5015009|SNOMEDCT_CORE|Economic problem|Economic problem
C0337664|T033|PT|77176002|SNOMEDCT_CORE|Smoker|Smoker
C0337664|T033|FN|77176002|SNOMEDCT_CORE|Smoker|Smoker
C0337664|T033|OF|77176002|SNOMEDCT_CORE|Smoker|Smoker
C0337664|T033|IS|77176002|SNOMEDCT_CORE|Smoker, NOS|Smoker
C0337667|T033|FN|65568007|SNOMEDCT_CORE|Cigarette smoker|Cigarette smoker
C0337667|T033|PT|65568007|SNOMEDCT_CORE|Cigarette smoker|Cigarette smoker
C0337667|T033|OF|65568007|SNOMEDCT_CORE|Cigarette smoker|Cigarette smoker
C0337667|T033|IS|65568007|SNOMEDCT_CORE|Cigarette smoker, NOS|Cigarette smoker
C0337671|T033|SY|8517006|SNOMEDCT_CORE|Cessation of smoking|Ex-smoker
C0337671|T033|PT|8517006|SNOMEDCT_CORE|Ex-smoker|Ex-smoker
C0337671|T033|FN|8517006|SNOMEDCT_CORE|Ex-smoker|Ex-smoker
C0337671|T033|OF|8517006|SNOMEDCT_CORE|Ex-smoker|Ex-smoker
C0337671|T033|IS|8517006|SNOMEDCT_CORE|Former smoker|Ex-smoker
C0337671|T033|SY|8517006|SNOMEDCT_CORE|Past tobacco smoker|Ex-smoker
C0337681|T033|PT|70545002|SNOMEDCT_CORE|Narcotic drug user|Narcotic drug user
C0337681|T033|FN|70545002|SNOMEDCT_CORE|Narcotic drug user|Narcotic drug user
C0337681|T033|OF|70545002|SNOMEDCT_CORE|Narcotic drug user|Narcotic drug user
C0338078|T191|PT|254962005|SNOMEDCT_CORE|Functionless pituitary adenoma|Functionless pituitary adenoma
C0338078|T191|FN|254962005|SNOMEDCT_CORE|Functionless pituitary adenoma|Functionless pituitary adenoma
C0338078|T191|SY|254962005|SNOMEDCT_CORE|Non-functioning pituitary adenoma|Functionless pituitary adenoma
C0338078|T191|IS|254962005|SNOMEDCT_CORE|Non-functioning pituitary tumor|Functionless pituitary adenoma
C0338078|T191|IS|254962005|SNOMEDCT_CORE|Non-functioning pituitary tumour|Functionless pituitary adenoma
C0338078|T191|SY|254962005|SNOMEDCT_CORE|Null cell pituitary adenoma|Functionless pituitary adenoma
C0338451|T047|PT|230270009|SNOMEDCT_CORE|Frontotemporal dementia|Frontotemporal dementia
C0338451|T047|FN|230270009|SNOMEDCT_CORE|Frontotemporal dementia|Frontotemporal dementia
C0338451|T047|SY|230270009|SNOMEDCT_CORE|Pick's disease|Frontotemporal dementia
C0338451|T047|SY|230270009|SNOMEDCT_CORE|Picks disease|Frontotemporal dementia
C0338480|T047|SY|56097005|SNOMEDCT_CORE|Atypical migraine|Migraine without aura
C0338480|T047|SY|56097005|SNOMEDCT_CORE|Common migraine|Migraine without aura
C0338480|T047|PT|56097005|SNOMEDCT_CORE|Migraine without aura|Migraine without aura
C0338480|T047|FN|56097005|SNOMEDCT_CORE|Migraine without aura|Migraine without aura
C0338480|T047|IS|56097005|SNOMEDCT_CORE|Sick headache|Migraine without aura
C0338481|T047|SY|95655001|SNOMEDCT_CORE|Ocular migraine|Ophthalmic migraine
C0338481|T047|PT|95655001|SNOMEDCT_CORE|Ophthalmic migraine|Ophthalmic migraine
C0338481|T047|FN|95655001|SNOMEDCT_CORE|Ophthalmic migraine|Ophthalmic migraine
C0338483|T047|SY|193039006|SNOMEDCT_CORE|Complex migraine|Complicated migraine
C0338483|T047|PT|193039006|SNOMEDCT_CORE|Complicated migraine|Complicated migraine
C0338483|T047|FN|193039006|SNOMEDCT_CORE|Complicated migraine|Complicated migraine
C0338486|T047|SY|230465000|SNOMEDCT_CORE|Acephalgic migraine|Migraine aura without headache
C0338486|T047|SY|230465000|SNOMEDCT_CORE|Migraine accompaniment|Migraine aura without headache
C0338486|T047|PT|230465000|SNOMEDCT_CORE|Migraine aura without headache|Migraine aura without headache
C0338486|T047|FN|230465000|SNOMEDCT_CORE|Migraine aura without headache|Migraine aura without headache
C0338502|T047|SY|95499004|SNOMEDCT_CORE|Hypoplasia of optic nerve|Hypoplasia of the optic nerve
C0338502|T047|PT|95499004|SNOMEDCT_CORE|Hypoplasia of the optic nerve|Hypoplasia of the optic nerve
C0338502|T047|FN|95499004|SNOMEDCT_CORE|Hypoplasia of the optic nerve|Hypoplasia of the optic nerve
C0338502|T047|SY|95499004|SNOMEDCT_CORE|ONH - Optic nerve hypoplasia|Hypoplasia of the optic nerve
C0338502|T047|SY|95499004|SNOMEDCT_CORE|Optic nerve hypoplasia|Hypoplasia of the optic nerve
C0338538|T047|PT|95675005|SNOMEDCT_CORE|Ulnar neuritis|Ulnar neuritis
C0338538|T047|FN|95675005|SNOMEDCT_CORE|Ulnar neuritis|Ulnar neuritis
C0338573|T047|PT|192759008|SNOMEDCT_CORE|Cerebral venous sinus thrombosis|Cerebral venous sinus thrombosis
C0338573|T047|FN|192759008|SNOMEDCT_CORE|Cerebral venous sinus thrombosis|Cerebral venous sinus thrombosis
C0338573|T047|SY|192759008|SNOMEDCT_CORE|Thrombosis of intracranial venous sinus|Cerebral venous sinus thrombosis
C0338585|T047|OAP|230729006|SNOMEDCT_CORE|Carotid artery dissection|Dissection of carotid artery
C0338585|T047|OAF|230729006|SNOMEDCT_CORE|Carotid artery dissection|Dissection of carotid artery
C0338585|T047|OAS|230729006|SNOMEDCT_CORE|Dissection of carotid artery|Dissection of carotid artery
C0338591|T048|SY|230736007|SNOMEDCT_CORE|TGA - Transient global amnesia|Transient global amnesia
C0338591|T048|PT|230736007|SNOMEDCT_CORE|Transient global amnesia|Transient global amnesia
C0338591|T048|FN|230736007|SNOMEDCT_CORE|Transient global amnesia|Transient global amnesia
C0338596|T019|SY|230773005|SNOMEDCT_CORE|Congenital spastic cerebral palsy|Spastic cerebral palsy
C0338596|T047|SY|230773005|SNOMEDCT_CORE|Congenital spastic cerebral palsy|Spastic cerebral palsy
C0338596|T019|SY|230773005|SNOMEDCT_CORE|Congenital spastic paralysis|Spastic cerebral palsy
C0338596|T047|SY|230773005|SNOMEDCT_CORE|Congenital spastic paralysis|Spastic cerebral palsy
C0338596|T019|SY|230773005|SNOMEDCT_CORE|Infantile spastic cerebral palsy|Spastic cerebral palsy
C0338596|T047|SY|230773005|SNOMEDCT_CORE|Infantile spastic cerebral palsy|Spastic cerebral palsy
C0338596|T019|SY|230773005|SNOMEDCT_CORE|Little's disease|Spastic cerebral palsy
C0338596|T047|SY|230773005|SNOMEDCT_CORE|Little's disease|Spastic cerebral palsy
C0338596|T019|SY|230773005|SNOMEDCT_CORE|Pyramidal cerebral palsy|Spastic cerebral palsy
C0338596|T047|SY|230773005|SNOMEDCT_CORE|Pyramidal cerebral palsy|Spastic cerebral palsy
C0338596|T019|PT|230773005|SNOMEDCT_CORE|Spastic cerebral palsy|Spastic cerebral palsy
C0338596|T047|PT|230773005|SNOMEDCT_CORE|Spastic cerebral palsy|Spastic cerebral palsy
C0338596|T019|FN|230773005|SNOMEDCT_CORE|Spastic cerebral palsy|Spastic cerebral palsy
C0338596|T047|FN|230773005|SNOMEDCT_CORE|Spastic cerebral palsy|Spastic cerebral palsy
C0338596|T019|SY|230773005|SNOMEDCT_CORE|Spastic infantile paralysis|Spastic cerebral palsy
C0338596|T047|SY|230773005|SNOMEDCT_CORE|Spastic infantile paralysis|Spastic cerebral palsy
C0338632|T048|PT|191519005|SNOMEDCT_CORE|Dementia associated with another disease|Dementia associated with another disease
C0338632|T048|FN|191519005|SNOMEDCT_CORE|Dementia associated with another disease|Dementia associated with another disease
C0338632|T048|IS|191519005|SNOMEDCT_CORE|Dementia in conditions EC|Dementia associated with another disease
C0338632|T048|OF|191519005|SNOMEDCT_CORE|Dementia in conditions EC|Dementia associated with another disease
C0338656|T048|SY|386806002|SNOMEDCT_CORE|Cognitive decline|Impaired cognition
C0338656|T048|SY|386806002|SNOMEDCT_CORE|Cognitive deficit|Impaired cognition
C0338656|T048|SY|386806002|SNOMEDCT_CORE|Cognitive disturbance|Impaired cognition
C0338656|T048|SY|386806002|SNOMEDCT_CORE|Cognitive dysfunction|Impaired cognition
C0338656|T048|SY|386806002|SNOMEDCT_CORE|Cognitive impairment|Impaired cognition
C0338656|T048|PT|386806002|SNOMEDCT_CORE|Impaired cognition|Impaired cognition
C0338656|T048|FN|386806002|SNOMEDCT_CORE|Impaired cognition|Impaired cognition
C0338676|T048|PT|191938005|SNOMEDCT_CORE|Nondependent mixed drug abuse in remission|Nondependent mixed drug abuse in remission
C0338676|T048|FN|191938005|SNOMEDCT_CORE|Nondependent mixed drug abuse in remission|Nondependent mixed drug abuse in remission
C0338687|T048|PT|191918009|SNOMEDCT_CORE|Nondependent cocaine abuse, continuous|Nondependent cocaine abuse, continuous
C0338687|T048|FN|191918009|SNOMEDCT_CORE|Nondependent cocaine abuse, continuous|Nondependent cocaine abuse, continuous
C0338688|T048|PT|191919001|SNOMEDCT_CORE|Nondependent cocaine abuse, episodic|Nondependent cocaine abuse, episodic
C0338688|T048|FN|191919001|SNOMEDCT_CORE|Nondependent cocaine abuse, episodic|Nondependent cocaine abuse, episodic
C0338689|T048|PT|191920007|SNOMEDCT_CORE|Nondependent cocaine abuse in remission|Nondependent cocaine abuse in remission
C0338689|T048|FN|191920007|SNOMEDCT_CORE|Nondependent cocaine abuse in remission|Nondependent cocaine abuse in remission
C0338693|T048|PT|191914006|SNOMEDCT_CORE|Nondependent opioid abuse in remission|Nondependent opioid abuse in remission
C0338693|T048|FN|191914006|SNOMEDCT_CORE|Nondependent opioid abuse in remission|Nondependent opioid abuse in remission
C0338707|T048|PT|191894006|SNOMEDCT_CORE|Nondependent cannabis abuse, episodic|Nondependent cannabis abuse, episodic
C0338707|T048|FN|191894006|SNOMEDCT_CORE|Nondependent cannabis abuse, episodic|Nondependent cannabis abuse, episodic
C0338708|T048|PT|191895007|SNOMEDCT_CORE|Nondependent cannabis abuse in remission|Nondependent cannabis abuse in remission
C0338708|T048|FN|191895007|SNOMEDCT_CORE|Nondependent cannabis abuse in remission|Nondependent cannabis abuse in remission
C0338710|T048|PT|191882002|SNOMEDCT_CORE|Nondependent alcohol abuse, continuous|Nondependent alcohol abuse, continuous
C0338710|T048|FN|191882002|SNOMEDCT_CORE|Nondependent alcohol abuse, continuous|Nondependent alcohol abuse, continuous
C0338711|T048|PT|191883007|SNOMEDCT_CORE|Nondependent alcohol abuse, episodic|Nondependent alcohol abuse, episodic
C0338711|T048|FN|191883007|SNOMEDCT_CORE|Nondependent alcohol abuse, episodic|Nondependent alcohol abuse, episodic
C0338712|T048|PT|191884001|SNOMEDCT_CORE|Nondependent alcohol abuse in remission|Nondependent alcohol abuse in remission
C0338712|T048|FN|191884001|SNOMEDCT_CORE|Nondependent alcohol abuse in remission|Nondependent alcohol abuse in remission
C0338726|T048|PT|191889006|SNOMEDCT_CORE|Tobacco dependence in remission|Tobacco dependence in remission
C0338726|T048|FN|191889006|SNOMEDCT_CORE|Tobacco dependence in remission|Tobacco dependence in remission
C0338726|T048|SY|191889006|SNOMEDCT_CORE|Tobacco dependence, in remission|Tobacco dependence in remission
C0338728|T048|PT|191871005|SNOMEDCT_CORE|Combined drug dependence, excluding opioids|Combined drug dependence, excluding opioids
C0338728|T048|FN|191871005|SNOMEDCT_CORE|Combined drug dependence, excluding opioids|Combined drug dependence, excluding opioids
C0338732|T047|PT|191875001|SNOMEDCT_CORE|Combined drug dependence, excluding opioid, in remission|Combined drug dependence, excluding opioid, in remission
C0338732|T047|FN|191875001|SNOMEDCT_CORE|Combined drug dependence, excluding opioid, in remission|Combined drug dependence, excluding opioid, in remission
C0338734|T048|FN|191865004|SNOMEDCT_CORE|Combined opioid with non-opioid drug dependence|Combined opioid with other drug dependence
C0338734|T048|SY|191865004|SNOMEDCT_CORE|Combined opioid with non-opioid drug dependence|Combined opioid with other drug dependence
C0338734|T048|PT|191865004|SNOMEDCT_CORE|Combined opioid with other drug dependence|Combined opioid with other drug dependence
C0338734|T048|OF|191865004|SNOMEDCT_CORE|Combined opioid with other drug dependence|Combined opioid with other drug dependence
C0338755|T048|SY|191845006|SNOMEDCT_CORE|Amfetamine or psychostimulant dependence in remission|Amphetamine or psychostimulant dependence in remission
C0338755|T048|PT|191845006|SNOMEDCT_CORE|Amphetamine or psychostimulant dependence in remission|Amphetamine or psychostimulant dependence in remission
C0338755|T048|FN|191845006|SNOMEDCT_CORE|Amphetamine or psychostimulant dependence in remission|Amphetamine or psychostimulant dependence in remission
C0338757|T048|PT|191837001|SNOMEDCT_CORE|Cannabis dependence, continuous|Cannabis dependence, continuous
C0338757|T048|FN|191837001|SNOMEDCT_CORE|Cannabis dependence, continuous|Cannabis dependence, continuous
C0338762|T048|PT|191831000|SNOMEDCT_CORE|Cocaine dependence, continuous|Cocaine dependence, continuous
C0338762|T048|FN|191831000|SNOMEDCT_CORE|Cocaine dependence, continuous|Cocaine dependence, continuous
C0338763|T048|PT|191832007|SNOMEDCT_CORE|Cocaine dependence, episodic|Cocaine dependence, episodic
C0338763|T048|FN|191832007|SNOMEDCT_CORE|Cocaine dependence, episodic|Cocaine dependence, episodic
C0338771|T048|SY|268640002|SNOMEDCT_CORE|Dependent sedative or hypnotic drug abuse|Hypnotic or anxiolytic dependence
C0338771|T048|PT|268640002|SNOMEDCT_CORE|Hypnotic or anxiolytic dependence|Hypnotic or anxiolytic dependence
C0338771|T048|FN|268640002|SNOMEDCT_CORE|Hypnotic or anxiolytic dependence|Hypnotic or anxiolytic dependence
C0338779|T047|PT|191819002|SNOMEDCT_CORE|Continuous opioid dependence|Continuous opioid dependence
C0338779|T047|FN|191819002|SNOMEDCT_CORE|Continuous opioid dependence|Continuous opioid dependence
C0338781|T047|PT|191821007|SNOMEDCT_CORE|Opioid dependence in remission|Opioid dependence in remission
C0338781|T047|FN|191821007|SNOMEDCT_CORE|Opioid dependence in remission|Opioid dependence in remission
C0338783|T047|PT|191813001|SNOMEDCT_CORE|Chronic alcoholism in remission|Chronic alcoholism in remission
C0338783|T047|FN|191813001|SNOMEDCT_CORE|Chronic alcoholism in remission|Chronic alcoholism in remission
C0338784|T048|PT|191812006|SNOMEDCT_CORE|Episodic chronic alcoholism|Episodic chronic alcoholism
C0338784|T048|FN|191812006|SNOMEDCT_CORE|Episodic chronic alcoholism|Episodic chronic alcoholism
C0338785|T048|PT|191811004|SNOMEDCT_CORE|Continuous chronic alcoholism|Continuous chronic alcoholism
C0338785|T048|FN|191811004|SNOMEDCT_CORE|Continuous chronic alcoholism|Continuous chronic alcoholism
C0338828|T048|PT|191574005|SNOMEDCT_CORE|Schizoaffective schizophrenia in remission|Schizoaffective schizophrenia in remission
C0338828|T048|FN|191574005|SNOMEDCT_CORE|Schizoaffective schizophrenia in remission|Schizoaffective schizophrenia in remission
C0338828|T048|SY|191574005|SNOMEDCT_CORE|Schizoaffective schizophrenia, in remission|Schizoaffective schizophrenia in remission
C0338828|T048|SY|191574005|SNOMEDCT_CORE|Schizophrenia, schizoaffective, in remission|Schizoaffective schizophrenia in remission
C0338831|T048|PT|231494001|SNOMEDCT_CORE|Mania|Mania
C0338831|T048|FN|231494001|SNOMEDCT_CORE|Mania|Mania
C0338831|T048|SY|231494001|SNOMEDCT_CORE|Manic|Mania
C0338873|T048|PT|191618007|SNOMEDCT_CORE|Bipolar affective disorder, current episode manic|Bipolar affective disorder, current episode manic
C0338873|T048|FN|191618007|SNOMEDCT_CORE|Bipolar affective disorder, current episode manic|Bipolar affective disorder, current episode manic
C0338873|T048|SY|191618007|SNOMEDCT_CORE|Manic-depressive - now manic|Bipolar affective disorder, current episode manic
C0338878|T048|PT|191623007|SNOMEDCT_CORE|Bipolar affective disorder, currently manic, severe, with psychosis|Bipolar affective disorder, currently manic, severe, with psychosis
C0338878|T048|FN|191623007|SNOMEDCT_CORE|Bipolar affective disorder, currently manic, severe, with psychosis|Bipolar affective disorder, currently manic, severe, with psychosis
C0338885|T048|PT|191604000|SNOMEDCT_CORE|Single major depressive episode, severe, with psychosis|Single major depressive episode, severe, with psychosis
C0338885|T048|FN|191604000|SNOMEDCT_CORE|Single major depressive episode, severe, with psychosis|Single major depressive episode, severe, with psychosis
C0338908|T048|SY|231504006|SNOMEDCT_CORE|Anxiety depression|Mixed anxiety and depressive disorder
C0338908|T048|PT|231504006|SNOMEDCT_CORE|Mixed anxiety and depressive disorder|Mixed anxiety and depressive disorder
C0338908|T048|FN|231504006|SNOMEDCT_CORE|Mixed anxiety and depressive disorder|Mixed anxiety and depressive disorder
C0338970|T048|PT|191765005|SNOMEDCT_CORE|Emotionally unstable personality disorder|Emotionally unstable personality disorder
C0338970|T048|FN|191765005|SNOMEDCT_CORE|Emotionally unstable personality disorder|Emotionally unstable personality disorder
C0338985|T048|PT|191689008|SNOMEDCT_CORE|Active infantile autism|Active infantile autism
C0338985|T048|FN|191689008|SNOMEDCT_CORE|Active infantile autism|Active infantile autism
C0339002|T048|SY|35253001|SNOMEDCT_CORE|ADD - Attention deficit disorder|Attention deficit hyperactivity disorder, predominantly inattentive type
C0339002|T048|SY|35253001|SNOMEDCT_CORE|ADD - Attention deficit disorder without hyperactivity|Attention deficit hyperactivity disorder, predominantly inattentive type
C0339002|T048|SY|35253001|SNOMEDCT_CORE|Attention deficit disorder|Attention deficit hyperactivity disorder, predominantly inattentive type
C0339002|T048|IS|35253001|SNOMEDCT_CORE|Attention deficit disorder|Attention deficit hyperactivity disorder, predominantly inattentive type
C0339002|T048|SY|35253001|SNOMEDCT_CORE|Attention deficit disorder without hyperactivity|Attention deficit hyperactivity disorder, predominantly inattentive type
C0339002|T048|PT|35253001|SNOMEDCT_CORE|Attention deficit hyperactivity disorder, predominantly inattentive type|Attention deficit hyperactivity disorder, predominantly inattentive type
C0339002|T048|FN|35253001|SNOMEDCT_CORE|Attention deficit hyperactivity disorder, predominantly inattentive type|Attention deficit hyperactivity disorder, predominantly inattentive type
C0339002|T048|SY|35253001|SNOMEDCT_CORE|Attention deficit without hyperactivity|Attention deficit hyperactivity disorder, predominantly inattentive type
C0339052|T037|PT|231791008|SNOMEDCT_CORE|Rupture of globe|Rupture of globe
C0339052|T037|FN|231791008|SNOMEDCT_CORE|Rupture of globe|Rupture of globe
C0339094|T037|FN|231816006|SNOMEDCT_CORE|Laceration of eyelid|Laceration of eyelid
C0339094|T037|PT|231816006|SNOMEDCT_CORE|Laceration of eyelid|Laceration of eyelid
C0339107|T191|PT|231824001|SNOMEDCT_CORE|Benign tumor of eyelid|Benign tumor of eyelid
C0339107|T191|FN|231824001|SNOMEDCT_CORE|Benign tumor of eyelid|Benign tumor of eyelid
C0339107|T191|PTGB|231824001|SNOMEDCT_CORE|Benign tumour of eyelid|Benign tumor of eyelid
C0339114|T191|PT|231832009|SNOMEDCT_CORE|Basal cell carcinoma of eyelid|Basal cell carcinoma of eyelid
C0339114|T191|FN|231832009|SNOMEDCT_CORE|Basal cell carcinoma of eyelid|Basal cell carcinoma of eyelid
C0339114|T191|SY|231832009|SNOMEDCT_CORE|Rodent ulcer of eyelid|Basal cell carcinoma of eyelid
C0339127|T047|SY|231839000|SNOMEDCT_CORE|Blocked tear duct|Complete obstruction of lacrimal canaliculus
C0339127|T047|PT|231839000|SNOMEDCT_CORE|Complete obstruction of lacrimal canaliculus|Complete obstruction of lacrimal canaliculus
C0339127|T047|FN|231839000|SNOMEDCT_CORE|Complete obstruction of lacrimal canaliculus|Complete obstruction of lacrimal canaliculus
C0339127|T047|SY|231839000|SNOMEDCT_CORE|Plugged tear duct|Complete obstruction of lacrimal canaliculus
C0339143|T047|IS|276177000|SNOMEDCT_CORE|Dysthroid orbitopathy|Thyroid eye disease
C0339143|T047|SY|276177000|SNOMEDCT_CORE|Dysthyroid eye disease|Thyroid eye disease
C0339143|T047|SY|276177000|SNOMEDCT_CORE|Dysthyroid orbitopathy|Thyroid eye disease
C0339143|T047|SY|276177000|SNOMEDCT_CORE|Endocrine ophthalmopathy|Thyroid eye disease
C0339143|T047|SY|276177000|SNOMEDCT_CORE|Endocrine orbitopathy|Thyroid eye disease
C0339143|T047|SY|276177000|SNOMEDCT_CORE|Graves eye disease|Thyroid eye disease
C0339143|T047|SY|276177000|SNOMEDCT_CORE|Graves ophthalmopathy|Thyroid eye disease
C0339143|T047|SY|276177000|SNOMEDCT_CORE|Graves' eye disease|Thyroid eye disease
C0339143|T047|SY|276177000|SNOMEDCT_CORE|Graves' ophthalmopathy|Thyroid eye disease
C0339143|T047|SY|276177000|SNOMEDCT_CORE|Ophthalmic Graves disease|Thyroid eye disease
C0339143|T047|PT|276177000|SNOMEDCT_CORE|Thyroid eye disease|Thyroid eye disease
C0339143|T047|FN|276177000|SNOMEDCT_CORE|Thyroid eye disease|Thyroid eye disease
C0339143|T047|SY|276177000|SNOMEDCT_CORE|Thyroid ophthalmopathy|Thyroid eye disease
C0339143|T047|SY|276177000|SNOMEDCT_CORE|Thyroid orbitopathy|Thyroid eye disease
C0339143|T047|SY|276177000|SNOMEDCT_CORE|Thyroid-associated ophthalmopathy|Thyroid eye disease
C0339150|T037|SY|49346003|SNOMEDCT_CORE|Closed blow-out fracture orbit|Closed blow-out fracture orbit
C0339150|T037|SY|49346003|SNOMEDCT_CORE|Closed orbital blow-out fracture|Closed blow-out fracture orbit
C0339164|T047|SY|231855007|SNOMEDCT_CORE|Hay fever conjunctivitis|Seasonal allergic conjunctivitis
C0339164|T047|PT|231855007|SNOMEDCT_CORE|Seasonal allergic conjunctivitis|Seasonal allergic conjunctivitis
C0339164|T047|FN|231855007|SNOMEDCT_CORE|Seasonal allergic conjunctivitis|Seasonal allergic conjunctivitis
C0339177|T037|PT|231866000|SNOMEDCT_CORE|Conjunctival foreign body|Conjunctival foreign body
C0339177|T037|FN|231866000|SNOMEDCT_CORE|Conjunctival foreign body|Conjunctival foreign body
C0339295|T047|SY|14366000|SNOMEDCT_CORE|Exposure keratitis|Exposure keratoconjunctivitis
C0339295|T047|PT|14366000|SNOMEDCT_CORE|Exposure keratoconjunctivitis|Exposure keratoconjunctivitis
C0339295|T047|FN|14366000|SNOMEDCT_CORE|Exposure keratoconjunctivitis|Exposure keratoconjunctivitis
C0339295|T047|SY|14366000|SNOMEDCT_CORE|Exposure keratopathy|Exposure keratoconjunctivitis
C0339295|T047|SY|14366000|SNOMEDCT_CORE|Lagophthalmic keratitis|Exposure keratoconjunctivitis
C0339295|T047|IS|14366000|SNOMEDCT_CORE|lagophthalmic keratitis|Exposure keratoconjunctivitis
C0339303|T047|PT|95742008|SNOMEDCT_CORE|Corneal graft rejection|Corneal graft rejection
C0339303|T047|FN|95742008|SNOMEDCT_CORE|Corneal graft rejection|Corneal graft rejection
C0339352|T047|FN|204125003|SNOMEDCT_CORE|Capsular cataract|Capsular cataract
C0339352|T047|PT|204125003|SNOMEDCT_CORE|Capsular cataract|Capsular cataract
C0339403|T047|OAS|240740001|SNOMEDCT_CORE|Ocular classical histoplasmosis|Presumed ocular histoplasmosis syndrome
C0339403|T047|OP|240740001|SNOMEDCT_CORE|Ocular histoplasmosis syndrome|Presumed ocular histoplasmosis syndrome
C0339403|T047|OAS|240740001|SNOMEDCT_CORE|POHS - Presumed ocular histoplasmosis syndrome|Presumed ocular histoplasmosis syndrome
C0339403|T047|OAP|240740001|SNOMEDCT_CORE|Presumed ocular histoplasmosis syndrome|Presumed ocular histoplasmosis syndrome
C0339403|T047|OAF|240740001|SNOMEDCT_CORE|Presumed ocular histoplasmosis syndrome|Presumed ocular histoplasmosis syndrome
C0339468|T047|PT|232017001|SNOMEDCT_CORE|Anterior proliferative vitreoretinopathy|Anterior proliferative vitreoretinopathy
C0339468|T047|FN|232017001|SNOMEDCT_CORE|Anterior proliferative vitreoretinopathy|Anterior proliferative vitreoretinopathy
C0339469|T047|PT|232018006|SNOMEDCT_CORE|Posterior proliferative vitreoretinopathy|Posterior proliferative vitreoretinopathy
C0339469|T047|FN|232018006|SNOMEDCT_CORE|Posterior proliferative vitreoretinopathy|Posterior proliferative vitreoretinopathy
C0339473|T047|IS|312905005|SNOMEDCT_CORE|Preproliferative diabetic retinopathy|Preproliferative diabetic retinopathy
C0339473|T047|IS|312905005|SNOMEDCT_CORE|Preproliferative retinopathy|Preproliferative diabetic retinopathy
C0339483|T046|PT|95221007|SNOMEDCT_CORE|Radiation retinopathy|Radiation retinopathy
C0339483|T046|FN|95221007|SNOMEDCT_CORE|Radiation retinopathy|Radiation retinopathy
C0339505|T046|SY|24596005|SNOMEDCT_CORE|Branch retinal vein occlusion|Venous retinal branch occlusion
C0339505|T046|SY|24596005|SNOMEDCT_CORE|Branch retinal vein thrombosis|Venous retinal branch occlusion
C0339505|T046|SY|24596005|SNOMEDCT_CORE|BRVO - Branch retinal vein occlusion|Venous retinal branch occlusion
C0339505|T046|SY|24596005|SNOMEDCT_CORE|BRVT - Branch retinal vein thrombosis|Venous retinal branch occlusion
C0339505|T046|SY|24596005|SNOMEDCT_CORE|BVO - Branch retinal occlusion|Venous retinal branch occlusion
C0339505|T046|PT|24596005|SNOMEDCT_CORE|Venous retinal branch occlusion|Venous retinal branch occlusion
C0339505|T046|FN|24596005|SNOMEDCT_CORE|Venous retinal branch occlusion|Venous retinal branch occlusion
C0339505|T046|SY|24596005|SNOMEDCT_CORE|Venous retinal tributary occlusion|Venous retinal branch occlusion
C0339543|T020|SY|367649002|SNOMEDCT_CORE|Cellophane maculopathy|Epiretinal membrane
C0339543|T020|PT|367649002|SNOMEDCT_CORE|Epiretinal membrane|Epiretinal membrane
C0339543|T020|FN|367649002|SNOMEDCT_CORE|Epiretinal membrane|Epiretinal membrane
C0339543|T020|SY|367649002|SNOMEDCT_CORE|ERM - Epiretinal membrane|Epiretinal membrane
C0339543|T020|SY|367649002|SNOMEDCT_CORE|Macular pucker|Epiretinal membrane
C0339543|T020|SY|367649002|SNOMEDCT_CORE|Macular retinal puckering|Epiretinal membrane
C0339543|T020|SY|367649002|SNOMEDCT_CORE|Preretinal fibrosis|Epiretinal membrane
C0339543|T020|SY|367649002|SNOMEDCT_CORE|Preretinal membrane|Epiretinal membrane
C0339555|T019|IS|232074003|SNOMEDCT_CORE|CHRPE - Congenital hypertophy of retinal pigment epithelium|Congenital hypertrophy of retinal pigment epithelium
C0339555|T019|SY|232074003|SNOMEDCT_CORE|CHRPE - Congenital hypertrophy of retinal pigment epithelium|Congenital hypertrophy of retinal pigment epithelium
C0339555|T019|SY|232074003|SNOMEDCT_CORE|Congenital hyperplasia of retinal pigment epithelium|Congenital hypertrophy of retinal pigment epithelium
C0339555|T019|PT|232074003|SNOMEDCT_CORE|Congenital hypertrophy of retinal pigment epithelium|Congenital hypertrophy of retinal pigment epithelium
C0339555|T019|FN|232074003|SNOMEDCT_CORE|Congenital hypertrophy of retinal pigment epithelium|Congenital hypertrophy of retinal pigment epithelium
C0339570|T047|PT|193533000|SNOMEDCT_CORE|Open-angle glaucoma - borderline|Open-angle glaucoma - borderline
C0339570|T047|FN|193533000|SNOMEDCT_CORE|Open-angle glaucoma - borderline|Open-angle glaucoma - borderline
C0339571|T047|PT|193534006|SNOMEDCT_CORE|Angle-closure glaucoma - borderline|Angle-closure glaucoma - borderline
C0339571|T047|FN|193534006|SNOMEDCT_CORE|Angle-closure glaucoma - borderline|Angle-closure glaucoma - borderline
C0339571|T047|SY|193534006|SNOMEDCT_CORE|Borderline angle closure glaucoma|Angle-closure glaucoma - borderline
C0339573|T047|SY|77075001|SNOMEDCT_CORE|Chronic simple glaucoma|Primary open angle glaucoma
C0339573|T047|SY|77075001|SNOMEDCT_CORE|COAG - Chronic open-angle glaucoma|Primary open angle glaucoma
C0339573|T047|SY|77075001|SNOMEDCT_CORE|CSG - Chronic simple glaucoma|Primary open angle glaucoma
C0339573|T047|SY|77075001|SNOMEDCT_CORE|POAG - Primary open-angle glaucoma|Primary open angle glaucoma
C0339573|T047|PT|77075001|SNOMEDCT_CORE|Primary open angle glaucoma|Primary open angle glaucoma
C0339573|T047|FN|77075001|SNOMEDCT_CORE|Primary open angle glaucoma|Primary open angle glaucoma
C0339573|T047|SY|77075001|SNOMEDCT_CORE|Primary open-angle glaucoma|Primary open angle glaucoma
C0339590|T047|SY|392300000|SNOMEDCT_CORE|Lens induced angle closure glaucoma|Phacomorphic glaucoma
C0339590|T047|SY|392300000|SNOMEDCT_CORE|Lens swelling glaucoma|Phacomorphic glaucoma
C0339590|T047|PT|392300000|SNOMEDCT_CORE|Phacomorphic glaucoma|Phacomorphic glaucoma
C0339590|T047|FN|392300000|SNOMEDCT_CORE|Phacomorphic glaucoma|Phacomorphic glaucoma
C0339593|T047|PT|37155002|SNOMEDCT_CORE|Glaucoma associated with ocular inflammation|Glaucoma associated with ocular inflammation
C0339593|T047|FN|37155002|SNOMEDCT_CORE|Glaucoma associated with ocular inflammation|Glaucoma associated with ocular inflammation
C0339593|T047|IS|37155002|SNOMEDCT_CORE|Glaucoma associated with ocular inflammations|Glaucoma associated with ocular inflammation
C0339593|T047|OF|37155002|SNOMEDCT_CORE|Glaucoma associated with ocular inflammations|Glaucoma associated with ocular inflammation
C0339593|T047|SY|37155002|SNOMEDCT_CORE|Glaucoma with ocular inflammation|Glaucoma associated with ocular inflammation
C0339594|T047|PT|68241007|SNOMEDCT_CORE|Glaucoma associated with ocular trauma|Glaucoma associated with ocular trauma
C0339594|T047|FN|68241007|SNOMEDCT_CORE|Glaucoma associated with ocular trauma|Glaucoma associated with ocular trauma
C0339594|T047|SY|68241007|SNOMEDCT_CORE|Glaucoma due to ocular trauma|Glaucoma associated with ocular trauma
C0339594|T047|SY|68241007|SNOMEDCT_CORE|Traumatic glaucoma|Glaucoma associated with ocular trauma
C0339670|T047|SY|72128008|SNOMEDCT_CORE|Disorder of refraction and accommodation|Disorder of refraction AND/OR accommodation
C0339670|T047|IS|72128008|SNOMEDCT_CORE|Disorder of refraction and accommodation, NOS|Disorder of refraction AND/OR accommodation
C0339670|T047|PT|72128008|SNOMEDCT_CORE|Disorder of refraction AND/OR accommodation|Disorder of refraction AND/OR accommodation
C0339670|T047|FN|72128008|SNOMEDCT_CORE|Disorder of refraction AND/OR accommodation|Disorder of refraction AND/OR accommodation
C0339696|T047|PT|232147001|SNOMEDCT_CORE|Anisometropic amblyopia|Anisometropic amblyopia
C0339696|T047|FN|232147001|SNOMEDCT_CORE|Anisometropic amblyopia|Anisometropic amblyopia
C0339711|T033|PT|193731001|SNOMEDCT_CORE|Legal blindness USA|Legal blindness USA
C0339711|T033|OF|193731001|SNOMEDCT_CORE|Legal blindness USA|Legal blindness USA
C0339753|T047|OAP|95806007|SNOMEDCT_CORE|Cellulitis of external ear|Cellulitis of external ear
C0339753|T047|OAF|95806007|SNOMEDCT_CORE|Cellulitis of external ear|Cellulitis of external ear
C0339767|T047|SY|38394007|SNOMEDCT_CORE|Chronic otitis media with perforation|Chronic otitis media with perforation
C0339804|T047|SY|232345000|SNOMEDCT_CORE|NINA - Non-infective non-allergic rhinitis|Non-infective non-allergic rhinitis
C0339804|T047|PT|232345000|SNOMEDCT_CORE|Non-infective non-allergic rhinitis|Non-infective non-allergic rhinitis
C0339804|T047|FN|232345000|SNOMEDCT_CORE|Non-infective non-allergic rhinitis|Non-infective non-allergic rhinitis
C0339808|T047|PT|232350006|SNOMEDCT_CORE|Allergy to dust mite protein|Allergy to dust mite protein
C0339808|T047|FN|232350006|SNOMEDCT_CORE|Allergy to dust mite protein|Allergy to dust mite protein
C0339808|T047|SY|232350006|SNOMEDCT_CORE|Allergy to house dust mite|Allergy to dust mite protein
C0339808|T047|OF|232350006|SNOMEDCT_CORE|Allergy to house dust mite|Allergy to dust mite protein
C0339808|T047|SY|232350006|SNOMEDCT_CORE|House dust mite allergy|Allergy to dust mite protein
C0339808|T047|OF|232350006|SNOMEDCT_CORE|House dust mite allergy|Allergy to dust mite protein
C0339820|T047|PT|232340005|SNOMEDCT_CORE|Disorder of nasal cavity|Disorder of nasal cavity
C0339820|T047|FN|232340005|SNOMEDCT_CORE|Disorder of nasal cavity|Disorder of nasal cavity
C0339825|T047|PT|23714000|SNOMEDCT_CORE|Nasal vestibulitis|Nasal vestibulitis
C0339825|T047|FN|23714000|SNOMEDCT_CORE|Nasal vestibulitis|Nasal vestibulitis
C0339825|T047|IS|23714000|SNOMEDCT_CORE|Nasal vestibulitis, NOS|Nasal vestibulitis
C0339848|T037|SY|263171005|SNOMEDCT_CORE|Broken nose|Fractured nasal bones
C0339848|T037|SY|263171005|SNOMEDCT_CORE|Fracture of nasal bones|Fractured nasal bones
C0339848|T037|SY|263171005|SNOMEDCT_CORE|Fracture of nasal complex|Fractured nasal bones
C0339848|T037|SY|263171005|SNOMEDCT_CORE|Fracture of nose|Fractured nasal bones
C0339848|T037|PT|263171005|SNOMEDCT_CORE|Fractured nasal bones|Fractured nasal bones
C0339848|T037|FN|263171005|SNOMEDCT_CORE|Fractured nasal bones|Fractured nasal bones
C0339848|T037|SY|263171005|SNOMEDCT_CORE|Fractured nose|Fractured nasal bones
C0339868|T047|SY|195677001|SNOMEDCT_CORE|RAT - Recurrent acute tonsillitis|Recurrent acute tonsillitis
C0339868|T047|PT|195677001|SNOMEDCT_CORE|Recurrent acute tonsillitis|Recurrent acute tonsillitis
C0339868|T047|FN|195677001|SNOMEDCT_CORE|Recurrent acute tonsillitis|Recurrent acute tonsillitis
C0339982|T047|PT|195984007|SNOMEDCT_CORE|Recurrent bronchiectasis|Recurrent bronchiectasis
C0339982|T047|FN|195984007|SNOMEDCT_CORE|Recurrent bronchiectasis|Recurrent bronchiectasis
C0340025|T047|PT|233659006|SNOMEDCT_CORE|Asbestos-induced pleural plaque|Asbestos-induced pleural plaque
C0340025|T047|FN|233659006|SNOMEDCT_CORE|Asbestos-induced pleural plaque|Asbestos-induced pleural plaque
C0340025|T047|IS|233659006|SNOMEDCT_CORE|Pleural plaque disease due to asbestosis|Asbestos-induced pleural plaque
C0340044|T047|PT|195951007|SNOMEDCT_CORE|Acute exacerbation of chronic obstructive airways disease|Acute exacerbation of chronic obstructive airways disease
C0340044|T047|FN|195951007|SNOMEDCT_CORE|Acute exacerbation of chronic obstructive airways disease|Acute exacerbation of chronic obstructive airways disease
C0340044|T047|SY|195951007|SNOMEDCT_CORE|Acute exacerbation of chronic obstructive pulmonary disease|Acute exacerbation of chronic obstructive airways disease
C0340044|T047|SY|195951007|SNOMEDCT_CORE|Acute exacerbation of COPD|Acute exacerbation of chronic obstructive airways disease
C0340050|T047|PT|233674008|SNOMEDCT_CORE|Pulmonary emphysema in alpha-1 PI deficiency|Pulmonary emphysema in alpha-1 PI deficiency
C0340050|T047|OF|233674008|SNOMEDCT_CORE|Pulmonary emphysema in alpha-1 PI deficiency|Pulmonary emphysema in alpha-1 PI deficiency
C0340050|T047|FN|233674008|SNOMEDCT_CORE|Pulmonary emphysema in alpha-1 primary immunodeficiency deficiency|Pulmonary emphysema in alpha-1 PI deficiency
C0340050|T047|SY|233674008|SNOMEDCT_CORE|Pulmonary emphysema in alpha-1 primary immunodeficiency deficiency|Pulmonary emphysema in alpha-1 PI deficiency
C0340062|T047|SY|195967001|SNOMEDCT_CORE|Hyperreactive airway disease|Hyperreactive airway disease
C0340145|T047|SY|196033004|SNOMEDCT_CORE|Pneumonitis caused by inhalation of regurgitated food|Pneumonitis due to inhalation of regurgitated food
C0340145|T047|FN|196033004|SNOMEDCT_CORE|Pneumonitis caused by inhalation of regurgitated food|Pneumonitis due to inhalation of regurgitated food
C0340145|T047|PT|196033004|SNOMEDCT_CORE|Pneumonitis due to inhalation of regurgitated food|Pneumonitis due to inhalation of regurgitated food
C0340145|T047|OF|196033004|SNOMEDCT_CORE|Pneumonitis due to inhalation of regurgitated food|Pneumonitis due to inhalation of regurgitated food
C0340194|T047|IS|233765002|SNOMEDCT_CORE|Hypoxemic respiratory failure|Respiratory failure without hypercapnia
C0340194|T047|PT|233765002|SNOMEDCT_CORE|Respiratory failure without hypercapnia|Respiratory failure without hypercapnia
C0340194|T047|FN|233765002|SNOMEDCT_CORE|Respiratory failure without hypercapnia|Respiratory failure without hypercapnia
C0340194|T047|SY|233765002|SNOMEDCT_CORE|Type 1 respiratory failure|Respiratory failure without hypercapnia
C0340194|T047|SY|233765002|SNOMEDCT_CORE|Type I respiratory failure|Respiratory failure without hypercapnia
C0340276|T046|PT|233816003|SNOMEDCT_CORE|Postoperative cardiac complication|Postoperative cardiac complication
C0340276|T046|FN|233816003|SNOMEDCT_CORE|Postoperative cardiac complication|Postoperative cardiac complication
C0340279|T047|PT|266249003|SNOMEDCT_CORE|Ventricular hypertrophy|Ventricular hypertrophy
C0340279|T047|FN|266249003|SNOMEDCT_CORE|Ventricular hypertrophy|Ventricular hypertrophy
C0340285|T047|SY|233817007|SNOMEDCT_CORE|Triple vessel coronary artery disease|Triple vessel disease of the heart
C0340285|T047|PT|233817007|SNOMEDCT_CORE|Triple vessel disease of the heart|Triple vessel disease of the heart
C0340285|T047|FN|233817007|SNOMEDCT_CORE|Triple vessel disease of the heart|Triple vessel disease of the heart
C0340288|T047|PT|233819005|SNOMEDCT_CORE|Stable angina|Stable angina
C0340288|T047|FN|233819005|SNOMEDCT_CORE|Stable angina|Stable angina
C0340311|T047|SY|58612006|SNOMEDCT_CORE|Acute lateral myocardial infarction|Acute myocardial infarction of lateral wall
C0340311|T047|PT|58612006|SNOMEDCT_CORE|Acute myocardial infarction of lateral wall|Acute myocardial infarction of lateral wall
C0340311|T047|FN|58612006|SNOMEDCT_CORE|Acute myocardial infarction of lateral wall|Acute myocardial infarction of lateral wall
C0340318|T047|PT|233838001|SNOMEDCT_CORE|Acute posterior myocardial infarction|Acute posterior myocardial infarction
C0340318|T047|FN|233838001|SNOMEDCT_CORE|Acute posterior myocardial infarction|Acute posterior myocardial infarction
C0340320|T047|PT|233839009|SNOMEDCT_CORE|Old anterior myocardial infarction|Old anterior myocardial infarction
C0340320|T047|FN|233839009|SNOMEDCT_CORE|Old anterior myocardial infarction|Old anterior myocardial infarction
C0340326|T047|PT|233844002|SNOMEDCT_CORE|Accelerated coronary artery disease in transplanted heart|Accelerated coronary artery disease in transplanted heart
C0340326|T047|FN|233844002|SNOMEDCT_CORE|Accelerated coronary artery disease in transplanted heart|Accelerated coronary artery disease in transplanted heart
C0340362|T047|SY|194978002|SNOMEDCT_CORE|Mitral incompetence, non-rheumatic|Non-rheumatic mitral regurgitation
C0340362|T047|PT|194978002|SNOMEDCT_CORE|Non-rheumatic mitral regurgitation|Non-rheumatic mitral regurgitation
C0340362|T047|FN|194978002|SNOMEDCT_CORE|Non-rheumatic mitral regurgitation|Non-rheumatic mitral regurgitation
C0340372|T047|PT|194984004|SNOMEDCT_CORE|Aortic stenosis, non-rheumatic|Aortic stenosis, non-rheumatic
C0340372|T047|FN|194984004|SNOMEDCT_CORE|Aortic stenosis, non-rheumatic|Aortic stenosis, non-rheumatic
C0340377|T047|PT|194983005|SNOMEDCT_CORE|Aortic incompetence, non-rheumatic|Aortic incompetence, non-rheumatic
C0340377|T047|FN|194983005|SNOMEDCT_CORE|Aortic incompetence, non-rheumatic|Aortic incompetence, non-rheumatic
C0340377|T047|SY|194983005|SNOMEDCT_CORE|Aortic insufficiency, non-rheumatic|Aortic incompetence, non-rheumatic
C0340377|T047|SY|194983005|SNOMEDCT_CORE|Aortic regurgitation, non-rheumatic|Aortic incompetence, non-rheumatic
C0340377|T047|SY|194983005|SNOMEDCT_CORE|Aortic valve regurgitation, nonrheumatic|Aortic incompetence, non-rheumatic
C0340389|T047|PT|194990000|SNOMEDCT_CORE|Tricuspid incompetence, non-rheumatic|Tricuspid incompetence, non-rheumatic
C0340389|T047|FN|194990000|SNOMEDCT_CORE|Tricuspid incompetence, non-rheumatic|Tricuspid incompetence, non-rheumatic
C0340389|T047|SY|194990000|SNOMEDCT_CORE|Tricuspid insufficiency, non-rheumatic|Tricuspid incompetence, non-rheumatic
C0340389|T047|SY|194990000|SNOMEDCT_CORE|Tricuspid regurgitation, non-rheumatic|Tricuspid incompetence, non-rheumatic
C0340389|T047|SY|194990000|SNOMEDCT_CORE|Tricuspid valve regurgitation, nonrheumatic|Tricuspid incompetence, non-rheumatic
C0340395|T047|PT|194997002|SNOMEDCT_CORE|Pulmonary stenosis, non-rheumatic|Pulmonary stenosis, non-rheumatic
C0340395|T047|FN|194997002|SNOMEDCT_CORE|Pulmonary stenosis, non-rheumatic|Pulmonary stenosis, non-rheumatic
C0340395|T047|SY|194997002|SNOMEDCT_CORE|Pulmonary valve stenosis, nonrheumatic|Pulmonary stenosis, non-rheumatic
C0340464|T047|IS|29717002|SNOMEDCT_CORE|Ectopic beats|Ectopic beats
C0340464|T047|PT|33413000|SNOMEDCT_CORE|Ectopic beats|Ectopic beats
C0340464|T047|FN|33413000|SNOMEDCT_CORE|Ectopic beats|Ectopic beats
C0340464|T047|SY|29717002|SNOMEDCT_CORE|Ectopics|Ectopic beats
C0340464|T047|SY|29717002|SNOMEDCT_CORE|Extrasystoles|Ectopic beats
C0340464|T047|SY|29717002|SNOMEDCT_CORE|Extrasystolic arrhythmia|Ectopic beats
C0340464|T047|PT|29717002|SNOMEDCT_CORE|Premature beats|Ectopic beats
C0340464|T047|FN|29717002|SNOMEDCT_CORE|Premature beats|Ectopic beats
C0340464|T047|IS|29717002|SNOMEDCT_CORE|Premature beats, NOS|Ectopic beats
C0340514|T047|PT|233927002|SNOMEDCT_CORE|Cardiac arrest with successful resuscitation|Cardiac arrest with successful resuscitation
C0340514|T047|FN|233927002|SNOMEDCT_CORE|Cardiac arrest with successful resuscitation|Cardiac arrest with successful resuscitation
C0340517|T047|PT|195147006|SNOMEDCT_CORE|Atrial thrombosis|Atrial thrombosis
C0340517|T047|FN|195147006|SNOMEDCT_CORE|Atrial thrombosis|Atrial thrombosis
C0340557|T047|SY|302910002|SNOMEDCT_CORE|ARAS - Atherosclerotic renal artery stenosis|Atherosclerotic renal artery stenosis
C0340557|T047|PT|302910002|SNOMEDCT_CORE|Atherosclerotic renal artery stenosis|Atherosclerotic renal artery stenosis
C0340557|T047|FN|302910002|SNOMEDCT_CORE|Atherosclerotic renal artery stenosis|Atherosclerotic renal artery stenosis
C0340566|T047|PTGB|233962007|SNOMEDCT_CORE|Critical lower limb ischaemia|Critical lower limb ischemia
C0340566|T047|PT|233962007|SNOMEDCT_CORE|Critical lower limb ischemia|Critical lower limb ischemia
C0340566|T047|FN|233962007|SNOMEDCT_CORE|Critical lower limb ischemia|Critical lower limb ischemia
C0340630|T047|PT|233984007|SNOMEDCT_CORE|Thoracoabdominal aortic aneurysm|Thoracoabdominal aortic aneurysm
C0340630|T047|FN|233984007|SNOMEDCT_CORE|Thoracoabdominal aortic aneurysm|Thoracoabdominal aortic aneurysm
C0340639|T047|SY|233988005|SNOMEDCT_CORE|Aneurysm of carotid artery|Carotid artery aneurysm
C0340639|T047|PT|233988005|SNOMEDCT_CORE|Carotid artery aneurysm|Carotid artery aneurysm
C0340639|T047|FN|233988005|SNOMEDCT_CORE|Carotid artery aneurysm|Carotid artery aneurysm
C0340643|T047|IS|308546005|SNOMEDCT_CORE|Dissecting aneurysm of aorta|Dissection of aorta
C0340643|T047|PT|308546005|SNOMEDCT_CORE|Dissection of aorta|Dissection of aorta
C0340643|T047|FN|308546005|SNOMEDCT_CORE|Dissection of aorta|Dissection of aorta
C0340644|T047|IS|233994002|SNOMEDCT_CORE|Dissecting aneurysm of thoracic aorta|Dissection of thoracic aorta
C0340644|T047|PT|233994002|SNOMEDCT_CORE|Dissection of thoracic aorta|Dissection of thoracic aorta
C0340644|T047|FN|233994002|SNOMEDCT_CORE|Dissection of thoracic aorta|Dissection of thoracic aorta
C0340704|T047|SY|197001004|SNOMEDCT_CORE|Deep venous thrombosis of the superior mesenteric vein|Superior mesenteric vein thrombosis
C0340704|T047|PT|197001004|SNOMEDCT_CORE|Superior mesenteric vein thrombosis|Superior mesenteric vein thrombosis
C0340704|T047|FN|197001004|SNOMEDCT_CORE|Superior mesenteric vein thrombosis|Superior mesenteric vein thrombosis
C0340708|T047|SY|404223003|SNOMEDCT_CORE|Deep vein thrombosis of lower limb|Deep venous thrombosis of lower extremity
C0340708|T047|SY|404223003|SNOMEDCT_CORE|Deep venous thrombosis of leg|Deep venous thrombosis of lower extremity
C0340708|T047|PT|404223003|SNOMEDCT_CORE|Deep venous thrombosis of lower extremity|Deep venous thrombosis of lower extremity
C0340708|T047|FN|404223003|SNOMEDCT_CORE|Deep venous thrombosis of lower extremity|Deep venous thrombosis of lower extremity
C0340708|T047|SY|404223003|SNOMEDCT_CORE|Deep venous thrombosis of lower limb|Deep venous thrombosis of lower extremity
C0340708|T047|SY|404223003|SNOMEDCT_CORE|DVT - Deep vein thrombosis of lower limb|Deep venous thrombosis of lower extremity
C0340858|T046|PT|234171009|SNOMEDCT_CORE|Drug-induced hypotension|Drug-induced hypotension
C0340858|T046|FN|234171009|SNOMEDCT_CORE|Drug-induced hypotension|Drug-induced hypotension
C0340858|T046|SY|234171009|SNOMEDCT_CORE|Hypotension due to drugs|Drug-induced hypotension
C0340914|T047|PT|271983002|SNOMEDCT_CORE|Disorder of cardiac pacemaker system|Disorder of cardiac pacemaker system
C0340914|T047|FN|271983002|SNOMEDCT_CORE|Disorder of cardiac pacemaker system|Disorder of cardiac pacemaker system
C0340933|T047|SY|234228008|SNOMEDCT_CORE|Disorder of implantable cardiovertor|Disorder of implantable defibrillator
C0340933|T047|PT|234228008|SNOMEDCT_CORE|Disorder of implantable defibrillator|Disorder of implantable defibrillator
C0340933|T047|FN|234228008|SNOMEDCT_CORE|Disorder of implantable defibrillator|Disorder of implantable defibrillator
C0340933|T047|SY|234228008|SNOMEDCT_CORE|ICD - Disorder of implantable cardiac defibrillator|Disorder of implantable defibrillator
C0341106|T047|PT|235599003|SNOMEDCT_CORE|Eosinophilic esophagitis|Eosinophilic esophagitis
C0341106|T047|FN|235599003|SNOMEDCT_CORE|Eosinophilic esophagitis|Eosinophilic esophagitis
C0341106|T047|PTGB|235599003|SNOMEDCT_CORE|Eosinophilic oesophagitis|Eosinophilic esophagitis
C0341164|T047|SY|15902003|SNOMEDCT_CORE|Bleeding gastric ulcer|Gastric ulcer with hemorrhage
C0341164|T047|PTGB|15902003|SNOMEDCT_CORE|Gastric ulcer with haemorrhage|Gastric ulcer with hemorrhage
C0341164|T047|PT|15902003|SNOMEDCT_CORE|Gastric ulcer with hemorrhage|Gastric ulcer with hemorrhage
C0341164|T047|FN|15902003|SNOMEDCT_CORE|Gastric ulcer with hemorrhage|Gastric ulcer with hemorrhage
C0341164|T047|IS|15902003|SNOMEDCT_CORE|Gastric ulcer, NOS with hemorrhage|Gastric ulcer with hemorrhage
C0341165|T047|PT|95529005|SNOMEDCT_CORE|Acute gastric ulcer|Acute gastric ulcer
C0341165|T047|FN|95529005|SNOMEDCT_CORE|Acute gastric ulcer|Acute gastric ulcer
C0341165|T047|IS|95529005|SNOMEDCT_CORE|Acute gastric ulcer, NOS|Acute gastric ulcer
C0341165|T047|SY|95529005|SNOMEDCT_CORE|Acute ulcer of stomach|Acute gastric ulcer
C0341165|T047|IS|95529005|SNOMEDCT_CORE|Acute ulcer of stomach, NOS|Acute gastric ulcer
C0341168|T047|SY|95529005|SNOMEDCT_CORE|Acute peptic ulcer of stomach|Acute peptic ulcer of stomach
C0341172|T047|PT|95530000|SNOMEDCT_CORE|Chronic gastric ulcer|Chronic gastric ulcer
C0341172|T047|FN|95530000|SNOMEDCT_CORE|Chronic gastric ulcer|Chronic gastric ulcer
C0341172|T047|IS|95530000|SNOMEDCT_CORE|Chronic gastric ulcer, NOS|Chronic gastric ulcer
C0341172|T047|SY|95530000|SNOMEDCT_CORE|Chronic ulcer of stomach|Chronic gastric ulcer
C0341172|T047|IS|95530000|SNOMEDCT_CORE|Chronic ulcer of stomach, NOS|Chronic gastric ulcer
C0341175|T047|SY|95530000|SNOMEDCT_CORE|Chronic peptic ulcer of stomach|Chronic peptic ulcer of stomach
C0341201|T047|PT|196757008|SNOMEDCT_CORE|Drug-induced gastrointestinal disturbance|Drug-induced gastrointestinal disturbance
C0341201|T047|FN|196757008|SNOMEDCT_CORE|Drug-induced gastrointestinal disturbance|Drug-induced gastrointestinal disturbance
C0341217|T047|SY|109558001|SNOMEDCT_CORE|Caliber persistent artery|Dieulafoy's vascular malformation
C0341217|T047|SYGB|109558001|SNOMEDCT_CORE|Calibre persistent artery|Dieulafoy's vascular malformation
C0341217|T047|SY|109558001|SNOMEDCT_CORE|Dieulafoy disease|Dieulafoy's vascular malformation
C0341217|T047|SY|109558001|SNOMEDCT_CORE|Dieulafoy vascular malformation|Dieulafoy's vascular malformation
C0341217|T047|PT|109558001|SNOMEDCT_CORE|Dieulafoy's vascular malformation|Dieulafoy's vascular malformation
C0341217|T047|FN|109558001|SNOMEDCT_CORE|Dieulafoy's vascular malformation|Dieulafoy's vascular malformation
C0341233|T047|PT|196652006|SNOMEDCT_CORE|Acute duodenal ulcer|Acute duodenal ulcer
C0341233|T047|FN|196652006|SNOMEDCT_CORE|Acute duodenal ulcer|Acute duodenal ulcer
C0341233|T047|SY|196652006|SNOMEDCT_CORE|ADU - Acute duodenal ulcer|Acute duodenal ulcer
C0341236|T047|SY|196652006|SNOMEDCT_CORE|Acute peptic ulcer of duodenum|Acute peptic ulcer of duodenum
C0341240|T047|PT|128286008|SNOMEDCT_CORE|Chronic duodenal ulcer|Chronic duodenal ulcer
C0341240|T047|FN|128286008|SNOMEDCT_CORE|Chronic duodenal ulcer|Chronic duodenal ulcer
C0341243|T047|SY|128286008|SNOMEDCT_CORE|Chronic peptic ulcer of duodenum|Chronic peptic ulcer of duodenum
C0341245|T047|IS|95531001|SNOMEDCT_CORE|Acute duodenitis|Hemorrhagic duodenitis
C0341245|T047|SY|95531001|SNOMEDCT_CORE|Erosive duodenitis|Hemorrhagic duodenitis
C0341245|T047|PTGB|95531001|SNOMEDCT_CORE|Haemorrhagic duodenitis|Hemorrhagic duodenitis
C0341245|T047|PT|95531001|SNOMEDCT_CORE|Hemorrhagic duodenitis|Hemorrhagic duodenitis
C0341245|T047|FN|95531001|SNOMEDCT_CORE|Hemorrhagic duodenitis|Hemorrhagic duodenitis
C0341247|T033|SY|95531001|SNOMEDCT_CORE|Multiple duodenal erosions|Multiple duodenal erosions
C0341318|T190|SY|197247001|SNOMEDCT_CORE|Enteric cutaneous fistula|Enterocutaneous fistula
C0341318|T190|PT|197247001|SNOMEDCT_CORE|Enterocutaneous fistula|Enterocutaneous fistula
C0341318|T190|FN|197247001|SNOMEDCT_CORE|Enterocutaneous fistula|Enterocutaneous fistula
C0341379|T190|PT|197155003|SNOMEDCT_CORE|Intersphincteric fistula|Intersphincteric fistula
C0341379|T190|FN|197155003|SNOMEDCT_CORE|Intersphincteric fistula|Intersphincteric fistula
C0341379|T190|SY|197155003|SNOMEDCT_CORE|Submucosal anal fistula|Intersphincteric fistula
C0341379|T190|SY|197155003|SNOMEDCT_CORE|Superficial anal fistula|Intersphincteric fistula
C0341395|T047|SY|235796008|SNOMEDCT_CORE|Perianal Crohn disease|Perianal Crohn's disease
C0341395|T047|PT|235796008|SNOMEDCT_CORE|Perianal Crohn's disease|Perianal Crohn's disease
C0341395|T047|FN|235796008|SNOMEDCT_CORE|Perianal Crohn's disease|Perianal Crohn's disease
C0341539|T020|PT|236048007|SNOMEDCT_CORE|Parastomal hernia|Parastomal hernia
C0341539|T020|FN|236048007|SNOMEDCT_CORE|Parastomal hernia|Parastomal hernia
C0341582|T047|PT|236104004|SNOMEDCT_CORE|Gastrointestinal anastomotic stricture|Gastrointestinal anastomotic stricture
C0341582|T047|FN|236104004|SNOMEDCT_CORE|Gastrointestinal anastomotic stricture|Gastrointestinal anastomotic stricture
C0341591|T046|PT|302918009|SNOMEDCT_CORE|Disorder of stoma|Disorder of stoma
C0341591|T046|FN|302918009|SNOMEDCT_CORE|Disorder of stoma|Disorder of stoma
C0341594|T047|SY|236117001|SNOMEDCT_CORE|Recession of stoma|Retraction of stoma
C0341594|T047|PT|236117001|SNOMEDCT_CORE|Retraction of stoma|Retraction of stoma
C0341594|T047|FN|236117001|SNOMEDCT_CORE|Retraction of stoma|Retraction of stoma
C0341601|T047|PT|236125004|SNOMEDCT_CORE|Peristomal dermatitis|Peristomal dermatitis
C0341601|T047|FN|236125004|SNOMEDCT_CORE|Peristomal dermatitis|Peristomal dermatitis
C0341601|T047|SY|236125004|SNOMEDCT_CORE|Peristomal eczema|Peristomal dermatitis
C0341677|T047|PT|197663003|SNOMEDCT_CORE|Impaired renal function disorder|Impaired renal function disorder
C0341677|T047|FN|197663003|SNOMEDCT_CORE|Impaired renal function disorder|Impaired renal function disorder
C0341687|T047|PT|197604006|SNOMEDCT_CORE|Nephrotic syndrome in amyloidosis|Nephrotic syndrome in amyloidosis
C0341687|T047|FN|197604006|SNOMEDCT_CORE|Nephrotic syndrome in amyloidosis|Nephrotic syndrome in amyloidosis
C0341698|T047|PT|197659005|SNOMEDCT_CORE|Atrophy of kidney|Atrophy of kidney
C0341698|T047|FN|197659005|SNOMEDCT_CORE|Atrophy of kidney|Atrophy of kidney
C0341698|T047|SY|197659005|SNOMEDCT_CORE|Renal atrophy|Atrophy of kidney
C0341740|T191|IS|236646007|SNOMEDCT_CORE|Benign prostatic hypertroph with outflow obstruction|Benign prostatic hypertrophy with outflow obstruction
C0341740|T191|OF|236646007|SNOMEDCT_CORE|Benign prostatic hypertroph with outflow obstruction|Benign prostatic hypertrophy with outflow obstruction
C0341740|T191|PT|236646007|SNOMEDCT_CORE|Benign prostatic hypertrophy with outflow obstruction|Benign prostatic hypertrophy with outflow obstruction
C0341740|T191|FN|236646007|SNOMEDCT_CORE|Benign prostatic hypertrophy with outflow obstruction|Benign prostatic hypertrophy with outflow obstruction
C0341741|T019|SY|268236002|SNOMEDCT_CORE|Bladder neck stenosis|Congenital bladder neck stenosis
C0341741|T019|SY|268236002|SNOMEDCT_CORE|BNS - Bladder neck stenosis|Congenital bladder neck stenosis
C0341741|T019|PT|268236002|SNOMEDCT_CORE|Congenital bladder neck stenosis|Congenital bladder neck stenosis
C0341741|T019|FN|268236002|SNOMEDCT_CORE|Congenital bladder neck stenosis|Congenital bladder neck stenosis
C0341741|T019|IS|268236002|SNOMEDCT_CORE|Contracture of bladder neck|Congenital bladder neck stenosis
C0341742|T184|PT|236648008|SNOMEDCT_CORE|Acute retention of urine|Acute retention of urine
C0341742|T184|FN|236648008|SNOMEDCT_CORE|Acute retention of urine|Acute retention of urine
C0341742|T184|SY|236648008|SNOMEDCT_CORE|Acute urinary retention|Acute retention of urine
C0341742|T184|SY|236648008|SNOMEDCT_CORE|ARU - Acute retention of urine|Acute retention of urine
C0341743|T046|PT|236650000|SNOMEDCT_CORE|Chronic retention of urine|Chronic retention of urine
C0341743|T046|FN|236650000|SNOMEDCT_CORE|Chronic retention of urine|Chronic retention of urine
C0341743|T046|SY|236650000|SNOMEDCT_CORE|CRU - Chronic retention of urine|Chronic retention of urine
C0341834|T047|PT|237084006|SNOMEDCT_CORE|Chlamydial cervicitis|Chlamydial cervicitis
C0341834|T047|FN|237084006|SNOMEDCT_CORE|Chlamydial cervicitis|Chlamydial cervicitis
C0341858|T047|IS|76376003|SNOMEDCT_CORE|Adenomyosis|Endometriosis of uterus
C0341858|T047|IS|76376003|SNOMEDCT_CORE|Adenomyosis uteri|Endometriosis of uterus
C0341858|T047|IS|76376003|SNOMEDCT_CORE|Endometriosis of myometrium|Endometriosis of uterus
C0341858|T047|PT|76376003|SNOMEDCT_CORE|Endometriosis of uterus|Endometriosis of uterus
C0341858|T047|FN|76376003|SNOMEDCT_CORE|Endometriosis of uterus|Endometriosis of uterus
C0341858|T047|IS|76376003|SNOMEDCT_CORE|Endometriosis of uterus, NOS|Endometriosis of uterus
C0341858|T047|SY|76376003|SNOMEDCT_CORE|Internal endometriosis|Endometriosis of uterus
C0341863|T046|SY|266601003|SNOMEDCT_CORE|Epimenorrhagia|Excessive and frequent menstruation
C0341863|T046|PT|266601003|SNOMEDCT_CORE|Excessive and frequent menstruation|Excessive and frequent menstruation
C0341863|T046|FN|266601003|SNOMEDCT_CORE|Excessive and frequent menstruation|Excessive and frequent menstruation
C0341863|T046|SY|266601003|SNOMEDCT_CORE|Frequent heavy periods|Excessive and frequent menstruation
C0341863|T046|SY|266601003|SNOMEDCT_CORE|Hyperpolymenorrhea|Excessive and frequent menstruation
C0341863|T046|SY|266601003|SNOMEDCT_CORE|Hyperpolymenorrhoea|Excessive and frequent menstruation
C0341863|T046|SY|266601003|SNOMEDCT_CORE|Polymenorrhagia|Excessive and frequent menstruation
C0341868|T047|PT|237138004|SNOMEDCT_CORE|Menopause ovarian failure|Menopause ovarian failure
C0341868|T047|FN|237138004|SNOMEDCT_CORE|Menopause ovarian failure|Menopause ovarian failure
C0341934|T046|PT|237279007|SNOMEDCT_CORE|Transient hypertension of pregnancy|Transient hypertension of pregnancy
C0341934|T046|FN|237279007|SNOMEDCT_CORE|Transient hypertension of pregnancy|Transient hypertension of pregnancy
C0341950|T046|SYGB|46764007|SNOMEDCT_CORE|PET - Severe pre-eclamptic toxaemia|Severe pre-eclampsia
C0341950|T046|SY|46764007|SNOMEDCT_CORE|PET - Severe pre-eclamptic toxemia|Severe pre-eclampsia
C0341950|T046|IS|46764007|SNOMEDCT_CORE|Severe edema|Severe pre-eclampsia
C0341950|T046|IS|46764007|SNOMEDCT_CORE|Severe oedema|Severe pre-eclampsia
C0341950|T046|PT|46764007|SNOMEDCT_CORE|Severe pre-eclampsia|Severe pre-eclampsia
C0341950|T046|FN|46764007|SNOMEDCT_CORE|Severe pre-eclampsia|Severe pre-eclampsia
C0341950|T046|SYGB|46764007|SNOMEDCT_CORE|Severe pre-eclamptic toxaemia|Severe pre-eclampsia
C0341950|T046|SY|46764007|SNOMEDCT_CORE|Severe pre-eclamptic toxemia|Severe pre-eclampsia
C0341950|T046|SY|46764007|SNOMEDCT_CORE|Severe proteinuric hypertension of pregnancy|Severe pre-eclampsia
C0341950|T046|IS|46764007|SNOMEDCT_CORE|Severe proteinuric hypertension of pregnancy|Severe pre-eclampsia
C0341973|T046|SY|267340006|SNOMEDCT_CORE|Maternal pyrexia during labor|Maternal pyrexia in labor
C0341973|T046|SYGB|267340006|SNOMEDCT_CORE|Maternal pyrexia during labour|Maternal pyrexia in labor
C0341973|T046|PT|267340006|SNOMEDCT_CORE|Maternal pyrexia in labor|Maternal pyrexia in labor
C0341973|T046|FN|267340006|SNOMEDCT_CORE|Maternal pyrexia in labor|Maternal pyrexia in labor
C0341973|T046|PTGB|267340006|SNOMEDCT_CORE|Maternal pyrexia in labour|Maternal pyrexia in labor
C0342115|T047|SY|190237002|SNOMEDCT_CORE|Non-toxic single thyroid nodule|Non-toxic uninodular goiter
C0342115|T047|FN|190237002|SNOMEDCT_CORE|Non-toxic uninodular goiter|Non-toxic uninodular goiter
C0342115|T047|PT|190237002|SNOMEDCT_CORE|Non-toxic uninodular goiter|Non-toxic uninodular goiter
C0342115|T047|PTGB|190237002|SNOMEDCT_CORE|Non-toxic uninodular goitre|Non-toxic uninodular goiter
C0342115|T047|SY|190237002|SNOMEDCT_CORE|Nontoxic uninodular thyroid goiter|Non-toxic uninodular goiter
C0342115|T047|SYGB|190237002|SNOMEDCT_CORE|Nontoxic uninodular thyroid goitre|Non-toxic uninodular goiter
C0342117|T020|SY|237496006|SNOMEDCT_CORE|Colloid nodule|Thyroid colloid nodule
C0342117|T020|PT|237496006|SNOMEDCT_CORE|Thyroid colloid nodule|Thyroid colloid nodule
C0342117|T020|FN|237496006|SNOMEDCT_CORE|Thyroid colloid nodule|Thyroid colloid nodule
C0342122|T047|SY|267374005|SNOMEDCT_CORE|Diffuse toxic goiter|Toxic diffuse goiter
C0342122|T047|SYGB|267374005|SNOMEDCT_CORE|Diffuse toxic goitre|Toxic diffuse goiter
C0342122|T047|SY|267374005|SNOMEDCT_CORE|Thyrotoxicosis with diffuse goiter|Toxic diffuse goiter
C0342122|T047|SYGB|267374005|SNOMEDCT_CORE|Thyrotoxicosis with diffuse goitre|Toxic diffuse goiter
C0342122|T047|PT|267374005|SNOMEDCT_CORE|Toxic diffuse goiter|Toxic diffuse goiter
C0342122|T047|FN|267374005|SNOMEDCT_CORE|Toxic diffuse goiter|Toxic diffuse goiter
C0342122|T047|PTGB|267374005|SNOMEDCT_CORE|Toxic diffuse goitre|Toxic diffuse goiter
C0342122|T047|SY|267374005|SNOMEDCT_CORE|Toxic diffuse thyroid goiter|Toxic diffuse goiter
C0342122|T047|SYGB|267374005|SNOMEDCT_CORE|Toxic diffuse thyroid goitre|Toxic diffuse goiter
C0342122|T047|SY|267374005|SNOMEDCT_CORE|Toxic primary thyroid hyperplasia|Toxic diffuse goiter
C0342165|T047|PT|237527007|SNOMEDCT_CORE|Postablative hypothyroidism|Postablative hypothyroidism
C0342165|T047|FN|237527007|SNOMEDCT_CORE|Postablative hypothyroidism|Postablative hypothyroidism
C0342168|T047|PT|40539002|SNOMEDCT_CORE|Hypothyroidism following radioiodine therapy|Hypothyroidism following radioiodine therapy
C0342168|T047|FN|40539002|SNOMEDCT_CORE|Hypothyroidism following radioiodine therapy|Hypothyroidism following radioiodine therapy
C0342168|T047|SY|40539002|SNOMEDCT_CORE|Hypothyroidism, postradioiodine therapy|Hypothyroidism following radioiodine therapy
C0342168|T047|SY|40539002|SNOMEDCT_CORE|Radioactive iodine-induced hypothyroidism|Hypothyroidism following radioiodine therapy
C0342200|T047|IS|217710005|SNOMEDCT_CORE|Endemic cretinism|Endemic cretinism
C0342205|T047|PT|237569006|SNOMEDCT_CORE|Uninodular goiter|Uninodular goiter
C0342205|T047|FN|237569006|SNOMEDCT_CORE|Uninodular goiter|Uninodular goiter
C0342205|T047|PTGB|237569006|SNOMEDCT_CORE|Uninodular goitre|Uninodular goiter
C0342208|T047|PT|237570007|SNOMEDCT_CORE|Multinodular goiter|Multinodular goiter
C0342208|T047|FN|237570007|SNOMEDCT_CORE|Multinodular goiter|Multinodular goiter
C0342208|T047|PTGB|237570007|SNOMEDCT_CORE|Multinodular goitre|Multinodular goiter
C0342208|T047|SY|237570007|SNOMEDCT_CORE|Multiple thyroid nodules|Multinodular goiter
C0342208|T047|SY|237570007|SNOMEDCT_CORE|Thyroid goiter multinodular|Multinodular goiter
C0342208|T047|SYGB|237570007|SNOMEDCT_CORE|Thyroid goitre multinodular|Multinodular goiter
C0342245|T047|SY|25093002|SNOMEDCT_CORE|Diabetic eye disease|Disorder of eye due to diabetes mellitus
C0342245|T047|IS|25093002|SNOMEDCT_CORE|Diabetic eye disease, NOS|Disorder of eye due to diabetes mellitus
C0342245|T047|SY|25093002|SNOMEDCT_CORE|Diabetic oculopathy|Disorder of eye due to diabetes mellitus
C0342245|T047|OF|25093002|SNOMEDCT_CORE|Diabetic oculopathy|Disorder of eye due to diabetes mellitus
C0342245|T047|IS|25093002|SNOMEDCT_CORE|Diabetic oculopathy, NOS|Disorder of eye due to diabetes mellitus
C0342245|T047|IS|25093002|SNOMEDCT_CORE|Disorder of eye co-occurrent and due to diabetes mellitus|Disorder of eye due to diabetes mellitus
C0342245|T047|OF|25093002|SNOMEDCT_CORE|Disorder of eye co-occurrent and due to diabetes mellitus|Disorder of eye due to diabetes mellitus
C0342245|T047|PT|25093002|SNOMEDCT_CORE|Disorder of eye due to diabetes mellitus|Disorder of eye due to diabetes mellitus
C0342245|T047|FN|25093002|SNOMEDCT_CORE|Disorder of eye due to diabetes mellitus|Disorder of eye due to diabetes mellitus
C0342245|T047|SY|25093002|SNOMEDCT_CORE|Eye disorder due to diabetes mellitus|Disorder of eye due to diabetes mellitus
C0342245|T047|SY|25093002|SNOMEDCT_CORE|Ophthalmic manifestations of diabetes|Disorder of eye due to diabetes mellitus
C0342257|T047|FN|74627003|SNOMEDCT_CORE|Complication due to diabetes mellitus|Complication due to diabetes mellitus
C0342257|T047|PT|74627003|SNOMEDCT_CORE|Complication due to diabetes mellitus|Complication due to diabetes mellitus
C0342257|T047|SY|74627003|SNOMEDCT_CORE|Diabetic complication|Complication due to diabetes mellitus
C0342257|T047|OF|74627003|SNOMEDCT_CORE|Diabetic complication|Complication due to diabetes mellitus
C0342257|T047|IS|74627003|SNOMEDCT_CORE|Diabetic complication, NOS|Complication due to diabetes mellitus
C0342257|T047|SY|74627003|SNOMEDCT_CORE|Disorder associated with diabetes mellitus|Complication due to diabetes mellitus
C0342266|T047|SY|237599002|SNOMEDCT_CORE|Diabetes type 2 on insulin|Insulin treated type 2 diabetes mellitus
C0342266|T047|IS|237599002|SNOMEDCT_CORE|Insulin treated non-insulin dependent diabetes mellitus|Insulin treated type 2 diabetes mellitus
C0342266|T047|PT|237599002|SNOMEDCT_CORE|Insulin treated type 2 diabetes mellitus|Insulin treated type 2 diabetes mellitus
C0342266|T047|FN|237599002|SNOMEDCT_CORE|Insulin treated type 2 diabetes mellitus|Insulin treated type 2 diabetes mellitus
C0342266|T047|SY|237599002|SNOMEDCT_CORE|Insulin treated Type II diabetes mellitus|Insulin treated type 2 diabetes mellitus
C0342266|T047|IS|237599002|SNOMEDCT_CORE|Insulin-treated non-insulin-dependent diabetes mellitus|Insulin treated type 2 diabetes mellitus
C0342266|T047|OF|237599002|SNOMEDCT_CORE|Insulin-treated non-insulin-dependent diabetes mellitus|Insulin treated type 2 diabetes mellitus
C0342266|T047|IS|237599002|SNOMEDCT_CORE|NIDDM - Insulin-treated non-insulin-dependent diabetes mellitus|Insulin treated type 2 diabetes mellitus
C0342269|T047|PT|190447002|SNOMEDCT_CORE|Steroid-induced diabetes|Steroid-induced diabetes
C0342269|T047|FN|190447002|SNOMEDCT_CORE|Steroid-induced diabetes|Steroid-induced diabetes
C0342294|T047|SY|420270002|SNOMEDCT_CORE|Diabetes type 1 with ketoacidosis|Ketoacidosis due to type 1 diabetes mellitus
C0342294|T047|PT|420270002|SNOMEDCT_CORE|Ketoacidosis due to type 1 diabetes mellitus|Ketoacidosis due to type 1 diabetes mellitus
C0342294|T047|FN|420270002|SNOMEDCT_CORE|Ketoacidosis due to type 1 diabetes mellitus|Ketoacidosis due to type 1 diabetes mellitus
C0342294|T047|IS|420270002|SNOMEDCT_CORE|Ketoacidosis in insulin-dependent diabetes mellitus|Ketoacidosis due to type 1 diabetes mellitus
C0342294|T047|IS|420270002|SNOMEDCT_CORE|Ketoacidosis in juvenile-onset type diabetes mellitus|Ketoacidosis due to type 1 diabetes mellitus
C0342294|T047|SY|420270002|SNOMEDCT_CORE|Ketoacidosis in type 1 diabetes mellitus|Ketoacidosis due to type 1 diabetes mellitus
C0342294|T047|SY|420270002|SNOMEDCT_CORE|Ketoacidosis in type I diabetes mellitus|Ketoacidosis due to type 1 diabetes mellitus
C0342294|T047|OF|420270002|SNOMEDCT_CORE|Ketoacidosis in type I diabetes mellitus|Ketoacidosis due to type 1 diabetes mellitus
C0342295|T047|SY|421750000|SNOMEDCT_CORE|Diabetes type 2 with ketoacidosis|Ketoacidosis due to type 2 diabetes mellitus
C0342295|T047|PT|421750000|SNOMEDCT_CORE|Ketoacidosis due to type 2 diabetes mellitus|Ketoacidosis due to type 2 diabetes mellitus
C0342295|T047|FN|421750000|SNOMEDCT_CORE|Ketoacidosis due to type 2 diabetes mellitus|Ketoacidosis due to type 2 diabetes mellitus
C0342295|T047|IS|421750000|SNOMEDCT_CORE|Ketoacidosis in adult-onset type diabetes mellitus|Ketoacidosis due to type 2 diabetes mellitus
C0342295|T047|IS|421750000|SNOMEDCT_CORE|Ketoacidosis in non-insulin-dependent diabetes mellitus|Ketoacidosis due to type 2 diabetes mellitus
C0342295|T047|SY|421750000|SNOMEDCT_CORE|Ketoacidosis in type 2 diabetes mellitus|Ketoacidosis due to type 2 diabetes mellitus
C0342295|T047|SY|421750000|SNOMEDCT_CORE|Ketoacidosis in type II diabetes mellitus|Ketoacidosis due to type 2 diabetes mellitus
C0342295|T047|OF|421750000|SNOMEDCT_CORE|Ketoacidosis in type II diabetes mellitus|Ketoacidosis due to type 2 diabetes mellitus
C0342297|T047|OP|190331003|SNOMEDCT_CORE|Diabetes mellitus, adult onset, with hyperosmolar coma|Hyperosmolar coma due to type 2 diabetes mellitus
C0342297|T047|OF|190331003|SNOMEDCT_CORE|Diabetes mellitus, adult onset, with hyperosmolar coma|Hyperosmolar coma due to type 2 diabetes mellitus
C0342297|T047|PT|190331003|SNOMEDCT_CORE|Hyperosmolar coma due to type 2 diabetes mellitus|Hyperosmolar coma due to type 2 diabetes mellitus
C0342297|T047|FN|190331003|SNOMEDCT_CORE|Hyperosmolar coma due to type 2 diabetes mellitus|Hyperosmolar coma due to type 2 diabetes mellitus
C0342297|T047|SY|190331003|SNOMEDCT_CORE|Type 2 diabetes mellitus with hyperosmolar coma|Hyperosmolar coma due to type 2 diabetes mellitus
C0342297|T047|OF|190331003|SNOMEDCT_CORE|Type 2 diabetes mellitus with hyperosmolar coma|Hyperosmolar coma due to type 2 diabetes mellitus
C0342302|T047|SY|11530004|SNOMEDCT_CORE|Brittle diabetes|Brittle diabetes mellitus
C0342302|T047|OF|11530004|SNOMEDCT_CORE|Brittle diabetes|Brittle diabetes mellitus
C0342302|T047|PT|11530004|SNOMEDCT_CORE|Brittle diabetes mellitus|Brittle diabetes mellitus
C0342302|T047|OF|11530004|SNOMEDCT_CORE|Brittle diabetes mellitus|Brittle diabetes mellitus
C0342302|T047|FN|11530004|SNOMEDCT_CORE|Brittle diabetes mellitus|Brittle diabetes mellitus
C0342302|T047|SY|11530004|SNOMEDCT_CORE|Labile diabetes|Brittle diabetes mellitus
C0342302|T047|OAP|275918005|SNOMEDCT_CORE|Unstable diabetes|Brittle diabetes mellitus
C0342302|T047|OF|275918005|SNOMEDCT_CORE|Unstable diabetes|Brittle diabetes mellitus
C0342302|T047|OAF|275918005|SNOMEDCT_CORE|Unstable diabetes mellitus|Brittle diabetes mellitus
C0342302|T047|OAS|275918005|SNOMEDCT_CORE|Unstable diabetes mellitus|Brittle diabetes mellitus
C0342302|T047|SY|11530004|SNOMEDCT_CORE|Unstable diabetes mellitus|Brittle diabetes mellitus
C0342305|T047|OAS|237626009|SNOMEDCT_CORE|Pregnancy and IDDM|Pregnancy and IDDM
C0342305|T047|OAP|237626009|SNOMEDCT_CORE|Pregnancy and insulin-dependent diabetes mellitus|Pregnancy and IDDM
C0342305|T047|OAF|237626009|SNOMEDCT_CORE|Pregnancy and insulin-dependent diabetes mellitus|Pregnancy and IDDM
C0342307|T047|SY|237628005|SNOMEDCT_CORE|IGT - Impaired glucose tolerance in pregnancy|Impaired glucose tolerance in pregnancy
C0342307|T047|PT|237628005|SNOMEDCT_CORE|Impaired glucose tolerance in pregnancy|Impaired glucose tolerance in pregnancy
C0342307|T047|FN|237628005|SNOMEDCT_CORE|Impaired glucose tolerance in pregnancy|Impaired glucose tolerance in pregnancy
C0342307|T047|SY|237628005|SNOMEDCT_CORE|Pregnancy and impaired glucose tolerance|Impaired glucose tolerance in pregnancy
C0342312|T047|PTGB|237632004|SNOMEDCT_CORE|Hypoglycaemic event due to diabetes|Hypoglycemic event due to diabetes
C0342312|T047|SYGB|237632004|SNOMEDCT_CORE|Hypoglycaemic event in diabetes|Hypoglycemic event due to diabetes
C0342312|T047|PT|237632004|SNOMEDCT_CORE|Hypoglycemic event due to diabetes|Hypoglycemic event due to diabetes
C0342312|T047|FN|237632004|SNOMEDCT_CORE|Hypoglycemic event due to diabetes|Hypoglycemic event due to diabetes
C0342312|T047|SY|237632004|SNOMEDCT_CORE|Hypoglycemic event in diabetes|Hypoglycemic event due to diabetes
C0342312|T047|OF|237632004|SNOMEDCT_CORE|Hypoglycemic event in diabetes|Hypoglycemic event due to diabetes
C0342317|T047|SYGB|170766006|SNOMEDCT_CORE|Hypoglycaemia unawareness|Loss of hypoglycemic warning due to diabetes mellitus
C0342317|T047|SY|170766006|SNOMEDCT_CORE|Hypoglycemia unawareness|Loss of hypoglycemic warning due to diabetes mellitus
C0342317|T047|SYGB|170766006|SNOMEDCT_CORE|Loss of hypoglycaemic warning|Loss of hypoglycemic warning due to diabetes mellitus
C0342317|T047|PTGB|170766006|SNOMEDCT_CORE|Loss of hypoglycaemic warning due to diabetes mellitus|Loss of hypoglycemic warning due to diabetes mellitus
C0342317|T047|SY|170766006|SNOMEDCT_CORE|Loss of hypoglycemic warning|Loss of hypoglycemic warning due to diabetes mellitus
C0342317|T047|OF|170766006|SNOMEDCT_CORE|Loss of hypoglycemic warning|Loss of hypoglycemic warning due to diabetes mellitus
C0342317|T047|PT|170766006|SNOMEDCT_CORE|Loss of hypoglycemic warning due to diabetes mellitus|Loss of hypoglycemic warning due to diabetes mellitus
C0342317|T047|FN|170766006|SNOMEDCT_CORE|Loss of hypoglycemic warning due to diabetes mellitus|Loss of hypoglycemic warning due to diabetes mellitus
C0342321|T046|PTGB|237640005|SNOMEDCT_CORE|Drug-induced hypoglycaemia|Drug-induced hypoglycemia
C0342321|T046|PT|237640005|SNOMEDCT_CORE|Drug-induced hypoglycemia|Drug-induced hypoglycemia
C0342321|T046|FN|237640005|SNOMEDCT_CORE|Drug-induced hypoglycemia|Drug-induced hypoglycemia
C0342388|T047|PT|237692001|SNOMEDCT_CORE|ACTH deficiency|ACTH deficiency
C0342388|T047|OF|237692001|SNOMEDCT_CORE|ACTH deficiency|ACTH deficiency
C0342388|T047|OF|237692001|SNOMEDCT_CORE|Adrenocorticotropic hormone deficiency|ACTH deficiency
C0342388|T047|FN|237692001|SNOMEDCT_CORE|Adrenocorticotropic hormone deficiency|ACTH deficiency
C0342388|T047|SY|237692001|SNOMEDCT_CORE|Adrenocorticotropic hormone deficiency|ACTH deficiency
C0342388|T047|SY|237692001|SNOMEDCT_CORE|Secondary hypoadrenalism|ACTH deficiency
C0342399|T033|PT|14900002|SNOMEDCT_CORE|Hypopituitarism due to radiotherapy|Hypopituitarism due to radiotherapy
C0342399|T033|SY|14900002|SNOMEDCT_CORE|Post-radiotherapy hypopituitarism|Hypopituitarism due to radiotherapy
C0342399|T033|SY|14900002|SNOMEDCT_CORE|Radiotherapy-induced hypopituitarism|Hypopituitarism due to radiotherapy
C0342399|T033|FN|14900002|SNOMEDCT_CORE|Radiotherapy-induced hypopituitarism|Hypopituitarism due to radiotherapy
C0342419|T190|SY|237715007|SNOMEDCT_CORE|Mass of pituitary|Pituitary mass
C0342419|T190|FN|237715007|SNOMEDCT_CORE|Mass of pituitary|Pituitary mass
C0342419|T190|PT|237715007|SNOMEDCT_CORE|Pituitary mass|Pituitary mass
C0342419|T190|OF|237715007|SNOMEDCT_CORE|Pituitary mass|Pituitary mass
C0342500|T047|PT|237783006|SNOMEDCT_CORE|Adrenal mass|Adrenal mass
C0342500|T047|OF|237783006|SNOMEDCT_CORE|Adrenal mass|Adrenal mass
C0342500|T047|SY|237783006|SNOMEDCT_CORE|Mass of adrenal gland|Adrenal mass
C0342500|T047|FN|237783006|SNOMEDCT_CORE|Mass of adrenal gland|Adrenal mass
C0342579|T046|PT|105593004|SNOMEDCT_CORE|Electrolyte imbalance|Electrolyte imbalance
C0342579|T046|FN|105593004|SNOMEDCT_CORE|Electrolyte imbalance|Electrolyte imbalance
C0342634|T047|PTGB|268846006|SNOMEDCT_CORE|Neonatal hypocalcaemia|Neonatal hypocalcemia
C0342634|T047|PT|268846006|SNOMEDCT_CORE|Neonatal hypocalcemia|Neonatal hypocalcemia
C0342634|T047|FN|268846006|SNOMEDCT_CORE|Neonatal hypocalcemia|Neonatal hypocalcemia
C0343020|T047|PT|238389005|SNOMEDCT_CORE|Boils of multiple sites|Boils of multiple sites
C0343020|T047|FN|238389005|SNOMEDCT_CORE|Boils of multiple sites|Boils of multiple sites
C0343021|T047|PT|200586004|SNOMEDCT_CORE|Carbuncle of back|Carbuncle of back
C0343021|T047|FN|200586004|SNOMEDCT_CORE|Carbuncle of back|Carbuncle of back
C0343024|T047|OAP|238402004|SNOMEDCT_CORE|Cellulitis of leg|Cellulitis of leg
C0343024|T047|OAF|238402004|SNOMEDCT_CORE|Cellulitis of leg|Cellulitis of leg
C0343024|T047|OAS|238402004|SNOMEDCT_CORE|Cellulitis of lower limb|Cellulitis of leg
C0343047|T047|SY|7297005|SNOMEDCT_CORE|Erythroderma desquamativum|Generalized seborrheic dermatitis of infants
C0343047|T047|PTGB|7297005|SNOMEDCT_CORE|Generalised seborrhoeic dermatitis of infants|Generalized seborrheic dermatitis of infants
C0343047|T047|PT|7297005|SNOMEDCT_CORE|Generalized seborrheic dermatitis of infants|Generalized seborrheic dermatitis of infants
C0343047|T047|FN|7297005|SNOMEDCT_CORE|Generalized seborrheic dermatitis of infants|Generalized seborrheic dermatitis of infants
C0343047|T047|OAP|200776003|SNOMEDCT_CORE|Infantile seborrheic dermatitis|Generalized seborrheic dermatitis of infants
C0343047|T047|SY|7297005|SNOMEDCT_CORE|Infantile seborrheic dermatitis|Generalized seborrheic dermatitis of infants
C0343047|T047|OAF|200776003|SNOMEDCT_CORE|Infantile seborrheic dermatitis|Generalized seborrheic dermatitis of infants
C0343047|T047|OAP|200776003|SNOMEDCT_CORE|Infantile seborrhoeic dermatitis|Generalized seborrheic dermatitis of infants
C0343047|T047|SYGB|7297005|SNOMEDCT_CORE|Infantile seborrhoeic dermatitis|Generalized seborrheic dermatitis of infants
C0343047|T047|SY|7297005|SNOMEDCT_CORE|Leiner's disease|Generalized seborrheic dermatitis of infants
C0343052|T047|PT|37042000|SNOMEDCT_CORE|Guttate psoriasis|Guttate psoriasis
C0343052|T047|FN|37042000|SNOMEDCT_CORE|Guttate psoriasis|Guttate psoriasis
C0343052|T047|SY|37042000|SNOMEDCT_CORE|Psoriasis guttata|Guttate psoriasis
C0343065|T047|PT|402410006|SNOMEDCT_CORE|Symptomatic dermographism|Symptomatic dermographism
C0343065|T047|FN|402410006|SNOMEDCT_CORE|Symptomatic dermographism|Symptomatic dermographism
C0343082|T191|SY|5050001|SNOMEDCT_CORE|Blood spots on skin|Senile angioma
C0343082|T191|SY|5050001|SNOMEDCT_CORE|Campbell de Morgan angioma|Senile angioma
C0343082|T191|SY|5050001|SNOMEDCT_CORE|Campbell de Morgan spot|Senile angioma
C0343082|T191|SY|5050001|SNOMEDCT_CORE|Cherry angioma|Senile angioma
C0343082|T191|SY|5050001|SNOMEDCT_CORE|De Morgan's spots|Senile angioma
C0343082|T191|PT|5050001|SNOMEDCT_CORE|Senile angioma|Senile angioma
C0343082|T191|FN|5050001|SNOMEDCT_CORE|Senile angioma|Senile angioma
C0343082|T191|SY|5050001|SNOMEDCT_CORE|Senile ectasia|Senile angioma
C0343082|T191|SYGB|5050001|SNOMEDCT_CORE|Senile naevus of skin|Senile angioma
C0343082|T191|SY|5050001|SNOMEDCT_CORE|Senile nevus of skin|Senile angioma
C0343140|T047|SY|111222003|SNOMEDCT_CORE|Derangement medial meniscus|Derangement of medial meniscus
C0343140|T047|PT|111222003|SNOMEDCT_CORE|Derangement of medial meniscus|Derangement of medial meniscus
C0343140|T047|FN|111222003|SNOMEDCT_CORE|Derangement of medial meniscus|Derangement of medial meniscus
C0343145|T020|PT|239735004|SNOMEDCT_CORE|Contracture of wrist joint|Contracture of wrist joint
C0343145|T020|FN|239735004|SNOMEDCT_CORE|Contracture of wrist joint|Contracture of wrist joint
C0343145|T020|SY|239735004|SNOMEDCT_CORE|Wrist joint contracture|Contracture of wrist joint
C0343146|T020|PT|239737007|SNOMEDCT_CORE|Contracture of joint of finger|Contracture of joint of finger
C0343146|T020|FN|239737007|SNOMEDCT_CORE|Contracture of joint of finger|Contracture of joint of finger
C0343147|T020|PT|239739005|SNOMEDCT_CORE|Contracture of knee joint|Contracture of knee joint
C0343147|T020|FN|239739005|SNOMEDCT_CORE|Contracture of knee joint|Contracture of knee joint
C0343147|T020|SY|239739005|SNOMEDCT_CORE|Knee joint contracture|Contracture of knee joint
C0343161|T020|OAP|239769003|SNOMEDCT_CORE|Joint mice in knee|Loose body in knee
C0343161|T020|OAF|239769003|SNOMEDCT_CORE|Joint mice in knee|Loose body in knee
C0343161|T020|SY|81512004|SNOMEDCT_CORE|Joint mice of knee|Loose body in knee
C0343161|T020|PT|81512004|SNOMEDCT_CORE|Loose body in knee|Loose body in knee
C0343161|T020|FN|81512004|SNOMEDCT_CORE|Loose body in knee|Loose body in knee
C0343161|T020|IS|81512004|SNOMEDCT_CORE|Loose body in knee, NOS|Loose body in knee
C0343166|T033|SY|202381003|SNOMEDCT_CORE|Effusion of knee|Knee joint effusion
C0343166|T033|PT|202381003|SNOMEDCT_CORE|Knee joint effusion|Knee joint effusion
C0343166|T033|FN|202381003|SNOMEDCT_CORE|Knee joint effusion|Knee joint effusion
C0343170|T046|PTGB|202413005|SNOMEDCT_CORE|Haemarthrosis of knee|Hemarthrosis of knee
C0343170|T046|PT|202413005|SNOMEDCT_CORE|Hemarthrosis of knee|Hemarthrosis of knee
C0343170|T046|FN|202413005|SNOMEDCT_CORE|Hemarthrosis of knee|Hemarthrosis of knee
C0343178|T046|SY|201724008|SNOMEDCT_CORE|Diabetic Charcot's arthropathy|Neuropathic arthropathy due to diabetes mellitus
C0343178|T046|SY|201724008|SNOMEDCT_CORE|Diabetic neuropathic arthropathy|Neuropathic arthropathy due to diabetes mellitus
C0343178|T046|OF|201724008|SNOMEDCT_CORE|Diabetic neuropathic arthropathy|Neuropathic arthropathy due to diabetes mellitus
C0343178|T046|FN|201724008|SNOMEDCT_CORE|Neuropathic arthropathy due to diabetes mellitus|Neuropathic arthropathy due to diabetes mellitus
C0343178|T046|PT|201724008|SNOMEDCT_CORE|Neuropathic arthropathy due to diabetes mellitus|Neuropathic arthropathy due to diabetes mellitus
C0343179|T047|SY|202924004|SNOMEDCT_CORE|Toxic synovitis|Transient synovitis
C0343179|T047|PT|202924004|SNOMEDCT_CORE|Transient synovitis|Transient synovitis
C0343179|T047|FN|202924004|SNOMEDCT_CORE|Transient synovitis|Transient synovitis
C0343216|T046|IS|302938005|SNOMEDCT_CORE|Tendinitis and tenosynovitis of the ankle region|Tendinitis AND/OR tenosynovitis of the ankle region
C0343216|T046|OF|302938005|SNOMEDCT_CORE|Tendinitis and tenosynovitis of the ankle region|Tendinitis AND/OR tenosynovitis of the ankle region
C0343216|T046|OAF|302938005|SNOMEDCT_CORE|Tendinitis AND/OR tenosynovitis of the ankle region|Tendinitis AND/OR tenosynovitis of the ankle region
C0343216|T046|OF|302938005|SNOMEDCT_CORE|Tendinitis and/or tenosynovitis of the ankle region|Tendinitis AND/OR tenosynovitis of the ankle region
C0343216|T046|OAP|302938005|SNOMEDCT_CORE|Tendinitis AND/OR tenosynovitis of the ankle region|Tendinitis AND/OR tenosynovitis of the ankle region
C0343216|T046|IS|302938005|SNOMEDCT_CORE|Tendinitis and/or tenosynovitis of the ankle region|Tendinitis AND/OR tenosynovitis of the ankle region
C0343216|T046|OAS|302938005|SNOMEDCT_CORE|Tendonitis AND/OR tenosynovitis of the ankle region|Tendinitis AND/OR tenosynovitis of the ankle region
C0343230|T047|IS|240008008|SNOMEDCT_CORE|Ganglion of knee|Ganglion of knee
C0343231|T047|SY|202942009|SNOMEDCT_CORE|Ganglion cyst of wrist|Ganglion of wrist
C0343231|T047|PT|202942009|SNOMEDCT_CORE|Ganglion of wrist|Ganglion of wrist
C0343231|T047|FN|202942009|SNOMEDCT_CORE|Ganglion of wrist|Ganglion of wrist
C0343238|T047|SY|193253000|SNOMEDCT_CORE|Myopathy due to Sjögren disease|Myopathy due to Sjögren's disease
C0343238|T047|PT|193253000|SNOMEDCT_CORE|Myopathy due to Sjögren's disease|Myopathy due to Sjögren's disease
C0343238|T047|SY|193253000|SNOMEDCT_CORE|Myopathy due to Sjogren's disease|Myopathy due to Sjögren's disease
C0343238|T047|FN|193253000|SNOMEDCT_CORE|Myopathy due to Sjögren's disease|Myopathy due to Sjögren's disease
C0343238|T047|OF|193253000|SNOMEDCT_CORE|Myopathy due to Sjogren's disease|Myopathy due to Sjögren's disease
C0343238|T047|SY|193253000|SNOMEDCT_CORE|Myopathy due to Sjogrens disease|Myopathy due to Sjögren's disease
C0343314|T047|PT|206356004|SNOMEDCT_CORE|Neonatal candidiasis of perineum|Neonatal candidiasis of perineum
C0343314|T047|FN|206356004|SNOMEDCT_CORE|Neonatal candidiasis of perineum|Neonatal candidiasis of perineum
C0343378|T047|IS|89538001|SNOMEDCT_CORE|Helicobacter pylori-associated gastritis|Helicobacter-associated gastritis
C0343378|T047|PT|89538001|SNOMEDCT_CORE|Helicobacter-associated gastritis|Helicobacter-associated gastritis
C0343378|T047|FN|89538001|SNOMEDCT_CORE|Helicobacter-associated gastritis|Helicobacter-associated gastritis
C0343386|T047|SY|186431008|SNOMEDCT_CORE|Clostridioides difficile gastrointestinal tract infection|Clostridioides difficile infection
C0343386|T047|FN|186431008|SNOMEDCT_CORE|Clostridioides difficile infection|Clostridioides difficile infection
C0343386|T047|PT|186431008|SNOMEDCT_CORE|Clostridioides difficile infection|Clostridioides difficile infection
C0343386|T047|SY|186431008|SNOMEDCT_CORE|Clostridium difficile gastrointestinal tract infection|Clostridioides difficile infection
C0343386|T047|SY|186431008|SNOMEDCT_CORE|Clostridium difficile infection|Clostridioides difficile infection
C0343386|T047|OF|186431008|SNOMEDCT_CORE|Clostridium difficile infection|Clostridioides difficile infection
C0343401|T047|SY|266096002|SNOMEDCT_CORE|Infection due to Methicillin resistant Staphylococcus aureus|Methicillin resistant Staphylococcus aureus infection
C0343401|T047|PT|266096002|SNOMEDCT_CORE|Methicillin resistant Staphylococcus aureus infection|Methicillin resistant Staphylococcus aureus infection
C0343401|T047|FN|266096002|SNOMEDCT_CORE|Methicillin resistant Staphylococcus aureus infection|Methicillin resistant Staphylococcus aureus infection
C0343401|T047|IS|266096002|SNOMEDCT_CORE|Methicillin-resistant staphylococcus aureus|Methicillin resistant Staphylococcus aureus infection
C0343401|T047|IS|266096002|SNOMEDCT_CORE|Methicillin-resistant staphylococcus aureus infection|Methicillin resistant Staphylococcus aureus infection
C0343401|T047|OF|266096002|SNOMEDCT_CORE|Methicillin-resistant staphylococcus aureus infection|Methicillin resistant Staphylococcus aureus infection
C0343401|T047|IS|266096002|SNOMEDCT_CORE|MRSA - Methicillin-resistant staphylococcus aureus|Methicillin resistant Staphylococcus aureus infection
C0343401|T047|IS|266096002|SNOMEDCT_CORE|MRSA infection|Methicillin resistant Staphylococcus aureus infection
C0343413|T047|PT|187252008|SNOMEDCT_CORE|Late effects of respiratory tuberculosis|Late effects of respiratory tuberculosis
C0343413|T047|FN|187252008|SNOMEDCT_CORE|Late effects of respiratory tuberculosis|Late effects of respiratory tuberculosis
C0343495|T033|IS|76902006|SNOMEDCT_CORE|Lockjaw|Lockjaw
C0343495|T033|IS|76902006|SNOMEDCT_CORE|Tetanus with trismus|Lockjaw
C0343641|T047|PT|240532009|SNOMEDCT_CORE|Human papilloma virus infection|Human papilloma virus infection
C0343641|T047|OF|240532009|SNOMEDCT_CORE|Human papilloma virus infection|Human papilloma virus infection
C0343641|T047|SY|240532009|SNOMEDCT_CORE|Human papillomavirus infection|Human papilloma virus infection
C0343641|T047|FN|240532009|SNOMEDCT_CORE|Human papillomavirus infection|Human papilloma virus infection
C0343751|T047|SY|91947003|SNOMEDCT_CORE|Asymptomatic HIV infection|Asymptomatic human immunodeficiency virus infection
C0343751|T047|PT|91947003|SNOMEDCT_CORE|Asymptomatic human immunodeficiency virus infection|Asymptomatic human immunodeficiency virus infection
C0343751|T047|FN|91947003|SNOMEDCT_CORE|Asymptomatic human immunodeficiency virus infection|Asymptomatic human immunodeficiency virus infection
C0343874|T047|SYGB|240711004|SNOMEDCT_CORE|Candidal nappy rash|Diaper candidiasis
C0343874|T047|PT|240711004|SNOMEDCT_CORE|Diaper candidiasis|Diaper candidiasis
C0343874|T047|FN|240711004|SNOMEDCT_CORE|Diaper candidiasis|Diaper candidiasis
C0343874|T047|SY|240711004|SNOMEDCT_CORE|Diaper candidosis|Diaper candidiasis
C0343874|T047|SYGB|240711004|SNOMEDCT_CORE|Monilial nappy rash|Diaper candidiasis
C0343874|T047|PTGB|240711004|SNOMEDCT_CORE|Napkin candidiasis|Diaper candidiasis
C0343874|T047|OF|240711004|SNOMEDCT_CORE|Napkin candidiasis|Diaper candidiasis
C0343874|T047|SYGB|240711004|SNOMEDCT_CORE|Napkin candidosis|Diaper candidiasis
C0344125|T037|OAP|111757004|SNOMEDCT_CORE|Poisoning by aromatic analgesic|Poisoning caused by aromatic analgesic
C0344125|T037|OF|111757004|SNOMEDCT_CORE|Poisoning by aromatic analgesic|Poisoning caused by aromatic analgesic
C0344125|T037|OAF|111757004|SNOMEDCT_CORE|Poisoning caused by aromatic analgesic|Poisoning caused by aromatic analgesic
C0344125|T037|OAS|111757004|SNOMEDCT_CORE|Poisoning caused by aromatic analgesic|Poisoning caused by aromatic analgesic
C0344155|T037|SY|11196001|SNOMEDCT_CORE|Narcotic poisoning|Narcotic poisoning
C0344198|T033|SY|406137001|SNOMEDCT_CORE|Adult abuse|Adult victim of abuse
C0344198|T033|FN|406137001|SNOMEDCT_CORE|Adult victim of abuse|Adult victim of abuse
C0344198|T033|PT|406137001|SNOMEDCT_CORE|Adult victim of abuse|Adult victim of abuse
C0344221|T033|SY|312081001|SNOMEDCT_CORE|Coil contraception|IUD contraception
C0344221|T033|IS|312081001|SNOMEDCT_CORE|Contraceptive IUD in situ|IUD contraception
C0344221|T033|SY|312081001|SNOMEDCT_CORE|Intrauterine device contraception|IUD contraception
C0344221|T033|FN|312081001|SNOMEDCT_CORE|Intrauterine device contraception|IUD contraception
C0344221|T033|OF|312081001|SNOMEDCT_CORE|Intrauterine device contraception|IUD contraception
C0344221|T033|PT|312081001|SNOMEDCT_CORE|IUD contraception|IUD contraception
C0344221|T033|OF|312081001|SNOMEDCT_CORE|IUD contraception|IUD contraception
C0344221|T033|IS|312081001|SNOMEDCT_CORE|IUD in situ|IUD contraception
C0344226|T033|PT|275917000|SNOMEDCT_CORE|Lithium monitoring|Lithium monitoring
C0344226|T033|FN|275917000|SNOMEDCT_CORE|Lithium monitoring|Lithium monitoring
C0344232|T033|IS|111516008|SNOMEDCT_CORE|Blurred vision|Hazy vision
C0344232|T033|IS|246636008|SNOMEDCT_CORE|Blurred vision|Hazy vision
C0344232|T033|IS|246636008|SNOMEDCT_CORE|Blurred vision - hazy|Hazy vision
C0344232|T033|IS|111516008|SNOMEDCT_CORE|Blurred vision, NOS|Hazy vision
C0344232|T033|PT|111516008|SNOMEDCT_CORE|Blurring of visual image|Hazy vision
C0344232|T033|FN|111516008|SNOMEDCT_CORE|Blurring of visual image|Hazy vision
C0344232|T033|SY|246636008|SNOMEDCT_CORE|Cloudy vision|Hazy vision
C0344232|T033|SY|246636008|SNOMEDCT_CORE|Foggy vision|Hazy vision
C0344232|T033|PT|246636008|SNOMEDCT_CORE|Hazy vision|Hazy vision
C0344232|T033|FN|246636008|SNOMEDCT_CORE|Hazy vision|Hazy vision
C0344232|T033|SY|246636008|SNOMEDCT_CORE|Mist over eyes|Hazy vision
C0344232|T033|SY|246636008|SNOMEDCT_CORE|Misty vision|Hazy vision
C0344233|T033|SY|23388006|SNOMEDCT_CORE|Blind spot|Blind spot
C0344304|T184|SY|102614006|SNOMEDCT_CORE|General abdominal pain-symptom|Generalized abdominal pain
C0344304|T184|PTGB|102614006|SNOMEDCT_CORE|Generalised abdominal pain|Generalized abdominal pain
C0344304|T184|PT|102614006|SNOMEDCT_CORE|Generalized abdominal pain|Generalized abdominal pain
C0344304|T184|FN|102614006|SNOMEDCT_CORE|Generalized abdominal pain|Generalized abdominal pain
C0344306|T184|PT|247389006|SNOMEDCT_CORE|Intercostal neuralgia|Intercostal neuralgia
C0344306|T184|FN|247389006|SNOMEDCT_CORE|Intercostal neuralgia|Intercostal neuralgia
C0344306|T184|OF|247389006|SNOMEDCT_CORE|Intercostal neuralgia|Intercostal neuralgia
C0344315|T048|OAS|41006004|SNOMEDCT_CORE|Depressed|Depressed mood
C0344315|T048|SY|35489007|SNOMEDCT_CORE|Depressed|Depressed mood
C0344315|T048|IS|41006004|SNOMEDCT_CORE|Depressed mood|Depressed mood
C0344315|T048|IS|41006004|SNOMEDCT_CORE|Feeling low|Depressed mood
C0344315|T048|IS|41006004|SNOMEDCT_CORE|Low mood|Depressed mood
C0344315|T048|OAS|41006004|SNOMEDCT_CORE|Melancholic|Depressed mood
C0344315|T048|OAS|41006004|SNOMEDCT_CORE|Miserable|Depressed mood
C0344315|T048|OAS|41006004|SNOMEDCT_CORE|Morose mood|Depressed mood
C0344315|T048|OAS|41006004|SNOMEDCT_CORE|Morosity|Depressed mood
C0344365|T184|SY|249288007|SNOMEDCT_CORE|Incomplete bladder emptying|Incomplete emptying of bladder
C0344365|T184|PT|249288007|SNOMEDCT_CORE|Incomplete emptying of bladder|Incomplete emptying of bladder
C0344365|T184|FN|249288007|SNOMEDCT_CORE|Incomplete emptying of bladder|Incomplete emptying of bladder
C0344453|T191|PT|253011004|SNOMEDCT_CORE|Macroprolactinoma|Macroprolactinoma
C0344453|T191|FN|253011004|SNOMEDCT_CORE|Macroprolactinoma|Macroprolactinoma
C0344503|T019|PT|253212001|SNOMEDCT_CORE|Epiblepharon|Epiblepharon
C0344503|T019|FN|253212001|SNOMEDCT_CORE|Epiblepharon|Epiblepharon
C0344616|T019|SY|83799000|SNOMEDCT_CORE|Congenitally corrected transposition of great arteries|Corrected transposition of great vessels
C0344616|T019|PT|83799000|SNOMEDCT_CORE|Corrected transposition of great vessels|Corrected transposition of great vessels
C0344616|T019|FN|83799000|SNOMEDCT_CORE|Corrected transposition of great vessels|Corrected transposition of great vessels
C0344616|T019|SY|83799000|SNOMEDCT_CORE|Discordant ventriculoarterial connection with discordant atrioventricular connection|Corrected transposition of great vessels
C0344616|T019|SY|83799000|SNOMEDCT_CORE|Transposition of great vessels with ventricular inversion|Corrected transposition of great vessels
C0344787|T019|PT|253416000|SNOMEDCT_CORE|Atrioventricular septal defect: atrial and ventricular components|Atrioventricular septal defect: atrial and ventricular components
C0344787|T019|FN|253416000|SNOMEDCT_CORE|Atrioventricular septal defect: atrial and ventricular components|Atrioventricular septal defect: atrial and ventricular components
C0344787|T019|SY|253416000|SNOMEDCT_CORE|Complete atrioventricular septal defect|Atrioventricular septal defect: atrial and ventricular components
C0344925|T019|PT|109428005|SNOMEDCT_CORE|Perimembranous ventricular septal defect|Perimembranous ventricular septal defect
C0344925|T019|FN|109428005|SNOMEDCT_CORE|Perimembranous ventricular septal defect|Perimembranous ventricular septal defect
C0345160|T019|PT|253737007|SNOMEDCT_CORE|Congenital laryngomalacia|Congenital laryngomalacia
C0345160|T019|FN|253737007|SNOMEDCT_CORE|Congenital laryngomalacia|Congenital laryngomalacia
C0345247|T019|PTGB|253785008|SNOMEDCT_CORE|Generalised congenital intestinal dysmotility|Generalized congenital intestinal dysmotility
C0345247|T019|IS|253785008|SNOMEDCT_CORE|Generalised intestinal dysmotility|Generalized congenital intestinal dysmotility
C0345247|T019|PT|253785008|SNOMEDCT_CORE|Generalized congenital intestinal dysmotility|Generalized congenital intestinal dysmotility
C0345247|T019|FN|253785008|SNOMEDCT_CORE|Generalized congenital intestinal dysmotility|Generalized congenital intestinal dysmotility
C0345247|T019|IS|253785008|SNOMEDCT_CORE|Generalized intestinal dysmotility|Generalized congenital intestinal dysmotility
C0345247|T019|OF|253785008|SNOMEDCT_CORE|Generalized intestinal dysmotility|Generalized congenital intestinal dysmotility
C0345303|T019|PT|253826001|SNOMEDCT_CORE|Embryonic cyst of broad ligament|Embryonic cyst of broad ligament
C0345303|T019|FN|253826001|SNOMEDCT_CORE|Embryonic cyst of broad ligament|Embryonic cyst of broad ligament
C0345325|T019|SY|39526006|SNOMEDCT_CORE|Long foreskin|Redundant prepuce
C0345325|T019|SY|39526006|SNOMEDCT_CORE|Redundant foreskin|Redundant prepuce
C0345325|T019|PT|39526006|SNOMEDCT_CORE|Redundant prepuce|Redundant prepuce
C0345325|T019|FN|39526006|SNOMEDCT_CORE|Redundant prepuce|Redundant prepuce
C0345354|T019|SY|205135003|SNOMEDCT_CORE|Preaxial polydactyly|Radial polydactyly
C0345354|T019|PT|205135003|SNOMEDCT_CORE|Radial polydactyly|Radial polydactyly
C0345354|T019|FN|205135003|SNOMEDCT_CORE|Radial polydactyly|Radial polydactyly
C0345392|T019|PT|405772002|SNOMEDCT_CORE|Congenital kyphoscoliosis|Congenital kyphoscoliosis
C0345392|T019|FN|405772002|SNOMEDCT_CORE|Congenital kyphoscoliosis|Congenital kyphoscoliosis
C0345468|T046|PT|213148006|SNOMEDCT_CORE|Transplanted organ rejection|Transplanted organ rejection
C0345468|T046|FN|213148006|SNOMEDCT_CORE|Transplanted organ rejection|Transplanted organ rejection
C0345602|T191|PT|254462001|SNOMEDCT_CORE|Carcinoma of parotid gland|Carcinoma of parotid gland
C0345602|T191|FN|254462001|SNOMEDCT_CORE|Carcinoma of parotid gland|Carcinoma of parotid gland
C0345779|T191|PT|254547001|SNOMEDCT_CORE|Carcinoma of upper third of esophagus|Carcinoma of upper third of esophagus
C0345779|T191|FN|254547001|SNOMEDCT_CORE|Carcinoma of upper third of esophagus|Carcinoma of upper third of esophagus
C0345779|T191|PTGB|254547001|SNOMEDCT_CORE|Carcinoma of upper third of oesophagus|Carcinoma of upper third of esophagus
C0345794|T191|PT|254553001|SNOMEDCT_CORE|Carcinoma of cardia|Carcinoma of cardia
C0345794|T191|FN|254553001|SNOMEDCT_CORE|Carcinoma of cardia|Carcinoma of cardia
C0345804|T191|PT|254557000|SNOMEDCT_CORE|Carcinoma of body of stomach|Carcinoma of body of stomach
C0345804|T191|FN|254557000|SNOMEDCT_CORE|Carcinoma of body of stomach|Carcinoma of body of stomach
C0345809|T191|PT|254559002|SNOMEDCT_CORE|Carcinoma of pyloric antrum|Carcinoma of pyloric antrum
C0345809|T191|FN|254559002|SNOMEDCT_CORE|Carcinoma of pyloric antrum|Carcinoma of pyloric antrum
C0345814|T191|PT|254561006|SNOMEDCT_CORE|Carcinoma of pylorus|Carcinoma of pylorus
C0345814|T191|FN|254561006|SNOMEDCT_CORE|Carcinoma of pylorus|Carcinoma of pylorus
C0345832|T191|PT|126832004|SNOMEDCT_CORE|Neoplasm of small intestine|Neoplasm of small intestine
C0345832|T191|FN|126832004|SNOMEDCT_CORE|Neoplasm of small intestine|Neoplasm of small intestine
C0345832|T191|SY|126832004|SNOMEDCT_CORE|Tumor of small intestine|Neoplasm of small intestine
C0345832|T191|SYGB|126832004|SNOMEDCT_CORE|Tumour of small intestine|Neoplasm of small intestine
C0345903|T190|PT|195469007|SNOMEDCT_CORE|Anal skin tag|Anal skin tag
C0345903|T190|FN|195469007|SNOMEDCT_CORE|Anal skin tag|Anal skin tag
C0345903|T190|SY|195469007|SNOMEDCT_CORE|Anal tag|Anal skin tag
C0345903|T190|SY|195469007|SNOMEDCT_CORE|Fibrous polyp of anus|Anal skin tag
C0345904|T191|SY|93870000|SNOMEDCT_CORE|CA - Liver cancer|Malignant neoplasm of liver
C0345904|T191|SY|93870000|SNOMEDCT_CORE|Liver cancer|Malignant neoplasm of liver
C0345904|T191|PT|93870000|SNOMEDCT_CORE|Malignant neoplasm of liver|Malignant neoplasm of liver
C0345904|T191|FN|93870000|SNOMEDCT_CORE|Malignant neoplasm of liver|Malignant neoplasm of liver
C0345904|T191|IS|93870000|SNOMEDCT_CORE|Malignant neoplasm of liver, NOS|Malignant neoplasm of liver
C0345904|T191|SY|93870000|SNOMEDCT_CORE|Malignant tumor of liver|Malignant neoplasm of liver
C0345904|T191|SYGB|93870000|SNOMEDCT_CORE|Malignant tumour of liver|Malignant neoplasm of liver
C0345950|T191|IS|254622008|SNOMEDCT_CORE|Primary bronchial cancer|Primary bronchial cancer
C0345989|T047|SY|254671003|SNOMEDCT_CORE|Infected sebaceous cyst|Infection of sebaceous cyst
C0345989|T047|OF|254671003|SNOMEDCT_CORE|Infected sebaceous cyst|Infection of sebaceous cyst
C0345989|T047|SY|254671003|SNOMEDCT_CORE|Infected sebaceous cyst of skin|Infection of sebaceous cyst
C0345989|T047|PT|254671003|SNOMEDCT_CORE|Infection of sebaceous cyst|Infection of sebaceous cyst
C0345989|T047|FN|254671003|SNOMEDCT_CORE|Infection of sebaceous cyst|Infection of sebaceous cyst
C0345996|T190|PT|254679001|SNOMEDCT_CORE|Milia|Milia
C0345996|T190|FN|254679001|SNOMEDCT_CORE|Milia|Milia
C0345996|T190|OAP|254683001|SNOMEDCT_CORE|Milial cyst|Milia
C0345996|T190|OAF|254683001|SNOMEDCT_CORE|Milial cyst|Milia
C0346032|T191|SY|254727007|SNOMEDCT_CORE|Extramammary Paget disease of skin|Extramammary Paget's disease of skin
C0346032|T191|PT|254727007|SNOMEDCT_CORE|Extramammary Paget's disease of skin|Extramammary Paget's disease of skin
C0346032|T191|FN|254727007|SNOMEDCT_CORE|Extramammary Paget's disease of skin|Extramammary Paget's disease of skin
C0346032|T191|SY|254727007|SNOMEDCT_CORE|Extramammary Pagets disease of skin|Extramammary Paget's disease of skin
C0346040|T191|SY|109266006|SNOMEDCT_CORE|In situ malignant melanoma of skin|Melanoma in situ of skin
C0346040|T191|SY|109266006|SNOMEDCT_CORE|In situ melanoma of skin|Melanoma in situ of skin
C0346040|T191|SY|109266006|SNOMEDCT_CORE|ISM - In situ melanoma of skin|Melanoma in situ of skin
C0346040|T191|SY|109266006|SNOMEDCT_CORE|ISMM - In situ malignant melanoma of skin|Melanoma in situ of skin
C0346040|T191|SY|109266006|SNOMEDCT_CORE|Melanoma in situ of skin|Melanoma in situ of skin
C0346040|T191|PT|109266006|SNOMEDCT_CORE|Melanoma in situ of skin|Melanoma in situ of skin
C0346040|T191|FN|109266006|SNOMEDCT_CORE|Melanoma in situ of skin|Melanoma in situ of skin
C0346081|T191|PT|254794007|SNOMEDCT_CORE|Angiosarcoma of skin|Angiosarcoma of skin
C0346081|T191|FN|254794007|SNOMEDCT_CORE|Angiosarcoma of skin|Angiosarcoma of skin
C0346156|T191|SY|269485000|SNOMEDCT_CORE|Benign neoplasm of breast|Benign tumor of breast
C0346156|T191|PT|269485000|SNOMEDCT_CORE|Benign tumor of breast|Benign tumor of breast
C0346156|T191|FN|269485000|SNOMEDCT_CORE|Benign tumor of breast|Benign tumor of breast
C0346156|T191|PTGB|269485000|SNOMEDCT_CORE|Benign tumour of breast|Benign tumor of breast
C0346186|T191|PT|119423009|SNOMEDCT_CORE|Benign teratoma of ovary|Benign teratoma of ovary
C0346186|T191|FN|119423009|SNOMEDCT_CORE|Benign teratoma of ovary|Benign teratoma of ovary
C0346186|T191|SY|119423009|SNOMEDCT_CORE|Ovarian mature cystic teratoma|Benign teratoma of ovary
C0346215|T046|IS|254902007|SNOMEDCT_CORE|Benign prostatic hypertroph without outflow obstruction|Benign prostatic hypertrophy without outflow obstruction
C0346215|T046|OF|254902007|SNOMEDCT_CORE|Benign prostatic hypertroph without outflow obstruction|Benign prostatic hypertrophy without outflow obstruction
C0346215|T046|PT|254902007|SNOMEDCT_CORE|Benign prostatic hypertrophy without outflow obstruction|Benign prostatic hypertrophy without outflow obstruction
C0346215|T046|FN|254902007|SNOMEDCT_CORE|Benign prostatic hypertrophy without outflow obstruction|Benign prostatic hypertrophy without outflow obstruction
C0346376|T191|SY|95711003|SNOMEDCT_CORE|Benign melanoma of iris|Nevus of iris
C0346376|T191|SYGB|95711003|SNOMEDCT_CORE|Iris naevus|Nevus of iris
C0346376|T191|SY|95711003|SNOMEDCT_CORE|Iris nevus|Nevus of iris
C0346376|T191|PTGB|95711003|SNOMEDCT_CORE|Naevus of iris|Nevus of iris
C0346376|T191|PT|95711003|SNOMEDCT_CORE|Nevus of iris|Nevus of iris
C0346376|T191|FN|95711003|SNOMEDCT_CORE|Nevus of iris|Nevus of iris
C0346388|T191|PT|255021005|SNOMEDCT_CORE|Malignant melanoma of choroid|Malignant melanoma of choroid
C0346388|T191|FN|255021005|SNOMEDCT_CORE|Malignant melanoma of choroid|Malignant melanoma of choroid
C0346392|T191|SY|255024002|SNOMEDCT_CORE|Benign melanoma of choroid|Nevus of choroid
C0346392|T191|SYGB|255024002|SNOMEDCT_CORE|Choroidal naevus|Nevus of choroid
C0346392|T191|SY|255024002|SNOMEDCT_CORE|Choroidal nevus|Nevus of choroid
C0346392|T191|PTGB|255024002|SNOMEDCT_CORE|Naevus of choroid|Nevus of choroid
C0346392|T191|PT|255024002|SNOMEDCT_CORE|Nevus of choroid|Nevus of choroid
C0346392|T191|FN|255024002|SNOMEDCT_CORE|Nevus of choroid|Nevus of choroid
C0346421|T191|SYGB|128835008|SNOMEDCT_CORE|Chronic eosinophilic leukaemia|Chronic eosinophilic leukemia
C0346421|T191|SY|128835008|SNOMEDCT_CORE|Chronic eosinophilic leukemia|Chronic eosinophilic leukemia
C0346455|T191|PT|94989005|SNOMEDCT_CORE|Neoplasm of uncertain behavior of parotid gland|Neoplasm of uncertain behavior of parotid gland
C0346455|T191|FN|94989005|SNOMEDCT_CORE|Neoplasm of uncertain behavior of parotid gland|Neoplasm of uncertain behavior of parotid gland
C0346455|T191|PTGB|94989005|SNOMEDCT_CORE|Neoplasm of uncertain behaviour of parotid gland|Neoplasm of uncertain behavior of parotid gland
C0346545|T191|PT|94963005|SNOMEDCT_CORE|Neoplasm of uncertain behavior of nervous system|Neoplasm of uncertain behavior of nervous system
C0346545|T191|FN|94963005|SNOMEDCT_CORE|Neoplasm of uncertain behavior of nervous system|Neoplasm of uncertain behavior of nervous system
C0346545|T191|IS|94963005|SNOMEDCT_CORE|Neoplasm of uncertain behavior of nervous system, NOS|Neoplasm of uncertain behavior of nervous system
C0346545|T191|PTGB|94963005|SNOMEDCT_CORE|Neoplasm of uncertain behaviour of nervous system|Neoplasm of uncertain behavior of nervous system
C0346564|T191|PT|271943005|SNOMEDCT_CORE|Carcinoma of base of tongue|Carcinoma of base of tongue
C0346564|T191|FN|271943005|SNOMEDCT_CORE|Carcinoma of base of tongue|Carcinoma of base of tongue
C0346619|T191|SY|187734007|SNOMEDCT_CORE|Gastroesophageal cancer|Malignant neoplasm of cardio-esophageal junction of stomach
C0346619|T191|PT|187734007|SNOMEDCT_CORE|Malignant neoplasm of cardio-esophageal junction of stomach|Malignant neoplasm of cardio-esophageal junction of stomach
C0346619|T191|PTGB|187734007|SNOMEDCT_CORE|Malignant neoplasm of cardio-oesophageal junction of stomach|Malignant neoplasm of cardio-esophageal junction of stomach
C0346619|T191|SY|187734007|SNOMEDCT_CORE|Malignant neoplasm of cardioesophageal junction of stomach|Malignant neoplasm of cardio-esophageal junction of stomach
C0346619|T191|FN|187734007|SNOMEDCT_CORE|Malignant neoplasm of cardioesophageal junction of stomach|Malignant neoplasm of cardio-esophageal junction of stomach
C0346619|T191|SY|187734007|SNOMEDCT_CORE|Malignant neoplasm of gastro-esophageal junction|Malignant neoplasm of cardio-esophageal junction of stomach
C0346619|T191|SYGB|187734007|SNOMEDCT_CORE|Malignant neoplasm of gastro-oesophageal junction|Malignant neoplasm of cardio-esophageal junction of stomach
C0346619|T191|SY|187734007|SNOMEDCT_CORE|Malignant neoplasm of gastroesophageal junction|Malignant neoplasm of cardio-esophageal junction of stomach
C0346619|T191|SY|187734007|SNOMEDCT_CORE|Malignant neoplasm of gastroesophageal junction of stomach|Malignant neoplasm of cardio-esophageal junction of stomach
C0346629|T191|SY|363510005|SNOMEDCT_CORE|CA - Cancer of large bowel|Malignant tumor of large intestine
C0346629|T191|SY|363510005|SNOMEDCT_CORE|Cancer of large bowel|Malignant tumor of large intestine
C0346629|T191|SY|363510005|SNOMEDCT_CORE|Cancer of large intestine|Malignant tumor of large intestine
C0346629|T191|IS|363510005|SNOMEDCT_CORE|Colorectal cancer|Malignant tumor of large intestine
C0346629|T191|PT|363510005|SNOMEDCT_CORE|Malignant tumor of large intestine|Malignant tumor of large intestine
C0346629|T191|FN|363510005|SNOMEDCT_CORE|Malignant tumor of large intestine|Malignant tumor of large intestine
C0346629|T191|PTGB|363510005|SNOMEDCT_CORE|Malignant tumour of large intestine|Malignant tumor of large intestine
C0346647|T191|SY|363418001|SNOMEDCT_CORE|CA - Cancer of pancreas|Malignant tumor of pancreas
C0346647|T191|SY|363418001|SNOMEDCT_CORE|CA - Pancreatic cancer|Malignant tumor of pancreas
C0346647|T191|PT|363418001|SNOMEDCT_CORE|Malignant tumor of pancreas|Malignant tumor of pancreas
C0346647|T191|FN|363418001|SNOMEDCT_CORE|Malignant tumor of pancreas|Malignant tumor of pancreas
C0346647|T191|PTGB|363418001|SNOMEDCT_CORE|Malignant tumour of pancreas|Malignant tumor of pancreas
C0346647|T191|SY|363418001|SNOMEDCT_CORE|Pancreatic cancer|Malignant tumor of pancreas
C0346773|T191|IS|188032002|SNOMEDCT_CORE|Malignant melanoma of ear and external auricular canal|Malignant melanoma of ear and/or external auditory canal
C0346773|T191|OF|188032002|SNOMEDCT_CORE|Malignant melanoma of ear and external auricular canal|Malignant melanoma of ear and/or external auditory canal
C0346773|T191|PT|188032002|SNOMEDCT_CORE|Malignant melanoma of ear and/or external auditory canal|Malignant melanoma of ear and/or external auditory canal
C0346773|T191|FN|188032002|SNOMEDCT_CORE|Malignant melanoma of ear and/or external auditory canal|Malignant melanoma of ear and/or external auditory canal
C0346773|T191|OF|188032002|SNOMEDCT_CORE|Malignant melanoma of ear and/or external auricular canal|Malignant melanoma of ear and/or external auditory canal
C0346773|T191|SY|188032002|SNOMEDCT_CORE|Malignant melanoma of ear and/or external auricular canal|Malignant melanoma of ear and/or external auditory canal
C0346782|T191|IS|188044004|SNOMEDCT_CORE|Malignant melanoma of scalp and neck|Malignant melanoma of scalp and/or neck
C0346782|T191|OF|188044004|SNOMEDCT_CORE|Malignant melanoma of scalp and neck|Malignant melanoma of scalp and/or neck
C0346782|T191|PT|188044004|SNOMEDCT_CORE|Malignant melanoma of scalp and/or neck|Malignant melanoma of scalp and/or neck
C0346782|T191|FN|188044004|SNOMEDCT_CORE|Malignant melanoma of scalp and/or neck|Malignant melanoma of scalp and/or neck
C0346782|T191|OF|188044004|SNOMEDCT_CORE|Malignant melanoma of scalp AND/OR neck|Malignant melanoma of scalp and/or neck
C0346794|T191|PT|188060000|SNOMEDCT_CORE|Malignant melanoma of shoulder|Malignant melanoma of shoulder
C0346794|T191|FN|188060000|SNOMEDCT_CORE|Malignant melanoma of shoulder|Malignant melanoma of shoulder
C0346795|T191|PT|188061001|SNOMEDCT_CORE|Malignant melanoma of upper arm|Malignant melanoma of upper arm
C0346795|T191|FN|188061001|SNOMEDCT_CORE|Malignant melanoma of upper arm|Malignant melanoma of upper arm
C0346808|T191|PT|188075008|SNOMEDCT_CORE|Malignant melanoma of foot|Malignant melanoma of foot
C0346808|T191|FN|188075008|SNOMEDCT_CORE|Malignant melanoma of foot|Malignant melanoma of foot
C0346836|T191|PT|187999008|SNOMEDCT_CORE|Malignant neoplasm of connective and soft tissue of hip and lower limb|Malignant neoplasm of connective and soft tissue of hip and lower limb
C0346836|T191|FN|187999008|SNOMEDCT_CORE|Malignant neoplasm of connective and soft tissue of hip and lower limb|Malignant neoplasm of connective and soft tissue of hip and lower limb
C0346957|T191|SY|405843009|SNOMEDCT_CORE|CA - Disseminated cancer|Widespread metastatic malignant neoplastic disease
C0346957|T191|SY|405843009|SNOMEDCT_CORE|Disseminated cancer|Widespread metastatic malignant neoplastic disease
C0346957|T191|SY|405843009|SNOMEDCT_CORE|Disseminated malignancy|Widespread metastatic malignant neoplastic disease
C0346957|T191|SYGB|405843009|SNOMEDCT_CORE|Generalised cancer|Widespread metastatic malignant neoplastic disease
C0346957|T191|SYGB|405843009|SNOMEDCT_CORE|Generalised malignancy|Widespread metastatic malignant neoplastic disease
C0346957|T191|SY|405843009|SNOMEDCT_CORE|Generalized cancer|Widespread metastatic malignant neoplastic disease
C0346957|T191|SY|405843009|SNOMEDCT_CORE|Generalized malignancy|Widespread metastatic malignant neoplastic disease
C0346957|T191|SY|405843009|SNOMEDCT_CORE|Malignant neoplasm, disseminated|Widespread metastatic malignant neoplastic disease
C0346957|T191|FN|405843009|SNOMEDCT_CORE|Widespread metastatic malignant neoplastic disease|Widespread metastatic malignant neoplastic disease
C0346957|T191|PT|405843009|SNOMEDCT_CORE|Widespread metastatic malignant neoplastic disease|Widespread metastatic malignant neoplastic disease
C0346973|T191|SY|94365007|SNOMEDCT_CORE|Cancer metastatic to large intestine|Secondary malignant neoplasm of large intestine
C0346973|T191|SY|94365007|SNOMEDCT_CORE|Metastasis to large intestine|Secondary malignant neoplasm of large intestine
C0346973|T191|SY|94365007|SNOMEDCT_CORE|Metastatic malignant neoplasm to large intestine|Secondary malignant neoplasm of large intestine
C0346973|T191|IS|94365007|SNOMEDCT_CORE|Metastatic malignant neoplasm to large intestine, NOS|Secondary malignant neoplasm of large intestine
C0346973|T191|PT|94365007|SNOMEDCT_CORE|Secondary malignant neoplasm of large intestine|Secondary malignant neoplasm of large intestine
C0346973|T191|FN|94365007|SNOMEDCT_CORE|Secondary malignant neoplasm of large intestine|Secondary malignant neoplasm of large intestine
C0346973|T191|IS|94365007|SNOMEDCT_CORE|Secondary malignant neoplasm of large intestine, NOS|Secondary malignant neoplasm of large intestine
C0346974|T191|SY|94260004|SNOMEDCT_CORE|Metastatic malignant neoplasm to colon|Secondary malignant neoplasm of colon
C0346974|T191|IS|94260004|SNOMEDCT_CORE|Metastatic malignant neoplasm to colon, NOS|Secondary malignant neoplasm of colon
C0346974|T191|PT|94260004|SNOMEDCT_CORE|Secondary malignant neoplasm of colon|Secondary malignant neoplasm of colon
C0346974|T191|FN|94260004|SNOMEDCT_CORE|Secondary malignant neoplasm of colon|Secondary malignant neoplasm of colon
C0346974|T191|IS|94260004|SNOMEDCT_CORE|Secondary malignant neoplasm of colon, NOS|Secondary malignant neoplasm of colon
C0346975|T191|SY|94513006|SNOMEDCT_CORE|Cancer metastatic to rectum|Secondary malignant neoplasm of rectum
C0346975|T191|SY|94513006|SNOMEDCT_CORE|Metastatic malignant neoplasm to rectum|Secondary malignant neoplasm of rectum
C0346975|T191|PT|94513006|SNOMEDCT_CORE|Secondary malignant neoplasm of rectum|Secondary malignant neoplasm of rectum
C0346975|T191|FN|94513006|SNOMEDCT_CORE|Secondary malignant neoplasm of rectum|Secondary malignant neoplasm of rectum
C0346976|T191|SY|94459006|SNOMEDCT_CORE|Cancer metastatic to pancreas|Secondary malignant neoplasm of pancreas
C0346976|T191|SY|94459006|SNOMEDCT_CORE|Metastasis to pancreas|Secondary malignant neoplasm of pancreas
C0346976|T191|SY|94459006|SNOMEDCT_CORE|Metastatic malignant neoplasm to pancreas|Secondary malignant neoplasm of pancreas
C0346976|T191|IS|94459006|SNOMEDCT_CORE|Metastatic malignant neoplasm to pancreas, NOS|Secondary malignant neoplasm of pancreas
C0346976|T191|SY|94459006|SNOMEDCT_CORE|Pancreatic metastasis|Secondary malignant neoplasm of pancreas
C0346976|T191|SY|94459006|SNOMEDCT_CORE|Secondary malignant deposit in pancreas|Secondary malignant neoplasm of pancreas
C0346976|T191|PT|94459006|SNOMEDCT_CORE|Secondary malignant neoplasm of pancreas|Secondary malignant neoplasm of pancreas
C0346976|T191|FN|94459006|SNOMEDCT_CORE|Secondary malignant neoplasm of pancreas|Secondary malignant neoplasm of pancreas
C0346976|T191|IS|94459006|SNOMEDCT_CORE|Secondary malignant neoplasm of pancreas, NOS|Secondary malignant neoplasm of pancreas
C0346989|T191|SY|94627008|SNOMEDCT_CORE|Cancer metastatic to peritoneum|Secondary malignant neoplasm of peritoneum
C0346989|T191|SY|94627008|SNOMEDCT_CORE|Metastasis to peritoneum|Secondary malignant neoplasm of peritoneum
C0346989|T191|SY|94627008|SNOMEDCT_CORE|Metastatic malignant neoplasm to peritoneum|Secondary malignant neoplasm of peritoneum
C0346989|T191|IS|94627008|SNOMEDCT_CORE|Metastatic malignant neoplasm to the peritoneum|Secondary malignant neoplasm of peritoneum
C0346989|T191|IS|94627008|SNOMEDCT_CORE|Metastatic malignant neoplasm to the peritoneum, NOS|Secondary malignant neoplasm of peritoneum
C0346989|T191|SY|94627008|SNOMEDCT_CORE|Peritoneal seedling|Secondary malignant neoplasm of peritoneum
C0346989|T191|PT|94627008|SNOMEDCT_CORE|Secondary malignant neoplasm of peritoneum|Secondary malignant neoplasm of peritoneum
C0346989|T191|FN|94627008|SNOMEDCT_CORE|Secondary malignant neoplasm of peritoneum|Secondary malignant neoplasm of peritoneum
C0346989|T191|OP|94627008|SNOMEDCT_CORE|Secondary malignant neoplasm of the peritoneum|Secondary malignant neoplasm of peritoneum
C0346989|T191|OF|94627008|SNOMEDCT_CORE|Secondary malignant neoplasm of the peritoneum|Secondary malignant neoplasm of peritoneum
C0346989|T191|IS|94627008|SNOMEDCT_CORE|Secondary malignant neoplasm of the peritoneum, NOS|Secondary malignant neoplasm of peritoneum
C0346989|T191|SY|94627008|SNOMEDCT_CORE|Secondary malignant peritoneal deposit|Secondary malignant neoplasm of peritoneum
C0346992|T191|SY|94628003|SNOMEDCT_CORE|Metastasis to retroperitoneum|Secondary malignant neoplasm of retroperitoneum
C0346992|T191|SY|94628003|SNOMEDCT_CORE|Metastatic malignant neoplasm to the retroperitoneum|Secondary malignant neoplasm of retroperitoneum
C0346992|T191|SY|94628003|SNOMEDCT_CORE|Retroperitoneal metastasis|Secondary malignant neoplasm of retroperitoneum
C0346992|T191|PT|94628003|SNOMEDCT_CORE|Secondary malignant neoplasm of retroperitoneum|Secondary malignant neoplasm of retroperitoneum
C0346992|T191|FN|94628003|SNOMEDCT_CORE|Secondary malignant neoplasm of retroperitoneum|Secondary malignant neoplasm of retroperitoneum
C0346992|T191|SY|94628003|SNOMEDCT_CORE|Secondary malignant neoplasm of the retroperitoneum|Secondary malignant neoplasm of retroperitoneum
C0346992|T191|OF|94628003|SNOMEDCT_CORE|Secondary malignant neoplasm of the retroperitoneum|Secondary malignant neoplasm of retroperitoneum
C0346993|T191|SY|94297009|SNOMEDCT_CORE|Metastasis to breast|Secondary malignant neoplasm of female breast
C0346993|T191|SY|94297009|SNOMEDCT_CORE|Metastatic malignant neoplasm to female breast|Secondary malignant neoplasm of female breast
C0346993|T191|IS|94297009|SNOMEDCT_CORE|Metastatic malignant neoplasm to female breast, NOS|Secondary malignant neoplasm of female breast
C0346993|T191|SY|94297009|SNOMEDCT_CORE|Secondary malignant deposit to breast|Secondary malignant neoplasm of female breast
C0346993|T191|SY|94297009|SNOMEDCT_CORE|Secondary malignant neoplasm of breast|Secondary malignant neoplasm of female breast
C0346993|T191|PT|94297009|SNOMEDCT_CORE|Secondary malignant neoplasm of female breast|Secondary malignant neoplasm of female breast
C0346993|T191|FN|94297009|SNOMEDCT_CORE|Secondary malignant neoplasm of female breast|Secondary malignant neoplasm of female breast
C0346993|T191|IS|94297009|SNOMEDCT_CORE|Secondary malignant neoplasm of female breast, NOS|Secondary malignant neoplasm of female breast
C0347001|T191|SY|94503003|SNOMEDCT_CORE|Cancer metastatic to prostate|Secondary malignant neoplasm of prostate
C0347001|T191|SY|94503003|SNOMEDCT_CORE|Metastasis to prostate|Secondary malignant neoplasm of prostate
C0347001|T191|SY|94503003|SNOMEDCT_CORE|Metastatic malignant neoplasm to prostate|Secondary malignant neoplasm of prostate
C0347001|T191|SY|94503003|SNOMEDCT_CORE|Metastatic tumor to prostate|Secondary malignant neoplasm of prostate
C0347001|T191|SYGB|94503003|SNOMEDCT_CORE|Metastatic tumour to prostate|Secondary malignant neoplasm of prostate
C0347001|T191|PT|94503003|SNOMEDCT_CORE|Secondary malignant neoplasm of prostate|Secondary malignant neoplasm of prostate
C0347001|T191|FN|94503003|SNOMEDCT_CORE|Secondary malignant neoplasm of prostate|Secondary malignant neoplasm of prostate
C0347003|T191|SY|94623007|SNOMEDCT_CORE|Metastasis to testis|Secondary malignant neoplasm of testis
C0347003|T191|SY|94623007|SNOMEDCT_CORE|Metastatic malignant neoplasm to testis|Secondary malignant neoplasm of testis
C0347003|T191|IS|94623007|SNOMEDCT_CORE|Metastatic malignant neoplasm to testis, NOS|Secondary malignant neoplasm of testis
C0347003|T191|SY|94623007|SNOMEDCT_CORE|Metastatic tumor to testis|Secondary malignant neoplasm of testis
C0347003|T191|SYGB|94623007|SNOMEDCT_CORE|Metastatic tumour to testis|Secondary malignant neoplasm of testis
C0347003|T191|PT|94623007|SNOMEDCT_CORE|Secondary malignant neoplasm of testis|Secondary malignant neoplasm of testis
C0347003|T191|FN|94623007|SNOMEDCT_CORE|Secondary malignant neoplasm of testis|Secondary malignant neoplasm of testis
C0347003|T191|IS|94623007|SNOMEDCT_CORE|Secondary malignant neoplasm of testis, NOS|Secondary malignant neoplasm of testis
C0347011|T191|SY|94186002|SNOMEDCT_CORE|Cancer metastatic to urinary bladder|Secondary malignant neoplasm of bladder
C0347011|T191|SY|94186002|SNOMEDCT_CORE|Metastasis to bladder|Secondary malignant neoplasm of bladder
C0347011|T191|SY|94186002|SNOMEDCT_CORE|Metastatic malignant neoplasm to bladder|Secondary malignant neoplasm of bladder
C0347011|T191|IS|94186002|SNOMEDCT_CORE|Metastatic malignant neoplasm to bladder, NOS|Secondary malignant neoplasm of bladder
C0347011|T191|SY|94186002|SNOMEDCT_CORE|Metastatic tumor to bladder|Secondary malignant neoplasm of bladder
C0347011|T191|SYGB|94186002|SNOMEDCT_CORE|Metastatic tumour to bladder|Secondary malignant neoplasm of bladder
C0347011|T191|PT|94186002|SNOMEDCT_CORE|Secondary malignant neoplasm of bladder|Secondary malignant neoplasm of bladder
C0347011|T191|FN|94186002|SNOMEDCT_CORE|Secondary malignant neoplasm of bladder|Secondary malignant neoplasm of bladder
C0347011|T191|IS|94186002|SNOMEDCT_CORE|Secondary malignant neoplasm of bladder, NOS|Secondary malignant neoplasm of bladder
C0347021|T191|SY|94254004|SNOMEDCT_CORE|Cancer metastatic to choroid|Secondary malignant neoplasm of choroid
C0347021|T191|SY|94254004|SNOMEDCT_CORE|Metastasis to choroid|Secondary malignant neoplasm of choroid
C0347021|T191|SY|94254004|SNOMEDCT_CORE|Metastatic malignant neoplasm to choroid|Secondary malignant neoplasm of choroid
C0347021|T191|SY|94254004|SNOMEDCT_CORE|Secondary choroidal tumor|Secondary malignant neoplasm of choroid
C0347021|T191|SYGB|94254004|SNOMEDCT_CORE|Secondary choroidal tumour|Secondary malignant neoplasm of choroid
C0347021|T191|PT|94254004|SNOMEDCT_CORE|Secondary malignant neoplasm of choroid|Secondary malignant neoplasm of choroid
C0347021|T191|FN|94254004|SNOMEDCT_CORE|Secondary malignant neoplasm of choroid|Secondary malignant neoplasm of choroid
C0347197|T191|PT|419645003|SNOMEDCT_CORE|Benign neoplasm of oral cavity|Benign neoplasm of oral cavity
C0347197|T191|FN|419645003|SNOMEDCT_CORE|Benign neoplasm of oral cavity|Benign neoplasm of oral cavity
C0347197|T191|SY|419645003|SNOMEDCT_CORE|Benign tumor of oral cavity|Benign neoplasm of oral cavity
C0347197|T191|SYGB|419645003|SNOMEDCT_CORE|Benign tumour of oral cavity|Benign neoplasm of oral cavity
C0347197|T191|SY|419645003|SNOMEDCT_CORE|Oral benign tumor|Benign neoplasm of oral cavity
C0347197|T191|SYGB|419645003|SNOMEDCT_CORE|Oral benign tumour|Benign neoplasm of oral cavity
C0347210|T191|PT|271472001|SNOMEDCT_CORE|Benign neoplasm of nose, middle ear and accessory sinuses|Benign neoplasm of nose, middle ear and accessory sinuses
C0347210|T191|FN|271472001|SNOMEDCT_CORE|Benign neoplasm of nose, middle ear and accessory sinuses|Benign neoplasm of nose, middle ear and accessory sinuses
C0347266|T191|SY|73861008|SNOMEDCT_CORE|Duodenal polyp|Polyp of duodenum
C0347266|T191|PT|73861008|SNOMEDCT_CORE|Polyp of duodenum|Polyp of duodenum
C0347266|T191|FN|73861008|SNOMEDCT_CORE|Polyp of duodenum|Polyp of duodenum
C0347284|T191|PT|92264007|SNOMEDCT_CORE|Benign neoplasm of pancreas|Benign neoplasm of pancreas
C0347284|T191|FN|92264007|SNOMEDCT_CORE|Benign neoplasm of pancreas|Benign neoplasm of pancreas
C0347284|T191|IS|92264007|SNOMEDCT_CORE|Benign neoplasm of pancreas, NOS|Benign neoplasm of pancreas
C0347284|T191|SY|92264007|SNOMEDCT_CORE|Benign tumor of pancreas|Benign neoplasm of pancreas
C0347284|T191|SYGB|92264007|SNOMEDCT_CORE|Benign tumour of pancreas|Benign neoplasm of pancreas
C0347353|T191|OAP|271477007|SNOMEDCT_CORE|Benign neoplasm of skin of ear and external auditory meatus|Benign neoplasm of skin of ear and external auditory meatus
C0347353|T191|OAF|271477007|SNOMEDCT_CORE|Benign neoplasm of skin of ear and external auditory meatus|Benign neoplasm of skin of ear and external auditory meatus
C0347354|T191|PT|255181009|SNOMEDCT_CORE|Benign neoplasm of ear|Benign neoplasm of ear
C0347354|T191|FN|255181009|SNOMEDCT_CORE|Benign neoplasm of ear|Benign neoplasm of ear
C0347365|T191|PT|92359006|SNOMEDCT_CORE|Benign neoplasm of skin of face|Benign neoplasm of skin of face
C0347365|T191|FN|92359006|SNOMEDCT_CORE|Benign neoplasm of skin of face|Benign neoplasm of skin of face
C0347365|T191|IS|92359006|SNOMEDCT_CORE|Benign neoplasm of skin of face, NOS|Benign neoplasm of skin of face
C0347366|T191|SY|92375009|SNOMEDCT_CORE|Benign neoplasm of scalp|Benign neoplasm of skin of scalp
C0347366|T191|PT|92375009|SNOMEDCT_CORE|Benign neoplasm of skin of scalp|Benign neoplasm of skin of scalp
C0347366|T191|FN|92375009|SNOMEDCT_CORE|Benign neoplasm of skin of scalp|Benign neoplasm of skin of scalp
C0347367|T191|PT|92371000|SNOMEDCT_CORE|Benign neoplasm of skin of neck|Benign neoplasm of skin of neck
C0347367|T191|FN|92371000|SNOMEDCT_CORE|Benign neoplasm of skin of neck|Benign neoplasm of skin of neck
C0347378|T191|PT|92376005|SNOMEDCT_CORE|Benign neoplasm of skin of shoulder|Benign neoplasm of skin of shoulder
C0347378|T191|FN|92376005|SNOMEDCT_CORE|Benign neoplasm of skin of shoulder|Benign neoplasm of skin of shoulder
C0347382|T191|SY|92370004|SNOMEDCT_CORE|Benign neoplasm of skin of leg|Benign neoplasm of skin of lower limb
C0347382|T191|PT|92370004|SNOMEDCT_CORE|Benign neoplasm of skin of lower limb|Benign neoplasm of skin of lower limb
C0347382|T191|FN|92370004|SNOMEDCT_CORE|Benign neoplasm of skin of lower limb|Benign neoplasm of skin of lower limb
C0347382|T191|IS|92370004|SNOMEDCT_CORE|Benign neoplasm of skin of lower limb, NOS|Benign neoplasm of skin of lower limb
C0347390|T191|PT|255184001|SNOMEDCT_CORE|Papilloma of skin|Papilloma of skin
C0347390|T191|FN|255184001|SNOMEDCT_CORE|Papilloma of skin|Papilloma of skin
C0347394|T191|PT|255187008|SNOMEDCT_CORE|Lipoma of skin|Lipoma of skin
C0347394|T191|FN|255187008|SNOMEDCT_CORE|Lipoma of skin|Lipoma of skin
C0347426|T191|SY|93160004|SNOMEDCT_CORE|Lipoma of neck|Lipoma of skin and subcutaneous tissue of neck
C0347426|T191|PT|93160004|SNOMEDCT_CORE|Lipoma of skin and subcutaneous tissue of neck|Lipoma of skin and subcutaneous tissue of neck
C0347426|T191|FN|93160004|SNOMEDCT_CORE|Lipoma of skin and subcutaneous tissue of neck|Lipoma of skin and subcutaneous tissue of neck
C0347493|T191|SY|255196008|SNOMEDCT_CORE|Adenomatous polyp - cervix uteri|Adenomatous polyp of cervix
C0347493|T191|OF|255196008|SNOMEDCT_CORE|Adenomatous polyp - cervix uteri|Adenomatous polyp of cervix
C0347493|T191|OAP|60535003|SNOMEDCT_CORE|Adenomatous polyp of cervix|Adenomatous polyp of cervix
C0347493|T191|PT|255196008|SNOMEDCT_CORE|Adenomatous polyp of cervix|Adenomatous polyp of cervix
C0347493|T191|OAF|60535003|SNOMEDCT_CORE|Adenomatous polyp of cervix|Adenomatous polyp of cervix
C0347493|T191|SY|255196008|SNOMEDCT_CORE|Adenomatous polyp of cervix uteri|Adenomatous polyp of cervix
C0347493|T191|FN|255196008|SNOMEDCT_CORE|Adenomatous polyp of cervix uteri|Adenomatous polyp of cervix
C0347493|T191|OAS|60535003|SNOMEDCT_CORE|Cervical adenomatous polyp|Adenomatous polyp of cervix
C0347525|T191|PT|271479005|SNOMEDCT_CORE|Benign neoplasm of pituitary gland and craniopharyngeal duct|Benign neoplasm of pituitary gland and craniopharyngeal duct
C0347525|T191|FN|271479005|SNOMEDCT_CORE|Benign neoplasm of pituitary gland and craniopharyngeal duct|Benign neoplasm of pituitary gland and craniopharyngeal duct
C0347535|T037|PT|127296001|SNOMEDCT_CORE|Intracranial injury|Intracranial injury
C0347535|T037|FN|127296001|SNOMEDCT_CORE|Intracranial injury|Intracranial injury
C0347544|T037|PT|283033008|SNOMEDCT_CORE|Superficial injury of forearm|Superficial injury of forearm
C0347544|T037|FN|283033008|SNOMEDCT_CORE|Superficial injury of forearm|Superficial injury of forearm
C0347545|T037|PT|274192001|SNOMEDCT_CORE|Superficial injury of wrist|Superficial injury of wrist
C0347545|T037|FN|274192001|SNOMEDCT_CORE|Superficial injury of wrist|Superficial injury of wrist
C0347573|T037|PT|125663008|SNOMEDCT_CORE|Open wound of foot|Open wound of foot
C0347573|T037|FN|125663008|SNOMEDCT_CORE|Open wound of foot|Open wound of foot
C0347575|T037|PT|275320004|SNOMEDCT_CORE|Injury of nail|Injury of nail
C0347575|T037|FN|275320004|SNOMEDCT_CORE|Injury of nail|Injury of nail
C0347577|T037|SY|262581006|SNOMEDCT_CORE|Burn of head|Head burn
C0347577|T037|SY|262581006|SNOMEDCT_CORE|Head - burn|Head burn
C0347577|T037|PT|262581006|SNOMEDCT_CORE|Head burn|Head burn
C0347577|T037|FN|262581006|SNOMEDCT_CORE|Head burn|Head burn
C0347577|T037|IS|262581006|SNOMEDCT_CORE|Head burns|Head burn
C0347577|T037|OF|262581006|SNOMEDCT_CORE|Head burns|Head burn
C0347584|T037|PT|95855003|SNOMEDCT_CORE|Traumatic amputation of finger|Traumatic amputation of finger
C0347584|T037|FN|95855003|SNOMEDCT_CORE|Traumatic amputation of finger|Traumatic amputation of finger
C0347584|T037|IS|95855003|SNOMEDCT_CORE|Traumatic amputation of finger, NOS|Traumatic amputation of finger
C0347620|T037|SY|3903005|SNOMEDCT_CORE|Closed traumatic pneumothorax|Traumatic pneumothorax without open wound into thorax
C0347620|T037|PT|3903005|SNOMEDCT_CORE|Traumatic pneumothorax without open wound into thorax|Traumatic pneumothorax without open wound into thorax
C0347620|T037|FN|3903005|SNOMEDCT_CORE|Traumatic pneumothorax without open wound into thorax|Traumatic pneumothorax without open wound into thorax
C0347633|T037|SY|262802005|SNOMEDCT_CORE|Hepatic laceration|Laceration of liver
C0347633|T037|PT|262802005|SNOMEDCT_CORE|Laceration of liver|Laceration of liver
C0347633|T037|FN|262802005|SNOMEDCT_CORE|Laceration of liver|Laceration of liver
C0347656|T037|SY|110015006|SNOMEDCT_CORE|Injuries of penis|Injury of penis
C0347656|T037|OF|110015006|SNOMEDCT_CORE|Injuries of penis|Injury of penis
C0347656|T037|PT|110015006|SNOMEDCT_CORE|Injury of penis|Injury of penis
C0347656|T037|FN|110015006|SNOMEDCT_CORE|Injury of penis|Injury of penis
C0347721|T037|IS|262965006|SNOMEDCT_CORE|Back strain|Strain of back muscle
C0347721|T037|IS|262965006|SNOMEDCT_CORE|Strain of back|Strain of back muscle
C0347721|T037|PT|262965006|SNOMEDCT_CORE|Strain of back muscle|Strain of back muscle
C0347721|T037|FN|262965006|SNOMEDCT_CORE|Strain of back muscle|Strain of back muscle
C0347775|T037|PT|263167007|SNOMEDCT_CORE|Blow out fracture of orbit|Blow out fracture of orbit
C0347775|T037|FN|263167007|SNOMEDCT_CORE|Blow out fracture of orbit|Blow out fracture of orbit
C0347775|T037|SY|263167007|SNOMEDCT_CORE|Blowout fracture of orbit|Blow out fracture of orbit
C0347780|T037|PT|125607007|SNOMEDCT_CORE|Fracture of thoracic spine|Fracture of thoracic spine
C0347780|T037|FN|125607007|SNOMEDCT_CORE|Fracture of thoracic spine|Fracture of thoracic spine
C0347780|T037|SY|125607007|SNOMEDCT_CORE|Fracture of thoracic vertebra|Fracture of thoracic spine
C0347781|T037|PT|207938004|SNOMEDCT_CORE|Closed fracture thoracic vertebra|Closed fracture thoracic vertebra
C0347781|T037|FN|207938004|SNOMEDCT_CORE|Closed fracture thoracic vertebra|Closed fracture thoracic vertebra
C0347804|T037|PT|64455005|SNOMEDCT_CORE|Fracture of acetabulum|Fracture of acetabulum
C0347804|T037|FN|64455005|SNOMEDCT_CORE|Fracture of acetabulum|Fracture of acetabulum
C0347804|T037|IS|64455005|SNOMEDCT_CORE|Fracture of acetabulum, NOS|Fracture of acetabulum
C0347854|T047|FN|186150001|SNOMEDCT_CORE|Enteritis caused by rotavirus|Enteritis due to rotavirus
C0347854|T047|SY|186150001|SNOMEDCT_CORE|Enteritis caused by rotavirus|Enteritis due to rotavirus
C0347854|T047|PT|186150001|SNOMEDCT_CORE|Enteritis due to rotavirus|Enteritis due to rotavirus
C0347854|T047|OF|186150001|SNOMEDCT_CORE|Enteritis due to rotavirus|Enteritis due to rotavirus
C0347854|T047|SY|186150001|SNOMEDCT_CORE|Rotavirus enteritis|Enteritis due to rotavirus
C0347887|T047|PT|42861008|SNOMEDCT_CORE|Thrombophlebitis of iliac vein|Thrombophlebitis of iliac vein
C0347887|T047|FN|42861008|SNOMEDCT_CORE|Thrombophlebitis of iliac vein|Thrombophlebitis of iliac vein
C0347940|T033|PT|274739003|SNOMEDCT_CORE|Chest swelling|Chest swelling
C0347940|T033|FN|274739003|SNOMEDCT_CORE|Chest swelling|Chest swelling
C0347941|T033|SY|440299000|SNOMEDCT_CORE|Chest mass|Chest mass
C0347943|T033|IS|74285003|SNOMEDCT_CORE|Pelvic swelling|Pelvic swelling
C0347943|T033|IS|74285003|SNOMEDCT_CORE|Pelvic swelling, NOS|Pelvic swelling
C0347944|T033|FN|74285003|SNOMEDCT_CORE|Mass of pelvic structure|Pelvic mass
C0347944|T033|SY|74285003|SNOMEDCT_CORE|Mass of pelvic structure|Pelvic mass
C0347944|T033|SY|74285003|SNOMEDCT_CORE|Pelvic lump|Pelvic mass
C0347944|T033|IS|74285003|SNOMEDCT_CORE|Pelvic lump, NOS|Pelvic mass
C0347944|T033|PT|74285003|SNOMEDCT_CORE|Pelvic mass|Pelvic mass
C0347944|T033|OF|74285003|SNOMEDCT_CORE|Pelvic mass|Pelvic mass
C0347944|T033|IS|74285003|SNOMEDCT_CORE|Pelvic mass, NOS|Pelvic mass
C0347952|T037|SY|428883008|SNOMEDCT_CORE|Rupture biceps tendon|Rupture of tendon of biceps
C0347952|T037|SY|428883008|SNOMEDCT_CORE|Rupture of biceps tendon|Rupture of tendon of biceps
C0347952|T037|PT|428883008|SNOMEDCT_CORE|Rupture of tendon of biceps|Rupture of tendon of biceps
C0347952|T037|FN|428883008|SNOMEDCT_CORE|Rupture of tendon of biceps|Rupture of tendon of biceps
C0347952|T037|SY|428883008|SNOMEDCT_CORE|Tear of biceps tendon|Rupture of tendon of biceps
C0347971|T037|PT|309710005|SNOMEDCT_CORE|Lumbosacral strain|Lumbosacral strain
C0347971|T037|FN|309710005|SNOMEDCT_CORE|Lumbosacral strain|Lumbosacral strain
C0348024|T046|PT|264580006|SNOMEDCT_CORE|Thyroid dysfunction|Thyroid dysfunction
C0348024|T046|FN|264580006|SNOMEDCT_CORE|Thyroid dysfunction|Thyroid dysfunction
C0348083|T190|PT|261827001|SNOMEDCT_CORE|High anal fistula|High anal fistula
C0348083|T190|FN|261827001|SNOMEDCT_CORE|High anal fistula|High anal fistula
C0348426|T191|PT|109913001|SNOMEDCT_CORE|Benign neoplasm of meninges|Benign neoplasm of meninges
C0348426|T191|FN|109913001|SNOMEDCT_CORE|Benign neoplasm of meninges|Benign neoplasm of meninges
C0348426|T191|SY|109913001|SNOMEDCT_CORE|Benign tumor of meninges|Benign neoplasm of meninges
C0348426|T191|SYGB|109913001|SNOMEDCT_CORE|Benign tumour of meninges|Benign neoplasm of meninges
C0348593|T047|SY|194856005|SNOMEDCT_CORE|Reinfarction of myocardium|Subsequent myocardial infarction
C0348593|T047|PT|194856005|SNOMEDCT_CORE|Subsequent myocardial infarction|Subsequent myocardial infarction
C0348593|T047|FN|194856005|SNOMEDCT_CORE|Subsequent myocardial infarction|Subsequent myocardial infarction
C0348799|T047|FN|195739001|SNOMEDCT_CORE|Acute bronchiolitis caused by respiratory syncytial virus|Acute bronchiolitis due to respiratory syncytial virus
C0348799|T047|SY|195739001|SNOMEDCT_CORE|Acute bronchiolitis caused by respiratory syncytial virus|Acute bronchiolitis due to respiratory syncytial virus
C0348799|T047|PT|195739001|SNOMEDCT_CORE|Acute bronchiolitis due to respiratory syncytial virus|Acute bronchiolitis due to respiratory syncytial virus
C0348799|T047|OF|195739001|SNOMEDCT_CORE|Acute bronchiolitis due to respiratory syncytial virus|Acute bronchiolitis due to respiratory syncytial virus
C0348809|T047|PT|186193001|SNOMEDCT_CORE|Tuberculosis of lung, confirmed by sputum microscopy with or without culture|Tuberculosis of lung, confirmed by sputum microscopy with or without culture
C0348809|T047|FN|186193001|SNOMEDCT_CORE|Tuberculosis of lung, confirmed by sputum microscopy with or without culture|Tuberculosis of lung, confirmed by sputum microscopy with or without culture
C0348810|T047|PT|186194007|SNOMEDCT_CORE|Tuberculosis of lung, confirmed by culture only|Tuberculosis of lung, confirmed by culture only
C0348810|T047|FN|186194007|SNOMEDCT_CORE|Tuberculosis of lung, confirmed by culture only|Tuberculosis of lung, confirmed by culture only
C0348811|T047|PT|186195008|SNOMEDCT_CORE|Tuberculosis of lung, confirmed histologically|Tuberculosis of lung, confirmed histologically
C0348811|T047|FN|186195008|SNOMEDCT_CORE|Tuberculosis of lung, confirmed histologically|Tuberculosis of lung, confirmed histologically
C0348818|T047|PT|196001008|SNOMEDCT_CORE|Chronic obstructive pulmonary disease with acute lower respiratory infection|Chronic obstructive pulmonary disease with acute lower respiratory infection
C0348818|T047|FN|196001008|SNOMEDCT_CORE|Chronic obstructive pulmonary disease with acute lower respiratory infection|Chronic obstructive pulmonary disease with acute lower respiratory infection
C0348860|T047|OAP|194774006|SNOMEDCT_CORE|Hypertensive renal disease with renal failure|Hypertensive renal disease with renal failure
C0348860|T047|OAF|194774006|SNOMEDCT_CORE|Hypertensive renal disease with renal failure|Hypertensive renal disease with renal failure
C0348879|T047|PT|194780003|SNOMEDCT_CORE|Hypertensive heart and renal disease with renal failure|Hypertensive heart and renal disease with renal failure
C0348879|T047|FN|194780003|SNOMEDCT_CORE|Hypertensive heart and renal disease with renal failure|Hypertensive heart and renal disease with renal failure
C0348919|T047|SY|422099009|SNOMEDCT_CORE|Diabetic oculopathy associated with type 2 diabetes mellitus|Disorder of eye due to type 2 diabetes mellitus
C0348919|T047|OF|422099009|SNOMEDCT_CORE|Diabetic oculopathy associated with type II diabetes mellitus|Disorder of eye due to type 2 diabetes mellitus
C0348919|T047|SY|422099009|SNOMEDCT_CORE|Diabetic oculopathy associated with type II diabetes mellitus|Disorder of eye due to type 2 diabetes mellitus
C0348919|T047|OF|422099009|SNOMEDCT_CORE|Disorder of eye co-occurrent and due to type 2 diabetes mellitus|Disorder of eye due to type 2 diabetes mellitus
C0348919|T047|IS|422099009|SNOMEDCT_CORE|Disorder of eye co-occurrent and due to type 2 diabetes mellitus|Disorder of eye due to type 2 diabetes mellitus
C0348919|T047|PT|422099009|SNOMEDCT_CORE|Disorder of eye due to type 2 diabetes mellitus|Disorder of eye due to type 2 diabetes mellitus
C0348919|T047|FN|422099009|SNOMEDCT_CORE|Disorder of eye due to type 2 diabetes mellitus|Disorder of eye due to type 2 diabetes mellitus
C0348919|T047|SY|422099009|SNOMEDCT_CORE|Disorder of eye with type 2 diabetes mellitus|Disorder of eye due to type 2 diabetes mellitus
C0348919|T047|IS|422099009|SNOMEDCT_CORE|Ophthalmic complication of adult-onset type diabetes mellitus|Disorder of eye due to type 2 diabetes mellitus
C0348919|T047|IS|422099009|SNOMEDCT_CORE|Ophthalmic complication of non-insulin-dependent diabetes mellitus|Disorder of eye due to type 2 diabetes mellitus
C0348921|T047|OP|199230006|SNOMEDCT_CORE|Pre-existing diabetes mellitus, non-insulin-dependent|Pre-existing type 2 diabetes mellitus
C0348921|T047|OF|199230006|SNOMEDCT_CORE|Pre-existing diabetes mellitus, non-insulin-dependent|Pre-existing type 2 diabetes mellitus
C0348921|T047|FN|199230006|SNOMEDCT_CORE|Pre-existing type 2 diabetes mellitus|Pre-existing type 2 diabetes mellitus
C0348921|T047|PT|199230006|SNOMEDCT_CORE|Pre-existing type 2 diabetes mellitus|Pre-existing type 2 diabetes mellitus
C0349006|T047|OAP|186385009|SNOMEDCT_CORE|Septicaemia due to Staphylococcus aureus|Septicemia due to Staphylococcus aureus
C0349006|T047|OAP|186385009|SNOMEDCT_CORE|Septicemia due to Staphylococcus aureus|Septicemia due to Staphylococcus aureus
C0349006|T047|OAF|186385009|SNOMEDCT_CORE|Septicemia due to Staphylococcus aureus|Septicemia due to Staphylococcus aureus
C0349007|T047|OAP|186386005|SNOMEDCT_CORE|Septicaemia due to coagulase-negative staphylococcus|Septicaemia due to coagulase-negative staphylococcus
C0349007|T047|OAP|186386005|SNOMEDCT_CORE|Septicemia due to coagulase-negative staphylococcus|Septicaemia due to coagulase-negative staphylococcus
C0349007|T047|OAF|186386005|SNOMEDCT_CORE|Septicemia due to coagulase-negative staphylococcus|Septicaemia due to coagulase-negative staphylococcus
C0349043|T191|SY|109371002|SNOMEDCT_CORE|Malignant neoplasm of overlapping lesion of bronchus and lung|Overlapping malignant neoplasm of bronchus and lung
C0349043|T191|PT|109371002|SNOMEDCT_CORE|Overlapping malignant neoplasm of bronchus and lung|Overlapping malignant neoplasm of bronchus and lung
C0349043|T191|FN|109371002|SNOMEDCT_CORE|Overlapping malignant neoplasm of bronchus and lung|Overlapping malignant neoplasm of bronchus and lung
C0349075|T047|PT|194727002|SNOMEDCT_CORE|Non-rheumatic mitral valve stenosis|Non-rheumatic mitral valve stenosis
C0349075|T047|FN|194727002|SNOMEDCT_CORE|Non-rheumatic mitral valve stenosis|Non-rheumatic mitral valve stenosis
C0349198|T048|PT|231489001|SNOMEDCT_CORE|Acute transient psychotic disorder|Acute transient psychotic disorder
C0349198|T048|FN|231489001|SNOMEDCT_CORE|Acute transient psychotic disorder|Acute transient psychotic disorder
C0349199|T048|PT|271428004|SNOMEDCT_CORE|Schizoaffective disorder, manic type|Schizoaffective disorder, manic type
C0349199|T048|FN|271428004|SNOMEDCT_CORE|Schizoaffective disorder, manic type|Schizoaffective disorder, manic type
C0349199|T048|SY|271428004|SNOMEDCT_CORE|Schizophreniform psychosis, manic type|Schizoaffective disorder, manic type
C0349217|T048|SY|35489007|SNOMEDCT_CORE|Depressive episode|Depressive episode
C0349245|T048|PT|191714002|SNOMEDCT_CORE|Dissociative convulsions|Dissociative convulsions
C0349245|T048|FN|191714002|SNOMEDCT_CORE|Dissociative convulsions|Dissociative convulsions
C0349245|T048|SY|191714002|SNOMEDCT_CORE|Dissociative seizures|Dissociative convulsions
C0349245|T048|SY|191714002|SNOMEDCT_CORE|Factitious seizures|Dissociative convulsions
C0349245|T048|SY|191714002|SNOMEDCT_CORE|Hysterical fit|Dissociative convulsions
C0349245|T048|SY|191714002|SNOMEDCT_CORE|Hysterical seizures|Dissociative convulsions
C0349245|T048|SY|191714002|SNOMEDCT_CORE|Pseudoseizures|Dissociative convulsions
C0349245|T048|SY|191714002|SNOMEDCT_CORE|Sham seizures|Dissociative convulsions
C0349255|T047|PT|192454004|SNOMEDCT_CORE|Nonorganic insomnia|Nonorganic insomnia
C0349255|T047|FN|192454004|SNOMEDCT_CORE|Nonorganic insomnia|Nonorganic insomnia
C0349280|T048|SY|66347000|SNOMEDCT_CORE|Habit and impulse disorder|Habit and impulse disorder
C0349347|T048|PT|192630004|SNOMEDCT_CORE|Psychogenic feeding disorder of infancy and childhood|Psychogenic feeding disorder of infancy and childhood
C0349347|T048|FN|192630004|SNOMEDCT_CORE|Psychogenic feeding disorder of infancy and childhood|Psychogenic feeding disorder of infancy and childhood
C0349391|T048|OAP|361276003|SNOMEDCT_CORE|Verbal apraxia|Verbal apraxia
C0349391|T048|OAF|361276003|SNOMEDCT_CORE|Verbal apraxia|Verbal apraxia
C0349453|T191|PT|237557003|SNOMEDCT_CORE|Mass of thyroid gland|Mass of thyroid gland
C0349453|T191|FN|237557003|SNOMEDCT_CORE|Mass of thyroid gland|Mass of thyroid gland
C0349453|T191|SY|237557003|SNOMEDCT_CORE|Thyroid lump|Mass of thyroid gland
C0349453|T191|OF|237557003|SNOMEDCT_CORE|Thyroid lump|Mass of thyroid gland
C0349453|T191|SY|237557003|SNOMEDCT_CORE|Thyroid mass|Mass of thyroid gland
C0349458|T191|PT|285836003|SNOMEDCT_CORE|Cervical intraepithelial neoplasia grade 1|Cervical intraepithelial neoplasia grade 1
C0349458|T191|FN|285836003|SNOMEDCT_CORE|Cervical intraepithelial neoplasia grade 1|Cervical intraepithelial neoplasia grade 1
C0349458|T191|SY|285836003|SNOMEDCT_CORE|Cervical intraepithelial neoplasia grade I|Cervical intraepithelial neoplasia grade 1
C0349458|T191|SY|285836003|SNOMEDCT_CORE|CIN I - Cervical intraepithelial neoplasia 1|Cervical intraepithelial neoplasia grade 1
C0349458|T191|SY|285836003|SNOMEDCT_CORE|Mild cervical dysplasia|Cervical intraepithelial neoplasia grade 1
C0349458|T191|SY|285836003|SNOMEDCT_CORE|Mild dysplasia of cervix|Cervical intraepithelial neoplasia grade 1
C0349459|T191|PT|285838002|SNOMEDCT_CORE|Cervical intraepithelial neoplasia grade 2|Cervical intraepithelial neoplasia grade 2
C0349459|T191|FN|285838002|SNOMEDCT_CORE|Cervical intraepithelial neoplasia grade 2|Cervical intraepithelial neoplasia grade 2
C0349459|T191|SY|285838002|SNOMEDCT_CORE|Cervical intraepithelial neoplasia grade II|Cervical intraepithelial neoplasia grade 2
C0349459|T191|SY|285838002|SNOMEDCT_CORE|CIN 2 - Cervical intraepithelial neoplasia 2|Cervical intraepithelial neoplasia grade 2
C0349459|T191|SY|285838002|SNOMEDCT_CORE|Moderate cervical dysplasia|Cervical intraepithelial neoplasia grade 2
C0349459|T191|SY|285838002|SNOMEDCT_CORE|Moderate dysplasia of cervix|Cervical intraepithelial neoplasia grade 2
C0349482|T033|PT|276613009|SNOMEDCT_CORE|High birth weight|High birth weight
C0349482|T033|FN|276613009|SNOMEDCT_CORE|High birth weight|High birth weight
C0349482|T033|SY|276613009|SNOMEDCT_CORE|High birth weight baby|High birth weight
C0349482|T033|OP|276613009|SNOMEDCT_CORE|High birth weight infant|High birth weight
C0349482|T033|OF|276613009|SNOMEDCT_CORE|High birth weight infant|High birth weight
C0349506|T046|PT|90128006|SNOMEDCT_CORE|Photosensitivity|Photosensitivity
C0349506|T046|FN|90128006|SNOMEDCT_CORE|Photosensitivity|Photosensitivity
C0349506|T046|SY|90128006|SNOMEDCT_CORE|Photosensitivity of skin|Photosensitivity
C0349541|T191|PT|276826005|SNOMEDCT_CORE|Malignant glioma of brain|Malignant glioma of brain
C0349541|T191|FN|276826005|SNOMEDCT_CORE|Malignant glioma of brain|Malignant glioma of brain
C0349549|T191|PT|276851006|SNOMEDCT_CORE|Intraduct papilloma of pancreas|Intraduct papilloma of pancreas
C0349549|T191|FN|276851006|SNOMEDCT_CORE|Intraduct papilloma of pancreas|Intraduct papilloma of pancreas
C0349566|T191|SY|276952000|SNOMEDCT_CORE|SCC - Squamous cell carcinoma of tongue|Squamous cell carcinoma of tongue
C0349566|T191|PT|276952000|SNOMEDCT_CORE|Squamous cell carcinoma of tongue|Squamous cell carcinoma of tongue
C0349566|T191|FN|276952000|SNOMEDCT_CORE|Squamous cell carcinoma of tongue|Squamous cell carcinoma of tongue
C0349568|T191|SY|276962007|SNOMEDCT_CORE|SCC - Squamous cell carcinoma of palate|Squamous cell carcinoma of palate
C0349568|T191|PT|276962007|SNOMEDCT_CORE|Squamous cell carcinoma of palate|Squamous cell carcinoma of palate
C0349568|T191|FN|276962007|SNOMEDCT_CORE|Squamous cell carcinoma of palate|Squamous cell carcinoma of palate
C0349571|T191|SY|255155005|SNOMEDCT_CORE|Adenoma of parotid gland|Pleomorphic adenoma of parotid gland
C0349571|T191|PT|255155005|SNOMEDCT_CORE|Pleomorphic adenoma of parotid gland|Pleomorphic adenoma of parotid gland
C0349571|T191|FN|255155005|SNOMEDCT_CORE|Pleomorphic adenoma of parotid gland|Pleomorphic adenoma of parotid gland
C0349571|T191|SY|255155005|SNOMEDCT_CORE|PSA - Pleomorphic adenoma of parotid gland|Pleomorphic adenoma of parotid gland
C0349577|T191|PT|277157002|SNOMEDCT_CORE|Benign tumor of external ear|Benign tumor of external ear
C0349577|T191|FN|277157002|SNOMEDCT_CORE|Benign tumor of external ear|Benign tumor of external ear
C0349577|T191|PTGB|277157002|SNOMEDCT_CORE|Benign tumour of external ear|Benign tumor of external ear
C0349588|T033|SY|237836003|SNOMEDCT_CORE|Small stature|SS - Short stature
C0349588|T033|SY|237836003|SNOMEDCT_CORE|SS - Short stature|SS - Short stature
C0349604|T191|SY|302820008|SNOMEDCT_CORE|Cranial meningioma|Intracranial meningioma
C0349604|T191|PT|302820008|SNOMEDCT_CORE|Intracranial meningioma|Intracranial meningioma
C0349604|T191|FN|302820008|SNOMEDCT_CORE|Intracranial meningioma|Intracranial meningioma
C0349604|T191|SY|302820008|SNOMEDCT_CORE|Meningioma of brain|Intracranial meningioma
C0349650|T047|PT|277869007|SNOMEDCT_CORE|Non-tuberculous mycobacterial pneumonia|Non-tuberculous mycobacterial pneumonia
C0349650|T047|FN|277869007|SNOMEDCT_CORE|Non-tuberculous mycobacterial pneumonia|Non-tuberculous mycobacterial pneumonia
C0349661|T191|FN|254936001|SNOMEDCT_CORE|Glial tumor of brain|Glial tumor of brain
C0349661|T191|PT|254936001|SNOMEDCT_CORE|Glial tumor of brain|Glial tumor of brain
C0349661|T191|PTGB|254936001|SNOMEDCT_CORE|Glial tumour of brain|Glial tumor of brain
C0349702|T033|PT|95726001|SNOMEDCT_CORE|Corneal scar|Corneal scar
C0349702|T033|FN|95726001|SNOMEDCT_CORE|Corneal scar|Corneal scar
C0349702|T033|IS|95726001|SNOMEDCT_CORE|Corneal scar, NOS|Corneal scar
C0349702|T033|IS|64634000|SNOMEDCT_CORE|Corneal scar, NOS|Corneal scar
C0349709|T048|PT|278853003|SNOMEDCT_CORE|Acute schizophrenia-like psychotic disorder|Acute schizophrenia-like psychotic disorder
C0349709|T048|FN|278853003|SNOMEDCT_CORE|Acute schizophrenia-like psychotic disorder|Acute schizophrenia-like psychotic disorder
C0349712|T048|PT|40568001|SNOMEDCT_CORE|Recurrent brief depressive disorder|Recurrent brief depressive disorder
C0349712|T048|FN|40568001|SNOMEDCT_CORE|Recurrent brief depressive disorder|Recurrent brief depressive disorder
C0349757|T046|PT|280972008|SNOMEDCT_CORE|Arteriovenous graft thrombosis|Arteriovenous graft thrombosis
C0349757|T046|FN|280972008|SNOMEDCT_CORE|Arteriovenous graft thrombosis|Arteriovenous graft thrombosis
C0349782|T047|PTGB|194849004|SNOMEDCT_CORE|Generalised ischaemic myocardial dysfunction|Generalized ischemic myocardial dysfunction
C0349782|T047|PT|194849004|SNOMEDCT_CORE|Generalized ischemic myocardial dysfunction|Generalized ischemic myocardial dysfunction
C0349782|T047|FN|194849004|SNOMEDCT_CORE|Generalized ischemic myocardial dysfunction|Generalized ischemic myocardial dysfunction
C0349782|T047|SYGB|194849004|SNOMEDCT_CORE|Ischaemic cardiomyopathy|Generalized ischemic myocardial dysfunction
C0349782|T047|SY|194849004|SNOMEDCT_CORE|Ischemic cardiomyopathy|Generalized ischemic myocardial dysfunction
C0349790|T033|IS|281239006|SNOMEDCT_CORE|Acute exacerbation of asthma|Exacerbation of asthma
C0349790|T033|PT|281239006|SNOMEDCT_CORE|Exacerbation of asthma|Exacerbation of asthma
C0349790|T033|FN|281239006|SNOMEDCT_CORE|Exacerbation of asthma|Exacerbation of asthma
C0362046|T047|IS|9414007|SNOMEDCT_CORE|Prediabetes|Prediabetes
C0362050|T046|SY|110270004|SNOMEDCT_CORE|Late effects of acute poliomyelitis|Late effects of poliomyelitis
C0362050|T046|PT|110270004|SNOMEDCT_CORE|Late effects of poliomyelitis|Late effects of poliomyelitis
C0362050|T046|OF|110270004|SNOMEDCT_CORE|Late effects of poliomyelitis|Late effects of poliomyelitis
C0362050|T046|FN|110270004|SNOMEDCT_CORE|Sequela of infection caused by Human poliovirus|Late effects of poliomyelitis
C0362050|T046|SY|110270004|SNOMEDCT_CORE|Sequela of infection caused by Human poliovirus|Late effects of poliomyelitis
C0362060|T033|PT|22268004|SNOMEDCT_CORE|Legal problem|Legal problem
C0362060|T033|FN|22268004|SNOMEDCT_CORE|Legal problem|Legal problem
C0362060|T033|IS|22268004|SNOMEDCT_CORE|Legal problem, NOS|Legal problem
C0375071|T191|SY|363367000|SNOMEDCT_CORE|Cancer of vulva|Malignant tumor of vulva
C0375071|T191|PT|363367000|SNOMEDCT_CORE|Malignant tumor of vulva|Malignant tumor of vulva
C0375071|T191|FN|363367000|SNOMEDCT_CORE|Malignant tumor of vulva|Malignant tumor of vulva
C0375071|T191|PTGB|363367000|SNOMEDCT_CORE|Malignant tumour of vulva|Malignant tumor of vulva
C0375209|T184|PT|442077006|SNOMEDCT_CORE|Flaccid hemiplegia of nondominant side|Flaccid hemiplegia of nondominant side
C0375209|T184|FN|442077006|SNOMEDCT_CORE|Flaccid hemiplegia of nondominant side|Flaccid hemiplegia of nondominant side
C0375257|T046|PT|60331006|SNOMEDCT_CORE|Abnormal auditory perception|Abnormal auditory perception
C0375257|T046|OF|60331006|SNOMEDCT_CORE|Abnormal auditory perception|Abnormal auditory perception
C0375257|T046|FN|60331006|SNOMEDCT_CORE|Abnormal auditory perception|Abnormal auditory perception
C0375257|T046|IS|60331006|SNOMEDCT_CORE|Abnormal auditory perception, NOS|Abnormal auditory perception
C0375305|T047|OAP|444701000|SNOMEDCT_CORE|Dissecting aneurysm of thoracoabdominal aorta|Dissecting aneurysm of thoracoabdominal aorta
C0375305|T047|OAF|444701000|SNOMEDCT_CORE|Dissecting aneurysm of thoracoabdominal aorta|Dissecting aneurysm of thoracoabdominal aorta
C0375336|T047|PT|441536000|SNOMEDCT_CORE|Iatrogenic pneumothorax|Iatrogenic pneumothorax
C0375336|T047|FN|441536000|SNOMEDCT_CORE|Iatrogenic pneumothorax|Iatrogenic pneumothorax
C0375359|T047|PT|441971007|SNOMEDCT_CORE|Chronic left-sided ulcerative colitis|Chronic left-sided ulcerative colitis
C0375359|T047|FN|441971007|SNOMEDCT_CORE|Chronic left-sided ulcerative colitis|Chronic left-sided ulcerative colitis
C0375732|T046|OAS|403676009|SNOMEDCT_CORE|Non healing surgical wound|Non-healing surgical wound
C0375732|T046|OAF|403676009|SNOMEDCT_CORE|Non-healing surgical wound|Non-healing surgical wound
C0375732|T046|OAP|403676009|SNOMEDCT_CORE|Non-healing surgical wound|Non-healing surgical wound
C0375732|T046|PT|781187003|SNOMEDCT_CORE|Non-healing surgical wound|Non-healing surgical wound
C0375732|T046|OF|403676009|SNOMEDCT_CORE|Non-healing surgical wound|Non-healing surgical wound
C0375732|T046|FN|781187003|SNOMEDCT_CORE|Non-healing surgical wound|Non-healing surgical wound
C0375812|T033|PT|161635002|SNOMEDCT_CORE|H/O: asbestos exposure|H/O: asbestos exposure
C0375812|T033|IS|161635002|SNOMEDCT_CORE|History of - asbestos exposure|H/O: asbestos exposure
C0375812|T033|OF|161635002|SNOMEDCT_CORE|History of - asbestos exposure|H/O: asbestos exposure
C0375812|T033|SY|161635002|SNOMEDCT_CORE|History of asbestos exposure|H/O: asbestos exposure
C0375812|T033|FN|161635002|SNOMEDCT_CORE|History of asbestos exposure|H/O: asbestos exposure
C0376117|T191|PT|442348004|SNOMEDCT_CORE|Inflamed seborrheic keratosis|Inflamed seborrheic keratosis
C0376117|T191|FN|442348004|SNOMEDCT_CORE|Inflamed seborrheic keratosis|Inflamed seborrheic keratosis
C0376117|T191|PTGB|442348004|SNOMEDCT_CORE|Inflamed seborrhoeic keratosis|Inflamed seborrheic keratosis
C0376154|T020|PT|201040000|SNOMEDCT_CORE|Callosity|Callosity
C0376154|T020|FN|201040000|SNOMEDCT_CORE|Callosity|Callosity
C0376154|T020|SY|201040000|SNOMEDCT_CORE|Callus|Callosity
C0376175|T047|SY|193093009|SNOMEDCT_CORE|Bell palsy|Bell's palsy
C0376175|T047|PT|193093009|SNOMEDCT_CORE|Bell's palsy|Bell's palsy
C0376175|T047|FN|193093009|SNOMEDCT_CORE|Bell's palsy|Bell's palsy
C0376175|T047|SY|193093009|SNOMEDCT_CORE|Bells palsy|Bell's palsy
C0376175|T047|SY|193093009|SNOMEDCT_CORE|Idiopathic acute facial nerve palsy|Bell's palsy
C0376186|T047|SY|48277006|SNOMEDCT_CORE|Impetigo contagiosa|Impetigo contagiosa
C0376356|T047|SY|82639001|SNOMEDCT_CORE|PMT - Premenstrual tension|Premenstrual tension syndrome
C0376356|T047|SY|82639001|SNOMEDCT_CORE|Premenstrual tension|Premenstrual tension syndrome
C0376356|T047|PT|82639001|SNOMEDCT_CORE|Premenstrual tension syndrome|Premenstrual tension syndrome
C0376356|T047|FN|82639001|SNOMEDCT_CORE|Premenstrual tension syndrome|Premenstrual tension syndrome
C0376356|T047|IS|82639001|SNOMEDCT_CORE|Premenstrual tension syndrome, NOS|Premenstrual tension syndrome
C0376358|T191|SY|399068003|SNOMEDCT_CORE|CA - Cancer of prostate|Malignant tumor of prostate
C0376358|T191|SY|399068003|SNOMEDCT_CORE|Cancer of prostate|Malignant tumor of prostate
C0376358|T191|IS|93974005|SNOMEDCT_CORE|Malignant neoplasm of prostate|Malignant tumor of prostate
C0376358|T191|SY|399068003|SNOMEDCT_CORE|Malignant prostatic tumor|Malignant tumor of prostate
C0376358|T191|SYGB|399068003|SNOMEDCT_CORE|Malignant prostatic tumour|Malignant tumor of prostate
C0376358|T191|PT|399068003|SNOMEDCT_CORE|Malignant tumor of prostate|Malignant tumor of prostate
C0376358|T191|FN|399068003|SNOMEDCT_CORE|Malignant tumor of prostate|Malignant tumor of prostate
C0376358|T191|PTGB|399068003|SNOMEDCT_CORE|Malignant tumour of prostate|Malignant tumor of prostate
C0376379|T047|SY|57920007|SNOMEDCT_CORE|Herpes simplex gingivostomatitis|Herpetic gingivostomatitis
C0376379|T047|PT|57920007|SNOMEDCT_CORE|Herpetic gingivostomatitis|Herpetic gingivostomatitis
C0376379|T047|FN|57920007|SNOMEDCT_CORE|Herpetic gingivostomatitis|Herpetic gingivostomatitis
C0376379|T047|SY|57920007|SNOMEDCT_CORE|Primary herpetic gingivostomatitis|Herpetic gingivostomatitis
C0376545|T191|PTGB|129154003|SNOMEDCT_CORE|Haematologic neoplasm|Hematologic neoplasm
C0376545|T191|PT|129154003|SNOMEDCT_CORE|Hematologic neoplasm|Hematologic neoplasm
C0376545|T191|FN|129154003|SNOMEDCT_CORE|Hematologic neoplasm|Hematologic neoplasm
C0376685|T047|SY|239960007|SNOMEDCT_CORE|Impingement syndrome of shoulder|Impingement syndrome of shoulder region
C0376685|T047|PT|239960007|SNOMEDCT_CORE|Impingement syndrome of shoulder region|Impingement syndrome of shoulder region
C0376685|T047|FN|239960007|SNOMEDCT_CORE|Impingement syndrome of shoulder region|Impingement syndrome of shoulder region
C0376685|T047|SY|239960007|SNOMEDCT_CORE|Shoulder impingement syndrome|Impingement syndrome of shoulder region
C0376710|T047|SY|236053002|SNOMEDCT_CORE|Sliding diaphragmatic hernia|Sliding hiatus hernia
C0376710|T047|SY|236053002|SNOMEDCT_CORE|Sliding esophageal hiatus hernia|Sliding hiatus hernia
C0376710|T047|PT|236053002|SNOMEDCT_CORE|Sliding hiatus hernia|Sliding hiatus hernia
C0376710|T047|FN|236053002|SNOMEDCT_CORE|Sliding hiatus hernia|Sliding hiatus hernia
C0376710|T047|SYGB|236053002|SNOMEDCT_CORE|Sliding oesophageal hiatus hernia|Sliding hiatus hernia
C0391820|T047|SY|190829000|SNOMEDCT_CORE|Gouty nephropathy|Gouty nephropathy
C0391920|T190|IS|20018005|SNOMEDCT_CORE|Intrinsic ureteral obstruction|Intrinsic ureteral obstruction
C0391924|T019|SYGB|72100002|SNOMEDCT_CORE|Naevoid lentigo|Nevoid lentigo
C0391924|T019|SY|72100002|SNOMEDCT_CORE|Nevoid lentigo|Nevoid lentigo
C0391959|T047|OAP|12731000|SNOMEDCT_CORE|Cervical sympathetic dystrophy|Cervical sympathetic paralysis
C0391959|T047|OAF|12731000|SNOMEDCT_CORE|Cervical sympathetic dystrophy|Cervical sympathetic paralysis
C0391959|T047|IS|12731000|SNOMEDCT_CORE|Cervical sympathetic paralysis|Cervical sympathetic paralysis
C0391970|T191|PT|445238008|SNOMEDCT_CORE|Malignant carcinoid tumor|Malignant carcinoid tumor
C0391970|T191|FN|445238008|SNOMEDCT_CORE|Malignant carcinoid tumor|Malignant carcinoid tumor
C0391970|T191|PTGB|445238008|SNOMEDCT_CORE|Malignant carcinoid tumour|Malignant carcinoid tumor
C0391993|T047|PT|49176002|SNOMEDCT_CORE|Arteriosclerotic gangrene|Arteriosclerotic gangrene
C0391993|T047|FN|49176002|SNOMEDCT_CORE|Arteriosclerotic gangrene|Arteriosclerotic gangrene
C0392003|T047|PT|75817003|SNOMEDCT_CORE|Cellulitis of breast|Cellulitis of breast
C0392003|T047|FN|75817003|SNOMEDCT_CORE|Cellulitis of breast|Cellulitis of breast
C0392042|T046|PT|427769002|SNOMEDCT_CORE|Infection of amputation stump|Infection of amputation stump
C0392042|T046|FN|427769002|SNOMEDCT_CORE|Infection of amputation stump|Infection of amputation stump
C0392118|T037|PT|274170000|SNOMEDCT_CORE|Open wound of abdominal wall|Open wound of abdominal wall
C0392118|T037|FN|274170000|SNOMEDCT_CORE|Open wound of abdominal wall|Open wound of abdominal wall
C0392120|T037|PT|210323002|SNOMEDCT_CORE|Open wound of scalp|Open wound of scalp
C0392120|T037|FN|210323002|SNOMEDCT_CORE|Open wound of scalp|Open wound of scalp
C0392163|T047|PT|50792001|SNOMEDCT_CORE|Corneal erosion|Corneal erosion
C0392163|T047|FN|50792001|SNOMEDCT_CORE|Corneal erosion|Corneal erosion
C0392163|T047|IS|50792001|SNOMEDCT_CORE|Superficial corneal ulcer|Corneal erosion
C0392163|T047|SY|50792001|SNOMEDCT_CORE|Superficial ulcer of cornea|Corneal erosion
C0392164|T047|PT|86555001|SNOMEDCT_CORE|Cystic fibrosis of the lung|Cystic fibrosis of the lung
C0392164|T047|FN|86555001|SNOMEDCT_CORE|Cystic fibrosis of the lung|Cystic fibrosis of the lung
C0392164|T047|SY|86555001|SNOMEDCT_CORE|Mucoviscidosis involving the lung|Cystic fibrosis of the lung
C0392164|T047|SY|86555001|SNOMEDCT_CORE|Pulmonary cystic fibrosis|Cystic fibrosis of the lung
C0392171|T184|SY|95891005|SNOMEDCT_CORE|Flu-like symptoms|Flu-like symptoms
C0392176|T184|SY|3696007|SNOMEDCT_CORE|Gastric irritation|Gastric irritation
C0392322|T048|SY|111484002|SNOMEDCT_CORE|Atypical schizophrenia|Undifferentiated schizophrenia
C0392322|T048|PT|111484002|SNOMEDCT_CORE|Undifferentiated schizophrenia|Undifferentiated schizophrenia
C0392322|T048|FN|111484002|SNOMEDCT_CORE|Undifferentiated schizophrenia|Undifferentiated schizophrenia
C0392322|T048|IS|111484002|SNOMEDCT_CORE|Undifferentiated schizophrenia, NOS|Undifferentiated schizophrenia
C0392454|T033|PT|68372009|SNOMEDCT_CORE|Upper respiratory tract obstruction|Upper respiratory tract obstruction
C0392454|T033|FN|68372009|SNOMEDCT_CORE|Upper respiratory tract obstruction|Upper respiratory tract obstruction
C0392462|T047|OAP|194766005|SNOMEDCT_CORE|Benign hypertensive heart disease without congestive cardiac failure|Benign hypertensive heart disease without congestive heart failure
C0392462|T047|OAF|194766005|SNOMEDCT_CORE|Benign hypertensive heart disease without congestive cardiac failure|Benign hypertensive heart disease without congestive heart failure
C0392462|T047|PT|77970009|SNOMEDCT_CORE|Benign hypertensive heart disease without congestive heart failure|Benign hypertensive heart disease without congestive heart failure
C0392462|T047|FN|77970009|SNOMEDCT_CORE|Benign hypertensive heart disease without congestive heart failure|Benign hypertensive heart disease without congestive heart failure
C0392477|T019|SY|23407003|SNOMEDCT_CORE|Congenital flat foot|Congenital pes planus
C0392477|T019|PT|23407003|SNOMEDCT_CORE|Congenital pes planus|Congenital pes planus
C0392477|T019|FN|23407003|SNOMEDCT_CORE|Congenital pes planus|Congenital pes planus
C0392477|T019|IS|23407003|SNOMEDCT_CORE|Pes planovalgus|Congenital pes planus
C0392477|T019|IS|23407003|SNOMEDCT_CORE|Pes planus|Congenital pes planus
C0392498|T020|PTGB|34580000|SNOMEDCT_CORE|Duodenal ulcer without haemorrhage, without perforation AND without obstruction|Duodenal ulcer without hemorrhage, without perforation AND without obstruction
C0392498|T020|PT|34580000|SNOMEDCT_CORE|Duodenal ulcer without hemorrhage, without perforation AND without obstruction|Duodenal ulcer without hemorrhage, without perforation AND without obstruction
C0392498|T020|FN|34580000|SNOMEDCT_CORE|Duodenal ulcer without hemorrhage, without perforation AND without obstruction|Duodenal ulcer without hemorrhage, without perforation AND without obstruction
C0392498|T020|IS|34580000|SNOMEDCT_CORE|Duodenal ulcer, NOS without hemorrhage or perforation and without obstruction|Duodenal ulcer without hemorrhage, without perforation AND without obstruction
C0392531|T190|PT|198047009|SNOMEDCT_CORE|Torsion of appendix of testis|Torsion of appendix of testis
C0392531|T190|FN|198047009|SNOMEDCT_CORE|Torsion of appendix of testis|Torsion of appendix of testis
C0392531|T190|SY|198047009|SNOMEDCT_CORE|Torsion of hydatid of Morgagni - male|Torsion of appendix of testis
C0392531|T190|IS|198047009|SNOMEDCT_CORE|Torsion of hydatid of Morgani - male|Torsion of appendix of testis
C0392534|T046|SY|17433009|SNOMEDCT_CORE|Aborted ectopic pregnancy|Ruptured ectopic pregnancy
C0392534|T046|PT|17433009|SNOMEDCT_CORE|Ruptured ectopic pregnancy|Ruptured ectopic pregnancy
C0392534|T046|FN|17433009|SNOMEDCT_CORE|Ruptured ectopic pregnancy|Ruptured ectopic pregnancy
C0392543|T047|PT|17140000|SNOMEDCT_CORE|Neonatal jaundice due to delayed conjugation|Neonatal jaundice due to delayed conjugation
C0392543|T047|FN|17140000|SNOMEDCT_CORE|Neonatal jaundice due to delayed conjugation|Neonatal jaundice due to delayed conjugation
C0392543|T047|IS|17140000|SNOMEDCT_CORE|Neonatal jaundice due to delayed conjugation, NOS|Neonatal jaundice due to delayed conjugation
C0392548|T047|PT|192970008|SNOMEDCT_CORE|Cauda equina syndrome|Cauda equina syndrome
C0392548|T047|FN|192970008|SNOMEDCT_CORE|Cauda equina syndrome|Cauda equina syndrome
C0392549|T047|IS|1178005|SNOMEDCT_CORE|Infantile cerebral palsy, NOS|Infantile cerebral palsy, NOS
C0392553|T047|PT|65017003|SNOMEDCT_CORE|Hereditary peripheral neuropathy|Hereditary peripheral neuropathy
C0392553|T047|FN|65017003|SNOMEDCT_CORE|Hereditary peripheral neuropathy|Hereditary peripheral neuropathy
C0392553|T047|IS|65017003|SNOMEDCT_CORE|Hereditary peripheral neuropathy, NOS|Hereditary peripheral neuropathy
C0392557|T047|IS|53889007|SNOMEDCT_CORE|Lenticular sclerosis|Nuclear cataract
C0392557|T047|SY|53889007|SNOMEDCT_CORE|NS - Nuclear sclerosis|Nuclear cataract
C0392557|T047|PT|53889007|SNOMEDCT_CORE|Nuclear cataract|Nuclear cataract
C0392557|T047|FN|53889007|SNOMEDCT_CORE|Nuclear cataract|Nuclear cataract
C0392557|T047|IS|53889007|SNOMEDCT_CORE|Nuclear cataract, NOS|Nuclear cataract
C0392557|T047|IS|53889007|SNOMEDCT_CORE|Nuclear sclerosis|Nuclear cataract
C0392611|T037|PT|25899002|SNOMEDCT_CORE|Closed bimalleolar fracture|Closed bimalleolar fracture
C0392611|T037|FN|25899002|SNOMEDCT_CORE|Closed bimalleolar fracture|Closed bimalleolar fracture
C0392618|T046|PT|33910007|SNOMEDCT_CORE|Postoperative infection|Postoperative infection
C0392618|T046|FN|33910007|SNOMEDCT_CORE|Postoperative infection|Postoperative infection
C0392646|T047|IS|88594005|SNOMEDCT_CORE|Herpes simplex without mention of complication|Herpes simplex without mention of complication
C0392650|T047|IS|14189004|SNOMEDCT_CORE|Measles without mention of complication|Measles without mention of complication
C0392672|T033|SY|386702006|SNOMEDCT_CORE|Battered person syndrome|Battered person syndrome
C0392672|T033|IS|386702006|SNOMEDCT_CORE|Battered person syndrome, NOS|Battered person syndrome
C0392678|T184|SY|399122003|SNOMEDCT_CORE|Impaired swallowing|Swallowing problem
C0392678|T184|SY|399122003|SNOMEDCT_CORE|Swallowing impairment|Swallowing problem
C0392678|T184|PT|399122003|SNOMEDCT_CORE|Swallowing problem|Swallowing problem
C0392678|T184|FN|399122003|SNOMEDCT_CORE|Swallowing problem|Swallowing problem
C0392681|T184|SY|56018004|SNOMEDCT_CORE|Asthmatic breath sounds|Asthmatic breathing
C0392681|T184|SY|56018004|SNOMEDCT_CORE|Asthmatic breathing|Asthmatic breathing
C0392682|T033|SY|371622005|SNOMEDCT_CORE|Elevated blood pressure reading without diagnosis of hypertension|Elevated blood-pressure reading without diagnosis of hypertension
C0392682|T033|FN|371622005|SNOMEDCT_CORE|Elevated blood pressure reading without diagnosis of hypertension|Elevated blood-pressure reading without diagnosis of hypertension
C0392682|T033|PT|371622005|SNOMEDCT_CORE|Elevated blood-pressure reading without diagnosis of hypertension|Elevated blood-pressure reading without diagnosis of hypertension
C0392682|T033|OF|371622005|SNOMEDCT_CORE|Elevated blood-pressure reading without diagnosis of hypertension|Elevated blood-pressure reading without diagnosis of hypertension
C0392699|T047|SYGB|279079003|SNOMEDCT_CORE|Abnormal sensation of dysaesthesia|Dysesthesia
C0392699|T047|SY|279079003|SNOMEDCT_CORE|Abnormal sensation of dysesthesia|Dysesthesia
C0392699|T047|PTGB|279079003|SNOMEDCT_CORE|Dysaesthesia|Dysesthesia
C0392699|T047|IS|279079003|SNOMEDCT_CORE|Dysaesthesia|Dysesthesia
C0392699|T047|PT|279079003|SNOMEDCT_CORE|Dysesthesia|Dysesthesia
C0392699|T047|IS|279079003|SNOMEDCT_CORE|Dysesthesia|Dysesthesia
C0392699|T047|FN|279079003|SNOMEDCT_CORE|Dysesthesia|Dysesthesia
C0392702|T047|PT|260912008|SNOMEDCT_CORE|Abnormal involuntary movement|Abnormal involuntary movement
C0392702|T047|FN|260912008|SNOMEDCT_CORE|Abnormal involuntary movement|Abnormal involuntary movement
C0393386|T046|PT|212904005|SNOMEDCT_CORE|Radiation therapy complication|Radiation therapy complication
C0393386|T046|FN|212904005|SNOMEDCT_CORE|Radiation therapy complication|Radiation therapy complication
C0393485|T047|PT|230193008|SNOMEDCT_CORE|Neurosarcoidosis|Neurosarcoidosis
C0393485|T047|FN|230193008|SNOMEDCT_CORE|Neurosarcoidosis|Neurosarcoidosis
C0393560|T047|PT|230285003|SNOMEDCT_CORE|Vascular dementia of acute onset|Vascular dementia of acute onset
C0393560|T047|FN|230285003|SNOMEDCT_CORE|Vascular dementia of acute onset|Vascular dementia of acute onset
C0393570|T047|SY|18842008|SNOMEDCT_CORE|Cortical basal ganglionic degeneration|Corticobasal degeneration
C0393570|T047|PT|18842008|SNOMEDCT_CORE|Corticobasal degeneration|Corticobasal degeneration
C0393570|T047|FN|18842008|SNOMEDCT_CORE|Corticobasal degeneration|Corticobasal degeneration
C0393570|T047|SY|18842008|SNOMEDCT_CORE|Corticodentatonigral degeneration with neuronal achromasia|Corticobasal degeneration
C0393571|T046|SY|230297002|SNOMEDCT_CORE|MSA - Multiple system atrophy|Multiple system atrophy
C0393571|T046|PT|230297002|SNOMEDCT_CORE|Multiple system atrophy|Multiple system atrophy
C0393571|T046|FN|230297002|SNOMEDCT_CORE|Multiple system atrophy|Multiple system atrophy
C0393593|T047|FN|15802004|SNOMEDCT_CORE|Dystonia|Dystonia
C0393593|T047|PT|15802004|SNOMEDCT_CORE|Dystonia|Dystonia
C0393593|T047|SY|15802004|SNOMEDCT_CORE|Dystonia disorder|Dystonia
C0393615|T047|OAP|192840004|SNOMEDCT_CORE|Benign familial tremor|Hereditary essential tremor
C0393615|T047|OAF|192840004|SNOMEDCT_CORE|Benign familial tremor|Hereditary essential tremor
C0393615|T047|OAS|192840004|SNOMEDCT_CORE|Familial tremor|Hereditary essential tremor
C0393615|T047|OAS|192839001|SNOMEDCT_CORE|Hereditary essential tremor|Hereditary essential tremor
C0393615|T047|PT|609559001|SNOMEDCT_CORE|Hereditary essential tremor|Hereditary essential tremor
C0393615|T047|FN|609559001|SNOMEDCT_CORE|Hereditary essential tremor|Hereditary essential tremor
C0393615|T047|OAS|192839001|SNOMEDCT_CORE|Heredofamilial tremor|Hereditary essential tremor
C0393666|T047|OAS|230374002|SNOMEDCT_CORE|Multiple sclerosis remitting progressive|Multiple sclerosis remitting progressive
C0393666|T047|OAP|230374002|SNOMEDCT_CORE|Remittent-progressive multiple sclerosis|Multiple sclerosis remitting progressive
C0393666|T047|OAF|230374002|SNOMEDCT_CORE|Remittent-progressive multiple sclerosis|Multiple sclerosis remitting progressive
C0393736|T047|SY|398126006|SNOMEDCT_CORE|Muscle contraction headache|Muscular headache
C0393736|T047|PT|398126006|SNOMEDCT_CORE|Muscular headache|Muscular headache
C0393736|T047|FN|398126006|SNOMEDCT_CORE|Muscular headache|Muscular headache
C0393737|T047|PT|230470007|SNOMEDCT_CORE|Episodic tension-type headache|Episodic tension-type headache
C0393737|T047|FN|230470007|SNOMEDCT_CORE|Episodic tension-type headache|Episodic tension-type headache
C0393738|T047|PT|230471006|SNOMEDCT_CORE|Chronic tension-type headache|Chronic tension-type headache
C0393738|T047|FN|230471006|SNOMEDCT_CORE|Chronic tension-type headache|Chronic tension-type headache
C0393758|T047|FN|191997003|SNOMEDCT_CORE|Persistent insomnia|Persistent insomnia
C0393758|T047|PT|191997003|SNOMEDCT_CORE|Persistent insomnia|Persistent insomnia
C0393770|T047|SY|80623000|SNOMEDCT_CORE|Circadian rhythm sleep disorder, delayed sleep phase|Sleep-wake schedule disorder, delayed phase type
C0393770|T047|SY|80623000|SNOMEDCT_CORE|Circadian rhythm sleep disorder, delayed sleep phase type|Sleep-wake schedule disorder, delayed phase type
C0393770|T047|SY|80623000|SNOMEDCT_CORE|Delayed sleep phase syndrome|Sleep-wake schedule disorder, delayed phase type
C0393770|T047|SY|80623000|SNOMEDCT_CORE|Delayed sleep-wake phase disorder|Sleep-wake schedule disorder, delayed phase type
C0393770|T047|PT|80623000|SNOMEDCT_CORE|Sleep-wake schedule disorder, delayed phase type|Sleep-wake schedule disorder, delayed phase type
C0393770|T047|FN|80623000|SNOMEDCT_CORE|Sleep-wake schedule disorder, delayed phase type|Sleep-wake schedule disorder, delayed phase type
C0393819|T047|OP|444728005|SNOMEDCT_CORE|Chronic inflammatory demyelinating polyneuritis|Chronic inflammatory demyelinating polyradiculoneuropathy
C0393819|T047|OF|444728005|SNOMEDCT_CORE|Chronic inflammatory demyelinating polyneuritis|Chronic inflammatory demyelinating polyradiculoneuropathy
C0393819|T047|OAF|444728005|SNOMEDCT_CORE|Chronic inflammatory demyelinating polyneuropathy|Chronic inflammatory demyelinating polyradiculoneuropathy
C0393819|T047|OAP|444728005|SNOMEDCT_CORE|Chronic inflammatory demyelinating polyneuropathy|Chronic inflammatory demyelinating polyradiculoneuropathy
C0393819|T047|SY|128209004|SNOMEDCT_CORE|Chronic inflammatory demyelinating polyneuropathy|Chronic inflammatory demyelinating polyradiculoneuropathy
C0393819|T047|PT|128209004|SNOMEDCT_CORE|Chronic inflammatory demyelinating polyradiculoneuropathy|Chronic inflammatory demyelinating polyradiculoneuropathy
C0393819|T047|FN|128209004|SNOMEDCT_CORE|Chronic inflammatory demyelinating polyradiculoneuropathy|Chronic inflammatory demyelinating polyradiculoneuropathy
C0393819|T047|IS|128209004|SNOMEDCT_CORE|CIDP|Chronic inflammatory demyelinating polyradiculoneuropathy
C0393819|T047|SY|128209004|SNOMEDCT_CORE|CIDP - Chronic inflammatory demyelinating polyneuropathy|Chronic inflammatory demyelinating polyradiculoneuropathy
C0393819|T047|SY|128209004|SNOMEDCT_CORE|CIDP - Chronic inflammatory demyelinating polyradiculoneuropathy|Chronic inflammatory demyelinating polyradiculoneuropathy
C0393847|T047|SY|230591002|SNOMEDCT_CORE|MMN - Motor neuropathy with multiple conduction block|Motor neuropathy with multiple conduction block
C0393847|T047|PT|230591002|SNOMEDCT_CORE|Motor neuropathy with multiple conduction block|Motor neuropathy with multiple conduction block
C0393847|T047|FN|230591002|SNOMEDCT_CORE|Motor neuropathy with multiple conduction block|Motor neuropathy with multiple conduction block
C0393847|T047|SY|230591002|SNOMEDCT_CORE|Multifocal motor neuropathy|Motor neuropathy with multiple conduction block
C0393951|T047|OF|230691006|SNOMEDCT_CORE|Cerebrovascular accident due to cerebral artery occlusion|CVA - cerebrovascular accident due to cerebral artery occlusion
C0393951|T047|SY|230691006|SNOMEDCT_CORE|Cerebrovascular accident due to cerebral artery occlusion|CVA - cerebrovascular accident due to cerebral artery occlusion
C0393951|T047|FN|230691006|SNOMEDCT_CORE|Cerebrovascular accident due to occlusion of cerebral artery|CVA - cerebrovascular accident due to cerebral artery occlusion
C0393951|T047|SY|230691006|SNOMEDCT_CORE|Cerebrovascular accident due to occlusion of cerebral artery|CVA - cerebrovascular accident due to cerebral artery occlusion
C0393951|T047|PT|230691006|SNOMEDCT_CORE|CVA - cerebrovascular accident due to cerebral artery occlusion|CVA - cerebrovascular accident due to cerebral artery occlusion
C0393951|T047|OF|230691006|SNOMEDCT_CORE|CVA - cerebrovascular accident due to cerebral artery occlusion|CVA - cerebrovascular accident due to cerebral artery occlusion
C0393995|T047|SY|48721008|SNOMEDCT_CORE|Cerebral palsy with spastic tetraplegia|Tetraplegic cerebral palsy
C0393995|T047|SY|48721008|SNOMEDCT_CORE|Quadriplegic cerebral palsy|Tetraplegic cerebral palsy
C0393995|T047|FN|48721008|SNOMEDCT_CORE|Quadriplegic cerebral palsy|Tetraplegic cerebral palsy
C0393995|T047|SY|48721008|SNOMEDCT_CORE|Quadriplegic spastic cerebral palsy|Tetraplegic cerebral palsy
C0393995|T047|SY|48721008|SNOMEDCT_CORE|Spastic quadriplegic cerebral palsy|Tetraplegic cerebral palsy
C0393995|T047|PT|48721008|SNOMEDCT_CORE|Tetraplegic cerebral palsy|Tetraplegic cerebral palsy
C0393995|T047|SY|48721008|SNOMEDCT_CORE|Tetraplegic spastic cerebral palsy|Tetraplegic cerebral palsy
C0394006|T047|SY|230782004|SNOMEDCT_CORE|DES - Dysequilibrium syndrome|Dysequilibrium syndrome
C0394006|T047|SY|230782004|SNOMEDCT_CORE|Disequilibrium|Dysequilibrium syndrome
C0394006|T047|SY|230782004|SNOMEDCT_CORE|Dysequilibrium|Dysequilibrium syndrome
C0394006|T047|PT|230782004|SNOMEDCT_CORE|Dysequilibrium syndrome|Dysequilibrium syndrome
C0394006|T047|FN|230782004|SNOMEDCT_CORE|Dysequilibrium syndrome|Dysequilibrium syndrome
C0394019|T046|PT|230802007|SNOMEDCT_CORE|Brainstem death|Brainstem death
C0394019|T046|FN|230802007|SNOMEDCT_CORE|Brainstem death|Brainstem death
C0394032|T020|PT|230808006|SNOMEDCT_CORE|Brain ventricular shunt obstruction|Brain ventricular shunt obstruction
C0394032|T020|FN|230808006|SNOMEDCT_CORE|Brain ventricular shunt obstruction|Brain ventricular shunt obstruction
C0394996|T048|SY|25702006|SNOMEDCT_CORE|Acute alcohol intoxication|Acute alcohol intoxication
C0395016|T033|PT|267095009|SNOMEDCT_CORE|Speech problem|Speech problem
C0395016|T033|FN|267095009|SNOMEDCT_CORE|Speech problem|Speech problem
C0395803|T047|PT|232214001|SNOMEDCT_CORE|Cellulitis of pinna|Cellulitis of pinna
C0395803|T047|FN|232214001|SNOMEDCT_CORE|Cellulitis of pinna|Cellulitis of pinna
C0395862|T047|SY|86279000|SNOMEDCT_CORE|Acute suppurative otitis media - tympanic membrane ruptured|Acute suppurative otitis media with spontaneous rupture of ear drum
C0395862|T047|PT|86279000|SNOMEDCT_CORE|Acute suppurative otitis media with spontaneous rupture of ear drum|Acute suppurative otitis media with spontaneous rupture of ear drum
C0395862|T047|FN|86279000|SNOMEDCT_CORE|Acute suppurative otitis media with spontaneous rupture of ear drum|Acute suppurative otitis media with spontaneous rupture of ear drum
C0395866|T047|PT|194287004|SNOMEDCT_CORE|Recurrent acute otitis media|Recurrent acute otitis media
C0395866|T047|FN|194287004|SNOMEDCT_CORE|Recurrent acute otitis media|Recurrent acute otitis media
C0395869|T047|PT|232254004|SNOMEDCT_CORE|Chronic non-suppurative otitis media|Chronic non-suppurative otitis media
C0395869|T047|FN|232254004|SNOMEDCT_CORE|Chronic non-suppurative otitis media|Chronic non-suppurative otitis media
C0396000|T047|PT|195662009|SNOMEDCT_CORE|Acute viral pharyngitis|Acute viral pharyngitis
C0396000|T047|FN|195662009|SNOMEDCT_CORE|Acute viral pharyngitis|Acute viral pharyngitis
C0396024|T047|PT|195798007|SNOMEDCT_CORE|Chronic adenotonsillitis|Chronic adenotonsillitis
C0396024|T047|FN|195798007|SNOMEDCT_CORE|Chronic adenotonsillitis|Chronic adenotonsillitis
C0396053|T033|OAP|195853009|SNOMEDCT_CORE|Singers' chorditis|Singers' chorditis
C0396053|T033|OAF|195853009|SNOMEDCT_CORE|Singers' chorditis|Singers' chorditis
C0398350|T047|PT|360371003|SNOMEDCT_CORE|Acute cardiac pulmonary edema|Acute cardiac pulmonary edema
C0398350|T047|FN|360371003|SNOMEDCT_CORE|Acute cardiac pulmonary edema|Acute cardiac pulmonary edema
C0398350|T047|PTGB|360371003|SNOMEDCT_CORE|Acute cardiac pulmonary oedema|Acute cardiac pulmonary edema
C0398350|T047|SY|360371003|SNOMEDCT_CORE|Acute cardiogenic pulmonary edema|Acute cardiac pulmonary edema
C0398350|T047|SYGB|360371003|SNOMEDCT_CORE|Acute cardiogenic pulmonary oedema|Acute cardiac pulmonary edema
C0398350|T047|SY|360371003|SNOMEDCT_CORE|Cardiogenic pulmonary edema|Acute cardiac pulmonary edema
C0398350|T047|SYGB|360371003|SNOMEDCT_CORE|Cardiogenic pulmonary oedema|Acute cardiac pulmonary edema
C0398353|T046|IS|15993004|SNOMEDCT_CORE|Hypercapnic respiratory failure|Hypercapnic respiratory failure
C0398353|T046|IS|15993004|SNOMEDCT_CORE|Type 2 respiratory failure|Hypercapnic respiratory failure
C0398353|T046|IS|15993004|SNOMEDCT_CORE|Ventilatory failure|Hypercapnic respiratory failure
C0398623|T047|SY|76612001|SNOMEDCT_CORE|Hypercoagulability|Thrombophilia
C0398623|T047|PT|76612001|SNOMEDCT_CORE|Hypercoagulability state|Thrombophilia
C0398623|T047|FN|76612001|SNOMEDCT_CORE|Hypercoagulability state|Thrombophilia
C0398623|T047|IS|76612001|SNOMEDCT_CORE|Hypercoagulability state, NOS|Thrombophilia
C0398623|T047|SY|76612001|SNOMEDCT_CORE|Hypercoagulable state|Thrombophilia
C0398623|T047|PT|234467004|SNOMEDCT_CORE|Thrombophilia|Thrombophilia
C0398623|T047|FN|234467004|SNOMEDCT_CORE|Thrombophilia|Thrombophilia
C0398650|T047|SY|32273002|SNOMEDCT_CORE|Idiopathic purpura|Idiopathic thrombocytopenic purpura
C0398650|T047|IS|32273002|SNOMEDCT_CORE|Idiopathic purpura, NOS|Idiopathic thrombocytopenic purpura
C0398650|T047|PT|32273002|SNOMEDCT_CORE|Idiopathic thrombocytopenic purpura|Idiopathic thrombocytopenic purpura
C0398650|T047|FN|32273002|SNOMEDCT_CORE|Idiopathic thrombocytopenic purpura|Idiopathic thrombocytopenic purpura
C0398650|T047|IS|32273002|SNOMEDCT_CORE|Idiopathic thrombocytopenic purpura, NOS|Idiopathic thrombocytopenic purpura
C0398650|T047|OAP|234490009|SNOMEDCT_CORE|Immune thrombocytopenic purpura|Idiopathic thrombocytopenic purpura
C0398650|T047|SY|32273002|SNOMEDCT_CORE|Immune thrombocytopenic purpura|Idiopathic thrombocytopenic purpura
C0398650|T047|OAF|234490009|SNOMEDCT_CORE|Immune thrombocytopenic purpura|Idiopathic thrombocytopenic purpura
C0398650|T047|IS|32273002|SNOMEDCT_CORE|ITP|Idiopathic thrombocytopenic purpura
C0398650|T047|SY|32273002|SNOMEDCT_CORE|ITP - idiopathic thrombocytopenic purpura|Idiopathic thrombocytopenic purpura
C0398650|T047|IS|32273002|SNOMEDCT_CORE|ITP - Idiopathic thrombocytopenic purpura|Idiopathic thrombocytopenic purpura
C0398650|T047|SY|32273002|SNOMEDCT_CORE|ITP - immune thrombocytopenic purpura|Idiopathic thrombocytopenic purpura
C0398650|T047|IS|32273002|SNOMEDCT_CORE|ITP, NOS|Idiopathic thrombocytopenic purpura
C0399396|T047|OAS|5170009|SNOMEDCT_CORE|Carious exposure of pulp|Carious exposure of pulp
C0399396|T047|PT|700046006|SNOMEDCT_CORE|Carious exposure of pulp|Carious exposure of pulp
C0399396|T047|FN|700046006|SNOMEDCT_CORE|Carious exposure of pulp|Carious exposure of pulp
C0399396|T047|OAP|5170009|SNOMEDCT_CORE|Complex dental caries|Carious exposure of pulp
C0399396|T047|OAF|5170009|SNOMEDCT_CORE|Complex dental caries|Carious exposure of pulp
C0399396|T047|OAS|5170009|SNOMEDCT_CORE|Complex dental cavity|Carious exposure of pulp
C0399396|T047|OAS|5170009|SNOMEDCT_CORE|Dental caries extending to pulp|Carious exposure of pulp
C0399396|T047|SY|700046006|SNOMEDCT_CORE|Dental caries extending to pulp|Carious exposure of pulp
C0399461|T047|PT|235019006|SNOMEDCT_CORE|Erosion of oral mucosa|Erosion of oral mucosa
C0399461|T047|FN|235019006|SNOMEDCT_CORE|Erosion of oral mucosa|Erosion of oral mucosa
C0399551|T046|SY|196417006|SNOMEDCT_CORE|Impacted 8|Impacted third molar tooth
C0399551|T046|PT|196417006|SNOMEDCT_CORE|Impacted third molar tooth|Impacted third molar tooth
C0399551|T046|FN|196417006|SNOMEDCT_CORE|Impacted third molar tooth|Impacted third molar tooth
C0399551|T046|SY|196417006|SNOMEDCT_CORE|Impacted wisdom tooth|Impacted third molar tooth
C0399561|T047|OAP|266423006|SNOMEDCT_CORE|Inflammatory disorder of jaw|Inflammatory disorder of jaw
C0399561|T047|OAF|266423006|SNOMEDCT_CORE|Inflammatory disorder of jaw|Inflammatory disorder of jaw
C0399586|T047|SY|196500001|SNOMEDCT_CORE|Submandibular calculus|Submandibular sialolithiasis
C0399586|T047|PT|196500001|SNOMEDCT_CORE|Submandibular sialolithiasis|Submandibular sialolithiasis
C0399586|T047|FN|196500001|SNOMEDCT_CORE|Submandibular sialolithiasis|Submandibular sialolithiasis
C0400821|T047|PT|235753003|SNOMEDCT_CORE|Microscopic colitis|Microscopic colitis
C0400821|T047|FN|235753003|SNOMEDCT_CORE|Microscopic colitis|Microscopic colitis
C0400822|T047|SY|31437008|SNOMEDCT_CORE|Lymphocytic colitis|Lymphocytic-plasmacytic colitis
C0400822|T047|PT|31437008|SNOMEDCT_CORE|Lymphocytic-plasmacytic colitis|Lymphocytic-plasmacytic colitis
C0400822|T047|FN|31437008|SNOMEDCT_CORE|Lymphocytic-plasmacytic colitis|Lymphocytic-plasmacytic colitis
C0400827|T046|SY|235760009|SNOMEDCT_CORE|Radiation induced proctitis|Radiation proctitis
C0400827|T046|PT|235760009|SNOMEDCT_CORE|Radiation proctitis|Radiation proctitis
C0400827|T046|FN|235760009|SNOMEDCT_CORE|Radiation proctitis|Radiation proctitis
C0400839|T047|SY|54609002|SNOMEDCT_CORE|Rectal ulcer|Ulcer of rectum
C0400839|T047|SY|54609002|SNOMEDCT_CORE|Solitary rectal ulcer|Ulcer of rectum
C0400839|T047|SY|54609002|SNOMEDCT_CORE|Solitary ulcer of rectum|Ulcer of rectum
C0400839|T047|PT|54609002|SNOMEDCT_CORE|Ulcer of rectum|Ulcer of rectum
C0400839|T047|FN|54609002|SNOMEDCT_CORE|Ulcer of rectum|Ulcer of rectum
C0400851|T020|PT|235810006|SNOMEDCT_CORE|Bolus obstruction of intestine|Bolus obstruction of intestine
C0400851|T020|FN|235810006|SNOMEDCT_CORE|Bolus obstruction of intestine|Bolus obstruction of intestine
C0400865|T047|SY|235823004|SNOMEDCT_CORE|Bowel dyskinesia|Motility disorder of intestine
C0400865|T047|PT|235823004|SNOMEDCT_CORE|Motility disorder of intestine|Motility disorder of intestine
C0400865|T047|FN|235823004|SNOMEDCT_CORE|Motility disorder of intestine|Motility disorder of intestine
C0400914|T047|PT|235866006|SNOMEDCT_CORE|Acute hepatitis C|Acute hepatitis C
C0400914|T047|FN|235866006|SNOMEDCT_CORE|Acute hepatitis C|Acute hepatitis C
C0400920|T033|FN|235872006|SNOMEDCT_CORE|Hepatitis C carrier|Hepatitis C carrier
C0400920|T033|PT|235872006|SNOMEDCT_CORE|Hepatitis C carrier|Hepatitis C carrier
C0400943|T047|PT|266468003|SNOMEDCT_CORE|Cirrhosis - non-alcoholic|Cirrhosis - non-alcoholic
C0400943|T047|FN|266468003|SNOMEDCT_CORE|Cirrhosis - non-alcoholic|Cirrhosis - non-alcoholic
C0400943|T047|SY|266468003|SNOMEDCT_CORE|Cirrhosis of liver not due to alcohol|Cirrhosis - non-alcoholic
C0400943|T047|OAF|111370006|SNOMEDCT_CORE|Cirrhosis of liver not due to alcohol|Cirrhosis - non-alcoholic
C0400943|T047|OAP|111370006|SNOMEDCT_CORE|Cirrhosis of liver not due to alcohol|Cirrhosis - non-alcoholic
C0400943|T047|SY|266468003|SNOMEDCT_CORE|Cirrhosis, nonalcoholic|Cirrhosis - non-alcoholic
C0400966|T047|SY|197315008|SNOMEDCT_CORE|NAFLD - Nonalcoholic fatty liver disease|Non-alcoholic fatty liver
C0400966|T047|PT|197315008|SNOMEDCT_CORE|Non-alcoholic fatty liver|Non-alcoholic fatty liver
C0400966|T047|FN|197315008|SNOMEDCT_CORE|Non-alcoholic fatty liver|Non-alcoholic fatty liver
C0400968|T046|PT|235911006|SNOMEDCT_CORE|Liver transplant rejection|Liver transplant rejection
C0400968|T046|FN|235911006|SNOMEDCT_CORE|Liver transplant rejection|Liver transplant rejection
C0400979|T047|PT|235918000|SNOMEDCT_CORE|Obstruction of biliary tree|Obstruction of biliary tree
C0400979|T047|FN|235918000|SNOMEDCT_CORE|Obstruction of biliary tree|Obstruction of biliary tree
C0400985|T047|SY|197377009|SNOMEDCT_CORE|Cholelithiasis AND acute cholecystitis without obstruction|Gallbladder calculus with acute cholecystitis and no obstruction
C0400985|T047|PT|197377009|SNOMEDCT_CORE|Gallbladder calculus with acute cholecystitis and no obstruction|Gallbladder calculus with acute cholecystitis and no obstruction
C0400985|T047|FN|197377009|SNOMEDCT_CORE|Gallbladder calculus with acute cholecystitis and no obstruction|Gallbladder calculus with acute cholecystitis and no obstruction
C0401066|T020|OAP|62120000|SNOMEDCT_CORE|Unilateral recurrent inguinal hernia|Unilateral recurrent inguinal hernia
C0401066|T020|OF|62120000|SNOMEDCT_CORE|Unilateral recurrent inguinal hernia|Unilateral recurrent inguinal hernia
C0401066|T020|OAF|62120000|SNOMEDCT_CORE|Unilateral recurrent inguinal hernia|Unilateral recurrent inguinal hernia
C0401067|T020|OAP|52278004|SNOMEDCT_CORE|Unilateral inguinal hernia|Unilateral inguinal hernia
C0401067|T020|OF|52278004|SNOMEDCT_CORE|Unilateral inguinal hernia|Unilateral inguinal hernia
C0401067|T020|OAF|52278004|SNOMEDCT_CORE|Unilateral inguinal hernia|Unilateral inguinal hernia
C0401096|T020|OF|60016005|SNOMEDCT_CORE|Unilateral femoral hernia without obstruction AND without gangrene|Unilateral femoral hernia without obstruction AND without gangrene
C0401096|T020|OAP|60016005|SNOMEDCT_CORE|Unilateral femoral hernia without obstruction AND without gangrene|Unilateral femoral hernia without obstruction AND without gangrene
C0401096|T020|OAF|60016005|SNOMEDCT_CORE|Unilateral femoral hernia without obstruction AND without gangrene|Unilateral femoral hernia without obstruction AND without gangrene
C0401096|T020|IS|60016005|SNOMEDCT_CORE|Unilateral femoral hernia without obstruction or gangrene|Unilateral femoral hernia without obstruction AND without gangrene
C0401096|T020|OAS|60016005|SNOMEDCT_CORE|Unilateral simple femoral hernia|Unilateral femoral hernia without obstruction AND without gangrene
C0401103|T020|OAP|38897008|SNOMEDCT_CORE|Unilateral femoral hernia with obstruction but no gangrene|Unilateral femoral hernia with obstruction but no gangrene
C0401103|T020|OF|38897008|SNOMEDCT_CORE|Unilateral femoral hernia with obstruction but no gangrene|Unilateral femoral hernia with obstruction but no gangrene
C0401103|T020|OAF|38897008|SNOMEDCT_CORE|Unilateral femoral hernia with obstruction but no gangrene|Unilateral femoral hernia with obstruction but no gangrene
C0401103|T020|OAS|38897008|SNOMEDCT_CORE|Unilateral obstructed femoral hernia|Unilateral femoral hernia with obstruction but no gangrene
C0401115|T020|PT|236042008|SNOMEDCT_CORE|Obstructed internal hernia|Obstructed internal hernia
C0401115|T020|FN|236042008|SNOMEDCT_CORE|Obstructed internal hernia|Obstructed internal hernia
C0401146|T047|PT|197118003|SNOMEDCT_CORE|Constipation - functional|Constipation - functional
C0401146|T047|FN|197118003|SNOMEDCT_CORE|Constipation - functional|Constipation - functional
C0401146|T047|SY|197118003|SNOMEDCT_CORE|Constipation-functional|Constipation - functional
C0401146|T047|SY|197118003|SNOMEDCT_CORE|Functional constipation|Constipation - functional
C0401149|T184|PT|236069009|SNOMEDCT_CORE|Chronic constipation|Chronic constipation
C0401149|T184|OF|236069009|SNOMEDCT_CORE|Chronic constipation|Chronic constipation
C0401149|T184|FN|236069009|SNOMEDCT_CORE|Chronic constipation|Chronic constipation
C0401151|T047|PT|236071009|SNOMEDCT_CORE|Chronic diarrhea|Chronic diarrhea
C0401151|T047|FN|236071009|SNOMEDCT_CORE|Chronic diarrhea|Chronic diarrhea
C0401151|T047|PTGB|236071009|SNOMEDCT_CORE|Chronic diarrhoea|Chronic diarrhea
C0403419|T047|PT|197618004|SNOMEDCT_CORE|Chronic focal glomerulonephritis|Chronic focal glomerulonephritis
C0403419|T047|FN|197618004|SNOMEDCT_CORE|Chronic focal glomerulonephritis|Chronic focal glomerulonephritis
C0403447|T047|OAP|236425005|SNOMEDCT_CORE|Chronic renal impairment|Chronic renal impairment
C0403447|T047|SY|709044004|SNOMEDCT_CORE|Chronic renal impairment|Chronic renal impairment
C0403447|T047|OAF|236425005|SNOMEDCT_CORE|Chronic renal impairment|Chronic renal impairment
C0403462|T047|SY|236433006|SNOMEDCT_CORE|Acute on chronic renal failure|Acute-on-chronic renal failure
C0403462|T047|PT|236433006|SNOMEDCT_CORE|Acute-on-chronic renal failure|Acute-on-chronic renal failure
C0403462|T047|FN|236433006|SNOMEDCT_CORE|Acute-on-chronic renal failure|Acute-on-chronic renal failure
C0403464|T047|PT|236435004|SNOMEDCT_CORE|End stage renal failure on dialysis|End stage renal failure on dialysis
C0403464|T047|FN|236435004|SNOMEDCT_CORE|End stage renal failure on dialysis|End stage renal failure on dialysis
C0403496|T047|SY|199132007|SNOMEDCT_CORE|Glycosuria during pregnancy|Pregnancy-related glycosuria
C0403496|T047|PT|199132007|SNOMEDCT_CORE|Pregnancy-related glycosuria|Pregnancy-related glycosuria
C0403496|T047|FN|199132007|SNOMEDCT_CORE|Pregnancy-related glycosuria|Pregnancy-related glycosuria
C0403571|T047|SY|236557008|SNOMEDCT_CORE|Peritoneal dialysis cannula exit site infection|Peritoneal dialysis catheter exit site infection
C0403571|T047|PT|236557008|SNOMEDCT_CORE|Peritoneal dialysis catheter exit site infection|Peritoneal dialysis catheter exit site infection
C0403571|T047|FN|236557008|SNOMEDCT_CORE|Peritoneal dialysis catheter exit site infection|Peritoneal dialysis catheter exit site infection
C0403576|T033|SY|236562009|SNOMEDCT_CORE|Blockage of peritoneal dialysis catheter|Obstruction of peritoneal dialysis catheter
C0403576|T033|PT|236562009|SNOMEDCT_CORE|Obstruction of peritoneal dialysis catheter|Obstruction of peritoneal dialysis catheter
C0403576|T033|FN|236562009|SNOMEDCT_CORE|Obstruction of peritoneal dialysis catheter|Obstruction of peritoneal dialysis catheter
C0403641|T047|PT|236632007|SNOMEDCT_CORE|Functional disorder of bladder|Functional disorder of bladder
C0403641|T047|FN|236632007|SNOMEDCT_CORE|Functional disorder of bladder|Functional disorder of bladder
C0403641|T047|SY|236632007|SNOMEDCT_CORE|Functional voiding disorder|Functional disorder of bladder
C0403643|T047|OAP|236633002|SNOMEDCT_CORE|Bladder muscle dysfunction - overactive|Bladder muscle dysfunction - overactive
C0403643|T047|OAF|236633002|SNOMEDCT_CORE|Bladder muscle dysfunction - overactive|Bladder muscle dysfunction - overactive
C0403645|T033|PT|197870000|SNOMEDCT_CORE|Acontractile detrusor|Acontractile detrusor
C0403645|T033|FN|197870000|SNOMEDCT_CORE|Acontractile detrusor|Acontractile detrusor
C0403645|T033|SY|197870000|SNOMEDCT_CORE|Atonic bladder|Acontractile detrusor
C0403645|T033|SY|197870000|SNOMEDCT_CORE|Atonic urinary bladder|Acontractile detrusor
C0403645|T033|SY|197870000|SNOMEDCT_CORE|Atony of bladder|Acontractile detrusor
C0403647|T047|FN|197871001|SNOMEDCT_CORE|Hypotonic bladder|Hypotonic bladder
C0403647|T047|PT|197871001|SNOMEDCT_CORE|Hypotonic bladder|Hypotonic bladder
C0403647|T047|SY|197871001|SNOMEDCT_CORE|Hypotonicity of bladder|Hypotonic bladder
C0403654|T020|PT|236645006|SNOMEDCT_CORE|Bladder outflow obstruction|Bladder outflow obstruction
C0403654|T020|FN|236645006|SNOMEDCT_CORE|Bladder outflow obstruction|Bladder outflow obstruction
C0403654|T020|SY|236645006|SNOMEDCT_CORE|BOO - Bladder outflow obstruction|Bladder outflow obstruction
C0403668|T033|SY|236664000|SNOMEDCT_CORE|PMD - Post-micturition dribbling|Post-micturition incontinence
C0403668|T033|SY|236664000|SNOMEDCT_CORE|Post-micturition dribbling|Post-micturition incontinence
C0403668|T033|PT|236664000|SNOMEDCT_CORE|Post-micturition incontinence|Post-micturition incontinence
C0403668|T033|FN|236664000|SNOMEDCT_CORE|Post-micturition incontinence|Post-micturition incontinence
C0403698|T037|SY|86347007|SNOMEDCT_CORE|Post-traumatic urethral stricture|Traumatic urethral stricture
C0403698|T037|PT|86347007|SNOMEDCT_CORE|Traumatic urethral stricture|Traumatic urethral stricture
C0403698|T037|FN|86347007|SNOMEDCT_CORE|Traumatic urethral stricture|Traumatic urethral stricture
C0403709|T047|PT|197926005|SNOMEDCT_CORE|Postoperative urinary tract infection|Postoperative urinary tract infection
C0403709|T047|FN|197926005|SNOMEDCT_CORE|Postoperative urinary tract infection|Postoperative urinary tract infection
C0403714|T047|PT|236708007|SNOMEDCT_CORE|Calyceal renal calculus|Calyceal renal calculus
C0403714|T047|FN|236708007|SNOMEDCT_CORE|Calyceal renal calculus|Calyceal renal calculus
C0403714|T047|SY|236708007|SNOMEDCT_CORE|Calyceal stone|Calyceal renal calculus
C0403717|T047|PT|236711008|SNOMEDCT_CORE|Calculus in pelviureteric junction|Calculus in pelviureteric junction
C0403717|T047|FN|236711008|SNOMEDCT_CORE|Calculus in pelviureteric junction|Calculus in pelviureteric junction
C0403717|T047|SY|236711008|SNOMEDCT_CORE|Stone in pelviureteric junction|Calculus in pelviureteric junction
C0403717|T047|SY|236711008|SNOMEDCT_CORE|Stone in PUJ - pelviureteric junction|Calculus in pelviureteric junction
C0403719|T047|IS|267441009|SNOMEDCT_CORE|Uric acid nephrolithiasis|Uric acid urolithiasis
C0403719|T047|PT|267441009|SNOMEDCT_CORE|Uric acid urolithiasis|Uric acid urolithiasis
C0403719|T047|FN|267441009|SNOMEDCT_CORE|Uric acid urolithiasis|Uric acid urolithiasis
C0404478|T047|SY|95598005|SNOMEDCT_CORE|Rupture of ovarian cyst|Ruptured cyst of ovary
C0404478|T047|PT|95598005|SNOMEDCT_CORE|Ruptured cyst of ovary|Ruptured cyst of ovary
C0404478|T047|FN|95598005|SNOMEDCT_CORE|Ruptured cyst of ovary|Ruptured cyst of ovary
C0404478|T047|SY|95598005|SNOMEDCT_CORE|Ruptured ovarian cyst|Ruptured cyst of ovary
C0404478|T047|IS|95598005|SNOMEDCT_CORE|Ruptured ovarian cyst, NOS|Ruptured cyst of ovary
C0404484|T184|FN|237067000|SNOMEDCT_CORE|Chronic pain in female pelvis|Chronic pelvic pain of female
C0404484|T184|SY|237067000|SNOMEDCT_CORE|Chronic pain in female pelvis|Chronic pelvic pain of female
C0404484|T184|IS|237067000|SNOMEDCT_CORE|Chronic pelvic pain|Chronic pelvic pain of female
C0404484|T184|PT|237067000|SNOMEDCT_CORE|Chronic pelvic pain of female|Chronic pelvic pain of female
C0404484|T184|OF|237067000|SNOMEDCT_CORE|Chronic pelvic pain of female|Chronic pelvic pain of female
C0404532|T020|PT|198279007|SNOMEDCT_CORE|Lax vaginal introitus|Lax vaginal introitus
C0404532|T020|FN|198279007|SNOMEDCT_CORE|Lax vaginal introitus|Lax vaginal introitus
C0404532|T020|OF|198279007|SNOMEDCT_CORE|Lax vaginal introitus|Lax vaginal introitus
C0404532|T020|SY|198279007|SNOMEDCT_CORE|Relaxation of vaginal outlet|Lax vaginal introitus
C0404559|T047|PT|266607004|SNOMEDCT_CORE|Perimenopausal disorder|Perimenopausal disorder
C0404559|T047|FN|266607004|SNOMEDCT_CORE|Perimenopausal disorder|Perimenopausal disorder
C0404572|T047|SY|266609001|SNOMEDCT_CORE|Anovulatory infertility|Female infertility of anovulatory origin
C0404572|T047|PT|266609001|SNOMEDCT_CORE|Female infertility of anovulatory origin|Female infertility of anovulatory origin
C0404572|T047|FN|266609001|SNOMEDCT_CORE|Female infertility of anovulatory origin|Female infertility of anovulatory origin
C0404596|T019|OAP|199516000|SNOMEDCT_CORE|Known or suspected fetal abnormality|Known or suspected fetal abnormality
C0404596|T019|OAP|609414006|SNOMEDCT_CORE|Known or suspected fetal abnormality|Known or suspected fetal abnormality
C0404596|T019|OAF|609414006|SNOMEDCT_CORE|Known or suspected fetal abnormality|Known or suspected fetal abnormality
C0404596|T019|OAF|199516000|SNOMEDCT_CORE|Known or suspected fetal abnormality|Known or suspected fetal abnormality
C0404596|T019|OAP|609414006|SNOMEDCT_CORE|Known or suspected foetal abnormality|Known or suspected fetal abnormality
C0404734|T033|PT|372054004|SNOMEDCT_CORE|Abnormal glucose tolerance test during pregnancy - baby not yet delivered|Abnormal glucose tolerance test during pregnancy - baby not yet delivered
C0404734|T033|FN|372054004|SNOMEDCT_CORE|Abnormal glucose tolerance test during pregnancy - baby not yet delivered|Abnormal glucose tolerance test during pregnancy - baby not yet delivered
C0404753|T048|PT|199257008|SNOMEDCT_CORE|Mental disorders during pregnancy, childbirth and the puerperium|Mental disorders during pregnancy, childbirth and the puerperium
C0404753|T048|FN|199257008|SNOMEDCT_CORE|Mental disorders during pregnancy, childbirth and the puerperium|Mental disorders during pregnancy, childbirth and the puerperium
C0404831|T033|PT|102876002|SNOMEDCT_CORE|Multigravida|Multigravida
C0404831|T033|FN|102876002|SNOMEDCT_CORE|Multigravida|Multigravida
C0404831|T033|SY|102876002|SNOMEDCT_CORE|Multip|Multigravida
C0404831|T033|IS|102876002|SNOMEDCT_CORE|Multiple previous pregnancies|Multigravida
C0404831|T033|IS|102876002|SNOMEDCT_CORE|Multiple previous pregnancies, NOS|Multigravida
C0404889|T033|SY|199088001|SNOMEDCT_CORE|Habitual aborter - not delivered|History of recurrent miscarriage - not delivered
C0404889|T033|FN|199088001|SNOMEDCT_CORE|Habitual aborter - not delivered|History of recurrent miscarriage - not delivered
C0404889|T033|PT|199088001|SNOMEDCT_CORE|History of recurrent miscarriage - not delivered|History of recurrent miscarriage - not delivered
C0405092|T046|PT|199064003|SNOMEDCT_CORE|Post-term pregnancy - not delivered|Post-term pregnancy - not delivered
C0405092|T046|FN|199064003|SNOMEDCT_CORE|Post-term pregnancy - not delivered|Post-term pregnancy - not delivered
C0406072|T047|OAP|200665006|SNOMEDCT_CORE|Cellulitis and abscess of arm|Cellulitis and abscess of arm
C0406072|T047|OAF|200665006|SNOMEDCT_CORE|Cellulitis and abscess of arm|Cellulitis and abscess of arm
C0406078|T047|PT|267780000|SNOMEDCT_CORE|Cellulitis and abscess of hand excluding digits|Cellulitis and abscess of hand excluding digits
C0406078|T047|FN|267780000|SNOMEDCT_CORE|Cellulitis and abscess of hand excluding digits|Cellulitis and abscess of hand excluding digits
C0406085|T047|PT|200681001|SNOMEDCT_CORE|Cellulitis and abscess of lower leg|Cellulitis and abscess of lower leg
C0406085|T047|FN|200681001|SNOMEDCT_CORE|Cellulitis and abscess of lower leg|Cellulitis and abscess of lower leg
C0406086|T047|PT|200682008|SNOMEDCT_CORE|Cellulitis and abscess of ankle|Cellulitis and abscess of ankle
C0406086|T047|FN|200682008|SNOMEDCT_CORE|Cellulitis and abscess of ankle|Cellulitis and abscess of ankle
C0406087|T047|OAP|267782008|SNOMEDCT_CORE|Cellulitis and abscess of leg|Cellulitis and abscess of leg
C0406087|T047|OAF|267782008|SNOMEDCT_CORE|Cellulitis and abscess of leg|Cellulitis and abscess of leg
C0406087|T047|OAS|267782008|SNOMEDCT_CORE|Leg cellulitis/abscess|Cellulitis and abscess of leg
C0406089|T047|PT|267783003|SNOMEDCT_CORE|Cellulitis and abscess of foot excluding toe|Cellulitis and abscess of foot excluding toe
C0406089|T047|FN|267783003|SNOMEDCT_CORE|Cellulitis and abscess of foot excluding toe|Cellulitis and abscess of foot excluding toe
C0406169|T047|SY|201040000|SNOMEDCT_CORE|Hyperkeratotic callus|Hyperkeratotic callus
C0406252|T047|PT|201201000|SNOMEDCT_CORE|Podopompholyx|Podopompholyx
C0406252|T047|FN|201201000|SNOMEDCT_CORE|Podopompholyx|Podopompholyx
C0406252|T047|SY|201201000|SNOMEDCT_CORE|Vesicular eczema of feet|Podopompholyx
C0406319|T047|PT|238602009|SNOMEDCT_CORE|Psoriasis-eczema overlap condition|Psoriasis-eczema overlap condition
C0406319|T047|FN|238602009|SNOMEDCT_CORE|Psoriasis-eczema overlap condition|Psoriasis-eczema overlap condition
C0406319|T047|IS|238602009|SNOMEDCT_CORE|Sebopsoriasis|Psoriasis-eczema overlap condition
C0406481|T047|PT|238744006|SNOMEDCT_CORE|Comedonal acne|Comedonal acne
C0406481|T047|FN|238744006|SNOMEDCT_CORE|Comedonal acne|Comedonal acne
C0406484|T047|SY|238748009|SNOMEDCT_CORE|Benign seborrheic hyperplasia|Sebaceous hyperplasia
C0406484|T047|SYGB|238748009|SNOMEDCT_CORE|Benign seborrhoeic hyperplasia|Sebaceous hyperplasia
C0406484|T047|SY|238748009|SNOMEDCT_CORE|Sebaceous gland hyperplasia|Sebaceous hyperplasia
C0406484|T047|PT|238748009|SNOMEDCT_CORE|Sebaceous hyperplasia|Sebaceous hyperplasia
C0406484|T047|FN|238748009|SNOMEDCT_CORE|Sebaceous hyperplasia|Sebaceous hyperplasia
C0406486|T047|PT|200933006|SNOMEDCT_CORE|Ocular rosacea|Ocular rosacea
C0406486|T047|FN|200933006|SNOMEDCT_CORE|Ocular rosacea|Ocular rosacea
C0406500|T047|PT|410016009|SNOMEDCT_CORE|Lipodermatosclerosis|Lipodermatosclerosis
C0406500|T047|FN|410016009|SNOMEDCT_CORE|Lipodermatosclerosis|Lipodermatosclerosis
C0406524|T047|SY|35222003|SNOMEDCT_CORE|Chronic neurogenic ulcer of leg|Chronic neurogenic ulcer of lower limb
C0406524|T047|IS|35222003|SNOMEDCT_CORE|Chronic neurogenic ulcer of leg, NOS|Chronic neurogenic ulcer of lower limb
C0406524|T047|PT|35222003|SNOMEDCT_CORE|Chronic neurogenic ulcer of lower limb|Chronic neurogenic ulcer of lower limb
C0406524|T047|FN|35222003|SNOMEDCT_CORE|Chronic neurogenic ulcer of lower limb|Chronic neurogenic ulcer of lower limb
C0406524|T047|SY|35222003|SNOMEDCT_CORE|Neurogenic leg ulcer|Chronic neurogenic ulcer of lower limb
C0406524|T047|SY|35222003|SNOMEDCT_CORE|Neuropathic leg ulcer|Chronic neurogenic ulcer of lower limb
C0406524|T047|IS|35222003|SNOMEDCT_CORE|Trophic leg ulcer|Chronic neurogenic ulcer of lower limb
C0406670|T047|IS|238968009|SNOMEDCT_CORE|Burning vulva|Vulvodynia
C0406670|T047|SY|162145001|SNOMEDCT_CORE|Pain of vulva|Vulvodynia
C0406670|T047|PT|162145001|SNOMEDCT_CORE|Vulval pain|Vulvodynia
C0406670|T047|FN|162145001|SNOMEDCT_CORE|Vulval pain|Vulvodynia
C0406670|T047|PT|238968009|SNOMEDCT_CORE|Vulvodynia|Vulvodynia
C0406670|T047|FN|238968009|SNOMEDCT_CORE|Vulvodynia|Vulvodynia
C0409204|T047|SY|442246002|SNOMEDCT_CORE|Arthropathy of ankle and/or foot|Disorder of joint of ankle and/or foot
C0409204|T047|PT|442246002|SNOMEDCT_CORE|Disorder of joint of ankle and/or foot|Disorder of joint of ankle and/or foot
C0409204|T047|FN|442246002|SNOMEDCT_CORE|Disorder of joint of ankle and/or foot|Disorder of joint of ankle and/or foot
C0409212|T047|PT|439656005|SNOMEDCT_CORE|Arthritis of elbow|Arthritis of elbow
C0409212|T047|FN|439656005|SNOMEDCT_CORE|Arthritis of elbow|Arthritis of elbow
C0409310|T037|SY|239724009|SNOMEDCT_CORE|ACL - Anterior cruciate ligament deficiency|Deficiency of anterior cruciate ligament
C0409310|T037|PT|239724009|SNOMEDCT_CORE|Deficiency of anterior cruciate ligament|Deficiency of anterior cruciate ligament
C0409310|T037|FN|239724009|SNOMEDCT_CORE|Deficiency of anterior cruciate ligament|Deficiency of anterior cruciate ligament
C0409312|T037|SY|239725005|SNOMEDCT_CORE|ACL - Anterior cruciate ligament rupture|Rupture of anterior cruciate ligament
C0409312|T037|SY|239725005|SNOMEDCT_CORE|Anterior cruciate ligament rupture|Rupture of anterior cruciate ligament
C0409312|T037|PT|239725005|SNOMEDCT_CORE|Rupture of anterior cruciate ligament|Rupture of anterior cruciate ligament
C0409312|T037|FN|239725005|SNOMEDCT_CORE|Rupture of anterior cruciate ligament|Rupture of anterior cruciate ligament
C0409312|T037|SY|239725005|SNOMEDCT_CORE|Tear of anterior cruciate ligament|Rupture of anterior cruciate ligament
C0409316|T037|SY|239727002|SNOMEDCT_CORE|PCL - Posterior cruciate ligament rupture|Rupture of posterior cruciate ligament
C0409316|T037|PT|239727002|SNOMEDCT_CORE|Rupture of posterior cruciate ligament|Rupture of posterior cruciate ligament
C0409316|T037|FN|239727002|SNOMEDCT_CORE|Rupture of posterior cruciate ligament|Rupture of posterior cruciate ligament
C0409316|T037|SY|239727002|SNOMEDCT_CORE|Tear of posterior cruciate ligament|Rupture of posterior cruciate ligament
C0409320|T037|SY|239729004|SNOMEDCT_CORE|MCL - Medial collateral ligament rupture of the knee|Rupture of medial collateral ligament of knee
C0409320|T037|PT|239729004|SNOMEDCT_CORE|Rupture of medial collateral ligament of knee|Rupture of medial collateral ligament of knee
C0409320|T037|FN|239729004|SNOMEDCT_CORE|Rupture of medial collateral ligament of knee|Rupture of medial collateral ligament of knee
C0409320|T037|SY|239729004|SNOMEDCT_CORE|Tear of medial collateral ligament of knee joint|Rupture of medial collateral ligament of knee
C0409377|T037|PT|202248001|SNOMEDCT_CORE|Recurrent subluxation of the patella|Recurrent subluxation of the patella
C0409377|T037|FN|202248001|SNOMEDCT_CORE|Recurrent subluxation of the patella|Recurrent subluxation of the patella
C0409415|T037|IS|30556007|SNOMEDCT_CORE|Recurrent dislocation of shoulder|Recurrent dislocation of shoulder
C0409415|T037|IS|30556007|SNOMEDCT_CORE|Recurrent dislocation of the shoulder joint|Recurrent dislocation of shoulder
C0409542|T047|PT|239777004|SNOMEDCT_CORE|Knee pyogenic arthritis|Knee pyogenic arthritis
C0409542|T047|FN|239777004|SNOMEDCT_CORE|Knee pyogenic arthritis|Knee pyogenic arthritis
C0409651|T047|PT|239791005|SNOMEDCT_CORE|Seropositive rheumatoid arthritis|Seropositive rheumatoid arthritis
C0409651|T047|FN|239791005|SNOMEDCT_CORE|Seropositive rheumatoid arthritis|Seropositive rheumatoid arthritis
C0409652|T047|PT|239792003|SNOMEDCT_CORE|Seronegative rheumatoid arthritis|Seronegative rheumatoid arthritis
C0409652|T047|FN|239792003|SNOMEDCT_CORE|Seronegative rheumatoid arthritis|Seronegative rheumatoid arthritis
C0409738|T037|SY|201954006|SNOMEDCT_CORE|Traumatic arthropathy of ankle|Traumatic arthropathy-ankle
C0409738|T037|FN|201954006|SNOMEDCT_CORE|Traumatic arthropathy of ankle|Traumatic arthropathy-ankle
C0409738|T037|PT|201954006|SNOMEDCT_CORE|Traumatic arthropathy-ankle|Traumatic arthropathy-ankle
C0409738|T037|OF|201954006|SNOMEDCT_CORE|Traumatic arthropathy-ankle|Traumatic arthropathy-ankle
C0409754|T037|SY|201938008|SNOMEDCT_CORE|Traumatic arthropathy of the ankle and foot|Traumatic arthropathy of the ankle and/or foot
C0409754|T037|OF|201938008|SNOMEDCT_CORE|Traumatic arthropathy of the ankle and foot|Traumatic arthropathy of the ankle and/or foot
C0409754|T037|PT|201938008|SNOMEDCT_CORE|Traumatic arthropathy of the ankle and/or foot|Traumatic arthropathy of the ankle and/or foot
C0409754|T037|FN|201938008|SNOMEDCT_CORE|Traumatic arthropathy of the ankle and/or foot|Traumatic arthropathy of the ankle and/or foot
C0409755|T037|OAP|201937003|SNOMEDCT_CORE|Traumatic arthropathy of the lower leg|Traumatic arthropathy of the lower leg
C0409755|T037|OAF|201937003|SNOMEDCT_CORE|Traumatic arthropathy of the lower leg|Traumatic arthropathy of the lower leg
C0409860|T047|IS|415352004|SNOMEDCT_CORE|Milwaukee shoulder|Rotator cuff tear arthropathy
C0409860|T047|PT|415352004|SNOMEDCT_CORE|Rotator cuff tear arthropathy|Rotator cuff tear arthropathy
C0409860|T047|FN|415352004|SNOMEDCT_CORE|Rotator cuff tear arthropathy|Rotator cuff tear arthropathy
C0409895|T047|OAS|60782007|SNOMEDCT_CORE|Idiopathic articular chondrocalcinosis|Idiopathic articular chondrocalcinosis
C0409931|T047|SY|239874001|SNOMEDCT_CORE|Degenerative joint disease of ankle|Osteoarthritis of ankle
C0409931|T047|SY|239874001|SNOMEDCT_CORE|OA - Osteoarthritis of ankle|Osteoarthritis of ankle
C0409931|T047|PT|239874001|SNOMEDCT_CORE|Osteoarthritis of ankle|Osteoarthritis of ankle
C0409931|T047|FN|239874001|SNOMEDCT_CORE|Osteoarthritis of ankle|Osteoarthritis of ankle
C0409936|T047|SY|239868001|SNOMEDCT_CORE|Degenerative joint disease of finger|Osteoarthritis of finger joint
C0409936|T047|SY|239868001|SNOMEDCT_CORE|OA - Osteoarthritis of joint of finger|Osteoarthritis of finger joint
C0409936|T047|SY|239868001|SNOMEDCT_CORE|Osteoarthritis of finger|Osteoarthritis of finger joint
C0409936|T047|PT|239868001|SNOMEDCT_CORE|Osteoarthritis of finger joint|Osteoarthritis of finger joint
C0409936|T047|FN|239868001|SNOMEDCT_CORE|Osteoarthritis of finger joint|Osteoarthritis of finger joint
C0409939|T047|SY|373623009|SNOMEDCT_CORE|Degenerative joint disease of glenohumeral joint|Osteoarthritis of glenohumeral joint
C0409939|T047|PT|67315001|SNOMEDCT_CORE|Degenerative joint disease of shoulder region|Osteoarthritis of glenohumeral joint
C0409939|T047|FN|67315001|SNOMEDCT_CORE|Degenerative joint disease of shoulder region|Osteoarthritis of glenohumeral joint
C0409939|T047|SY|67315001|SNOMEDCT_CORE|OA - Osteoarthritis of shoulder|Osteoarthritis of glenohumeral joint
C0409939|T047|PT|373623009|SNOMEDCT_CORE|Osteoarthritis of glenohumeral joint|Osteoarthritis of glenohumeral joint
C0409939|T047|FN|373623009|SNOMEDCT_CORE|Osteoarthritis of glenohumeral joint|Osteoarthritis of glenohumeral joint
C0409939|T047|SY|67315001|SNOMEDCT_CORE|Osteoarthritis of shoulder|Osteoarthritis of glenohumeral joint
C0409939|T047|SY|67315001|SNOMEDCT_CORE|Osteoarthritis of shoulder joint|Osteoarthritis of glenohumeral joint
C0409939|T047|SY|67315001|SNOMEDCT_CORE|Osteoarthritis of shoulder region|Osteoarthritis of glenohumeral joint
C0409954|T047|IS|239866002|SNOMEDCT_CORE|Degenerative joint diease of elbow|Osteoarthritis of elbow
C0409954|T047|SY|239866002|SNOMEDCT_CORE|Degenerative joint disease of elbow|Osteoarthritis of elbow
C0409954|T047|SY|239866002|SNOMEDCT_CORE|OA - Osteoarthritis of elbow|Osteoarthritis of elbow
C0409954|T047|PT|239866002|SNOMEDCT_CORE|Osteoarthritis of elbow|Osteoarthritis of elbow
C0409954|T047|FN|239866002|SNOMEDCT_CORE|Osteoarthritis of elbow|Osteoarthritis of elbow
C0409955|T047|SY|239867006|SNOMEDCT_CORE|Degenerative joint disease of wrist|Osteoarthritis of wrist
C0409955|T047|SY|239867006|SNOMEDCT_CORE|OA - Osteoarthritis of wrist|Osteoarthritis of wrist
C0409955|T047|PT|239867006|SNOMEDCT_CORE|Osteoarthritis of wrist|Osteoarthritis of wrist
C0409955|T047|FN|239867006|SNOMEDCT_CORE|Osteoarthritis of wrist|Osteoarthritis of wrist
C0409956|T047|SY|37895003|SNOMEDCT_CORE|Osteoarthritis basilar joint of thumb|Osteoarthrosis of the carpometacarpal joint of the thumb
C0409956|T047|SY|37895003|SNOMEDCT_CORE|Osteoarthritis of first carpometacarpal joint|Osteoarthrosis of the carpometacarpal joint of the thumb
C0409956|T047|PT|37895003|SNOMEDCT_CORE|Osteoarthrosis of the carpometacarpal joint of the thumb|Osteoarthrosis of the carpometacarpal joint of the thumb
C0409956|T047|FN|37895003|SNOMEDCT_CORE|Osteoarthrosis of the carpometacarpal joint of the thumb|Osteoarthrosis of the carpometacarpal joint of the thumb
C0409959|T047|SY|239873007|SNOMEDCT_CORE|Degenerative joint disease of knee|Osteoarthritis of knee
C0409959|T047|SY|239873007|SNOMEDCT_CORE|Gonarthrosis|Osteoarthritis of knee
C0409959|T047|SY|239873007|SNOMEDCT_CORE|Knee DJD|Osteoarthritis of knee
C0409959|T047|IS|239873007|SNOMEDCT_CORE|Knee DJD|Osteoarthritis of knee
C0409959|T047|SY|239873007|SNOMEDCT_CORE|OA - Osteoarthritis of knee|Osteoarthritis of knee
C0409959|T047|PT|239873007|SNOMEDCT_CORE|Osteoarthritis of knee|Osteoarthritis of knee
C0409959|T047|FN|239873007|SNOMEDCT_CORE|Osteoarthritis of knee|Osteoarthritis of knee
C0409961|T047|PT|1679003|SNOMEDCT_CORE|Arthritis associated with another disorder|Arthritis associated with another disorder
C0409961|T047|FN|1679003|SNOMEDCT_CORE|Arthritis associated with another disorder|Arthritis associated with another disorder
C0409961|T047|IS|1679003|SNOMEDCT_CORE|Arthritis associated with disorder classified elsewhere|Arthritis associated with another disorder
C0409963|T047|SY|239865003|SNOMEDCT_CORE|Degenerative joint disease of acromioclavicular joint|Osteoarthritis of acromioclavicular joint
C0409963|T047|SY|239865003|SNOMEDCT_CORE|OA - Osteoarthritis of acromioclavicular joint|Osteoarthritis of acromioclavicular joint
C0409963|T047|PT|239865003|SNOMEDCT_CORE|Osteoarthritis of acromioclavicular joint|Osteoarthritis of acromioclavicular joint
C0409963|T047|FN|239865003|SNOMEDCT_CORE|Osteoarthritis of acromioclavicular joint|Osteoarthritis of acromioclavicular joint
C0409974|T047|SY|200936003|SNOMEDCT_CORE|LE - Lupus erythematosus|Lupus erythematosus
C0409974|T047|SY|200936003|SNOMEDCT_CORE|Lupus|Lupus erythematosus
C0409974|T047|PT|200936003|SNOMEDCT_CORE|Lupus erythematosus|Lupus erythematosus
C0409974|T047|FN|200936003|SNOMEDCT_CORE|Lupus erythematosus|Lupus erythematosus
C0409999|T047|PT|239918008|SNOMEDCT_CORE|Undifferentiated connective tissue disease|Undifferentiated connective tissue disease
C0409999|T047|FN|239918008|SNOMEDCT_CORE|Undifferentiated connective tissue disease|Undifferentiated connective tissue disease
C0410017|T037|SY|202843000|SNOMEDCT_CORE|Complete rupture of rotator cuff|Full thickness rotator cuff tear
C0410017|T037|PT|202843000|SNOMEDCT_CORE|Full thickness rotator cuff tear|Full thickness rotator cuff tear
C0410017|T037|FN|202843000|SNOMEDCT_CORE|Full thickness rotator cuff tear|Full thickness rotator cuff tear
C0410031|T047|IS|239965002|SNOMEDCT_CORE|Tendinitis and tenosynovitis of the elbow region|Tendinitis AND/OR tenosynovitis of the elbow region
C0410031|T047|OF|239965002|SNOMEDCT_CORE|Tendinitis and tenosynovitis of the elbow region|Tendinitis AND/OR tenosynovitis of the elbow region
C0410031|T047|OAF|239965002|SNOMEDCT_CORE|Tendinitis AND/OR tenosynovitis of the elbow region|Tendinitis AND/OR tenosynovitis of the elbow region
C0410031|T047|OAP|239965002|SNOMEDCT_CORE|Tendinitis AND/OR tenosynovitis of the elbow region|Tendinitis AND/OR tenosynovitis of the elbow region
C0410031|T047|OAS|239965002|SNOMEDCT_CORE|Tendonitis AND/OR tenosynovitis of the elbow region|Tendinitis AND/OR tenosynovitis of the elbow region
C0410039|T047|IS|239973006|SNOMEDCT_CORE|Tendinitis and tenosynovitis of the wrist and hand|Tendinitis AND/OR tenosynovitis of wrist AND/OR hand
C0410039|T047|OF|239973006|SNOMEDCT_CORE|Tendinitis and tenosynovitis of the wrist and hand|Tendinitis AND/OR tenosynovitis of wrist AND/OR hand
C0410039|T047|OF|239973006|SNOMEDCT_CORE|Tendinitis AND/OR tenosynovitis of the wrist AND/OR hand|Tendinitis AND/OR tenosynovitis of wrist AND/OR hand
C0410039|T047|OAS|239973006|SNOMEDCT_CORE|Tendinitis AND/OR tenosynovitis of the wrist AND/OR hand|Tendinitis AND/OR tenosynovitis of wrist AND/OR hand
C0410039|T047|OAF|239973006|SNOMEDCT_CORE|Tendinitis AND/OR tenosynovitis of wrist AND/OR hand|Tendinitis AND/OR tenosynovitis of wrist AND/OR hand
C0410039|T047|OAP|239973006|SNOMEDCT_CORE|Tendinitis AND/OR tenosynovitis of wrist AND/OR hand|Tendinitis AND/OR tenosynovitis of wrist AND/OR hand
C0410043|T047|PT|202912006|SNOMEDCT_CORE|Flexor tenosynovitis of finger|Flexor tenosynovitis of finger
C0410043|T047|FN|202912006|SNOMEDCT_CORE|Flexor tenosynovitis of finger|Flexor tenosynovitis of finger
C0410055|T046|SY|302936009|SNOMEDCT_CORE|Enthesopathy of wrist and hand|Enthesopathy of wrist and/or hand
C0410055|T046|OF|302936009|SNOMEDCT_CORE|Enthesopathy of wrist and hand|Enthesopathy of wrist and/or hand
C0410055|T046|PT|302936009|SNOMEDCT_CORE|Enthesopathy of wrist and/or hand|Enthesopathy of wrist and/or hand
C0410055|T046|FN|302936009|SNOMEDCT_CORE|Enthesopathy of wrist and/or hand|Enthesopathy of wrist and/or hand
C0410060|T020|SY|42786005|SNOMEDCT_CORE|Clicking thumb|Snapping thumb syndrome
C0410060|T020|SY|42786005|SNOMEDCT_CORE|Nodular tendinous disease of thumb|Snapping thumb syndrome
C0410060|T020|PT|42786005|SNOMEDCT_CORE|Snapping thumb syndrome|Snapping thumb syndrome
C0410060|T020|FN|42786005|SNOMEDCT_CORE|Snapping thumb syndrome|Snapping thumb syndrome
C0410060|T020|SY|42786005|SNOMEDCT_CORE|Trigger thumb|Snapping thumb syndrome
C0410060|T020|SY|42786005|SNOMEDCT_CORE|Trigger thumb - acquired|Snapping thumb syndrome
C0410060|T020|SY|42786005|SNOMEDCT_CORE|Triggering of thumb|Snapping thumb syndrome
C0410061|T019|PT|205274004|SNOMEDCT_CORE|Congenital trigger thumb|Congenital trigger thumb
C0410061|T019|FN|205274004|SNOMEDCT_CORE|Congenital trigger thumb|Congenital trigger thumb
C0410076|T047|PT|239993003|SNOMEDCT_CORE|Ischial bursitis|Ischial bursitis
C0410076|T047|FN|239993003|SNOMEDCT_CORE|Ischial bursitis|Ischial bursitis
C0410092|T047|PT|240004005|SNOMEDCT_CORE|Semimembranosus bursitis|Semimembranosus bursitis
C0410092|T047|FN|240004005|SNOMEDCT_CORE|Semimembranosus bursitis|Semimembranosus bursitis
C0410118|T047|PT|240027002|SNOMEDCT_CORE|Bursitis of foot region|Bursitis of foot region
C0410118|T047|FN|240027002|SNOMEDCT_CORE|Bursitis of foot region|Bursitis of foot region
C0410119|T047|PT|240028007|SNOMEDCT_CORE|Enthesopathy of foot region|Enthesopathy of foot region
C0410119|T047|FN|240028007|SNOMEDCT_CORE|Enthesopathy of foot region|Enthesopathy of foot region
C0410132|T037|PT|202888004|SNOMEDCT_CORE|Anterior shin splints|Anterior shin splints
C0410132|T037|FN|202888004|SNOMEDCT_CORE|Anterior shin splints|Anterior shin splints
C0410139|T047|PT|240036003|SNOMEDCT_CORE|Tenosynovitis of fingers|Tenosynovitis of fingers
C0410139|T047|FN|240036003|SNOMEDCT_CORE|Tenosynovitis of fingers|Tenosynovitis of fingers
C0410264|T190|SY|203076007|SNOMEDCT_CORE|Achilles tendon contracture|Contracture of Achilles tendon
C0410264|T190|PT|203076007|SNOMEDCT_CORE|Contracture of Achilles tendon|Contracture of Achilles tendon
C0410264|T190|FN|203076007|SNOMEDCT_CORE|Contracture of Achilles tendon|Contracture of Achilles tendon
C0410264|T190|OP|203076007|SNOMEDCT_CORE|Contracture of tendo achilles|Contracture of Achilles tendon
C0410264|T190|SY|203076007|SNOMEDCT_CORE|Contracture of tendo Achilles|Contracture of Achilles tendon
C0410264|T190|OF|203076007|SNOMEDCT_CORE|Contracture of tendo achilles|Contracture of Achilles tendon
C0410340|T037|PT|202332000|SNOMEDCT_CORE|Glenoid labrum tear|Glenoid labrum tear
C0410340|T037|FN|202332000|SNOMEDCT_CORE|Glenoid labrum tear|Glenoid labrum tear
C0410340|T037|SY|202332000|SNOMEDCT_CORE|Tear of glenoid labrum|Glenoid labrum tear
C0410480|T047|PT|203476003|SNOMEDCT_CORE|Avascular necrosis of the head of femur|Avascular necrosis of the head of femur
C0410480|T047|FN|203476003|SNOMEDCT_CORE|Avascular necrosis of the head of femur|Avascular necrosis of the head of femur
C0410549|T033|SY|240198002|SNOMEDCT_CORE|Collapse of vertebra due to osteoporosis|Osteoporotic vertebral collapse
C0410549|T033|PT|240198002|SNOMEDCT_CORE|Osteoporotic vertebral collapse|Osteoporotic vertebral collapse
C0410549|T033|FN|240198002|SNOMEDCT_CORE|Osteoporotic vertebral collapse|Osteoporotic vertebral collapse
C0410550|T047|PT|84138006|SNOMEDCT_CORE|Collapse of vertebra|Collapse of vertebra
C0410550|T047|FN|84138006|SNOMEDCT_CORE|Collapse of vertebra|Collapse of vertebra
C0410550|T047|IS|84138006|SNOMEDCT_CORE|Collapse of vertebra, NOS|Collapse of vertebra
C0410550|T047|SY|84138006|SNOMEDCT_CORE|Collapsed vertebra|Collapse of vertebra
C0410550|T047|SY|84138006|SNOMEDCT_CORE|Spondylomalacia|Collapse of vertebra
C0410601|T047|PT|202717005|SNOMEDCT_CORE|Cervical disc disorder with myelopathy|Cervical disc disorder with myelopathy
C0410601|T047|FN|202717005|SNOMEDCT_CORE|Cervical disc disorder with myelopathy|Cervical disc disorder with myelopathy
C0410619|T020|PT|240215009|SNOMEDCT_CORE|Prolapsed cervical intervertebral disc|Prolapsed cervical intervertebral disc
C0410619|T020|FN|240215009|SNOMEDCT_CORE|Prolapsed cervical intervertebral disc|Prolapsed cervical intervertebral disc
C0410629|T047|PT|202735001|SNOMEDCT_CORE|Lumbar disc prolapse with radiculopathy|Lumbar disc prolapse with radiculopathy
C0410629|T047|FN|202735001|SNOMEDCT_CORE|Lumbar disc prolapse with radiculopathy|Lumbar disc prolapse with radiculopathy
C0410629|T047|SY|202735001|SNOMEDCT_CORE|Lumbar disc prolapse with root compression|Lumbar disc prolapse with radiculopathy
C0410807|T033|SY|213082003|SNOMEDCT_CORE|Dislocation of joint prosthesis|Prosthetic joint dislocation
C0410807|T033|PT|213082003|SNOMEDCT_CORE|Prosthetic joint dislocation|Prosthetic joint dislocation
C0410807|T033|FN|213082003|SNOMEDCT_CORE|Prosthetic joint dislocation|Prosthetic joint dislocation
C0410808|T047|SY|213121005|SNOMEDCT_CORE|Infected arthroplasty|Prosthetic joint infection
C0410808|T047|SY|213121005|SNOMEDCT_CORE|Infected joint prosthesis|Prosthetic joint infection
C0410808|T047|PT|213121005|SNOMEDCT_CORE|Prosthetic joint infection|Prosthetic joint infection
C0410808|T047|FN|213121005|SNOMEDCT_CORE|Prosthetic joint infection|Prosthetic joint infection
C0410816|T184|PT|240271006|SNOMEDCT_CORE|Persistent prosthetic joint pain|Persistent prosthetic joint pain
C0410816|T184|FN|240271006|SNOMEDCT_CORE|Persistent prosthetic joint pain|Persistent prosthetic joint pain
C0410928|T033|IS|240301009|SNOMEDCT_CORE|Breast-feeding problem in the newborn|Breastfeeding problem in the newborn
C0410928|T033|OF|240301009|SNOMEDCT_CORE|Breast-feeding problem in the newborn|Breastfeeding problem in the newborn
C0410928|T033|PT|240301009|SNOMEDCT_CORE|Breastfeeding problem in the newborn|Breastfeeding problem in the newborn
C0410928|T033|FN|240301009|SNOMEDCT_CORE|Breastfeeding problem in the newborn|Breastfeeding problem in the newborn
C0410988|T047|PT|206439006|SNOMEDCT_CORE|Neonatal jaundice due to glucose-6-phosphate dehydrogenase deficiency|Neonatal jaundice due to glucose-6-phosphate dehydrogenase deficiency
C0410988|T047|FN|206439006|SNOMEDCT_CORE|Neonatal jaundice due to glucose-6-phosphate dehydrogenase deficiency|Neonatal jaundice due to glucose-6-phosphate dehydrogenase deficiency
C0410988|T047|SY|206439006|SNOMEDCT_CORE|Neonatal jaundice with glucose-6-phosphate dehydrogenase deficiency|Neonatal jaundice due to glucose-6-phosphate dehydrogenase deficiency
C0410988|T047|OF|206439006|SNOMEDCT_CORE|Neonatal jaundice with glucose-6-phosphate dehydrogenase deficiency|Neonatal jaundice due to glucose-6-phosphate dehydrogenase deficiency
C0411160|T046|PT|206037001|SNOMEDCT_CORE|Fetal or neonatal effect of maternal premature rupture of membrane|Fetal or neonatal effect of maternal premature rupture of membrane
C0411160|T046|FN|206037001|SNOMEDCT_CORE|Fetal or neonatal effect of maternal premature rupture of membrane|Fetal or neonatal effect of maternal premature rupture of membrane
C0411160|T046|OP|206037001|SNOMEDCT_CORE|Fetus or neonate affected by maternal premature rupture of membrane|Fetal or neonatal effect of maternal premature rupture of membrane
C0411160|T046|OF|206037001|SNOMEDCT_CORE|Fetus or neonate affected by maternal premature rupture of membrane|Fetal or neonatal effect of maternal premature rupture of membrane
C0411160|T046|IS|38511004|SNOMEDCT_CORE|Fetus or newborn affected by premature rupture of membranes|Fetal or neonatal effect of maternal premature rupture of membrane
C0411160|T046|OAP|38511004|SNOMEDCT_CORE|Fetus OR newborn affected by premature rupture of membranes|Fetal or neonatal effect of maternal premature rupture of membrane
C0411160|T046|OAF|38511004|SNOMEDCT_CORE|Fetus OR newborn affected by premature rupture of membranes|Fetal or neonatal effect of maternal premature rupture of membrane
C0411160|T046|SY|206037001|SNOMEDCT_CORE|Foetal or neonatal effect of maternal premature rupture of membrane|Fetal or neonatal effect of maternal premature rupture of membrane
C0411160|T046|OP|206037001|SNOMEDCT_CORE|Foetus or neonate affected by maternal premature rupture of membrane|Fetal or neonatal effect of maternal premature rupture of membrane
C0411161|T047|PT|206038006|SNOMEDCT_CORE|Fetal or neonatal effect of maternal oligohydramnios|Fetal or neonatal effect of maternal oligohydramnios
C0411161|T047|FN|206038006|SNOMEDCT_CORE|Fetal or neonatal effect of maternal oligohydramnios|Fetal or neonatal effect of maternal oligohydramnios
C0411161|T047|OAP|65599008|SNOMEDCT_CORE|Fetal or neonatal effect of oligohydramnios|Fetal or neonatal effect of maternal oligohydramnios
C0411161|T047|SY|206038006|SNOMEDCT_CORE|Fetal or neonatal effect of oligohydramnios|Fetal or neonatal effect of maternal oligohydramnios
C0411161|T047|OAF|65599008|SNOMEDCT_CORE|Fetal or neonatal effect of oligohydramnios|Fetal or neonatal effect of maternal oligohydramnios
C0411161|T047|OP|206038006|SNOMEDCT_CORE|Fetus or neonate affected by maternal oligohydramnios|Fetal or neonatal effect of maternal oligohydramnios
C0411161|T047|OF|206038006|SNOMEDCT_CORE|Fetus or neonate affected by maternal oligohydramnios|Fetal or neonatal effect of maternal oligohydramnios
C0411161|T047|SY|206038006|SNOMEDCT_CORE|Foetal or neonatal effect of maternal oligohydramnios|Fetal or neonatal effect of maternal oligohydramnios
C0411161|T047|SY|206038006|SNOMEDCT_CORE|Foetal or neonatal effect of oligohydramnios|Fetal or neonatal effect of maternal oligohydramnios
C0411162|T047|IS|268798004|SNOMEDCT_CORE|Fetus affected by hydramnios|Fetus affected by hydramnios
C0411162|T047|OP|268798004|SNOMEDCT_CORE|Fetus or neonate affected by maternal polyhydramnios|Fetus affected by hydramnios
C0411162|T047|OF|268798004|SNOMEDCT_CORE|Fetus or neonate affected by maternal polyhydramnios|Fetus affected by hydramnios
C0411169|T046|OP|206046007|SNOMEDCT_CORE|Fetus or neonate affected by multiple pregnancy|Fetus or neonate affected by multiple pregnancy
C0411169|T046|OF|206046007|SNOMEDCT_CORE|Fetus or neonate affected by multiple pregnancy|Fetus or neonate affected by multiple pregnancy
C0411169|T046|OP|18001006|SNOMEDCT_CORE|Fetus OR newborn affected by multiple pregnancy|Fetus or neonate affected by multiple pregnancy
C0411169|T046|OF|18001006|SNOMEDCT_CORE|Fetus OR newborn affected by multiple pregnancy|Fetus or neonate affected by multiple pregnancy
C0411169|T046|IS|18001006|SNOMEDCT_CORE|Fetus or newborn affected by multiple pregnancy, NOS|Fetus or neonate affected by multiple pregnancy
C0411169|T046|IS|18001006|SNOMEDCT_CORE|Foetus or newborn affected by multiple pregnancy, NOS|Fetus or neonate affected by multiple pregnancy
C0411175|T047|PT|206002004|SNOMEDCT_CORE|Fetal or neonatal effect of maternal medical problem|Fetal or neonatal effect of maternal medical problem
C0411175|T047|FN|206002004|SNOMEDCT_CORE|Fetal or neonatal effect of maternal medical problem|Fetal or neonatal effect of maternal medical problem
C0411175|T047|OP|206002004|SNOMEDCT_CORE|Fetus or neonate affected by maternal medical problem|Fetal or neonatal effect of maternal medical problem
C0411175|T047|OF|206002004|SNOMEDCT_CORE|Fetus or neonate affected by maternal medical problem|Fetal or neonatal effect of maternal medical problem
C0411175|T047|IS|206002004|SNOMEDCT_CORE|Fetus or neonate affected by maternal medical problems|Fetal or neonatal effect of maternal medical problem
C0411175|T047|OF|206002004|SNOMEDCT_CORE|Fetus or neonate affected by maternal medical problems|Fetal or neonatal effect of maternal medical problem
C0411175|T047|IS|206002004|SNOMEDCT_CORE|Fetus OR newborn affected by maternal condition|Fetal or neonatal effect of maternal medical problem
C0411175|T047|SY|206002004|SNOMEDCT_CORE|Foetal or neonatal effect of maternal medical problem|Fetal or neonatal effect of maternal medical problem
C0411178|T046|PT|206005002|SNOMEDCT_CORE|Fetal or neonatal effect of maternal infection|Fetal or neonatal effect of maternal infection
C0411178|T046|FN|206005002|SNOMEDCT_CORE|Fetal or neonatal effect of maternal infection|Fetal or neonatal effect of maternal infection
C0411178|T046|SY|206005002|SNOMEDCT_CORE|Fetal or neonatal effect of maternal infectious disease|Fetal or neonatal effect of maternal infection
C0411178|T046|OP|206005002|SNOMEDCT_CORE|Fetus or neonate affected by maternal infection|Fetal or neonatal effect of maternal infection
C0411178|T046|OF|206005002|SNOMEDCT_CORE|Fetus or neonate affected by maternal infection|Fetal or neonatal effect of maternal infection
C0411178|T046|IS|206005002|SNOMEDCT_CORE|Fetus or neonate affected by maternal infections|Fetal or neonatal effect of maternal infection
C0411178|T046|OF|206005002|SNOMEDCT_CORE|Fetus or neonate affected by maternal infections|Fetal or neonatal effect of maternal infection
C0411178|T046|IS|206005002|SNOMEDCT_CORE|Fetus OR newborn affected by maternal infection|Fetal or neonatal effect of maternal infection
C0411178|T046|IS|206005002|SNOMEDCT_CORE|Fetus OR newborn affected by maternal infectious disease|Fetal or neonatal effect of maternal infection
C0411178|T046|SY|206005002|SNOMEDCT_CORE|Foetal or neonatal effect of maternal infection|Fetal or neonatal effect of maternal infection
C0411178|T046|SY|206005002|SNOMEDCT_CORE|Foetal or neonatal effect of maternal infectious disease|Fetal or neonatal effect of maternal infection
C0412849|T037|PT|241748001|SNOMEDCT_CORE|Poisoning by analgesic drug|Poisoning by analgesic drug
C0412849|T037|OF|241748001|SNOMEDCT_CORE|Poisoning by analgesic drug|Poisoning by analgesic drug
C0412849|T037|SY|241748001|SNOMEDCT_CORE|Poisoning caused by analgesic drug|Poisoning by analgesic drug
C0412849|T037|FN|241748001|SNOMEDCT_CORE|Poisoning caused by analgesic drug|Poisoning by analgesic drug
C0412877|T037|SY|56951005|SNOMEDCT_CORE|Poisoning by cardiac glycoside|Poisoning by cardiotonic glycoside
C0412877|T037|PT|56951005|SNOMEDCT_CORE|Poisoning by cardiotonic glycoside|Poisoning by cardiotonic glycoside
C0412877|T037|OF|56951005|SNOMEDCT_CORE|Poisoning by cardiotonic glycoside|Poisoning by cardiotonic glycoside
C0412877|T037|IS|56951005|SNOMEDCT_CORE|Poisoning by cardiotonic glycoside, NOS|Poisoning by cardiotonic glycoside
C0412877|T037|SY|56951005|SNOMEDCT_CORE|Poisoning caused by cardiac glycoside|Poisoning by cardiotonic glycoside
C0412877|T037|SY|56951005|SNOMEDCT_CORE|Poisoning caused by cardiotonic glycoside|Poisoning by cardiotonic glycoside
C0412877|T037|FN|56951005|SNOMEDCT_CORE|Poisoning caused by cardiotonic glycoside|Poisoning by cardiotonic glycoside
C0413120|T037|PT|241820008|SNOMEDCT_CORE|Bee sting|Bee sting
C0413120|T037|FN|241820008|SNOMEDCT_CORE|Bee sting|Bee sting
C0413671|T046|SY|293331003|SNOMEDCT_CORE|Adverse reaction to anticoagulants|Anticoagulant adverse reaction
C0413671|T046|PT|293331003|SNOMEDCT_CORE|Anticoagulant adverse reaction|Anticoagulant adverse reaction
C0413671|T046|FN|293331003|SNOMEDCT_CORE|Anticoagulant adverse reaction|Anticoagulant adverse reaction
C0414592|T037|PT|214206004|SNOMEDCT_CORE|Motor vehicle on road in collision with pedestrian|Motor vehicle on road in collision with pedestrian
C0414592|T037|OF|214206004|SNOMEDCT_CORE|Motor vehicle on road in collision with pedestrian|Motor vehicle on road in collision with pedestrian
C0414592|T037|FN|214206004|SNOMEDCT_CORE|Motor vehicle on road in collision with pedestrian|Motor vehicle on road in collision with pedestrian
C0416591|T037|OAP|433086005|SNOMEDCT_CORE|Accidental poisoning by aromatic analgesic|Accidental poisoning caused by aromatic analgesic
C0416591|T037|OF|433086005|SNOMEDCT_CORE|Accidental poisoning by aromatic analgesic|Accidental poisoning caused by aromatic analgesic
C0416591|T037|OAS|433086005|SNOMEDCT_CORE|Accidental poisoning caused by aromatic analgesic|Accidental poisoning caused by aromatic analgesic
C0416591|T037|OAF|433086005|SNOMEDCT_CORE|Accidental poisoning caused by aromatic analgesic|Accidental poisoning caused by aromatic analgesic
C0416892|T037|PT|242374007|SNOMEDCT_CORE|Accidental exposure to metallic lead|Accidental exposure to metallic lead
C0416892|T037|OF|242374007|SNOMEDCT_CORE|Accidental exposure to metallic lead|Accidental exposure to metallic lead
C0416892|T037|FN|242374007|SNOMEDCT_CORE|Accidental exposure to metallic lead|Accidental exposure to metallic lead
C0416987|T037|PT|217155007|SNOMEDCT_CORE|Fall on same level from slipping|Fall on same level from slipping
C0416987|T037|OF|217155007|SNOMEDCT_CORE|Fall on same level from slipping|Fall on same level from slipping
C0416987|T037|FN|217155007|SNOMEDCT_CORE|Fall on same level from slipping|Fall on same level from slipping
C0416999|T037|PT|217157004|SNOMEDCT_CORE|Fall on same level from stumbling|Fall on same level from stumbling
C0416999|T037|OF|217157004|SNOMEDCT_CORE|Fall on same level from stumbling|Fall on same level from stumbling
C0416999|T037|FN|217157004|SNOMEDCT_CORE|Fall on same level from stumbling|Fall on same level from stumbling
C0417006|T037|PT|274919008|SNOMEDCT_CORE|Fall on same level due to impact against another person|Fall on same level due to impact against another person
C0417006|T037|OF|274919008|SNOMEDCT_CORE|Fall on same level due to impact against another person|Fall on same level due to impact against another person
C0417006|T037|FN|274919008|SNOMEDCT_CORE|Fall on same level due to impact against another person|Fall on same level due to impact against another person
C0417023|T037|SY|217094006|SNOMEDCT_CORE|Fall down steps|Fall from steps
C0417023|T037|PT|217094006|SNOMEDCT_CORE|Fall from steps|Fall from steps
C0417023|T037|OF|217094006|SNOMEDCT_CORE|Fall from steps|Fall from steps
C0417023|T037|FN|217094006|SNOMEDCT_CORE|Fall from steps|Fall from steps
C0417024|T037|PT|242408008|SNOMEDCT_CORE|Fall from one level to another|Fall from one level to another
C0417024|T037|OF|242408008|SNOMEDCT_CORE|Fall from one level to another|Fall from one level to another
C0417024|T037|FN|242408008|SNOMEDCT_CORE|Fall from one level to another|Fall from one level to another
C0417508|T037|PT|242489002|SNOMEDCT_CORE|Accident due to contact with hot or corrosive substance|Accident due to contact with hot or corrosive substance
C0417508|T037|OF|242489002|SNOMEDCT_CORE|Accident due to contact with hot or corrosive substance|Accident due to contact with hot or corrosive substance
C0417508|T037|FN|242489002|SNOMEDCT_CORE|Accident due to contact with hot or corrosive substance|Accident due to contact with hot or corrosive substance
C0417950|T037|SY|269716005|SNOMEDCT_CORE|Industrial machinery accident|Industrial machinery accident
C0418294|T037|PT|242840004|SNOMEDCT_CORE|Self poisoning by carbon monoxide|Self poisoning by carbon monoxide
C0418294|T037|OF|242840004|SNOMEDCT_CORE|Self poisoning by carbon monoxide|Self poisoning by carbon monoxide
C0418294|T037|SY|242840004|SNOMEDCT_CORE|Self poisoning caused by carbon monoxide|Self poisoning by carbon monoxide
C0418294|T037|FN|242840004|SNOMEDCT_CORE|Self poisoning caused by carbon monoxide|Self poisoning by carbon monoxide
C0418384|T037|PT|219218005|SNOMEDCT_CORE|Assault by cutting and stabbing instruments|Assault by cutting and stabbing instruments
C0418384|T037|OF|219218005|SNOMEDCT_CORE|Assault by cutting and stabbing instruments|Assault by cutting and stabbing instruments
C0418384|T037|FN|219218005|SNOMEDCT_CORE|Assault by cutting and stabbing instruments|Assault by cutting and stabbing instruments
C0418570|T037|PT|219346009|SNOMEDCT_CORE|Injury of unknown intent due to fall from height|Injury of unknown intent due to fall from height
C0418570|T037|OF|219346009|SNOMEDCT_CORE|Injury of unknown intent due to fall from height|Injury of unknown intent due to fall from height
C0418570|T037|FN|219346009|SNOMEDCT_CORE|Injury of unknown intent due to fall from height|Injury of unknown intent due to fall from height
C0419373|T033|PT|281050002|SNOMEDCT_CORE|Livebirth|Livebirth
C0419373|T033|FN|281050002|SNOMEDCT_CORE|Livebirth|Livebirth
C0419530|T033|PT|268464009|SNOMEDCT_CORE|Contraception using injectable contraceptive medication|Contraception using injectable contraceptive medication
C0419530|T033|SY|268464009|SNOMEDCT_CORE|Depot contraception|Contraception using injectable contraceptive medication
C0419530|T033|FN|268464009|SNOMEDCT_CORE|Depot contraception|Contraception using injectable contraceptive medication
C0419530|T033|SY|268464009|SNOMEDCT_CORE|Depot contraceptive|Contraception using injectable contraceptive medication
C0419551|T033|PT|169582001|SNOMEDCT_CORE|A/N care: H/O stillbirth|A/N care: H/O stillbirth
C0419551|T033|OF|169582001|SNOMEDCT_CORE|Antenatal care: H/O stillbirth|A/N care: H/O stillbirth
C0419551|T033|FN|169582001|SNOMEDCT_CORE|Antenatal care: history of stillbirth|A/N care: H/O stillbirth
C0419551|T033|SY|169582001|SNOMEDCT_CORE|Antenatal care: history of stillbirth|A/N care: H/O stillbirth
C0419552|T033|PT|169583006|SNOMEDCT_CORE|A/N care: H/O perinatal death|A/N care: H/O perinatal death
C0419552|T033|OF|169583006|SNOMEDCT_CORE|Antenatal care: H/O perinatal death|A/N care: H/O perinatal death
C0419552|T033|FN|169583006|SNOMEDCT_CORE|Antenatal care: history of perinatal death|A/N care: H/O perinatal death
C0419552|T033|SY|169583006|SNOMEDCT_CORE|Antenatal care: history of perinatal death|A/N care: H/O perinatal death
C0419553|T033|PT|169584000|SNOMEDCT_CORE|A/N care: poor obstetric history|A/N care: poor obstetric history
C0419553|T033|OF|169584000|SNOMEDCT_CORE|Antenatal care: poor obstetric history|A/N care: poor obstetric history
C0419553|T033|FN|169584000|SNOMEDCT_CORE|Antenatal care: poor obstetric history|A/N care: poor obstetric history
C0419553|T033|SY|169584000|SNOMEDCT_CORE|Antenatal care: poor obstetric history|A/N care: poor obstetric history
C0420948|T033|SY|169665005|SNOMEDCT_CORE|A/N U/S scan abnormal|Antenatal ultrasound scan abnormal
C0420948|T033|SY|169665005|SNOMEDCT_CORE|Abnormal ultrasonic finding on antenatal screening of mother|Antenatal ultrasound scan abnormal
C0420948|T033|PT|169665005|SNOMEDCT_CORE|Antenatal ultrasound scan abnormal|Antenatal ultrasound scan abnormal
C0420948|T033|FN|169665005|SNOMEDCT_CORE|Antenatal ultrasound scan abnormal|Antenatal ultrasound scan abnormal
C0420968|T033|PT|169696001|SNOMEDCT_CORE|Rubella status not known|Rubella status not known
C0420968|T033|FN|169696001|SNOMEDCT_CORE|Rubella status not known|Rubella status not known
C0421373|T033|PTGB|171259000|SNOMEDCT_CORE|Not up to date with immunisations|Not up to date with immunizations
C0421373|T033|PT|171259000|SNOMEDCT_CORE|Not up to date with immunizations|Not up to date with immunizations
C0421373|T033|FN|171259000|SNOMEDCT_CORE|Not up to date with immunizations|Not up to date with immunizations
C0421373|T033|IS|171259000|SNOMEDCT_CORE|Not up-to-date with immunisation|Not up to date with immunizations
C0421373|T033|OP|171259000|SNOMEDCT_CORE|Not up-to-date with immunisations|Not up to date with immunizations
C0421373|T033|IS|171259000|SNOMEDCT_CORE|Not up-to-date with immunization|Not up to date with immunizations
C0421373|T033|OF|171259000|SNOMEDCT_CORE|Not up-to-date with immunization|Not up to date with immunizations
C0421373|T033|OP|171259000|SNOMEDCT_CORE|Not up-to-date with immunizations|Not up to date with immunizations
C0421373|T033|OF|171259000|SNOMEDCT_CORE|Not up-to-date with immunizations|Not up to date with immunizations
C0421565|T033|PT|184238003|SNOMEDCT_CORE|Repeat prescription card duplicate issue|Repeat prescription card duplicate issue
C0421565|T033|FN|184238003|SNOMEDCT_CORE|Repeat prescription card duplicate issue|Repeat prescription card duplicate issue
C0422987|T033|PT|246656009|SNOMEDCT_CORE|Loss of part of visual field|Loss of part of visual field
C0422987|T033|FN|246656009|SNOMEDCT_CORE|Loss of part of visual field|Loss of part of visual field
C0423004|T184|OAP|246676003|SNOMEDCT_CORE|Hyperaemia of surface of eye|Hyperaemia of surface of eye
C0423004|T184|OAP|246676003|SNOMEDCT_CORE|Hyperemia of surface of eye|Hyperaemia of surface of eye
C0423004|T184|OAS|246676003|SNOMEDCT_CORE|Injection of surface of eye|Hyperaemia of surface of eye
C0423004|T184|OAF|246676003|SNOMEDCT_CORE|Injection of surface of eye|Hyperaemia of surface of eye
C0423062|T047|SY|63988001|SNOMEDCT_CORE|Intermittent comitant exotropia|Intermittent exotropia
C0423062|T047|SY|63988001|SNOMEDCT_CORE|Intermittent divergent squint|Intermittent exotropia
C0423062|T047|PT|63988001|SNOMEDCT_CORE|Intermittent exotropia|Intermittent exotropia
C0423062|T047|FN|63988001|SNOMEDCT_CORE|Intermittent exotropia|Intermittent exotropia
C0423062|T047|IS|63988001|SNOMEDCT_CORE|Intermittent exotropia, NOS|Intermittent exotropia
C0423062|T047|SY|63988001|SNOMEDCT_CORE|X - Intermittent exotropia|Intermittent exotropia
C0423086|T047|SY|103262002|SNOMEDCT_CORE|Gazing fixedly|Staring
C0423086|T047|PT|103262002|SNOMEDCT_CORE|Staring|Staring
C0423086|T047|FN|103262002|SNOMEDCT_CORE|Staring|Staring
C0423122|T047|SY|246813002|SNOMEDCT_CORE|Brow ptosis|Ptosis of eyebrow
C0423122|T047|IS|246813002|SNOMEDCT_CORE|Eyebow ptosis|Ptosis of eyebrow
C0423122|T047|SY|246813002|SNOMEDCT_CORE|Eyebrow ptosis|Ptosis of eyebrow
C0423122|T047|SY|246813002|SNOMEDCT_CORE|Ptosis brow|Ptosis of eyebrow
C0423122|T047|PT|246813002|SNOMEDCT_CORE|Ptosis of eyebrow|Ptosis of eyebrow
C0423122|T047|FN|246813002|SNOMEDCT_CORE|Ptosis of eyebrow|Ptosis of eyebrow
C0423124|T033|SY|246815009|SNOMEDCT_CORE|Dermatochalasis|Excess skin of eyelid
C0423124|T033|PT|246815009|SNOMEDCT_CORE|Excess skin of eyelid|Excess skin of eyelid
C0423124|T033|FN|246815009|SNOMEDCT_CORE|Excess skin of eyelid|Excess skin of eyelid
C0423361|T047|PT|247081001|SNOMEDCT_CORE|Posterior vitreous detachment|Posterior vitreous detachment
C0423361|T047|FN|247081001|SNOMEDCT_CORE|Posterior vitreous detachment|Posterior vitreous detachment
C0423361|T047|SY|247081001|SNOMEDCT_CORE|PVD - Posterior vitreous detachment|Posterior vitreous detachment
C0423422|T033|PT|247146001|SNOMEDCT_CORE|Macular pigment deposit|Macular pigment deposit
C0423422|T033|OF|247146001|SNOMEDCT_CORE|Macular pigment deposit|Macular pigment deposit
C0423422|T033|FN|247146001|SNOMEDCT_CORE|Macular pigment deposit|Macular pigment deposit
C0423428|T020|SY|18410006|SNOMEDCT_CORE|Macular scar|Scarred macula
C0423428|T020|PT|18410006|SNOMEDCT_CORE|Scarred macula|Scarred macula
C0423428|T020|FN|18410006|SNOMEDCT_CORE|Scarred macula|Scarred macula
C0423433|T033|OAS|23911001|SNOMEDCT_CORE|CNV-Choroidal neovascularisation|Subretinal neovascularization
C0423433|T033|OAS|23911001|SNOMEDCT_CORE|CNV-Choroidal neovascularization|Subretinal neovascularization
C0423433|T033|OAS|23911001|SNOMEDCT_CORE|NVM - Subretinal neovascular membrane|Subretinal neovascularization
C0423433|T033|OAS|23911001|SNOMEDCT_CORE|Presumed subretinal neovascular membrane|Subretinal neovascularization
C0423433|T033|OAS|23911001|SNOMEDCT_CORE|SRNV-Subretinal neovascularisation|Subretinal neovascularization
C0423433|T033|OAS|23911001|SNOMEDCT_CORE|SRNV-Subretinal neovascularization|Subretinal neovascularization
C0423433|T033|OAS|23911001|SNOMEDCT_CORE|Subretinal neovascular membrane|Subretinal neovascularization
C0423433|T033|OAP|23911001|SNOMEDCT_CORE|Subretinal neovascularisation|Subretinal neovascularization
C0423433|T033|OAP|23911001|SNOMEDCT_CORE|Subretinal neovascularization|Subretinal neovascularization
C0423433|T033|OF|23911001|SNOMEDCT_CORE|Subretinal neovascularization|Subretinal neovascularization
C0423433|T033|OAF|23911001|SNOMEDCT_CORE|Subretinal neovascularization|Subretinal neovascularization
C0423572|T184|PT|62507009|SNOMEDCT_CORE|Pins and needles|Pins and needles
C0423572|T184|FN|62507009|SNOMEDCT_CORE|Pins and needles|Pins and needles
C0423572|T184|SY|62507009|SNOMEDCT_CORE|Pins and needles sensation|Pins and needles
C0423610|T184|SY|162143008|SNOMEDCT_CORE|Female genital pain|Pain in female genitalia
C0423610|T184|PT|162143008|SNOMEDCT_CORE|Pain in female genitalia|Pain in female genitalia
C0423610|T184|FN|162143008|SNOMEDCT_CORE|Pain in female genitalia|Pain in female genitalia
C0423632|T184|SY|2237002|SNOMEDCT_CORE|Painful breathing -pleurodynia|Painful breathing -pleurodynia
C0423658|T184|SY|267954009|SNOMEDCT_CORE|Ankle and/or foot joint pain|Arthralgia of the ankle and/or foot
C0423658|T184|SY|267954009|SNOMEDCT_CORE|Arthralgia of the ankle and foot|Arthralgia of the ankle and/or foot
C0423658|T184|OF|267954009|SNOMEDCT_CORE|Arthralgia of the ankle and foot|Arthralgia of the ankle and/or foot
C0423658|T184|PT|267954009|SNOMEDCT_CORE|Arthralgia of the ankle and/or foot|Arthralgia of the ankle and/or foot
C0423658|T184|FN|267954009|SNOMEDCT_CORE|Arthralgia of the ankle and/or foot|Arthralgia of the ankle and/or foot
C0423661|T184|OAP|267953003|SNOMEDCT_CORE|Arthralgia of the lower leg|Arthralgia of the lower leg
C0423661|T184|OAF|267953003|SNOMEDCT_CORE|Arthralgia of the lower leg|Arthralgia of the lower leg
C0423663|T184|PT|267952008|SNOMEDCT_CORE|Arthralgia of the pelvic region and thigh|Arthralgia of the pelvic region and thigh
C0423663|T184|FN|267952008|SNOMEDCT_CORE|Arthralgia of the pelvic region and thigh|Arthralgia of the pelvic region and thigh
C0423665|T184|SY|202472008|SNOMEDCT_CORE|Arthralgia of the hand|Hand joint pain
C0423665|T184|PT|202472008|SNOMEDCT_CORE|Hand joint pain|Hand joint pain
C0423665|T184|FN|202472008|SNOMEDCT_CORE|Hand joint pain|Hand joint pain
C0423668|T184|PT|267950000|SNOMEDCT_CORE|Arthralgia of the upper arm|Arthralgia of the upper arm
C0423668|T184|FN|267950000|SNOMEDCT_CORE|Arthralgia of the upper arm|Arthralgia of the upper arm
C0423669|T184|SY|202480001|SNOMEDCT_CORE|Arthralgia of elbow|Elbow joint pain
C0423669|T184|PT|202480001|SNOMEDCT_CORE|Elbow joint pain|Elbow joint pain
C0423669|T184|FN|202480001|SNOMEDCT_CORE|Elbow joint pain|Elbow joint pain
C0423670|T184|SY|267949000|SNOMEDCT_CORE|Arthralgia of shoulder|Shoulder joint pain
C0423670|T184|SY|267949000|SNOMEDCT_CORE|Arthralgia of the shoulder region|Shoulder joint pain
C0423670|T184|PT|267949000|SNOMEDCT_CORE|Shoulder joint pain|Shoulder joint pain
C0423670|T184|FN|267949000|SNOMEDCT_CORE|Shoulder joint pain|Shoulder joint pain
C0423674|T184|PT|279029001|SNOMEDCT_CORE|Pain in cervical spine|Pain in cervical spine
C0423674|T184|FN|279029001|SNOMEDCT_CORE|Pain in cervical spine|Pain in cervical spine
C0423675|T047|PT|202796002|SNOMEDCT_CORE|Thoracic and lumbosacral neuritis|Thoracic and lumbosacral neuritis
C0423675|T047|FN|202796002|SNOMEDCT_CORE|Thoracic and lumbosacral neuritis|Thoracic and lumbosacral neuritis
C0423676|T047|PT|62195001|SNOMEDCT_CORE|Lumbosacral neuritis|Lumbosacral neuritis
C0423676|T047|FN|62195001|SNOMEDCT_CORE|Lumbosacral neuritis|Lumbosacral neuritis
C0423676|T047|IS|62195001|SNOMEDCT_CORE|Lumbosacral neuritis, NOS|Lumbosacral neuritis
C0423682|T047|PT|279040009|SNOMEDCT_CORE|Mechanical low back pain|Mechanical low back pain
C0423682|T047|FN|279040009|SNOMEDCT_CORE|Mechanical low back pain|Mechanical low back pain
C0423682|T047|OF|279040009|SNOMEDCT_CORE|Mechanical low back pain|Mechanical low back pain
C0423684|T033|PT|279038004|SNOMEDCT_CORE|Thoracic back pain|Thoracic back pain
C0423684|T033|FN|279038004|SNOMEDCT_CORE|Thoracic back pain|Thoracic back pain
C0423684|T033|OF|279038004|SNOMEDCT_CORE|Thoracic back pain|Thoracic back pain
C0423690|T047|PT|247369005|SNOMEDCT_CORE|Facet joint pain|Facet joint pain
C0423690|T047|FN|247369005|SNOMEDCT_CORE|Facet joint pain|Facet joint pain
C0423690|T047|SY|247369005|SNOMEDCT_CORE|Facet joint syndrome|Facet joint pain
C0423736|T184|IS|58250006|SNOMEDCT_CORE|Burning on urination|Scalding pain on urination
C0423736|T184|SY|58250006|SNOMEDCT_CORE|Burning pain on urination|Scalding pain on urination
C0423736|T184|PT|58250006|SNOMEDCT_CORE|Scalding pain on urination|Scalding pain on urination
C0423736|T184|FN|58250006|SNOMEDCT_CORE|Scalding pain on urination|Scalding pain on urination
C0423775|T047|IS|200767005|SNOMEDCT_CORE|Dandruff|Pityriasis simplex
C0423775|T047|IS|200767005|SNOMEDCT_CORE|Furfuracea|Pityriasis simplex
C0423775|T047|OF|200767005|SNOMEDCT_CORE|Pityriasis simplex|Pityriasis simplex
C0423775|T047|PT|200767005|SNOMEDCT_CORE|Pityriasis simplex|Pityriasis simplex
C0423775|T047|FN|200767005|SNOMEDCT_CORE|Pityriasis simplex|Pityriasis simplex
C0423791|T033|PT|247471006|SNOMEDCT_CORE|Maculopapular eruption|Maculopapular eruption
C0423791|T033|FN|247471006|SNOMEDCT_CORE|Maculopapular eruption|Maculopapular eruption
C0423791|T033|SY|247471006|SNOMEDCT_CORE|Maculopapular exanthema|Maculopapular eruption
C0423791|T033|SY|247471006|SNOMEDCT_CORE|Maculopapular rash|Maculopapular eruption
C0423798|T033|PT|424131007|SNOMEDCT_CORE|Easy bruising|Easy bruising
C0423798|T033|FN|424131007|SNOMEDCT_CORE|Easy bruising|Easy bruising
C0423798|T033|SY|424131007|SNOMEDCT_CORE|Increased tendency to bruise|Easy bruising
C0423927|T048|PT|192071009|SNOMEDCT_CORE|Mild memory disturbance|Mild memory disturbance
C0423927|T048|FN|192071009|SNOMEDCT_CORE|Mild memory disturbance|Mild memory disturbance
C0424000|T033|FN|225457007|SNOMEDCT_CORE|Feeling suicidal|Suicidal thoughts
C0424000|T033|PT|225457007|SNOMEDCT_CORE|Feeling suicidal|Suicidal thoughts
C0424000|T033|SY|6471006|SNOMEDCT_CORE|Suicidal ideation|Suicidal thoughts
C0424000|T033|PT|6471006|SNOMEDCT_CORE|Suicidal thoughts|Suicidal thoughts
C0424000|T033|FN|6471006|SNOMEDCT_CORE|Suicidal thoughts|Suicidal thoughts
C0424101|T048|SY|22058002|SNOMEDCT_CORE|General inattentiveness|Inattention
C0424101|T048|PT|22058002|SNOMEDCT_CORE|Inattention|Inattention
C0424101|T048|FN|22058002|SNOMEDCT_CORE|Inattention|Inattention
C0424295|T048|SY|44548000|SNOMEDCT_CORE|HA - Hyperactivity|Hyperactive behavior
C0424295|T048|PT|44548000|SNOMEDCT_CORE|Hyperactive behavior|Hyperactive behavior
C0424295|T048|FN|44548000|SNOMEDCT_CORE|Hyperactive behavior|Hyperactive behavior
C0424295|T048|PTGB|44548000|SNOMEDCT_CORE|Hyperactive behaviour|Hyperactive behavior
C0424295|T048|IS|44548000|SNOMEDCT_CORE|Hyperactivity|Hyperactive behavior
C0424295|T048|IS|44548000|SNOMEDCT_CORE|Hyperactivity, NOS|Hyperactive behavior
C0424295|T048|SY|44548000|SNOMEDCT_CORE|Hyperkinesis|Hyperactive behavior
C0424295|T048|SY|44548000|SNOMEDCT_CORE|Increased purposeful goal-directed activity|Hyperactive behavior
C0424295|T048|IS|44548000|SNOMEDCT_CORE|Increased purposeful goal-directed activity, NOS|Hyperactive behavior
C0424366|T033|OAS|248061004|SNOMEDCT_CORE|Self-damage|Self-harm
C0424366|T033|OAP|248061004|SNOMEDCT_CORE|Self-harm|Self-harm
C0424366|T033|OAF|248061004|SNOMEDCT_CORE|Self-harm|Self-harm
C0424531|T033|SY|248228001|SNOMEDCT_CORE|Bad turn|Funny turn
C0424531|T033|SY|248228001|SNOMEDCT_CORE|Funny spell|Funny turn
C0424531|T033|FN|248228001|SNOMEDCT_CORE|Funny turn|Funny turn
C0424531|T033|PT|248228001|SNOMEDCT_CORE|Funny turn|Funny turn
C0424593|T033|PT|248278004|SNOMEDCT_CORE|Attacks of weakness|Attacks of weakness
C0424593|T033|FN|248278004|SNOMEDCT_CORE|Attacks of weakness|Attacks of weakness
C0424605|T048|FN|248290002|SNOMEDCT_CORE|Developmental delay|Developmental delay
C0424605|T048|PT|248290002|SNOMEDCT_CORE|Developmental delay|Developmental delay
C0424641|T033|PT|71781005|SNOMEDCT_CORE|Decrease in height|Decrease in height
C0424641|T033|FN|71781005|SNOMEDCT_CORE|Decrease in height|Decrease in height
C0424671|T033|SY|162864005|SNOMEDCT_CORE|BMI 30+ - obesity|Body mass index 30+ - obesity
C0424671|T033|PT|162864005|SNOMEDCT_CORE|Body mass index 30+ - obesity|Body mass index 30+ - obesity
C0424671|T033|FN|162864005|SNOMEDCT_CORE|Body mass index 30+ - obesity|Body mass index 30+ - obesity
C0424672|T033|SY|162863004|SNOMEDCT_CORE|BMI 25-29 - overweight|Body mass index 25-29 - overweight
C0424672|T033|PT|162863004|SNOMEDCT_CORE|Body mass index 25-29 - overweight|Body mass index 25-29 - overweight
C0424672|T033|FN|162863004|SNOMEDCT_CORE|Body mass index 25-29 - overweight|Body mass index 25-29 - overweight
C0424672|T033|IS|162863004|SNOMEDCT_CORE|Body mass index index 25-29 - overweight|Body mass index 25-29 - overweight
C0424672|T033|OF|162863004|SNOMEDCT_CORE|Body mass index index 25-29 - overweight|Body mass index 25-29 - overweight
C0424802|T033|IS|67162002|SNOMEDCT_CORE|Ammoniacal body odor|Smells of urine
C0424802|T033|PT|67162002|SNOMEDCT_CORE|Smells of urine|Smells of urine
C0424802|T033|FN|67162002|SNOMEDCT_CORE|Smells of urine|Smells of urine
C0424802|T033|SY|67162002|SNOMEDCT_CORE|Urinary body odor|Smells of urine
C0424802|T033|SYGB|67162002|SNOMEDCT_CORE|Urinary body odour|Smells of urine
C0424853|T184|PT|248521008|SNOMEDCT_CORE|Lump on finger|Lump on finger
C0424853|T184|FN|248521008|SNOMEDCT_CORE|Lump on finger|Lump on finger
C0424853|T184|SY|248521008|SNOMEDCT_CORE|Mass of finger|Lump on finger
C0424939|T033|SY|161129001|SNOMEDCT_CORE|LD - Learning difficulties|Learning difficulties
C0424939|T033|PT|161129001|SNOMEDCT_CORE|Learning difficulties|Learning difficulties
C0424939|T033|FN|161129001|SNOMEDCT_CORE|Learning difficulties|Learning difficulties
C0424960|T033|PT|248539004|SNOMEDCT_CORE|Family problems|Family problems
C0424960|T033|FN|248539004|SNOMEDCT_CORE|Family problems|Family problems
C0424961|T033|OAP|248540002|SNOMEDCT_CORE|Constantly crying baby|Constantly crying baby
C0424961|T033|OAF|248540002|SNOMEDCT_CORE|Constantly crying baby|Constantly crying baby
C0424964|T033|PT|270472006|SNOMEDCT_CORE|Maternal concern|Maternal concern
C0424964|T033|FN|270472006|SNOMEDCT_CORE|Maternal concern|Maternal concern
C0425043|T033|IS|398033008|SNOMEDCT_CORE|Death in family, NOS|Death of relative
C0425043|T033|SY|398033008|SNOMEDCT_CORE|Death of family member|Death of relative
C0425043|T033|PT|398033008|SNOMEDCT_CORE|Death of relative|Death of relative
C0425043|T033|FN|398033008|SNOMEDCT_CORE|Death of relative|Death of relative
C0425043|T033|SY|398033008|SNOMEDCT_CORE|Family members dead|Death of relative
C0425043|T033|SY|398033008|SNOMEDCT_CORE|Family members deceased|Death of relative
C0425043|T033|SY|398033008|SNOMEDCT_CORE|Relative died|Death of relative
C0425043|T033|SY|398033008|SNOMEDCT_CORE|Relatives dead|Death of relative
C0425043|T033|SY|398033008|SNOMEDCT_CORE|Relatives deceased|Death of relative
C0425043|T033|SY|398033008|SNOMEDCT_CORE|Relatives died|Death of relative
C0425043|T033|OF|398033008|SNOMEDCT_CORE|Relatives died|Death of relative
C0425168|T033|SY|160822004|SNOMEDCT_CORE|Relational problem|Relationship problems
C0425168|T033|FN|160822004|SNOMEDCT_CORE|Relationship problems|Relationship problems
C0425168|T033|PT|160822004|SNOMEDCT_CORE|Relationship problems|Relationship problems
C0425265|T033|IS|160656007|SNOMEDCT_CORE|Will donate kidney|Willing to be donor of kidney
C0425265|T033|OF|160656007|SNOMEDCT_CORE|Will donate kidney|Willing to be donor of kidney
C0425265|T033|PT|160656007|SNOMEDCT_CORE|Willing to be donor of kidney|Willing to be donor of kidney
C0425265|T033|FN|160656007|SNOMEDCT_CORE|Willing to be donor of kidney|Willing to be donor of kidney
C0425293|T033|SY|266919005|SNOMEDCT_CORE|Never smoked|Never smoked tobacco
C0425293|T033|PT|266919005|SNOMEDCT_CORE|Never smoked tobacco|Never smoked tobacco
C0425293|T033|FN|266919005|SNOMEDCT_CORE|Never smoked tobacco|Never smoked tobacco
C0425293|T033|OF|266919005|SNOMEDCT_CORE|Never smoked tobacco|Never smoked tobacco
C0425309|T033|SY|43381005|SNOMEDCT_CORE|ETS - Exposed to tobacco smoke|Passive smoker
C0425309|T033|SY|43381005|SNOMEDCT_CORE|Exposed to environmental tobacco smoke|Passive smoker
C0425309|T033|SY|43381005|SNOMEDCT_CORE|Exposed to second hand tobacco smoke|Passive smoker
C0425309|T033|SY|43381005|SNOMEDCT_CORE|Exposed to tobacco smoke|Passive smoker
C0425309|T033|SY|43381005|SNOMEDCT_CORE|Involuntary smoker|Passive smoker
C0425309|T033|PT|43381005|SNOMEDCT_CORE|Passive smoker|Passive smoker
C0425309|T033|FN|43381005|SNOMEDCT_CORE|Passive smoker|Passive smoker
C0425310|T033|PT|160617001|SNOMEDCT_CORE|Stopped smoking|Stopped smoking
C0425310|T033|FN|160617001|SNOMEDCT_CORE|Stopped smoking|Stopped smoking
C0425310|T033|OF|160617001|SNOMEDCT_CORE|Stopped smoking|Stopped smoking
C0425311|T033|PT|160618006|SNOMEDCT_CORE|Current non-smoker|Current non-smoker
C0425311|T033|FN|160618006|SNOMEDCT_CORE|Current non-smoker|Current non-smoker
C0425311|T033|OF|160618006|SNOMEDCT_CORE|Current non-smoker|Current non-smoker
C0425496|T033|PT|248589007|SNOMEDCT_CORE|Clearing throat - hawking|Clearing throat - hawking
C0425496|T033|FN|248589007|SNOMEDCT_CORE|Clearing throat - hawking|Clearing throat - hawking
C0425512|T184|PT|248596009|SNOMEDCT_CORE|Sputum - symptom|Sputum - symptom
C0425512|T184|FN|248596009|SNOMEDCT_CORE|Sputum - symptom|Sputum - symptom
C0425770|T033|PT|116339002|SNOMEDCT_CORE|Breast finding|Breast finding
C0425770|T033|FN|116339002|SNOMEDCT_CORE|Breast finding|Breast finding
C0425770|T033|SY|116339002|SNOMEDCT_CORE|Breast observations|Breast finding
C0425775|T033|FN|248802009|SNOMEDCT_CORE|Absence of breast|Absence of breast
C0425775|T033|PT|248802009|SNOMEDCT_CORE|Absence of breast|Absence of breast
C0425779|T033|PT|271691008|SNOMEDCT_CORE|Breasts asymmetrical|Breasts asymmetrical
C0425779|T033|FN|271691008|SNOMEDCT_CORE|Breasts asymmetrical|Breasts asymmetrical
C0426065|T046|PT|199363002|SNOMEDCT_CORE|Transverse lie with antenatal problem|Transverse lie with antenatal problem
C0426065|T046|FN|199363002|SNOMEDCT_CORE|Transverse lie with antenatal problem|Transverse lie with antenatal problem
C0426066|T033|SY|86356004|SNOMEDCT_CORE|Baby keeps changing position|Unstable lie
C0426066|T033|SY|86356004|SNOMEDCT_CORE|Fetus - unstable lie|Unstable lie
C0426066|T033|SY|86356004|SNOMEDCT_CORE|Foetus - unstable lie|Unstable lie
C0426066|T033|PT|86356004|SNOMEDCT_CORE|Unstable lie|Unstable lie
C0426066|T033|FN|86356004|SNOMEDCT_CORE|Unstable lie|Unstable lie
C0426066|T033|IS|86356004|SNOMEDCT_CORE|Unstable lie of fetus|Unstable lie
C0426093|T033|SY|90381008|SNOMEDCT_CORE|OA - Occipitoanterior position|Occipitoanterior position
C0426093|T033|PT|90381008|SNOMEDCT_CORE|Occipitoanterior position|Occipitoanterior position
C0426093|T033|FN|90381008|SNOMEDCT_CORE|Occipitoanterior position|Occipitoanterior position
C0426093|T033|IS|90381008|SNOMEDCT_CORE|Occiput anterior position|Occipitoanterior position
C0426147|T033|SY|249097002|SNOMEDCT_CORE|Fetal foot presenting|Footling breech presentation
C0426147|T033|SY|249097002|SNOMEDCT_CORE|Fetal leg presenting|Footling breech presentation
C0426147|T033|SY|249097002|SNOMEDCT_CORE|Foetal foot presenting|Footling breech presentation
C0426147|T033|SY|249097002|SNOMEDCT_CORE|Foetal leg presenting|Footling breech presentation
C0426147|T033|PT|249097002|SNOMEDCT_CORE|Footling breech presentation|Footling breech presentation
C0426147|T033|FN|249097002|SNOMEDCT_CORE|Footling breech presentation|Footling breech presentation
C0426196|T033|PT|268471004|SNOMEDCT_CORE|Vaginal show|Vaginal show
C0426196|T033|FN|268471004|SNOMEDCT_CORE|Vaginal show|Vaginal show
C0426209|T033|PT|168092006|SNOMEDCT_CORE|Amniotic fluid -meconium stain|Amniotic fluid -meconium stain
C0426209|T033|FN|168092006|SNOMEDCT_CORE|Amniotic fluid -meconium stain|Amniotic fluid -meconium stain
C0426209|T033|SY|168092006|SNOMEDCT_CORE|Meconium stained amniotic fluid|Amniotic fluid -meconium stain
C0426209|T033|SY|168092006|SNOMEDCT_CORE|Meconium stained liquor|Amniotic fluid -meconium stain
C0426270|T037|SY|249220002|SNOMEDCT_CORE|Vaginal tear during delivery|Vaginal tear resulting from childbirth
C0426270|T037|PT|249220002|SNOMEDCT_CORE|Vaginal tear resulting from childbirth|Vaginal tear resulting from childbirth
C0426270|T037|FN|249220002|SNOMEDCT_CORE|Vaginal tear resulting from childbirth|Vaginal tear resulting from childbirth
C0426317|T184|PT|267062003|SNOMEDCT_CORE|Genitourinary symptoms|Genitourinary symptoms
C0426317|T184|FN|267062003|SNOMEDCT_CORE|Genitourinary symptoms|Genitourinary symptoms
C0426317|T184|SY|267062003|SNOMEDCT_CORE|GU symptoms|Genitourinary symptoms
C0426317|T184|SY|267062003|SNOMEDCT_CORE|GUT symptoms|Genitourinary symptoms
C0426348|T033|PT|249263004|SNOMEDCT_CORE|Adhesions of foreskin|Adhesions of foreskin
C0426348|T033|FN|249263004|SNOMEDCT_CORE|Adhesions of foreskin|Adhesions of foreskin
C0426359|T184|PT|249274008|SNOMEDCT_CORE|Urinary symptoms|Urinary symptoms
C0426359|T184|FN|249274008|SNOMEDCT_CORE|Urinary symptoms|Urinary symptoms
C0426359|T184|SY|249274008|SNOMEDCT_CORE|Urinary system symptoms|Urinary symptoms
C0426390|T184|SY|249297006|SNOMEDCT_CORE|Bladder spasm|Spasm of bladder
C0426390|T184|PT|249297006|SNOMEDCT_CORE|Spasm of bladder|Spasm of bladder
C0426390|T184|FN|249297006|SNOMEDCT_CORE|Spasm of bladder|Spasm of bladder
C0426551|T020|PT|249444002|SNOMEDCT_CORE|Vocal cord cyst|Vocal cord cyst
C0426551|T020|FN|249444002|SNOMEDCT_CORE|Vocal cord cyst|Vocal cord cyst
C0426623|T184|PT|162076009|SNOMEDCT_CORE|Excessive upper gastrointestinal gas|Excessive upper gastrointestinal gas
C0426623|T184|FN|162076009|SNOMEDCT_CORE|Excessive upper gastrointestinal gas|Excessive upper gastrointestinal gas
C0426636|T184|SYGB|71820002|SNOMEDCT_CORE|Defaecation urgency|Urgent desire for stool
C0426636|T184|SY|71820002|SNOMEDCT_CORE|Defecation urgency|Urgent desire for stool
C0426636|T184|SY|71820002|SNOMEDCT_CORE|Fecal urgency|Urgent desire for stool
C0426636|T184|SYGB|71820002|SNOMEDCT_CORE|Precipitancy of defaecation|Urgent desire for stool
C0426636|T184|SY|71820002|SNOMEDCT_CORE|Precipitancy of defecation|Urgent desire for stool
C0426636|T184|IS|71820002|SNOMEDCT_CORE|Rectal urgency|Urgent desire for stool
C0426636|T184|PT|71820002|SNOMEDCT_CORE|Urgent desire for stool|Urgent desire for stool
C0426636|T184|FN|71820002|SNOMEDCT_CORE|Urgent desire for stool|Urgent desire for stool
C0426732|T033|SY|249607009|SNOMEDCT_CORE|Enlarged prostate|Large prostate
C0426732|T033|PT|249607009|SNOMEDCT_CORE|Large prostate|Large prostate
C0426732|T033|FN|249607009|SNOMEDCT_CORE|Large prostate|Large prostate
C0426732|T033|SY|249607009|SNOMEDCT_CORE|Prostatomegaly|Large prostate
C0426747|T046|PT|6072007|SNOMEDCT_CORE|Bleeding from anus|Bleeding from anus
C0426747|T046|FN|6072007|SNOMEDCT_CORE|Bleeding from anus|Bleeding from anus
C0426747|T046|IS|6072007|SNOMEDCT_CORE|Hemorrhage of anus|Bleeding from anus
C0426848|T033|PT|311897005|SNOMEDCT_CORE|Sacral dimple|Sacral dimple
C0426848|T033|FN|311897005|SNOMEDCT_CORE|Sacral dimple|Sacral dimple
C0426848|T033|OAP|249729002|SNOMEDCT_CORE|Sacral dimples|Sacral dimple
C0426848|T033|OAF|249729002|SNOMEDCT_CORE|Sacral dimples|Sacral dimple
C0426900|T033|PT|249785006|SNOMEDCT_CORE|Tibial torsion|Tibial torsion
C0426900|T033|FN|249785006|SNOMEDCT_CORE|Tibial torsion|Tibial torsion
C0427036|T033|PT|249915009|SNOMEDCT_CORE|Hand joint stiff|Hand joint stiff
C0427036|T033|FN|249915009|SNOMEDCT_CORE|Hand joint stiff|Hand joint stiff
C0427068|T033|PT|249945007|SNOMEDCT_CORE|Monoparesis - leg|Monoparesis - leg
C0427068|T033|FN|249945007|SNOMEDCT_CORE|Monoparesis - leg|Monoparesis - leg
C0427068|T033|SY|249945007|SNOMEDCT_CORE|Weakness of leg|Monoparesis - leg
C0427144|T033|SY|250018006|SNOMEDCT_CORE|Toe walking|Toe-walking gait
C0427144|T033|PT|250018006|SNOMEDCT_CORE|Toe-walking gait|Toe-walking gait
C0427144|T033|FN|250018006|SNOMEDCT_CORE|Toe-walking gait|Toe-walking gait
C0427262|T033|SY|250102002|SNOMEDCT_CORE|Instability of knee|Unstable knee
C0427262|T033|SY|250102002|SNOMEDCT_CORE|Instability of knee joint|Unstable knee
C0427262|T033|SY|250102002|SNOMEDCT_CORE|Knee gives way|Unstable knee
C0427262|T033|PT|250102002|SNOMEDCT_CORE|Unstable knee|Unstable knee
C0427262|T033|FN|250102002|SNOMEDCT_CORE|Unstable knee|Unstable knee
C0427285|T184|PT|202606004|SNOMEDCT_CORE|Clicking hip|Clicking hip
C0427285|T184|FN|202606004|SNOMEDCT_CORE|Clicking hip|Clicking hip
C0427792|T033|SY|249134008|SNOMEDCT_CORE|Bloodstained amniotic fluid|Bloodstained liquor
C0427792|T033|PT|249134008|SNOMEDCT_CORE|Bloodstained liquor|Bloodstained liquor
C0427792|T033|FN|249134008|SNOMEDCT_CORE|Bloodstained liquor|Bloodstained liquor
C0428047|T033|PT|302764009|SNOMEDCT_CORE|Rubella non-immune|Rubella non-immune
C0428047|T033|FN|302764009|SNOMEDCT_CORE|Rubella non-immune|Rubella non-immune
C0428468|T033|OAP|166829003|SNOMEDCT_CORE|Serum cholesterol borderline|Serum cholesterol borderline
C0428468|T033|OAF|166829003|SNOMEDCT_CORE|Serum cholesterol borderline|Serum cholesterol borderline
C0428796|T047|SY|67754003|SNOMEDCT_CORE|Senile sclerosis of aortic cusp|Senile sclerosis of aortic cusp
C0428908|T047|SY|60423000|SNOMEDCT_CORE|Coronary sinus rhythm disorder|Sinus node dysfunction
C0428908|T047|IS|60423000|SNOMEDCT_CORE|Sinoatrial node dysfunction|Sinus node dysfunction
C0428908|T047|FN|60423000|SNOMEDCT_CORE|Sinus node dysfunction|Sinus node dysfunction
C0428908|T047|PT|60423000|SNOMEDCT_CORE|Sinus node dysfunction|Sinus node dysfunction
C0428974|T047|PT|72654001|SNOMEDCT_CORE|Supraventricular arrhythmia|Supraventricular arrhythmia
C0428974|T047|FN|72654001|SNOMEDCT_CORE|Supraventricular arrhythmia|Supraventricular arrhythmia
C0428974|T047|IS|72654001|SNOMEDCT_CORE|Supraventricular arrhythmia, NOS|Supraventricular arrhythmia
C0428977|T033|PT|48867003|SNOMEDCT_CORE|Bradycardia|Bradycardia
C0428977|T033|FN|48867003|SNOMEDCT_CORE|Bradycardia|Bradycardia
C0428977|T033|OF|48867003|SNOMEDCT_CORE|Bradycardia|Bradycardia
C0428977|T033|IS|48867003|SNOMEDCT_CORE|Bradycardia, NOS|Bradycardia
C0428977|T033|SY|48867003|SNOMEDCT_CORE|Decreased heart rate|Bradycardia
C0428977|T033|SY|48867003|SNOMEDCT_CORE|Heart rate slow|Bradycardia
C0428977|T033|SY|48867003|SNOMEDCT_CORE|Slow heart beat|Bradycardia
C0429468|T047|SY|266609001|SNOMEDCT_CORE|Anovular cycle|Anovular cycle
C0429803|T190|PT|79184009|SNOMEDCT_CORE|Bladder trabeculation|Bladder trabeculation
C0429803|T190|FN|79184009|SNOMEDCT_CORE|Bladder trabeculation|Bladder trabeculation
C0429803|T190|SY|79184009|SNOMEDCT_CORE|Trabeculated bladder|Bladder trabeculation
C0429826|T033|SY|252030006|SNOMEDCT_CORE|Dysfunctional elimination of urine|Dysfunctional voiding of urine
C0429826|T033|PT|252030006|SNOMEDCT_CORE|Dysfunctional voiding of urine|Dysfunctional voiding of urine
C0429826|T033|FN|252030006|SNOMEDCT_CORE|Dysfunctional voiding of urine|Dysfunctional voiding of urine
C0429826|T033|SY|252030006|SNOMEDCT_CORE|Voiding dysfunction|Dysfunctional voiding of urine
C0431108|T191|SY|22217002|SNOMEDCT_CORE|Anaplastic oligoastrocytoma|Anaplastic oligoastrocytoma
C0431319|T019|PT|203936004|SNOMEDCT_CORE|Lumbar spina bifida with hydrocephalus|Lumbar spina bifida with hydrocephalus
C0431319|T019|FN|203936004|SNOMEDCT_CORE|Lumbar spina bifida with hydrocephalus|Lumbar spina bifida with hydrocephalus
C0431661|T019|SY|268228006|SNOMEDCT_CORE|Imperfectly descended testes - bilateral|Imperfectly descended testes - bilateral
C0431661|T019|SY|268228006|SNOMEDCT_CORE|Maldescent of testes - bilateral|Imperfectly descended testes - bilateral
C0431662|T019|SY|268227001|SNOMEDCT_CORE|IDT - Imperfectly descended testis - unilateral|IDT - Imperfectly descended testis - unilateral
C0431662|T019|SY|268227001|SNOMEDCT_CORE|Imperfectly descended testis - unilateral|IDT - Imperfectly descended testis - unilateral
C0431662|T019|SY|268227001|SNOMEDCT_CORE|Maldescent of testis - unilateral|IDT - Imperfectly descended testis - unilateral
C0431663|T019|SY|268228006|SNOMEDCT_CORE|Cryptorchidism, bilateral|Undescended testes - bilateral
C0431663|T019|SY|268228006|SNOMEDCT_CORE|UDT - Undescended testes bilateral|Undescended testes - bilateral
C0431663|T019|PT|268228006|SNOMEDCT_CORE|Undescended testes - bilateral|Undescended testes - bilateral
C0431663|T019|FN|268228006|SNOMEDCT_CORE|Undescended testes - bilateral|Undescended testes - bilateral
C0431663|T019|SY|268228006|SNOMEDCT_CORE|Undescended testis, bilateral|Undescended testes - bilateral
C0431664|T019|SY|268227001|SNOMEDCT_CORE|Cryptorchidism, unilateral|Unilateral undescended testis
C0431664|T019|SY|268227001|SNOMEDCT_CORE|UDT - Undescended testis unilateral|Unilateral undescended testis
C0431664|T019|SY|268227001|SNOMEDCT_CORE|Undescended testis, unilateral|Unilateral undescended testis
C0431664|T019|OF|268227001|SNOMEDCT_CORE|Undescended testis, unilateral|Unilateral undescended testis
C0431664|T019|PT|268227001|SNOMEDCT_CORE|Unilateral undescended testis|Unilateral undescended testis
C0431664|T019|FN|268227001|SNOMEDCT_CORE|Unilateral undescended testis|Unilateral undescended testis
C0431750|T047|SY|197919005|SNOMEDCT_CORE|Meatal stenosis|Stenosis of urinary meatus
C0431750|T047|PT|197919005|SNOMEDCT_CORE|Stenosis of urinary meatus|Stenosis of urinary meatus
C0431750|T047|FN|197919005|SNOMEDCT_CORE|Stenosis of urinary meatus|Stenosis of urinary meatus
C0432162|T019|SY|80712009|SNOMEDCT_CORE|Congenital lumbosacral spondylolysis|Congenital spondylolysis of lumbosacral region
C0432162|T019|PT|80712009|SNOMEDCT_CORE|Congenital spondylolysis of lumbosacral region|Congenital spondylolysis of lumbosacral region
C0432162|T019|FN|80712009|SNOMEDCT_CORE|Congenital spondylolysis of lumbosacral region|Congenital spondylolysis of lumbosacral region
C0432556|T191|PT|93195001|SNOMEDCT_CORE|Malignant lymphoma of lymph nodes of head, face AND/OR neck|Malignant lymphoma of lymph nodes of head, face AND/OR neck
C0432556|T191|FN|93195001|SNOMEDCT_CORE|Malignant lymphoma of lymph nodes of head, face AND/OR neck|Malignant lymphoma of lymph nodes of head, face AND/OR neck
C0432556|T191|IS|93195001|SNOMEDCT_CORE|Malignant lymphoma, NOS of lymph nodes of head, face, and neck|Malignant lymphoma of lymph nodes of head, face AND/OR neck
C0432563|T191|PT|93197009|SNOMEDCT_CORE|Malignant lymphoma of lymph nodes of multiple sites|Malignant lymphoma of lymph nodes of multiple sites
C0432563|T191|FN|93197009|SNOMEDCT_CORE|Malignant lymphoma of lymph nodes of multiple sites|Malignant lymphoma of lymph nodes of multiple sites
C0432563|T191|IS|93197009|SNOMEDCT_CORE|Malignant lymphoma, NOS of lymph nodes of multiple sites|Malignant lymphoma of lymph nodes of multiple sites
C0432750|T037|SY|125668004|SNOMEDCT_CORE|Bruise of face|Contusion of face
C0432750|T037|PT|125668004|SNOMEDCT_CORE|Contusion of face|Contusion of face
C0432750|T037|FN|125668004|SNOMEDCT_CORE|Contusion of face|Contusion of face
C0432750|T037|SY|125668004|SNOMEDCT_CORE|Superficial bruising of face|Contusion of face
C0432762|T037|PT|39812007|SNOMEDCT_CORE|Contusion of forearm|Contusion of forearm
C0432762|T037|FN|39812007|SNOMEDCT_CORE|Contusion of forearm|Contusion of forearm
C0432762|T037|SY|39812007|SNOMEDCT_CORE|Contusion, forearm area|Contusion of forearm
C0432762|T037|SY|39812007|SNOMEDCT_CORE|Superficial bruising of forearm|Contusion of forearm
C0432763|T037|PT|91613004|SNOMEDCT_CORE|Contusion of elbow|Contusion of elbow
C0432763|T037|FN|91613004|SNOMEDCT_CORE|Contusion of elbow|Contusion of elbow
C0432763|T037|SY|91613004|SNOMEDCT_CORE|Contusion, elbow area|Contusion of elbow
C0432763|T037|SY|91613004|SNOMEDCT_CORE|Superficial bruising of elbow|Contusion of elbow
C0432769|T037|PT|5662003|SNOMEDCT_CORE|Contusion of hand|Contusion of hand
C0432769|T037|FN|5662003|SNOMEDCT_CORE|Contusion of hand|Contusion of hand
C0432769|T037|SY|5662003|SNOMEDCT_CORE|Superficial bruising of hand|Contusion of hand
C0432773|T037|PT|69787006|SNOMEDCT_CORE|Contusion of finger|Contusion of finger
C0432773|T037|FN|69787006|SNOMEDCT_CORE|Contusion of finger|Contusion of finger
C0432773|T037|SY|69787006|SNOMEDCT_CORE|Contusion, finger|Contusion of finger
C0432773|T037|SY|69787006|SNOMEDCT_CORE|Superficial bruising of finger|Contusion of finger
C0432794|T037|PT|210987008|SNOMEDCT_CORE|Abrasion of face|Abrasion of face
C0432794|T037|FN|210987008|SNOMEDCT_CORE|Abrasion of face|Abrasion of face
C0432794|T037|SY|210987008|SNOMEDCT_CORE|Abrasion, face|Abrasion of face
C0432794|T037|SY|210987008|SNOMEDCT_CORE|Facial graze|Abrasion of face
C0432794|T037|SY|210987008|SNOMEDCT_CORE|Graze of face|Abrasion of face
C0432929|T037|PT|210456000|SNOMEDCT_CORE|Open wound of anterior abdominal wall|Open wound of anterior abdominal wall
C0432929|T037|FN|210456000|SNOMEDCT_CORE|Open wound of anterior abdominal wall|Open wound of anterior abdominal wall
C0432948|T037|PT|210339009|SNOMEDCT_CORE|Open wound of face|Open wound of face
C0432948|T037|FN|210339009|SNOMEDCT_CORE|Open wound of face|Open wound of face
C0432966|T037|PT|125651003|SNOMEDCT_CORE|Open wound of wrist|Open wound of wrist
C0432966|T037|FN|125651003|SNOMEDCT_CORE|Open wound of wrist|Open wound of wrist
C0432975|T037|PT|284549007|SNOMEDCT_CORE|Laceration of hand|Laceration of hand
C0432975|T037|FN|284549007|SNOMEDCT_CORE|Laceration of hand|Laceration of hand
C0432980|T037|PT|210565009|SNOMEDCT_CORE|Open wound of hand with complication|Open wound of hand with complication
C0432980|T037|FN|210565009|SNOMEDCT_CORE|Open wound of hand with complication|Open wound of hand with complication
C0432981|T037|PT|274172008|SNOMEDCT_CORE|Laceration of finger|Laceration of finger
C0432981|T037|FN|274172008|SNOMEDCT_CORE|Laceration of finger|Laceration of finger
C0432988|T037|PT|210682000|SNOMEDCT_CORE|Open wound of knee and/or leg and/or ankle|Open wound of knee and/or leg and/or ankle
C0432988|T037|FN|210682000|SNOMEDCT_CORE|Open wound of knee and/or leg and/or ankle|Open wound of knee and/or leg and/or ankle
C0432988|T037|SY|210682000|SNOMEDCT_CORE|Open wound of knee, leg and ankle|Open wound of knee and/or leg and/or ankle
C0432988|T037|OF|210682000|SNOMEDCT_CORE|Open wound of knee, leg and ankle|Open wound of knee and/or leg and/or ankle
C0433054|T037|PT|262555007|SNOMEDCT_CORE|Human bite - wound|Human bite - wound
C0433054|T037|FN|262555007|SNOMEDCT_CORE|Human bite - wound|Human bite - wound
C0433163|T037|PT|262582004|SNOMEDCT_CORE|Burn of face|Burn of face
C0433163|T037|FN|262582004|SNOMEDCT_CORE|Burn of face|Burn of face
C0433163|T037|SY|262582004|SNOMEDCT_CORE|Face burns|Burn of face
C0433163|T037|OF|262582004|SNOMEDCT_CORE|Face burns|Burn of face
C0433163|T037|SY|262582004|SNOMEDCT_CORE|Facial burn|Burn of face
C0433654|T037|PT|262599003|SNOMEDCT_CORE|Foreign body in respiratory tract|Foreign body in respiratory tract
C0433654|T037|FN|262599003|SNOMEDCT_CORE|Foreign body in respiratory tract|Foreign body in respiratory tract
C0434302|T037|PT|210566005|SNOMEDCT_CORE|Open wound of hand with tendon involvement|Open wound of hand with tendon involvement
C0434302|T037|FN|210566005|SNOMEDCT_CORE|Open wound of hand with tendon involvement|Open wound of hand with tendon involvement
C0434321|T037|IS|262975009|SNOMEDCT_CORE|Back strain|Strain of tendon of back
C0434321|T037|IS|262975009|SNOMEDCT_CORE|Strain of back|Strain of tendon of back
C0434321|T037|PT|262975009|SNOMEDCT_CORE|Strain of tendon of back|Strain of tendon of back
C0434321|T037|FN|262975009|SNOMEDCT_CORE|Strain of tendon of back|Strain of tendon of back
C0434322|T037|OAP|74779009|SNOMEDCT_CORE|Strain of rotator cuff capsule|Strain of rotator cuff of shoulder
C0434322|T037|OAF|74779009|SNOMEDCT_CORE|Strain of rotator cuff capsule|Strain of rotator cuff of shoulder
C0434322|T037|OAS|74779009|SNOMEDCT_CORE|Strain of rotator cuff of shoulder|Strain of rotator cuff of shoulder
C0434322|T037|PT|789758005|SNOMEDCT_CORE|Strain of rotator cuff of shoulder|Strain of rotator cuff of shoulder
C0434322|T037|FN|789758005|SNOMEDCT_CORE|Strain of rotator cuff of shoulder|Strain of rotator cuff of shoulder
C0434416|T037|SY|269134004|SNOMEDCT_CORE|Sprain elbow and forearm|Sprain of elbow and forearm
C0434416|T037|PT|269134004|SNOMEDCT_CORE|Sprain of elbow and forearm|Sprain of elbow and forearm
C0434416|T037|FN|269134004|SNOMEDCT_CORE|Sprain of elbow and forearm|Sprain of elbow and forearm
C0434421|T037|SY|17883008|SNOMEDCT_CORE|Sprain of hip and thigh|Sprain of hip and thigh
C0434423|T037|OAP|262992000|SNOMEDCT_CORE|Hamstring sprain|Hamstring sprain
C0434423|T037|OAF|262992000|SNOMEDCT_CORE|Hamstring sprain|Hamstring sprain
C0434425|T037|OAP|269137006|SNOMEDCT_CORE|Sprain of knee and leg|Sprain of knee and leg
C0434425|T037|OAF|269137006|SNOMEDCT_CORE|Sprain of knee and leg|Sprain of knee and leg
C0434480|T037|PT|262998001|SNOMEDCT_CORE|Sprain of toe joint|Sprain of toe joint
C0434480|T037|FN|262998001|SNOMEDCT_CORE|Sprain of toe joint|Sprain of toe joint
C0434480|T037|SY|262998001|SNOMEDCT_CORE|Sprained toe|Sprain of toe joint
C0434480|T037|SY|262998001|SNOMEDCT_CORE|Toe sprain|Sprain of toe joint
C0434482|T037|PT|263000005|SNOMEDCT_CORE|Joint capsule sprain|Joint capsule sprain
C0434482|T037|FN|263000005|SNOMEDCT_CORE|Joint capsule sprain|Joint capsule sprain
C0434579|T037|IS|125614009|SNOMEDCT_CORE|Closed dislocation of glenohumeral joint|Closed traumatic dislocation of glenohumeral joint
C0434579|T037|IS|125614009|SNOMEDCT_CORE|Closed dislocation of humerus|Closed traumatic dislocation of glenohumeral joint
C0434579|T037|IS|22911007|SNOMEDCT_CORE|Closed dislocation of humerus, NOS|Closed traumatic dislocation of glenohumeral joint
C0434579|T037|OP|22911007|SNOMEDCT_CORE|Closed dislocation of shoulder region|Closed traumatic dislocation of glenohumeral joint
C0434579|T037|IS|22911007|SNOMEDCT_CORE|Closed dislocation of shoulder, NOS|Closed traumatic dislocation of glenohumeral joint
C0434579|T037|PT|125614009|SNOMEDCT_CORE|Closed traumatic dislocation of glenohumeral joint|Closed traumatic dislocation of glenohumeral joint
C0434579|T037|FN|125614009|SNOMEDCT_CORE|Closed traumatic dislocation of glenohumeral joint|Closed traumatic dislocation of glenohumeral joint
C0434579|T037|FN|22911007|SNOMEDCT_CORE|Closed traumatic dislocation of joint of shoulder region|Closed traumatic dislocation of glenohumeral joint
C0434579|T037|PT|22911007|SNOMEDCT_CORE|Closed traumatic dislocation of joint of shoulder region|Closed traumatic dislocation of glenohumeral joint
C0434579|T037|SY|125614009|SNOMEDCT_CORE|Closed traumatic shoulder dislocation|Closed traumatic dislocation of glenohumeral joint
C0434599|T037|OP|2651006|SNOMEDCT_CORE|Closed dislocation of elbow|Closed traumatic dislocation of elbow joint
C0434599|T037|IS|2651006|SNOMEDCT_CORE|Closed dislocation of elbow, NOS|Closed traumatic dislocation of elbow joint
C0434599|T037|PT|2651006|SNOMEDCT_CORE|Closed traumatic dislocation of elbow joint|Closed traumatic dislocation of elbow joint
C0434599|T037|FN|2651006|SNOMEDCT_CORE|Closed traumatic dislocation of elbow joint|Closed traumatic dislocation of elbow joint
C0434662|T037|PT|208892001|SNOMEDCT_CORE|Closed traumatic dislocation of hip|Closed traumatic dislocation of hip
C0434662|T037|FN|208892001|SNOMEDCT_CORE|Closed traumatic dislocation of hip|Closed traumatic dislocation of hip
C0434662|T037|OAF|63079007|SNOMEDCT_CORE|Closed traumatic dislocation of hip joint|Closed traumatic dislocation of hip
C0434662|T037|OAS|63079007|SNOMEDCT_CORE|Closed traumatic dislocation of hip joint|Closed traumatic dislocation of hip
C0434662|T037|SY|208892001|SNOMEDCT_CORE|Closed traumatic dislocation of hip joint|Closed traumatic dislocation of hip
C0434685|T037|SY|208929003|SNOMEDCT_CORE|Closed traumatic dislocation of patella|Closed traumatic dislocation of patellofemoral joint
C0434685|T037|PT|208929003|SNOMEDCT_CORE|Closed traumatic dislocation of patellofemoral joint|Closed traumatic dislocation of patellofemoral joint
C0434685|T037|FN|208929003|SNOMEDCT_CORE|Closed traumatic dislocation of patellofemoral joint|Closed traumatic dislocation of patellofemoral joint
C0434692|T037|PT|208981003|SNOMEDCT_CORE|Closed traumatic dislocation ankle joint|Closed traumatic dislocation ankle joint
C0434692|T037|FN|208981003|SNOMEDCT_CORE|Closed traumatic dislocation ankle joint|Closed traumatic dislocation ankle joint
C0434984|T037|PT|269113006|SNOMEDCT_CORE|Acute meniscal tear, medial|Acute meniscal tear, medial
C0434984|T037|FN|269113006|SNOMEDCT_CORE|Acute meniscal tear, medial|Acute meniscal tear, medial
C0434993|T037|PT|208921000|SNOMEDCT_CORE|Acute meniscal tear, lateral|Acute meniscal tear, lateral
C0434993|T037|FN|208921000|SNOMEDCT_CORE|Acute meniscal tear, lateral|Acute meniscal tear, lateral
C0435002|T037|SY|398878007|SNOMEDCT_CORE|Ligament sprain|Sprain of ligament
C0435002|T037|PT|398878007|SNOMEDCT_CORE|Sprain of ligament|Sprain of ligament
C0435002|T037|FN|398878007|SNOMEDCT_CORE|Sprain of ligament|Sprain of ligament
C0435024|T037|SY|263128001|SNOMEDCT_CORE|Elbow sprain|Sprain of ligament of elbow
C0435024|T037|SY|263128001|SNOMEDCT_CORE|Sprain of elbow|Sprain of ligament of elbow
C0435024|T037|SY|263128001|SNOMEDCT_CORE|Sprain of elbow joint|Sprain of ligament of elbow
C0435024|T037|PT|263128001|SNOMEDCT_CORE|Sprain of ligament of elbow|Sprain of ligament of elbow
C0435024|T037|FN|263128001|SNOMEDCT_CORE|Sprain of ligament of elbow|Sprain of ligament of elbow
C0435128|T037|PT|209629006|SNOMEDCT_CORE|Complete tear, knee, anterior cruciate ligament|Complete tear, knee, anterior cruciate ligament
C0435128|T037|FN|209629006|SNOMEDCT_CORE|Complete tear, knee, anterior cruciate ligament|Complete tear, knee, anterior cruciate ligament
C0435236|T037|PT|207687004|SNOMEDCT_CORE|Closed fracture vault of skull with intracranial injury|Closed fracture vault of skull with intracranial injury
C0435236|T037|OF|207687004|SNOMEDCT_CORE|Closed fracture vault of skull with intracranial injury|Closed fracture vault of skull with intracranial injury
C0435236|T037|FN|207687004|SNOMEDCT_CORE|Intracranial injury co-occurrent and due to closed fracture of vault of skull|Closed fracture vault of skull with intracranial injury
C0435236|T037|SY|207687004|SNOMEDCT_CORE|Intracranial injury co-occurrent and due to closed fracture of vault of skull|Closed fracture vault of skull with intracranial injury
C0435352|T037|PT|269062008|SNOMEDCT_CORE|Closed fracture of cervical spine|Closed fracture of cervical spine
C0435352|T037|FN|269062008|SNOMEDCT_CORE|Closed fracture of cervical spine|Closed fracture of cervical spine
C0435522|T037|SY|1658003|SNOMEDCT_CORE|Closed fracture clavicle, lateral end|Closed fracture of acromial end of clavicle
C0435522|T037|PT|1658003|SNOMEDCT_CORE|Closed fracture of acromial end of clavicle|Closed fracture of acromial end of clavicle
C0435522|T037|FN|1658003|SNOMEDCT_CORE|Closed fracture of acromial end of clavicle|Closed fracture of acromial end of clavicle
C0435532|T037|SY|208241000|SNOMEDCT_CORE|Closed fracture of anatomical neck of humerus|Closed fracture of proximal humerus, anatomical neck
C0435532|T037|PT|208241000|SNOMEDCT_CORE|Closed fracture of proximal humerus, anatomical neck|Closed fracture of proximal humerus, anatomical neck
C0435532|T037|FN|208241000|SNOMEDCT_CORE|Closed fracture of proximal humerus, anatomical neck|Closed fracture of proximal humerus, anatomical neck
C0435533|T037|PT|208242007|SNOMEDCT_CORE|Closed fracture proximal humerus, greater tuberosity|Closed fracture proximal humerus, greater tuberosity
C0435533|T037|FN|208242007|SNOMEDCT_CORE|Closed fracture proximal humerus, greater tuberosity|Closed fracture proximal humerus, greater tuberosity
C0435552|T037|PT|208271008|SNOMEDCT_CORE|Closed fracture distal humerus, lateral epicondyle|Closed fracture distal humerus, lateral epicondyle
C0435552|T037|FN|208271008|SNOMEDCT_CORE|Closed fracture distal humerus, lateral epicondyle|Closed fracture distal humerus, lateral epicondyle
C0435553|T037|IS|21419000|SNOMEDCT_CORE|Closed fracture distal humerus, medial epicondyle|Closed fracture of medial condyle of humerus
C0435553|T037|IS|21419000|SNOMEDCT_CORE|Closed fracture of internal epicondyle of humerus|Closed fracture of medial condyle of humerus
C0435553|T037|PT|21419000|SNOMEDCT_CORE|Closed fracture of medial condyle of humerus|Closed fracture of medial condyle of humerus
C0435553|T037|FN|21419000|SNOMEDCT_CORE|Closed fracture of medial condyle of humerus|Closed fracture of medial condyle of humerus
C0435569|T037|SY|58580000|SNOMEDCT_CORE|Closed fracture distal humerus, supracondylar|Closed supracondylar fracture of humerus
C0435569|T037|PT|58580000|SNOMEDCT_CORE|Closed supracondylar fracture of humerus|Closed supracondylar fracture of humerus
C0435569|T037|FN|58580000|SNOMEDCT_CORE|Closed supracondylar fracture of humerus|Closed supracondylar fracture of humerus
C0435577|T037|PT|263196008|SNOMEDCT_CORE|Fracture of radial head|Fracture of radial head
C0435577|T037|FN|263196008|SNOMEDCT_CORE|Fracture of radial head|Fracture of radial head
C0435579|T037|PT|263197004|SNOMEDCT_CORE|Fracture of radial neck|Fracture of radial neck
C0435579|T037|FN|263197004|SNOMEDCT_CORE|Fracture of radial neck|Fracture of radial neck
C0435585|T037|PT|263199001|SNOMEDCT_CORE|Fracture of distal end of radius|Fracture of distal end of radius
C0435585|T037|FN|263199001|SNOMEDCT_CORE|Fracture of distal end of radius|Fracture of distal end of radius
C0435585|T037|SY|263199001|SNOMEDCT_CORE|Fracture of lower end of radius|Fracture of distal end of radius
C0435603|T037|PT|68819003|SNOMEDCT_CORE|Closed fracture of coronoid process of ulna|Closed fracture of coronoid process of ulna
C0435603|T037|FN|68819003|SNOMEDCT_CORE|Closed fracture of coronoid process of ulna|Closed fracture of coronoid process of ulna
C0435603|T037|SY|68819003|SNOMEDCT_CORE|Closed fracture of ulna, coronoid|Closed fracture of coronoid process of ulna
C0435612|T037|PT|53792000|SNOMEDCT_CORE|Closed fracture of shaft of ulna|Closed fracture of shaft of ulna
C0435612|T037|FN|53792000|SNOMEDCT_CORE|Closed fracture of shaft of ulna|Closed fracture of shaft of ulna
C0435612|T037|SY|53792000|SNOMEDCT_CORE|Closed fracture of the ulnar shaft|Closed fracture of shaft of ulna
C0435620|T037|PT|91419009|SNOMEDCT_CORE|Closed fracture of forearm|Closed fracture of forearm
C0435620|T037|FN|91419009|SNOMEDCT_CORE|Closed fracture of forearm|Closed fracture of forearm
C0435620|T037|IS|91419009|SNOMEDCT_CORE|Closed fracture of forearm, NOS|Closed fracture of forearm
C0435627|T037|SY|263207000|SNOMEDCT_CORE|Fracture of shaft of radius and ulna|Fracture of shaft of radius and/or ulna
C0435627|T037|OF|263207000|SNOMEDCT_CORE|Fracture of shaft of radius and ulna|Fracture of shaft of radius and/or ulna
C0435627|T037|PT|263207000|SNOMEDCT_CORE|Fracture of shaft of radius and/or ulna|Fracture of shaft of radius and/or ulna
C0435627|T037|FN|263207000|SNOMEDCT_CORE|Fracture of shaft of radius and/or ulna|Fracture of shaft of radius and/or ulna
C0435630|T037|PT|263208005|SNOMEDCT_CORE|Fracture of distal end of radius and ulna|Fracture of distal end of radius and ulna
C0435630|T037|FN|263208005|SNOMEDCT_CORE|Fracture of distal end of radius and ulna|Fracture of distal end of radius and ulna
C0435630|T037|SY|263208005|SNOMEDCT_CORE|Fracture of lower end of both ulna and radius|Fracture of distal end of radius and ulna
C0435630|T037|IS|263208005|SNOMEDCT_CORE|Fracture of wrist|Fracture of distal end of radius and ulna
C0435632|T037|SY|20511007|SNOMEDCT_CORE|Fracture of bone of hand|Fracture of hand
C0435632|T037|PT|20511007|SNOMEDCT_CORE|Fracture of hand|Fracture of hand
C0435632|T037|FN|20511007|SNOMEDCT_CORE|Fracture of hand|Fracture of hand
C0435632|T037|SY|20511007|SNOMEDCT_CORE|Fracture of hand bone|Fracture of hand
C0435632|T037|IS|20511007|SNOMEDCT_CORE|Fracture of hand bone, NOS|Fracture of hand
C0435632|T037|IS|20511007|SNOMEDCT_CORE|Fracture of hand, NOS|Fracture of hand
C0435644|T037|SY|42818005|SNOMEDCT_CORE|Closed fracture of navicular bone of wrist|Closed fracture of scaphoid bone of wrist
C0435644|T037|FN|42818005|SNOMEDCT_CORE|Closed fracture of navicular bone of wrist|Closed fracture of scaphoid bone of wrist
C0435644|T037|IS|42818005|SNOMEDCT_CORE|Closed fracture of of navicular bone of wrist|Closed fracture of scaphoid bone of wrist
C0435644|T037|OF|42818005|SNOMEDCT_CORE|Closed fracture of of navicular bone of wrist|Closed fracture of scaphoid bone of wrist
C0435644|T037|PT|42818005|SNOMEDCT_CORE|Closed fracture of scaphoid bone of wrist|Closed fracture of scaphoid bone of wrist
C0435644|T037|SY|42818005|SNOMEDCT_CORE|Closed fracture of the scaphoid|Closed fracture of scaphoid bone of wrist
C0435700|T037|PT|208444006|SNOMEDCT_CORE|Closed fracture finger proximal phalanx|Closed fracture finger proximal phalanx
C0435700|T037|FN|208444006|SNOMEDCT_CORE|Closed fracture finger proximal phalanx|Closed fracture finger proximal phalanx
C0435702|T037|PT|208446008|SNOMEDCT_CORE|Closed fracture finger proximal phalanx, shaft|Closed fracture finger proximal phalanx, shaft
C0435702|T037|FN|208446008|SNOMEDCT_CORE|Closed fracture finger proximal phalanx, shaft|Closed fracture finger proximal phalanx, shaft
C0435705|T037|PT|208449001|SNOMEDCT_CORE|Closed fracture finger proximal phalanx, multiple|Closed fracture finger proximal phalanx, multiple
C0435705|T037|FN|208449001|SNOMEDCT_CORE|Closed fracture finger proximal phalanx, multiple|Closed fracture finger proximal phalanx, multiple
C0435706|T037|PT|208450001|SNOMEDCT_CORE|Closed fracture finger middle phalanx|Closed fracture finger middle phalanx
C0435706|T037|FN|208450001|SNOMEDCT_CORE|Closed fracture finger middle phalanx|Closed fracture finger middle phalanx
C0435750|T037|PT|60667009|SNOMEDCT_CORE|Closed fracture of rib|Closed fracture of rib
C0435750|T037|FN|60667009|SNOMEDCT_CORE|Closed fracture of rib|Closed fracture of rib
C0435750|T037|IS|60667009|SNOMEDCT_CORE|Closed fracture of rib, NOS|Closed fracture of rib
C0435750|T037|SY|60667009|SNOMEDCT_CORE|Closed fracture rib|Closed fracture of rib
C0435805|T037|PT|263225007|SNOMEDCT_CORE|Fracture of proximal end of femur|Fracture of proximal end of femur
C0435805|T037|FN|263225007|SNOMEDCT_CORE|Fracture of proximal end of femur|Fracture of proximal end of femur
C0435844|T037|SY|30905007|SNOMEDCT_CORE|Closed fracture distal femur, supracondylar|Closed supracondylar fracture of femur
C0435844|T037|PT|30905007|SNOMEDCT_CORE|Closed supracondylar fracture of femur|Closed supracondylar fracture of femur
C0435844|T037|FN|30905007|SNOMEDCT_CORE|Closed supracondylar fracture of femur|Closed supracondylar fracture of femur
C0435884|T037|PT|208634001|SNOMEDCT_CORE|Closed fracture distal tibia|Closed fracture distal tibia
C0435884|T037|FN|208634001|SNOMEDCT_CORE|Closed fracture distal tibia|Closed fracture distal tibia
C0435890|T037|SY|15385006|SNOMEDCT_CORE|Closed fracture ankle, medial malleolus|Closed fracture of medial malleolus
C0435890|T037|PT|15385006|SNOMEDCT_CORE|Closed fracture of medial malleolus|Closed fracture of medial malleolus
C0435890|T037|FN|15385006|SNOMEDCT_CORE|Closed fracture of medial malleolus|Closed fracture of medial malleolus
C0435892|T037|SY|34268009|SNOMEDCT_CORE|Closed fracture ankle, lateral malleolus|Closed fracture of lateral malleolus
C0435892|T037|PT|34268009|SNOMEDCT_CORE|Closed fracture of lateral malleolus|Closed fracture of lateral malleolus
C0435892|T037|FN|34268009|SNOMEDCT_CORE|Closed fracture of lateral malleolus|Closed fracture of lateral malleolus
C0435908|T037|PT|263244000|SNOMEDCT_CORE|Bimalleolar fracture of ankle|Bimalleolar fracture of ankle
C0435908|T037|FN|263244000|SNOMEDCT_CORE|Bimalleolar fracture of ankle|Bimalleolar fracture of ankle
C0435908|T037|SY|263244000|SNOMEDCT_CORE|Fracture of medial and lateral malleoli|Bimalleolar fracture of ankle
C0435943|T037|SY|263251009|SNOMEDCT_CORE|Fracture of metatarsal bone|Metatarsal bone fracture
C0435943|T037|PT|263251009|SNOMEDCT_CORE|Metatarsal bone fracture|Metatarsal bone fracture
C0435943|T037|FN|263251009|SNOMEDCT_CORE|Metatarsal bone fracture|Metatarsal bone fracture
C0435944|T037|SY|36924003|SNOMEDCT_CORE|Closed fracture metatarsal|Closed fracture of metatarsal bone
C0435944|T037|PT|36924003|SNOMEDCT_CORE|Closed fracture of metatarsal bone|Closed fracture of metatarsal bone
C0435944|T037|FN|36924003|SNOMEDCT_CORE|Closed fracture of metatarsal bone|Closed fracture of metatarsal bone
C0435944|T037|IS|36924003|SNOMEDCT_CORE|Closed fracture of metatarsal bone, NOS|Closed fracture of metatarsal bone
C0435961|T037|PT|208713003|SNOMEDCT_CORE|Closed fracture multiple phalanges, toe|Closed fracture multiple phalanges, toe
C0435961|T037|FN|208713003|SNOMEDCT_CORE|Closed fracture multiple phalanges, toe|Closed fracture multiple phalanges, toe
C0436449|T033|PT|168749009|SNOMEDCT_CORE|Mammography normal|Mammography normal
C0436449|T033|FN|168749009|SNOMEDCT_CORE|Mammography normal|Mammography normal
C0436485|T033|PT|168501001|SNOMEDCT_CORE|Radiology result abnormal|Radiology result abnormal
C0436485|T033|FN|168501001|SNOMEDCT_CORE|Radiology result abnormal|Radiology result abnormal
C0436503|T033|PT|168734001|SNOMEDCT_CORE|Standard chest X-ray abnormal|Standard chest X-ray abnormal
C0436503|T033|FN|168734001|SNOMEDCT_CORE|Standard chest X-ray abnormal|Standard chest X-ray abnormal
C0436515|T033|PT|168840001|SNOMEDCT_CORE|Barium enema abnormal|Barium enema abnormal
C0436515|T033|FN|168840001|SNOMEDCT_CORE|Barium enema abnormal|Barium enema abnormal
C0436539|T033|IS|129679001|SNOMEDCT_CORE|Abnormal CT scan|Computed tomography result abnormal
C0436539|T033|OF|129679001|SNOMEDCT_CORE|Abnormal CT scan|Computed tomography result abnormal
C0436539|T033|IS|129679001|SNOMEDCT_CORE|CAT scan abnormal|Computed tomography result abnormal
C0436539|T033|PT|129679001|SNOMEDCT_CORE|Computed tomography result abnormal|Computed tomography result abnormal
C0436539|T033|FN|129679001|SNOMEDCT_CORE|Computed tomography result abnormal|Computed tomography result abnormal
C0436540|T033|FN|169083003|SNOMEDCT_CORE|Magnetic resonance imaging scan abnormal|MRI scan abnormal
C0436540|T033|SY|169083003|SNOMEDCT_CORE|Magnetic resonance imaging scan abnormal|MRI scan abnormal
C0436540|T033|PT|169083003|SNOMEDCT_CORE|MRI scan abnormal|MRI scan abnormal
C0436540|T033|IS|169083003|SNOMEDCT_CORE|Nuclear magn.reson. abnormal|MRI scan abnormal
C0436540|T033|OF|169083003|SNOMEDCT_CORE|Nuclear magnetic resonance abnormal|MRI scan abnormal
C0436540|T033|OP|169083003|SNOMEDCT_CORE|Nuclear magnetic resonance abnormal|MRI scan abnormal
C0438065|T033|PT|161800001|SNOMEDCT_CORE|H/O: hysterectomy|H/O: hysterectomy
C0438065|T033|OF|161800001|SNOMEDCT_CORE|History of - hysterectomy|H/O: hysterectomy
C0438065|T033|IS|161800001|SNOMEDCT_CORE|History of - hysterectomy|H/O: hysterectomy
C0438065|T033|FN|161800001|SNOMEDCT_CORE|History of hysterectomy|H/O: hysterectomy
C0438065|T033|SY|161800001|SNOMEDCT_CORE|History of hysterectomy|H/O: hysterectomy
C0438066|T033|PT|267020005|SNOMEDCT_CORE|H/O: tubal ligation|H/O: tubal ligation
C0438066|T033|OF|267020005|SNOMEDCT_CORE|History of - tubal ligation|H/O: tubal ligation
C0438066|T033|IS|267020005|SNOMEDCT_CORE|History of - tubal ligation|H/O: tubal ligation
C0438066|T033|FN|267020005|SNOMEDCT_CORE|History of tubal ligation|H/O: tubal ligation
C0438066|T033|SY|267020005|SNOMEDCT_CORE|History of tubal ligation|H/O: tubal ligation
C0438069|T033|OAP|161803004|SNOMEDCT_CORE|H/O: obstetric problem|H/O: obstetric problem
C0438069|T033|OF|161803004|SNOMEDCT_CORE|History of - obstetric problem|H/O: obstetric problem
C0438069|T033|IS|161803004|SNOMEDCT_CORE|History of - obstetric problem|H/O: obstetric problem
C0438069|T033|OAF|161803004|SNOMEDCT_CORE|History of obstetric problem|H/O: obstetric problem
C0438069|T033|OAS|161803004|SNOMEDCT_CORE|History of obstetric problem|H/O: obstetric problem
C0438076|T033|PT|161765003|SNOMEDCT_CORE|H/O: premature delivery|H/O: premature delivery
C0438076|T033|IS|161765003|SNOMEDCT_CORE|History of - premature delivery|H/O: premature delivery
C0438076|T033|OF|161765003|SNOMEDCT_CORE|History of - premature delivery|H/O: premature delivery
C0438076|T033|SY|161765003|SNOMEDCT_CORE|History of premature delivery|H/O: premature delivery
C0438076|T033|FN|161765003|SNOMEDCT_CORE|History of premature delivery|H/O: premature delivery
C0438076|T033|SY|161765003|SNOMEDCT_CORE|History of preterm delivery|H/O: premature delivery
C0438080|T033|PT|161744009|SNOMEDCT_CORE|H/O: miscarriage|H/O: miscarriage
C0438080|T033|OF|161744009|SNOMEDCT_CORE|History of - miscarriage|H/O: miscarriage
C0438080|T033|IS|161744009|SNOMEDCT_CORE|History of - miscarriage|H/O: miscarriage
C0438080|T033|FN|161744009|SNOMEDCT_CORE|History of miscarriage|H/O: miscarriage
C0438080|T033|SY|161744009|SNOMEDCT_CORE|History of miscarriage|H/O: miscarriage
C0438097|T033|SY|161811009|SNOMEDCT_CORE|H/O: perinatal death|H/O: perinatal fetal loss
C0438097|T033|PT|161811009|SNOMEDCT_CORE|H/O: perinatal fetal loss|H/O: perinatal fetal loss
C0438097|T033|SY|161811009|SNOMEDCT_CORE|H/O: perinatal foetal loss|H/O: perinatal fetal loss
C0438097|T033|OF|161811009|SNOMEDCT_CORE|History of - perinatal fetal loss|H/O: perinatal fetal loss
C0438097|T033|IS|161811009|SNOMEDCT_CORE|History of - perinatal fetal loss|H/O: perinatal fetal loss
C0438097|T033|SY|161811009|SNOMEDCT_CORE|History of - perinatal foetal loss|H/O: perinatal fetal loss
C0438097|T033|FN|161811009|SNOMEDCT_CORE|History of perinatal fetal loss|H/O: perinatal fetal loss
C0438097|T033|SY|161811009|SNOMEDCT_CORE|History of perinatal fetal loss|H/O: perinatal fetal loss
C0438142|T033|PT|171251002|SNOMEDCT_CORE|Urine screening abnormal|Urine screening abnormal
C0438142|T033|FN|171251002|SNOMEDCT_CORE|Urine screening abnormal|Urine screening abnormal
C0438228|T033|PT|165563002|SNOMEDCT_CORE|Coag./bleeding tests abnormal|Coag./bleeding tests abnormal
C0438228|T033|FN|165563002|SNOMEDCT_CORE|Coagulation/bleeding tests abnormal|Coag./bleeding tests abnormal
C0438228|T033|SY|165563002|SNOMEDCT_CORE|Coagulation/bleeding tests abnormal|Coag./bleeding tests abnormal
C0438237|T033|PT|166643006|SNOMEDCT_CORE|Liver enzymes abnormal|Liver enzymes abnormal
C0438237|T033|FN|166643006|SNOMEDCT_CORE|Liver enzymes abnormal|Liver enzymes abnormal
C0438258|T033|PT|166318006|SNOMEDCT_CORE|Blood chemistry abnormal|Blood chemistry abnormal
C0438258|T033|FN|166318006|SNOMEDCT_CORE|Blood chemistry abnormal|Blood chemistry abnormal
C0438623|T037|OAP|209410007|SNOMEDCT_CORE|Sprain of shoulder and upper arm|Sprain of shoulder and upper arm
C0438623|T037|OAF|209410007|SNOMEDCT_CORE|Sprain of shoulder and upper arm|Sprain of shoulder and upper arm
C0438623|T037|OAS|209410007|SNOMEDCT_CORE|Sprain shoulder and upper arm|Sprain of shoulder and upper arm
C0438624|T037|SY|367423000|SNOMEDCT_CORE|Bruise of eye|Contusion of eye
C0438624|T037|PT|367423000|SNOMEDCT_CORE|Contusion of eye|Contusion of eye
C0438624|T037|FN|367423000|SNOMEDCT_CORE|Contusion of eye|Contusion of eye
C0438624|T037|IS|367423000|SNOMEDCT_CORE|Contusion of eye, NOS|Contusion of eye
C0438638|T047|FN|282095007|SNOMEDCT_CORE|Allergic reaction caused by bee sting|Allergic reaction to bee sting
C0438638|T047|SY|282095007|SNOMEDCT_CORE|Allergic reaction caused by bee sting|Allergic reaction to bee sting
C0438638|T047|PT|282095007|SNOMEDCT_CORE|Allergic reaction to bee sting|Allergic reaction to bee sting
C0438638|T047|OF|282095007|SNOMEDCT_CORE|Allergic reaction to bee sting|Allergic reaction to bee sting
C0438716|T184|SY|23924001|SNOMEDCT_CORE|Pressure in chest|Pressure in chest
C0439032|T033|PT|272036004|SNOMEDCT_CORE|C/O - debility - malaise|C/O - debility - malaise
C0439032|T033|OF|272036004|SNOMEDCT_CORE|C/O - debility - malaise|C/O - debility - malaise
C0439032|T033|FN|272036004|SNOMEDCT_CORE|Complaining of debility and malaise|C/O - debility - malaise
C0439032|T033|SY|272036004|SNOMEDCT_CORE|Complaining of debility and malaise|C/O - debility - malaise
C0439044|T033|IS|105529008|SNOMEDCT_CORE|Home alone|Lives alone
C0439044|T033|PT|105529008|SNOMEDCT_CORE|Lives alone|Lives alone
C0439044|T033|FN|105529008|SNOMEDCT_CORE|Lives alone|Lives alone
C0439044|T033|IS|105529008|SNOMEDCT_CORE|Living alone|Lives alone
C0442874|T047|IS|42658009|SNOMEDCT_CORE|Neuropathy|Neuropathy
C0442874|T047|PT|386033004|SNOMEDCT_CORE|Neuropathy|Neuropathy
C0442874|T047|SY|386033004|SNOMEDCT_CORE|Neuropathy|Neuropathy
C0442874|T047|FN|386033004|SNOMEDCT_CORE|Neuropathy|Neuropathy
C0442874|T047|IS|42658009|SNOMEDCT_CORE|Neuropathy, NOS|Neuropathy
C0451641|T047|PT|95566004|SNOMEDCT_CORE|Urolithiasis|Urolithiasis
C0451641|T047|FN|95566004|SNOMEDCT_CORE|Urolithiasis|Urolithiasis
C0451641|T047|IS|95566004|SNOMEDCT_CORE|Urolithiasis, NOS|Urolithiasis
C0451664|T037|PT|212363007|SNOMEDCT_CORE|Injury of multiple nerves at shoulder and upper arm level|Injury of multiple nerves at shoulder and upper arm level
C0451664|T037|FN|212363007|SNOMEDCT_CORE|Injury of multiple nerves at shoulder and upper arm level|Injury of multiple nerves at shoulder and upper arm level
C0451674|T046|PT|195189003|SNOMEDCT_CORE|Cerebral infarction due to thrombosis of cerebral arteries|Cerebral infarction due to thrombosis of cerebral arteries
C0451674|T046|FN|195189003|SNOMEDCT_CORE|Cerebral infarction due to thrombosis of cerebral arteries|Cerebral infarction due to thrombosis of cerebral arteries
C0451675|T047|PT|195190007|SNOMEDCT_CORE|Cerebral infarction due to embolism of cerebral arteries|Cerebral infarction due to embolism of cerebral arteries
C0451675|T047|FN|195190007|SNOMEDCT_CORE|Cerebral infarction due to embolism of cerebral arteries|Cerebral infarction due to embolism of cerebral arteries
C0451718|T047|SY|197764002|SNOMEDCT_CORE|Chronic non-obstructive atrophic pyelonephritis|Non-obstructive reflux-associated chronic pyelonephritis
C0451718|T047|SY|197764002|SNOMEDCT_CORE|Nephropathy associated with vesicoureteral reflux|Non-obstructive reflux-associated chronic pyelonephritis
C0451718|T047|FN|197764002|SNOMEDCT_CORE|Non-obstructive reflux-associated chronic pyelonephritis|Non-obstructive reflux-associated chronic pyelonephritis
C0451718|T047|PT|197764002|SNOMEDCT_CORE|Non-obstructive reflux-associated chronic pyelonephritis|Non-obstructive reflux-associated chronic pyelonephritis
C0451718|T047|SY|197764002|SNOMEDCT_CORE|Reflux nephropathy|Non-obstructive reflux-associated chronic pyelonephritis
C0451718|T047|SY|197764002|SNOMEDCT_CORE|RN - Reflux nephropathy|Non-obstructive reflux-associated chronic pyelonephritis
C0451772|T046|SY|199111004|SNOMEDCT_CORE|Postpartum urinary tract infection|Urinary tract infection following delivery
C0451772|T046|PT|199111004|SNOMEDCT_CORE|Urinary tract infection following delivery|Urinary tract infection following delivery
C0451772|T046|FN|199111004|SNOMEDCT_CORE|Urinary tract infection following delivery|Urinary tract infection following delivery
C0451805|T033|PT|199734003|SNOMEDCT_CORE|Abnormal biochemical finding on antenatal screening of mother|Abnormal biochemical finding on antenatal screening of mother
C0451805|T033|OF|199734003|SNOMEDCT_CORE|Abnormal biochemical finding on antenatal screening of mother|Abnormal biochemical finding on antenatal screening of mother
C0451805|T033|FN|199734003|SNOMEDCT_CORE|Abnormal biochemical finding on antenatal screening of mother|Abnormal biochemical finding on antenatal screening of mother
C0451819|T047|SY|415530009|SNOMEDCT_CORE|Obesity due to excess calories|Simple obesity
C0451819|T047|PT|415530009|SNOMEDCT_CORE|Simple obesity|Simple obesity
C0451819|T047|FN|415530009|SNOMEDCT_CORE|Simple obesity|Simple obesity
C0451891|T037|PT|212454006|SNOMEDCT_CORE|Traumatic rupture of lumbar intervertebral disc|Traumatic rupture of lumbar intervertebral disc
C0451891|T037|FN|212454006|SNOMEDCT_CORE|Traumatic rupture of lumbar intervertebral disc|Traumatic rupture of lumbar intervertebral disc
C0451918|T037|PT|210773002|SNOMEDCT_CORE|Open wounds involving multiple regions of lower limb|Open wounds involving multiple regions of lower limb
C0451918|T037|FN|210773002|SNOMEDCT_CORE|Open wounds involving multiple regions of lower limb|Open wounds involving multiple regions of lower limb
C0452138|T047|PT|194424005|SNOMEDCT_CORE|Sensorineural hearing loss, bilateral|Sensorineural hearing loss, bilateral
C0452138|T047|OF|194424005|SNOMEDCT_CORE|Sensorineural hearing loss, bilateral|Sensorineural hearing loss, bilateral
C0452138|T047|FN|194424005|SNOMEDCT_CORE|Sensorineural hearing loss, bilateral|Sensorineural hearing loss, bilateral
C0452167|T046|PT|200125006|SNOMEDCT_CORE|Infection of obstetric surgical wound|Infection of obstetric surgical wound
C0452167|T046|FN|200125006|SNOMEDCT_CORE|Infection of obstetric surgical wound|Infection of obstetric surgical wound
C0452168|T019|PT|204891000|SNOMEDCT_CORE|Hypospadias, balanic|Hypospadias, balanic
C0452168|T019|FN|204891000|SNOMEDCT_CORE|Hypospadias, balanic|Hypospadias, balanic
C0452168|T019|SY|204891000|SNOMEDCT_CORE|Hypospadias, glandular|Hypospadias, balanic
C0452168|T019|IS|204891000|SNOMEDCT_CORE|Hypospadias, glanular|Hypospadias, balanic
C0452221|T047|PT|203241002|SNOMEDCT_CORE|Osteomyelitis of vertebra|Osteomyelitis of vertebra
C0452221|T047|FN|203241002|SNOMEDCT_CORE|Osteomyelitis of vertebra|Osteomyelitis of vertebra
C0454644|T033|PT|62415009|SNOMEDCT_CORE|Delayed articulatory and language development|Delayed articulatory and language development
C0454644|T033|FN|62415009|SNOMEDCT_CORE|Delayed articulatory and language development|Delayed articulatory and language development
C0454644|T033|SY|62415009|SNOMEDCT_CORE|Developmental language delay|Delayed articulatory and language development
C0455366|T033|OF|160302006|SNOMEDCT_CORE|Family history: Thyroid disorder|FH: Thyroid disorder
C0455366|T033|FN|160302006|SNOMEDCT_CORE|Family history: Thyroid disorder|FH: Thyroid disorder
C0455366|T033|SY|160302006|SNOMEDCT_CORE|Family history: Thyroid disorder|FH: Thyroid disorder
C0455366|T033|SY|160302006|SNOMEDCT_CORE|FH: Thyroid disease|FH: Thyroid disorder
C0455366|T033|PT|160302006|SNOMEDCT_CORE|FH: Thyroid disorder|FH: Thyroid disorder
C0455369|T033|OF|266887003|SNOMEDCT_CORE|Family history: Raised blood lipids|FH: Raised blood lipids
C0455369|T033|FN|266887003|SNOMEDCT_CORE|Family history: Raised blood lipids|FH: Raised blood lipids
C0455369|T033|SY|266887003|SNOMEDCT_CORE|Family history: Raised blood lipids|FH: Raised blood lipids
C0455369|T033|SY|266887003|SNOMEDCT_CORE|FH: Fats raised|FH: Raised blood lipids
C0455369|T033|PT|266887003|SNOMEDCT_CORE|FH: Raised blood lipids|FH: Raised blood lipids
C0455376|T033|SY|160316001|SNOMEDCT_CORE|Family history of blood disorder|FH: Blood disorder
C0455376|T033|SY|160316001|SNOMEDCT_CORE|Family history: Blood disorder|FH: Blood disorder
C0455376|T033|OF|160316001|SNOMEDCT_CORE|Family history: Blood disorder|FH: Blood disorder
C0455376|T033|FN|160316001|SNOMEDCT_CORE|Family history: Blood disorder|FH: Blood disorder
C0455376|T033|PT|160316001|SNOMEDCT_CORE|FH: Blood disorder|FH: Blood disorder
C0455397|T033|SY|160347007|SNOMEDCT_CORE|Family history of glaucoma|FH: Glaucoma
C0455397|T033|SY|160347007|SNOMEDCT_CORE|Family history: Glaucoma|FH: Glaucoma
C0455397|T033|OF|160347007|SNOMEDCT_CORE|Family history: Glaucoma|FH: Glaucoma
C0455397|T033|FN|160347007|SNOMEDCT_CORE|Family history: Glaucoma|FH: Glaucoma
C0455397|T033|PT|160347007|SNOMEDCT_CORE|FH: Glaucoma|FH: Glaucoma
C0455404|T033|SY|266894000|SNOMEDCT_CORE|Family history of cardiovascular disease|FH: Cardiovascular disease
C0455404|T033|SY|266894000|SNOMEDCT_CORE|Family history: Cardiovascular disease|FH: Cardiovascular disease
C0455404|T033|OF|266894000|SNOMEDCT_CORE|Family history: Cardiovascular disease|FH: Cardiovascular disease
C0455404|T033|FN|266894000|SNOMEDCT_CORE|Family history: Cardiovascular disease|FH: Cardiovascular disease
C0455404|T033|PT|266894000|SNOMEDCT_CORE|FH: Cardiovascular disease|FH: Cardiovascular disease
C0455404|T033|SY|266894000|SNOMEDCT_CORE|FH: CVS disorder|FH: Cardiovascular disease
C0455405|T033|SY|160357008|SNOMEDCT_CORE|Family history of hypertension|FH: Hypertension
C0455405|T033|SY|160357008|SNOMEDCT_CORE|Family history: Hypertension|FH: Hypertension
C0455405|T033|OF|160357008|SNOMEDCT_CORE|Family history: Hypertension|FH: Hypertension
C0455405|T033|FN|160357008|SNOMEDCT_CORE|Family history: Hypertension|FH: Hypertension
C0455405|T033|PT|160357008|SNOMEDCT_CORE|FH: Hypertension|FH: Hypertension
C0455420|T033|SY|160381001|SNOMEDCT_CORE|Family history of gastrointestinal disease|FH: Gastrointestinal disease
C0455420|T033|SY|160381001|SNOMEDCT_CORE|Family history: Gastrointestinal disease|FH: Gastrointestinal disease
C0455420|T033|OF|160381001|SNOMEDCT_CORE|Family history: Gastrointestinal disease|FH: Gastrointestinal disease
C0455420|T033|FN|160381001|SNOMEDCT_CORE|Family history: Gastrointestinal disease|FH: Gastrointestinal disease
C0455420|T033|PT|160381001|SNOMEDCT_CORE|FH: Gastrointestinal disease|FH: Gastrointestinal disease
C0455425|T033|SY|160392000|SNOMEDCT_CORE|Family history of breast disorder|FH: Breast disease
C0455425|T033|OF|160392000|SNOMEDCT_CORE|Family history: Breast disease|FH: Breast disease
C0455425|T033|FN|160392000|SNOMEDCT_CORE|Family history: Breast disease|FH: Breast disease
C0455425|T033|SY|160392000|SNOMEDCT_CORE|Family history: Breast disease|FH: Breast disease
C0455425|T033|PT|160392000|SNOMEDCT_CORE|FH: Breast disease|FH: Breast disease
C0455434|T033|OF|160402005|SNOMEDCT_CORE|Family history: Diabetes in pregnancy|FH: Diabetes in pregnancy
C0455434|T033|FN|160402005|SNOMEDCT_CORE|Family history: Diabetes in pregnancy|FH: Diabetes in pregnancy
C0455434|T033|SY|160402005|SNOMEDCT_CORE|Family history: Diabetes in pregnancy|FH: Diabetes in pregnancy
C0455434|T033|PT|160402005|SNOMEDCT_CORE|FH: Diabetes in pregnancy|FH: Diabetes in pregnancy
C0455453|T033|SY|160469004|SNOMEDCT_CORE|Family history of allergy|FH: Allergy
C0455453|T033|SY|160469004|SNOMEDCT_CORE|Family history: Allergy|FH: Allergy
C0455453|T033|OF|160469004|SNOMEDCT_CORE|Family history: Allergy|FH: Allergy
C0455453|T033|FN|160469004|SNOMEDCT_CORE|Family history: Allergy|FH: Allergy
C0455453|T033|PT|160469004|SNOMEDCT_CORE|FH: Allergy|FH: Allergy
C0455457|T033|OF|160474007|SNOMEDCT_CORE|Family history: Atopy|FH: Atopy
C0455457|T033|FN|160474007|SNOMEDCT_CORE|Family history: Atopy|FH: Atopy
C0455457|T033|SY|160474007|SNOMEDCT_CORE|Family history: Atopy|FH: Atopy
C0455457|T033|PT|160474007|SNOMEDCT_CORE|FH: Atopy|FH: Atopy
C0455460|T033|PT|161414005|SNOMEDCT_CORE|H/O: tuberculosis|H/O: tuberculosis
C0455460|T033|OF|161414005|SNOMEDCT_CORE|History of - tuberculosis|H/O: tuberculosis
C0455460|T033|IS|161414005|SNOMEDCT_CORE|History of - tuberculosis|H/O: tuberculosis
C0455460|T033|FN|161414005|SNOMEDCT_CORE|History of tuberculosis|H/O: tuberculosis
C0455460|T033|SY|161414005|SNOMEDCT_CORE|History of tuberculosis|H/O: tuberculosis
C0455461|T033|PT|161415006|SNOMEDCT_CORE|H/O: poliomyelitis|H/O: poliomyelitis
C0455461|T033|OF|161415006|SNOMEDCT_CORE|History of - poliomyelitis|H/O: poliomyelitis
C0455461|T033|IS|161415006|SNOMEDCT_CORE|History of - poliomyelitis|H/O: poliomyelitis
C0455461|T033|FN|161415006|SNOMEDCT_CORE|History of poliomyelitis|H/O: poliomyelitis
C0455461|T033|SY|161415006|SNOMEDCT_CORE|History of poliomyelitis|H/O: poliomyelitis
C0455462|T033|PT|161416007|SNOMEDCT_CORE|H/O: malaria|H/O: malaria
C0455462|T033|OF|161416007|SNOMEDCT_CORE|History of - malaria|H/O: malaria
C0455462|T033|IS|161416007|SNOMEDCT_CORE|History of - malaria|H/O: malaria
C0455462|T033|FN|161416007|SNOMEDCT_CORE|History of malaria|H/O: malaria
C0455462|T033|SY|161416007|SNOMEDCT_CORE|History of malaria|H/O: malaria
C0455469|T033|PT|161423008|SNOMEDCT_CORE|H/O: chickenpox|H/O: chickenpox
C0455469|T033|OF|161423008|SNOMEDCT_CORE|History of - chickenpox|H/O: chickenpox
C0455469|T033|IS|161423008|SNOMEDCT_CORE|History of - chickenpox|H/O: chickenpox
C0455469|T033|FN|161423008|SNOMEDCT_CORE|History of chickenpox|H/O: chickenpox
C0455469|T033|SY|161423008|SNOMEDCT_CORE|History of chickenpox|H/O: chickenpox
C0455486|T033|PT|161443002|SNOMEDCT_CORE|H/O: hypothyroidism|H/O: hypothyroidism
C0455486|T033|OF|161443002|SNOMEDCT_CORE|History of - hypothyroidism|H/O: hypothyroidism
C0455486|T033|IS|161443002|SNOMEDCT_CORE|History of - hypothyroidism|H/O: hypothyroidism
C0455486|T033|FN|161443002|SNOMEDCT_CORE|History of hypothyroidism|H/O: hypothyroidism
C0455486|T033|SY|161443002|SNOMEDCT_CORE|History of hypothyroidism|H/O: hypothyroidism
C0455488|T033|PT|161445009|SNOMEDCT_CORE|H/O: diabetes mellitus|H/O: diabetes mellitus
C0455488|T033|OF|161445009|SNOMEDCT_CORE|History of - diabetes mellitus|H/O: diabetes mellitus
C0455488|T033|IS|161445009|SNOMEDCT_CORE|History of - diabetes mellitus|H/O: diabetes mellitus
C0455488|T033|FN|161445009|SNOMEDCT_CORE|History of diabetes mellitus|H/O: diabetes mellitus
C0455488|T033|SY|161445009|SNOMEDCT_CORE|History of diabetes mellitus|H/O: diabetes mellitus
C0455488|T033|SY|161445009|SNOMEDCT_CORE|Pre-existing diabetes mellitus|H/O: diabetes mellitus
C0455491|T033|PT|161450003|SNOMEDCT_CORE|H/O: raised blood lipids|H/O: raised blood lipids
C0455491|T033|OF|161450003|SNOMEDCT_CORE|History of - raised blood lipids|H/O: raised blood lipids
C0455491|T033|IS|161450003|SNOMEDCT_CORE|History of - raised blood lipids|H/O: raised blood lipids
C0455491|T033|FN|161450003|SNOMEDCT_CORE|History of raised blood lipids|H/O: raised blood lipids
C0455491|T033|SY|161450003|SNOMEDCT_CORE|History of raised blood lipids|H/O: raised blood lipids
C0455492|T033|PT|161451004|SNOMEDCT_CORE|H/O: gout|H/O: gout
C0455492|T033|OF|161451004|SNOMEDCT_CORE|History of - gout|H/O: gout
C0455492|T033|IS|161451004|SNOMEDCT_CORE|History of - gout|H/O: gout
C0455492|T033|FN|161451004|SNOMEDCT_CORE|History of gout|H/O: gout
C0455492|T033|SY|161451004|SNOMEDCT_CORE|History of gout|H/O: gout
C0455500|T033|PT|161466001|SNOMEDCT_CORE|H/O: alcoholism|H/O: alcoholism
C0455500|T033|OF|161466001|SNOMEDCT_CORE|History of - alcoholism|H/O: alcoholism
C0455500|T033|IS|161466001|SNOMEDCT_CORE|History of - alcoholism|H/O: alcoholism
C0455500|T033|FN|161466001|SNOMEDCT_CORE|History of alcoholism|H/O: alcoholism
C0455500|T033|SY|161466001|SNOMEDCT_CORE|History of alcoholism|H/O: alcoholism
C0455502|T033|PT|161468000|SNOMEDCT_CORE|H/O: schizophrenia|H/O: schizophrenia
C0455502|T033|OF|161468000|SNOMEDCT_CORE|History of - schizophrenia|H/O: schizophrenia
C0455502|T033|IS|161468000|SNOMEDCT_CORE|History of - schizophrenia|H/O: schizophrenia
C0455502|T033|FN|161468000|SNOMEDCT_CORE|History of schizophrenia|H/O: schizophrenia
C0455502|T033|SY|161468000|SNOMEDCT_CORE|History of schizophrenia|H/O: schizophrenia
C0455503|T033|PT|161469008|SNOMEDCT_CORE|H/O: depression|H/O: depression
C0455503|T033|SY|161469008|SNOMEDCT_CORE|Has had depression|H/O: depression
C0455503|T033|OF|161469008|SNOMEDCT_CORE|History of - depression|H/O: depression
C0455503|T033|IS|161469008|SNOMEDCT_CORE|History of - depression|H/O: depression
C0455503|T033|FN|161469008|SNOMEDCT_CORE|History of depression|H/O: depression
C0455503|T033|SY|161469008|SNOMEDCT_CORE|History of depression|H/O: depression
C0455503|T033|SY|161469008|SNOMEDCT_CORE|History of depressive disorder|H/O: depression
C0455514|T033|PT|161483005|SNOMEDCT_CORE|H/O: Bell's palsy|H/O: Bell's palsy
C0455514|T033|IS|161483005|SNOMEDCT_CORE|History of - Bell palsy|H/O: Bell's palsy
C0455514|T033|OF|161483005|SNOMEDCT_CORE|History of - Bell's palsy|H/O: Bell's palsy
C0455514|T033|IS|161483005|SNOMEDCT_CORE|History of - Bell's palsy|H/O: Bell's palsy
C0455514|T033|SY|161483005|SNOMEDCT_CORE|History of Bell palsy|H/O: Bell's palsy
C0455514|T033|FN|161483005|SNOMEDCT_CORE|History of Bell's palsy|H/O: Bell's palsy
C0455514|T033|SY|161483005|SNOMEDCT_CORE|History of Bell's palsy|H/O: Bell's palsy
C0455527|T033|PT|161501007|SNOMEDCT_CORE|H/O: hypertension|H/O: hypertension
C0455527|T033|OF|161501007|SNOMEDCT_CORE|History of - hypertension|H/O: hypertension
C0455527|T033|IS|161501007|SNOMEDCT_CORE|History of - hypertension|H/O: hypertension
C0455527|T033|FN|161501007|SNOMEDCT_CORE|History of hypertension|H/O: hypertension
C0455527|T033|SY|161501007|SNOMEDCT_CORE|History of hypertension|H/O: hypertension
C0455531|T033|PT|161505003|SNOMEDCT_CORE|H/O: heart failure|H/O: heart failure
C0455531|T033|OF|161505003|SNOMEDCT_CORE|History of - heart failure|H/O: heart failure
C0455531|T033|IS|161505003|SNOMEDCT_CORE|History of - heart failure|H/O: heart failure
C0455531|T033|FN|161505003|SNOMEDCT_CORE|History of heart failure|H/O: heart failure
C0455531|T033|SY|161505003|SNOMEDCT_CORE|History of heart failure|H/O: heart failure
C0455536|T033|OP|161511000|SNOMEDCT_CORE|H/O: TIA|History of transient ischemic attack
C0455536|T033|OF|161511000|SNOMEDCT_CORE|History of - TIA|History of transient ischemic attack
C0455536|T033|IS|161511000|SNOMEDCT_CORE|History of - transient ischemic attack|History of transient ischemic attack
C0455536|T033|OF|161511000|SNOMEDCT_CORE|History of - transient ischemic attack|History of transient ischemic attack
C0455536|T033|PTGB|161511000|SNOMEDCT_CORE|History of transient ischaemic attack|History of transient ischemic attack
C0455536|T033|PT|161511000|SNOMEDCT_CORE|History of transient ischemic attack|History of transient ischemic attack
C0455536|T033|FN|161511000|SNOMEDCT_CORE|History of transient ischemic attack|History of transient ischemic attack
C0455537|T033|PT|161512007|SNOMEDCT_CORE|H/O: pulmonary embolus|H/O: pulmonary embolus
C0455537|T033|OF|161512007|SNOMEDCT_CORE|History of - pulmonary embolus|H/O: pulmonary embolus
C0455537|T033|IS|161512007|SNOMEDCT_CORE|History of - pulmonary embolus|H/O: pulmonary embolus
C0455537|T033|FN|161512007|SNOMEDCT_CORE|History of pulmonary embolus|H/O: pulmonary embolus
C0455537|T033|SY|161512007|SNOMEDCT_CORE|History of pulmonary embolus|H/O: pulmonary embolus
C0455539|T033|PT|266995000|SNOMEDCT_CORE|H/O: cardiovascular disease|H/O: cardiovascular disease
C0455539|T033|OF|266995000|SNOMEDCT_CORE|History of - cardiovascular disease|H/O: cardiovascular disease
C0455539|T033|IS|266995000|SNOMEDCT_CORE|History of - cardiovascular disease|H/O: cardiovascular disease
C0455539|T033|FN|266995000|SNOMEDCT_CORE|History of cardiovascular disease|H/O: cardiovascular disease
C0455539|T033|SY|266995000|SNOMEDCT_CORE|History of cardiovascular disease|H/O: cardiovascular disease
C0455539|T033|SY|266995000|SNOMEDCT_CORE|History of circulatory system disease|H/O: cardiovascular disease
C0455540|T033|PT|161523006|SNOMEDCT_CORE|H/O: respiratory disease|H/O: respiratory disease
C0455540|T033|IS|161523006|SNOMEDCT_CORE|History of - respiratory disease|H/O: respiratory disease
C0455540|T033|OF|161523006|SNOMEDCT_CORE|History of - respiratory disease|H/O: respiratory disease
C0455540|T033|SY|161523006|SNOMEDCT_CORE|History of respiratory disease|H/O: respiratory disease
C0455540|T033|FN|161523006|SNOMEDCT_CORE|History of respiratory disease|H/O: respiratory disease
C0455542|T033|PT|161525004|SNOMEDCT_CORE|H/O: pneumonia|H/O: pneumonia
C0455542|T033|OF|161525004|SNOMEDCT_CORE|History of - pneumonia|H/O: pneumonia
C0455542|T033|IS|161525004|SNOMEDCT_CORE|History of - pneumonia|H/O: pneumonia
C0455542|T033|FN|161525004|SNOMEDCT_CORE|History of pneumonia|H/O: pneumonia
C0455542|T033|SY|161525004|SNOMEDCT_CORE|History of pneumonia|H/O: pneumonia
C0455546|T033|PT|266998003|SNOMEDCT_CORE|H/O: peptic ulcer|H/O: peptic ulcer
C0455546|T033|OF|266998003|SNOMEDCT_CORE|History of - peptic ulcer|H/O: peptic ulcer
C0455546|T033|IS|266998003|SNOMEDCT_CORE|History of - peptic ulcer|H/O: peptic ulcer
C0455546|T033|FN|266998003|SNOMEDCT_CORE|History of peptic ulcer|H/O: peptic ulcer
C0455546|T033|SY|266998003|SNOMEDCT_CORE|History of peptic ulcer|H/O: peptic ulcer
C0455553|T033|PT|266997008|SNOMEDCT_CORE|H/O: gastrointestinal disease|H/O: gastrointestinal disease
C0455553|T033|OF|266997008|SNOMEDCT_CORE|History of - gastrointestinal disease|H/O: gastrointestinal disease
C0455553|T033|IS|266997008|SNOMEDCT_CORE|History of - gastrointestinal disease|H/O: gastrointestinal disease
C0455553|T033|FN|266997008|SNOMEDCT_CORE|History of gastrointestinal disease|H/O: gastrointestinal disease
C0455553|T033|SY|266997008|SNOMEDCT_CORE|History of gastrointestinal disease|H/O: gastrointestinal disease
C0455557|T033|PT|161548009|SNOMEDCT_CORE|H/O: urinary stone|H/O: urinary stone
C0455557|T033|OF|161548009|SNOMEDCT_CORE|History of - urinary stone|H/O: urinary stone
C0455557|T033|IS|161548009|SNOMEDCT_CORE|History of - urinary stone|H/O: urinary stone
C0455557|T033|FN|161548009|SNOMEDCT_CORE|History of urinary stone|H/O: urinary stone
C0455557|T033|SY|161548009|SNOMEDCT_CORE|History of urinary stone|H/O: urinary stone
C0455557|T033|SY|161548009|SNOMEDCT_CORE|History of urinary tract calculus|H/O: urinary stone
C0455564|T033|PT|161558008|SNOMEDCT_CORE|H/O: vasectomy|H/O: vasectomy
C0455564|T033|OF|161558008|SNOMEDCT_CORE|History of - vasectomy|H/O: vasectomy
C0455564|T033|IS|161558008|SNOMEDCT_CORE|History of - vasectomy|H/O: vasectomy
C0455564|T033|FN|161558008|SNOMEDCT_CORE|History of vasectomy|H/O: vasectomy
C0455564|T033|SY|161558008|SNOMEDCT_CORE|History of vasectomy|H/O: vasectomy
C0455581|T033|PT|161579008|SNOMEDCT_CORE|H/O: perinatal problem|H/O: perinatal problem
C0455581|T033|OF|161579008|SNOMEDCT_CORE|History of - perinatal problem|H/O: perinatal problem
C0455581|T033|IS|161579008|SNOMEDCT_CORE|History of - perinatal problem|H/O: perinatal problem
C0455581|T033|SY|161579008|SNOMEDCT_CORE|History of perinatal problem|H/O: perinatal problem
C0455581|T033|FN|161579008|SNOMEDCT_CORE|History of perinatal problem|H/O: perinatal problem
C0455586|T033|PT|161586000|SNOMEDCT_CORE|H/O: injury|H/O: injury
C0455586|T033|OF|161586000|SNOMEDCT_CORE|History of - injury|H/O: injury
C0455586|T033|IS|161586000|SNOMEDCT_CORE|History of - injury|H/O: injury
C0455586|T033|SY|161586000|SNOMEDCT_CORE|History of injury|H/O: injury
C0455586|T033|FN|161586000|SNOMEDCT_CORE|History of injury|H/O: injury
C0455587|T033|PT|161587009|SNOMEDCT_CORE|H/O: head injury|H/O: head injury
C0455587|T033|OF|161587009|SNOMEDCT_CORE|History of - head injury|H/O: head injury
C0455587|T033|IS|161587009|SNOMEDCT_CORE|History of - head injury|H/O: head injury
C0455587|T033|FN|161587009|SNOMEDCT_CORE|History of head injury|H/O: head injury
C0455587|T033|SY|161587009|SNOMEDCT_CORE|History of head injury|H/O: head injury
C0455589|T033|OAP|161590003|SNOMEDCT_CORE|H/O: drug allergy|H/O: drug allergy
C0455589|T033|OF|161590003|SNOMEDCT_CORE|History of - drug allergy|H/O: drug allergy
C0455589|T033|IS|161590003|SNOMEDCT_CORE|History of - drug allergy|H/O: drug allergy
C0455589|T033|OAS|161590003|SNOMEDCT_CORE|History of drug allergy|H/O: drug allergy
C0455589|T033|OAF|161590003|SNOMEDCT_CORE|History of drug allergy|H/O: drug allergy
C0455590|T033|OAP|161591004|SNOMEDCT_CORE|H/O: penicillin allergy|H/O: penicillin allergy
C0455590|T033|OF|161591004|SNOMEDCT_CORE|History of - penicillin allergy|H/O: penicillin allergy
C0455590|T033|IS|161591004|SNOMEDCT_CORE|History of - penicillin allergy|H/O: penicillin allergy
C0455590|T033|OAS|161591004|SNOMEDCT_CORE|History of penicillin allergy|H/O: penicillin allergy
C0455590|T033|OAF|161591004|SNOMEDCT_CORE|History of penicillin allergy|H/O: penicillin allergy
C0455607|T033|OAP|161612000|SNOMEDCT_CORE|H/O: food allergy|H/O: food allergy
C0455607|T033|IS|161612000|SNOMEDCT_CORE|History of - food allergy|H/O: food allergy
C0455607|T033|OF|161612000|SNOMEDCT_CORE|History of - food allergy|H/O: food allergy
C0455607|T033|OAS|161612000|SNOMEDCT_CORE|History of food allergy|H/O: food allergy
C0455607|T033|OAF|161612000|SNOMEDCT_CORE|History of food allergy|H/O: food allergy
C0455610|T033|SY|161615003|SNOMEDCT_CORE|H/O: operation|H/O: surgery
C0455610|T033|PT|161615003|SNOMEDCT_CORE|H/O: surgery|H/O: surgery
C0455610|T033|OF|161615003|SNOMEDCT_CORE|History of - surgery|H/O: surgery
C0455610|T033|SY|161615003|SNOMEDCT_CORE|History of - surgery|H/O: surgery
C0455610|T033|SY|161615003|SNOMEDCT_CORE|History of surgery|H/O: surgery
C0455610|T033|FN|161615003|SNOMEDCT_CORE|History of surgery|H/O: surgery
C0455610|T033|IS|161615003|SNOMEDCT_CORE|Past surgical history of|H/O: surgery
C0455616|T033|PT|161622006|SNOMEDCT_CORE|H/O: lower limb amputation|H/O: lower limb amputation
C0455616|T033|OF|161622006|SNOMEDCT_CORE|History of - lower limb amputation|H/O: lower limb amputation
C0455616|T033|IS|161622006|SNOMEDCT_CORE|History of - lower limb amputation|H/O: lower limb amputation
C0455616|T033|FN|161622006|SNOMEDCT_CORE|History of lower limb amputation|H/O: lower limb amputation
C0455616|T033|SY|161622006|SNOMEDCT_CORE|History of lower limb amputation|H/O: lower limb amputation
C0455620|T033|PT|161633009|SNOMEDCT_CORE|H/O: radiation exposure|H/O: radiation exposure
C0455620|T033|IS|161633009|SNOMEDCT_CORE|History of - radiation exposure|H/O: radiation exposure
C0455620|T033|OF|161633009|SNOMEDCT_CORE|History of - radiation exposure|H/O: radiation exposure
C0455620|T033|SY|161633009|SNOMEDCT_CORE|History of irradiation|H/O: radiation exposure
C0455620|T033|SY|161633009|SNOMEDCT_CORE|History of radiation exposure|H/O: radiation exposure
C0455620|T033|FN|161633009|SNOMEDCT_CORE|History of radiation exposure|H/O: radiation exposure
C0455636|T033|PT|161659007|SNOMEDCT_CORE|H/O: kidney donation|H/O: kidney donation
C0455636|T033|OF|161659007|SNOMEDCT_CORE|History of - kidney donation|H/O: kidney donation
C0455636|T033|IS|161659007|SNOMEDCT_CORE|History of - kidney donation|H/O: kidney donation
C0455636|T033|FN|161659007|SNOMEDCT_CORE|History of kidney donation|H/O: kidney donation
C0455636|T033|SY|161659007|SNOMEDCT_CORE|History of kidney donation|H/O: kidney donation
C0455641|T033|SY|161665007|SNOMEDCT_CORE|H/O: kidney recipient|History of renal transplant
C0455641|T033|OF|161665007|SNOMEDCT_CORE|History of - kidney recipient|History of renal transplant
C0455641|T033|SY|161665007|SNOMEDCT_CORE|History of - kidney recipient|History of renal transplant
C0455641|T033|PT|161665007|SNOMEDCT_CORE|History of renal transplant|History of renal transplant
C0455641|T033|FN|161665007|SNOMEDCT_CORE|History of renal transplant|History of renal transplant
C0455642|T033|PT|161666008|SNOMEDCT_CORE|H/O: heart recipient|H/O: heart recipient
C0455642|T033|OF|161666008|SNOMEDCT_CORE|History of - heart recipient|H/O: heart recipient
C0455642|T033|IS|161666008|SNOMEDCT_CORE|History of - heart recipient|H/O: heart recipient
C0455642|T033|FN|161666008|SNOMEDCT_CORE|History of heart recipient|H/O: heart recipient
C0455642|T033|SY|161666008|SNOMEDCT_CORE|History of heart recipient|H/O: heart recipient
C0455646|T033|PT|161670000|SNOMEDCT_CORE|H/O: cornea recipient|H/O: cornea recipient
C0455646|T033|OF|161670000|SNOMEDCT_CORE|History of - cornea recipient|H/O: cornea recipient
C0455646|T033|IS|161670000|SNOMEDCT_CORE|History of - cornea recipient|H/O: cornea recipient
C0455646|T033|FN|161670000|SNOMEDCT_CORE|History of cornea recipient|H/O: cornea recipient
C0455646|T033|SY|161670000|SNOMEDCT_CORE|History of cornea recipient|H/O: cornea recipient
C0455647|T033|PT|161671001|SNOMEDCT_CORE|H/O: liver recipient|H/O: liver recipient
C0455647|T033|IS|161671001|SNOMEDCT_CORE|History of - liver recipient|H/O: liver recipient
C0455647|T033|OF|161671001|SNOMEDCT_CORE|History of - liver recipient|H/O: liver recipient
C0455647|T033|SY|161671001|SNOMEDCT_CORE|History of liver recipient|H/O: liver recipient
C0455647|T033|FN|161671001|SNOMEDCT_CORE|History of liver recipient|H/O: liver recipient
C0455650|T033|PT|161675005|SNOMEDCT_CORE|H/O: artificial eyeglobe|H/O: artificial eyeglobe
C0455650|T033|OF|161675005|SNOMEDCT_CORE|History of - artificial eyeglobe|H/O: artificial eyeglobe
C0455650|T033|IS|161675005|SNOMEDCT_CORE|History of - artificial eyeglobe|H/O: artificial eyeglobe
C0455650|T033|FN|161675005|SNOMEDCT_CORE|History of artificial eyeglobe|H/O: artificial eyeglobe
C0455650|T033|SY|161675005|SNOMEDCT_CORE|History of artificial eyeglobe|H/O: artificial eyeglobe
C0455652|T033|PT|161677002|SNOMEDCT_CORE|H/O: artificial heart valve|H/O: artificial heart valve
C0455652|T033|OF|161677002|SNOMEDCT_CORE|History of - artificial heart valve|H/O: artificial heart valve
C0455652|T033|IS|161677002|SNOMEDCT_CORE|History of - artificial heart valve|H/O: artificial heart valve
C0455652|T033|FN|161677002|SNOMEDCT_CORE|History of artificial heart valve|H/O: artificial heart valve
C0455652|T033|SY|161677002|SNOMEDCT_CORE|History of artificial heart valve|H/O: artificial heart valve
C0455654|T033|PT|161679004|SNOMEDCT_CORE|H/O: artificial joint|H/O: artificial joint
C0455654|T033|OF|161679004|SNOMEDCT_CORE|History of - artificial joint|H/O: artificial joint
C0455654|T033|IS|161679004|SNOMEDCT_CORE|History of - artificial joint|H/O: artificial joint
C0455654|T033|FN|161679004|SNOMEDCT_CORE|History of artificial joint|H/O: artificial joint
C0455654|T033|SY|161679004|SNOMEDCT_CORE|History of artificial joint|H/O: artificial joint
C0455660|T033|PT|161685006|SNOMEDCT_CORE|H/O: tracheostomy|H/O: tracheostomy
C0455660|T033|OF|161685006|SNOMEDCT_CORE|History of - tracheostomy|H/O: tracheostomy
C0455660|T033|IS|161685006|SNOMEDCT_CORE|History of - tracheostomy|H/O: tracheostomy
C0455660|T033|FN|161685006|SNOMEDCT_CORE|History of tracheostomy|H/O: tracheostomy
C0455660|T033|SY|161685006|SNOMEDCT_CORE|History of tracheostomy|H/O: tracheostomy
C0455661|T033|PT|161686007|SNOMEDCT_CORE|H/O: ileostomy|H/O: ileostomy
C0455661|T033|OF|161686007|SNOMEDCT_CORE|History of - ileostomy|H/O: ileostomy
C0455661|T033|IS|161686007|SNOMEDCT_CORE|History of - ileostomy|H/O: ileostomy
C0455661|T033|FN|161686007|SNOMEDCT_CORE|History of ileostomy|H/O: ileostomy
C0455661|T033|SY|161686007|SNOMEDCT_CORE|History of ileostomy|H/O: ileostomy
C0455662|T033|PT|161687003|SNOMEDCT_CORE|H/O: colostomy|H/O: colostomy
C0455662|T033|OF|161687003|SNOMEDCT_CORE|History of - colostomy|H/O: colostomy
C0455662|T033|IS|161687003|SNOMEDCT_CORE|History of - colostomy|H/O: colostomy
C0455662|T033|FN|161687003|SNOMEDCT_CORE|History of colostomy|H/O: colostomy
C0455662|T033|SY|161687003|SNOMEDCT_CORE|History of colostomy|H/O: colostomy
C0455664|T033|PT|161689000|SNOMEDCT_CORE|H/O: gastrostomy|H/O: gastrostomy
C0455664|T033|OF|161689000|SNOMEDCT_CORE|History of - gastrostomy|H/O: gastrostomy
C0455664|T033|IS|161689000|SNOMEDCT_CORE|History of - gastrostomy|H/O: gastrostomy
C0455664|T033|FN|161689000|SNOMEDCT_CORE|History of gastrostomy|H/O: gastrostomy
C0455664|T033|SY|161689000|SNOMEDCT_CORE|History of gastrostomy|H/O: gastrostomy
C0455667|T033|SY|161693006|SNOMEDCT_CORE|H/O: kidney dialysis|H/O: renal dialysis
C0455667|T033|PT|161693006|SNOMEDCT_CORE|H/O: renal dialysis|H/O: renal dialysis
C0455667|T033|OF|161693006|SNOMEDCT_CORE|History of - renal dialysis|H/O: renal dialysis
C0455667|T033|IS|161693006|SNOMEDCT_CORE|History of - renal dialysis|H/O: renal dialysis
C0455667|T033|FN|161693006|SNOMEDCT_CORE|History of renal dialysis|H/O: renal dialysis
C0455667|T033|SY|161693006|SNOMEDCT_CORE|History of renal dialysis|H/O: renal dialysis
C0455669|T033|OP|267010000|SNOMEDCT_CORE|H/O: GIT bypass/anastomosis|History of gastrointestinal tract bypass
C0455669|T033|OF|267010000|SNOMEDCT_CORE|History of - gastrointestinal tract bypass/anastomosis|History of gastrointestinal tract bypass
C0455669|T033|IS|267010000|SNOMEDCT_CORE|History of - gastrointestinal tract bypass/anastomosis|History of gastrointestinal tract bypass
C0455669|T033|SY|267010000|SNOMEDCT_CORE|History of gastrointestinal tract anastomosis|History of gastrointestinal tract bypass
C0455669|T033|PT|267010000|SNOMEDCT_CORE|History of gastrointestinal tract bypass|History of gastrointestinal tract bypass
C0455669|T033|FN|267010000|SNOMEDCT_CORE|History of gastrointestinal tract bypass|History of gastrointestinal tract bypass
C0455669|T033|OF|267010000|SNOMEDCT_CORE|History of gastrointestinal tract bypass/anastomosis|History of gastrointestinal tract bypass
C0455669|T033|IS|267010000|SNOMEDCT_CORE|History of gastrointestinal tract bypass/anastomosis|History of gastrointestinal tract bypass
C0455693|T033|PT|275563002|SNOMEDCT_CORE|H/O: bone marrow donation|H/O: bone marrow donation
C0455693|T033|OF|275563002|SNOMEDCT_CORE|History of - bone marrow donation|H/O: bone marrow donation
C0455693|T033|IS|275563002|SNOMEDCT_CORE|History of - bone marrow donation|H/O: bone marrow donation
C0455693|T033|FN|275563002|SNOMEDCT_CORE|History of bone marrow donation|H/O: bone marrow donation
C0455693|T033|SY|275563002|SNOMEDCT_CORE|History of bone marrow donation|H/O: bone marrow donation
C0455899|T033|IS|126662008|SNOMEDCT_CORE|Erythema of mucous membrane of oropharynx|Red throat
C0455899|T033|PT|126662008|SNOMEDCT_CORE|Red throat|Red throat
C0455899|T033|FN|126662008|SNOMEDCT_CORE|Red throat|Red throat
C0456003|T047|PT|68550008|SNOMEDCT_CORE|Disturbance of temperature regulation of newborn|Disturbance of temperature regulation of newborn
C0456003|T047|FN|68550008|SNOMEDCT_CORE|Disturbance of temperature regulation of newborn|Disturbance of temperature regulation of newborn
C0456003|T047|IS|68550008|SNOMEDCT_CORE|Disturbance of temperature regulation of newborn, NOS|Disturbance of temperature regulation of newborn
C0456003|T047|SY|68550008|SNOMEDCT_CORE|Perinatal disorders of temperature regulation|Disturbance of temperature regulation of newborn
C0456058|T047|PT|276603001|SNOMEDCT_CORE|Perinatal disorder of growth and/or development|Perinatal disorder of growth and/or development
C0456058|T047|FN|276603001|SNOMEDCT_CORE|Perinatal disorder of growth and/or development|Perinatal disorder of growth and/or development
C0456058|T047|OP|276603001|SNOMEDCT_CORE|Perinatal disorders of growth and development|Perinatal disorder of growth and/or development
C0456058|T047|OF|276603001|SNOMEDCT_CORE|Perinatal disorders of growth and development|Perinatal disorder of growth and/or development
C0456070|T046|OAP|276617005|SNOMEDCT_CORE|Growth delay|Growth delay
C0456070|T046|OAF|276617005|SNOMEDCT_CORE|Growth delay|Growth delay
C0456091|T033|SY|199616008|SNOMEDCT_CORE|Accelerated fetal growth|Large for gestation age fetus
C0456091|T033|SY|199616008|SNOMEDCT_CORE|Accelerated foetal growth|Large for gestation age fetus
C0456091|T033|SY|199616008|SNOMEDCT_CORE|Fetal growth acceleration|Large for gestation age fetus
C0456091|T033|SY|199616008|SNOMEDCT_CORE|Foetal growth acceleration|Large for gestation age fetus
C0456091|T033|PT|199616008|SNOMEDCT_CORE|Large for gestation age fetus|Large for gestation age fetus
C0456091|T033|SY|199616008|SNOMEDCT_CORE|Large for gestation age foetus|Large for gestation age fetus
C0456091|T033|SY|199616008|SNOMEDCT_CORE|Large for gestational dates|Large for gestation age fetus
C0456091|T033|SY|199616008|SNOMEDCT_CORE|Large-for-dates fetus|Large for gestation age fetus
C0456091|T033|FN|199616008|SNOMEDCT_CORE|Large-for-dates fetus|Large for gestation age fetus
C0456091|T033|SY|199616008|SNOMEDCT_CORE|Large-for-dates foetus|Large for gestation age fetus
C0456091|T033|SY|199616008|SNOMEDCT_CORE|LFD - Fetus large for dates|Large for gestation age fetus
C0456091|T033|SY|199616008|SNOMEDCT_CORE|LFD - Foetus large for dates|Large for gestation age fetus
C0456091|T033|SY|199616008|SNOMEDCT_CORE|LGA - Large for gestational age fetus|Large for gestation age fetus
C0456091|T033|SY|199616008|SNOMEDCT_CORE|LGA - Large for gestational age foetus|Large for gestation age fetus
C0456128|T033|SY|57891003|SNOMEDCT_CORE|Baby full term maturity|Term infant
C0456128|T033|IS|57891003|SNOMEDCT_CORE|Term infancy|Term infant
C0456128|T033|FN|57891003|SNOMEDCT_CORE|Term infant|Term infant
C0456128|T033|PT|57891003|SNOMEDCT_CORE|Term infant|Term infant
C0456239|T047|PT|276883000|SNOMEDCT_CORE|Peritoneal dialysis-associated peritonitis|Peritoneal dialysis-associated peritonitis
C0456239|T047|FN|276883000|SNOMEDCT_CORE|Peritoneal dialysis-associated peritonitis|Peritoneal dialysis-associated peritonitis
C0456239|T047|SY|276883000|SNOMEDCT_CORE|Peritonitis secondary to peritoneal dialysis|Peritoneal dialysis-associated peritonitis
C0456537|T033|OAP|277213009|SNOMEDCT_CORE|Hearing aid worn|Hearing aid worn
C0456537|T033|OAF|277213009|SNOMEDCT_CORE|Hearing aid worn|Hearing aid worn
C0456541|T033|SY|249316004|SNOMEDCT_CORE|Crooked nose|Nasal deviation
C0456541|T033|PT|249316004|SNOMEDCT_CORE|Nasal deviation|Nasal deviation
C0456541|T033|FN|249316004|SNOMEDCT_CORE|Nasal deviation|Nasal deviation
C0456673|T033|PT|277357006|SNOMEDCT_CORE|Sputum retention|Sputum retention
C0456673|T033|FN|277357006|SNOMEDCT_CORE|Sputum retention|Sputum retention
C0456824|T037|PT|231466009|SNOMEDCT_CORE|Acute drug intoxication|Acute drug intoxication
C0456824|T037|FN|231466009|SNOMEDCT_CORE|Acute drug intoxication|Acute drug intoxication
C0456824|T037|SY|231466009|SNOMEDCT_CORE|Acute intoxication|Acute drug intoxication
C0456824|T037|SY|231466009|SNOMEDCT_CORE|Stoned|Acute drug intoxication
C0456909|T047|OAP|277675000|SNOMEDCT_CORE|Blind|Blind
C0456909|T047|OAF|277675000|SNOMEDCT_CORE|Blind|Blind
C0456973|T046|PT|87500009|SNOMEDCT_CORE|Hilar lymphadenopathy|Hilar lymphadenopathy
C0456973|T046|FN|87500009|SNOMEDCT_CORE|Hilar lymphadenopathy|Hilar lymphadenopathy
C0457084|T033|SY|277890004|SNOMEDCT_CORE|Swollen toe|Toe swelling
C0457084|T033|PT|277890004|SNOMEDCT_CORE|Toe swelling|Toe swelling
C0457084|T033|FN|277890004|SNOMEDCT_CORE|Toe swelling|Toe swelling
C0457205|T020|PT|197805009|SNOMEDCT_CORE|Postoperative ureteric constriction|Postoperative ureteric constriction
C0457205|T020|FN|197805009|SNOMEDCT_CORE|Postoperative ureteric constriction|Postoperative ureteric constriction
C0457205|T020|SY|197805009|SNOMEDCT_CORE|Postprocedural ureteric obstruction|Postoperative ureteric constriction
C0457238|T033|SY|278073009|SNOMEDCT_CORE|Technically poor CTG|Unsatisfactory CTG tracing
C0457238|T033|FN|278073009|SNOMEDCT_CORE|Unsatisfactory cardiotochogram tracing|Unsatisfactory CTG tracing
C0457238|T033|SY|278073009|SNOMEDCT_CORE|Unsatisfactory cardiotochogram tracing|Unsatisfactory CTG tracing
C0457238|T033|PT|278073009|SNOMEDCT_CORE|Unsatisfactory CTG tracing|Unsatisfactory CTG tracing
C0457238|T033|OF|278073009|SNOMEDCT_CORE|Unsatisfactory CTG tracing|Unsatisfactory CTG tracing
C0457798|T047|PT|93423006|SNOMEDCT_CORE|Dermatitis of eyelid|Dermatitis of eyelid
C0457798|T047|FN|93423006|SNOMEDCT_CORE|Dermatitis of eyelid|Dermatitis of eyelid
C0457798|T047|IS|93423006|SNOMEDCT_CORE|Dermatitis of eyelid, NOS|Dermatitis of eyelid
C0457949|T047|PT|278860009|SNOMEDCT_CORE|Chronic low back pain|Chronic low back pain
C0457949|T047|FN|278860009|SNOMEDCT_CORE|Chronic low back pain|Chronic low back pain
C0457949|T047|OF|278860009|SNOMEDCT_CORE|Chronic low back pain|Chronic low back pain
C0457949|T047|SY|278860009|SNOMEDCT_CORE|CLBP - Chronic low back pain|Chronic low back pain
C0457950|T184|SY|278862001|SNOMEDCT_CORE|Acute back pain - lumbar|Acute low back pain
C0457950|T184|PT|278862001|SNOMEDCT_CORE|Acute low back pain|Acute low back pain
C0457950|T184|FN|278862001|SNOMEDCT_CORE|Acute low back pain|Acute low back pain
C0457950|T184|OF|278862001|SNOMEDCT_CORE|Acute low back pain|Acute low back pain
C0457969|T033|PT|161432005|SNOMEDCT_CORE|H/O Malignant melanoma|H/O Malignant melanoma
C0457969|T033|OF|161432005|SNOMEDCT_CORE|History of - malignant melanoma|H/O Malignant melanoma
C0457969|T033|IS|161432005|SNOMEDCT_CORE|History of - malignant melanoma|H/O Malignant melanoma
C0457969|T033|FN|161432005|SNOMEDCT_CORE|History of malignant melanoma|H/O Malignant melanoma
C0457969|T033|SY|161432005|SNOMEDCT_CORE|History of malignant melanoma|H/O Malignant melanoma
C0457978|T020|SY|229811005|SNOMEDCT_CORE|Callosity on foot|Foot callus
C0457978|T020|PT|229811005|SNOMEDCT_CORE|Foot callus|Foot callus
C0457978|T020|FN|229811005|SNOMEDCT_CORE|Foot callus|Foot callus
C0458101|T047|PT|279016001|SNOMEDCT_CORE|Cervicogenic headache|Cervicogenic headache
C0458101|T047|FN|279016001|SNOMEDCT_CORE|Cervicogenic headache|Cervicogenic headache
C0458219|T047|SY|128200000|SNOMEDCT_CORE|Algodystrophy|Complex regional pain syndrome
C0458219|T047|PT|128200000|SNOMEDCT_CORE|Complex regional pain syndrome|Complex regional pain syndrome
C0458219|T047|IS|128200000|SNOMEDCT_CORE|Complex regional pain syndrome|Complex regional pain syndrome
C0458219|T047|FN|128200000|SNOMEDCT_CORE|Complex regional pain syndrome|Complex regional pain syndrome
C0458219|T047|OF|128200000|SNOMEDCT_CORE|Complex regional pain syndromes|Complex regional pain syndrome
C0458219|T047|IS|128200000|SNOMEDCT_CORE|Complex regional pain syndromes|Complex regional pain syndrome
C0458219|T047|SY|128200000|SNOMEDCT_CORE|CRPS - complex regional pain syndrome|Complex regional pain syndrome
C0458219|T047|IS|128200000|SNOMEDCT_CORE|Reflex sympathetic dystrophy|Complex regional pain syndrome
C0458219|T047|IS|128200000|SNOMEDCT_CORE|Sudek atrophy|Complex regional pain syndrome
C0458224|T047|SY|129179000|SNOMEDCT_CORE|Pelvic outlet syndrome|Piriformis syndrome
C0458224|T047|PT|129179000|SNOMEDCT_CORE|Piriformis syndrome|Piriformis syndrome
C0458224|T047|FN|129179000|SNOMEDCT_CORE|Piriformis syndrome|Piriformis syndrome
C0458224|T047|IS|129179000|SNOMEDCT_CORE|Sciatica due to compression of sciatic nerve at pelvic outlet|Piriformis syndrome
C0458228|T184|PT|202479004|SNOMEDCT_CORE|Acromioclavicular joint pain|Acromioclavicular joint pain
C0458228|T184|FN|202479004|SNOMEDCT_CORE|Acromioclavicular joint pain|Acromioclavicular joint pain
C0458228|T184|SY|202479004|SNOMEDCT_CORE|Arthralgia of acromioclavicular joint|Acromioclavicular joint pain
C0458232|T184|SY|202487003|SNOMEDCT_CORE|Arthralgia of sacroiliac joint|Sacroiliac joint pain
C0458232|T184|PT|202487003|SNOMEDCT_CORE|Sacroiliac joint pain|Sacroiliac joint pain
C0458232|T184|FN|202487003|SNOMEDCT_CORE|Sacroiliac joint pain|Sacroiliac joint pain
C0458233|T184|SY|202489000|SNOMEDCT_CORE|Arthralgia of tibiofibular joint|Tibiofibular joint pain
C0458233|T184|PT|202489000|SNOMEDCT_CORE|Tibiofibular joint pain|Tibiofibular joint pain
C0458233|T184|FN|202489000|SNOMEDCT_CORE|Tibiofibular joint pain|Tibiofibular joint pain
C0458239|T184|SY|279066007|SNOMEDCT_CORE|Arthralgia of foot|Foot joint pain
C0458239|T184|PT|279066007|SNOMEDCT_CORE|Foot joint pain|Foot joint pain
C0458239|T184|FN|279066007|SNOMEDCT_CORE|Foot joint pain|Foot joint pain
C0458990|T033|PT|279992002|SNOMEDCT_CORE|Recurrent falls|Recurrent falls
C0458990|T033|FN|279992002|SNOMEDCT_CORE|Recurrent falls|Recurrent falls
C0459830|T047|PT|195303005|SNOMEDCT_CORE|Gangrene of foot|Gangrene of foot
C0459830|T047|FN|195303005|SNOMEDCT_CORE|Gangrene of foot|Gangrene of foot
C0459853|T033|PT|161508001|SNOMEDCT_CORE|H/O: Deep vein thrombosis|H/O: Deep vein thrombosis
C0459853|T033|IS|161508001|SNOMEDCT_CORE|H/O: Deep Vein Thrombosis|H/O: Deep vein thrombosis
C0459853|T033|OF|161508001|SNOMEDCT_CORE|History of - deep vein thrombosis|H/O: Deep vein thrombosis
C0459853|T033|IS|161508001|SNOMEDCT_CORE|History of - deep vein thrombosis|H/O: Deep vein thrombosis
C0459853|T033|FN|161508001|SNOMEDCT_CORE|History of deep vein thrombosis|H/O: Deep vein thrombosis
C0459853|T033|SY|161508001|SNOMEDCT_CORE|History of deep vein thrombosis|H/O: Deep vein thrombosis
C0460098|T033|PT|281305005|SNOMEDCT_CORE|Unwanted fertility|Unwanted fertility
C0460098|T033|FN|281305005|SNOMEDCT_CORE|Unwanted fertility|Unwanted fertility
C0472692|T047|SY|33129002|SNOMEDCT_CORE|Elephantiasis due to mastectomy|Postmastectomy lymphedema syndrome
C0472692|T047|SY|33129002|SNOMEDCT_CORE|Obliteration of lymphatic vessel due to mastectomy|Postmastectomy lymphedema syndrome
C0472692|T047|SY|33129002|SNOMEDCT_CORE|Post-mastectomy secondary lymphedema|Postmastectomy lymphedema syndrome
C0472692|T047|SYGB|33129002|SNOMEDCT_CORE|Post-mastectomy secondary lymphoedema|Postmastectomy lymphedema syndrome
C0472692|T047|PT|33129002|SNOMEDCT_CORE|Postmastectomy lymphedema syndrome|Postmastectomy lymphedema syndrome
C0472692|T047|FN|33129002|SNOMEDCT_CORE|Postmastectomy lymphedema syndrome|Postmastectomy lymphedema syndrome
C0472692|T047|PTGB|33129002|SNOMEDCT_CORE|Postmastectomy lymphoedema syndrome|Postmastectomy lymphedema syndrome
C0472713|T047|PTGB|234348004|SNOMEDCT_CORE|Anaemia of renal disease|Anemia of renal disease
C0472713|T047|PT|234348004|SNOMEDCT_CORE|Anemia of renal disease|Anemia of renal disease
C0472713|T047|FN|234348004|SNOMEDCT_CORE|Anemia of renal disease|Anemia of renal disease
C0472713|T047|SYGB|234348004|SNOMEDCT_CORE|Nephrogenic anaemia|Anemia of renal disease
C0472713|T047|SY|234348004|SNOMEDCT_CORE|Nephrogenic anemia|Anemia of renal disease
C0472762|T047|SYGB|191187006|SNOMEDCT_CORE|Alpha thalassaemia trait|Alpha trait thalassemia
C0472762|T047|SY|191187006|SNOMEDCT_CORE|Alpha thalassemia trait|Alpha trait thalassemia
C0472762|T047|PTGB|191187006|SNOMEDCT_CORE|Alpha trait thalassaemia|Alpha trait thalassemia
C0472762|T047|PT|191187006|SNOMEDCT_CORE|Alpha trait thalassemia|Alpha trait thalassemia
C0472762|T047|FN|191187006|SNOMEDCT_CORE|Alpha trait thalassemia|Alpha trait thalassemia
C0472793|T047|PTGB|234413005|SNOMEDCT_CORE|Alpha/beta lipoproteinaemia|Alpha/beta lipoproteinemia
C0472793|T047|PT|234413005|SNOMEDCT_CORE|Alpha/beta lipoproteinemia|Alpha/beta lipoproteinemia
C0472793|T047|FN|234413005|SNOMEDCT_CORE|Alpha/beta lipoproteinemia|Alpha/beta lipoproteinemia
C0473119|T047|PTGB|235985005|SNOMEDCT_CORE|Faecal peritonitis|Fecal peritonitis
C0473119|T047|PT|235985005|SNOMEDCT_CORE|Fecal peritonitis|Fecal peritonitis
C0473119|T047|FN|235985005|SNOMEDCT_CORE|Fecal peritonitis|Fecal peritonitis
C0473237|T033|PTGB|197941005|SNOMEDCT_CORE|Frank haematuria|Frank hematuria
C0473237|T033|PT|197941005|SNOMEDCT_CORE|Frank hematuria|Frank hematuria
C0473237|T033|FN|197941005|SNOMEDCT_CORE|Frank hematuria|Frank hematuria
C0473237|T033|SY|197941005|SNOMEDCT_CORE|Gross hematuria|Frank hematuria
C0473237|T033|SYGB|197941005|SNOMEDCT_CORE|Macroscopic haematuria|Frank hematuria
C0473237|T033|SY|197941005|SNOMEDCT_CORE|Macroscopic hematuria|Frank hematuria
C0473313|T020|PTGB|237102006|SNOMEDCT_CORE|Vaginal vault haematoma|Vaginal vault hematoma
C0473313|T020|PT|237102006|SNOMEDCT_CORE|Vaginal vault hematoma|Vaginal vault hematoma
C0473313|T020|FN|237102006|SNOMEDCT_CORE|Vaginal vault hematoma|Vaginal vault hematoma
C0473326|T047|PTGB|199246003|SNOMEDCT_CORE|Anaemia during pregnancy - baby not yet delivered|Anemia during pregnancy - baby not yet delivered
C0473326|T047|PT|199246003|SNOMEDCT_CORE|Anemia during pregnancy - baby not yet delivered|Anemia during pregnancy - baby not yet delivered
C0473326|T047|FN|199246003|SNOMEDCT_CORE|Anemia during pregnancy - baby not yet delivered|Anemia during pregnancy - baby not yet delivered
C0473326|T047|SYGB|199246003|SNOMEDCT_CORE|Maternal anaemia in pregnancy, before birth|Anemia during pregnancy - baby not yet delivered
C0473326|T047|SY|199246003|SNOMEDCT_CORE|Maternal anemia in pregnancy, before birth|Anemia during pregnancy - baby not yet delivered
C0473389|T033|SY|199049003|SNOMEDCT_CORE|False premature labor|Threatened premature labor - not delivered
C0473389|T033|SYGB|199049003|SNOMEDCT_CORE|False premature labour|Threatened premature labor - not delivered
C0473389|T033|PT|199049003|SNOMEDCT_CORE|Threatened premature labor - not delivered|Threatened premature labor - not delivered
C0473389|T033|FN|199049003|SNOMEDCT_CORE|Threatened premature labor - not delivered|Threatened premature labor - not delivered
C0473389|T033|OF|199049003|SNOMEDCT_CORE|Threatened premature labor - not delivered|Threatened premature labor - not delivered
C0473389|T033|PTGB|199049003|SNOMEDCT_CORE|Threatened premature labour - not delivered|Threatened premature labor - not delivered
C0473390|T046|OAS|4946002|SNOMEDCT_CORE|Premature labor after 22 weeks but before 37 completed weeks of gestation without delivery|Threatened premature labor
C0473390|T046|OAS|4946002|SNOMEDCT_CORE|Premature labour after 22 weeks but before 37 completed weeks of gestation without delivery|Threatened premature labor
C0473390|T046|IS|199047001|SNOMEDCT_CORE|Threatened premature labor|Threatened premature labor
C0473390|T046|OAP|4946002|SNOMEDCT_CORE|Threatened premature labor|Threatened premature labor
C0473390|T046|OAF|4946002|SNOMEDCT_CORE|Threatened premature labor|Threatened premature labor
C0473390|T046|IS|199047001|SNOMEDCT_CORE|Threatened premature labour|Threatened premature labor
C0473390|T046|OAP|4946002|SNOMEDCT_CORE|Threatened premature labour|Threatened premature labor
C0473408|T047|PTGB|199583002|SNOMEDCT_CORE|Rhesus isoimmunisation with antenatal problem|Rhesus isoimmunization with antenatal problem
C0473408|T047|PT|199583002|SNOMEDCT_CORE|Rhesus isoimmunization with antenatal problem|Rhesus isoimmunization with antenatal problem
C0473408|T047|FN|199583002|SNOMEDCT_CORE|Rhesus isoimmunization with antenatal problem|Rhesus isoimmunization with antenatal problem
C0473508|T046|PTGB|23171006|SNOMEDCT_CORE|Delayed AND/OR secondary postpartum haemorrhage|Delayed AND/OR secondary postpartum hemorrhage
C0473508|T046|PT|23171006|SNOMEDCT_CORE|Delayed AND/OR secondary postpartum hemorrhage|Delayed AND/OR secondary postpartum hemorrhage
C0473508|T046|FN|23171006|SNOMEDCT_CORE|Delayed AND/OR secondary postpartum hemorrhage|Delayed AND/OR secondary postpartum hemorrhage
C0473508|T046|IS|23171006|SNOMEDCT_CORE|Delayed or secondary postpartum hemorrhage|Delayed AND/OR secondary postpartum hemorrhage
C0473508|T046|SYGB|23171006|SNOMEDCT_CORE|Delayed postpartum haemorrhage|Delayed AND/OR secondary postpartum hemorrhage
C0473508|T046|SY|23171006|SNOMEDCT_CORE|Delayed postpartum hemorrhage|Delayed AND/OR secondary postpartum hemorrhage
C0473508|T046|SYGB|23171006|SNOMEDCT_CORE|Haemorrhage after first 24 hours following delivery of placenta|Delayed AND/OR secondary postpartum hemorrhage
C0473508|T046|SY|23171006|SNOMEDCT_CORE|Hemorrhage after first 24 hours following delivery of placenta|Delayed AND/OR secondary postpartum hemorrhage
C0473508|T046|SYGB|23171006|SNOMEDCT_CORE|Postpartum haemorrhage specified as delayed or secondary|Delayed AND/OR secondary postpartum hemorrhage
C0473508|T046|SYGB|23171006|SNOMEDCT_CORE|Postpartum haemorrhage, delayed AND/OR secondary|Delayed AND/OR secondary postpartum hemorrhage
C0473508|T046|SY|23171006|SNOMEDCT_CORE|Postpartum hemorrhage specified as delayed or secondary|Delayed AND/OR secondary postpartum hemorrhage
C0473508|T046|SY|23171006|SNOMEDCT_CORE|Postpartum hemorrhage, delayed AND/OR secondary|Delayed AND/OR secondary postpartum hemorrhage
C0473527|T047|OAP|190784001|SNOMEDCT_CORE|High density lipoid deficiency|High density lipoid deficiency
C0473527|T047|OAF|190784001|SNOMEDCT_CORE|High density lipoid deficiency|High density lipoid deficiency
C0473557|T047|OAP|238793001|SNOMEDCT_CORE|Ischaemic leg ulcer|Ischemic leg ulcer
C0473557|T047|OAP|238793001|SNOMEDCT_CORE|Ischemic leg ulcer|Ischemic leg ulcer
C0473557|T047|OAF|238793001|SNOMEDCT_CORE|Ischemic leg ulcer|Ischemic leg ulcer
C0473748|T047|PTGB|201835007|SNOMEDCT_CORE|Localised, primary osteoarthritis of the pelvic region and thigh|Localized, primary osteoarthritis of the pelvic region and thigh
C0473748|T047|PT|201835007|SNOMEDCT_CORE|Localized, primary osteoarthritis of the pelvic region and thigh|Localized, primary osteoarthritis of the pelvic region and thigh
C0473748|T047|FN|201835007|SNOMEDCT_CORE|Localized, primary osteoarthritis of the pelvic region and thigh|Localized, primary osteoarthritis of the pelvic region and thigh
C0473762|T047|PTGB|201849003|SNOMEDCT_CORE|Localised, secondary osteoarthritis of the shoulder region|Localized, secondary osteoarthritis of the shoulder region
C0473762|T047|PT|201849003|SNOMEDCT_CORE|Localized, secondary osteoarthritis of the shoulder region|Localized, secondary osteoarthritis of the shoulder region
C0473762|T047|FN|201849003|SNOMEDCT_CORE|Localized, secondary osteoarthritis of the shoulder region|Localized, secondary osteoarthritis of the shoulder region
C0473762|T047|SYGB|201849003|SNOMEDCT_CORE|Secondary localised osteoarthrosis of shoulder region|Localized, secondary osteoarthritis of the shoulder region
C0473762|T047|SY|201849003|SNOMEDCT_CORE|Secondary localized osteoarthrosis of shoulder region|Localized, secondary osteoarthritis of the shoulder region
C0473785|T047|PTGB|206470003|SNOMEDCT_CORE|Perinatal jaundice due to galactosaemia|Perinatal jaundice due to galactosemia
C0473785|T047|PT|206470003|SNOMEDCT_CORE|Perinatal jaundice due to galactosemia|Perinatal jaundice due to galactosemia
C0473785|T047|FN|206470003|SNOMEDCT_CORE|Perinatal jaundice due to galactosemia|Perinatal jaundice due to galactosemia
C0473839|T033|PT|206116006|SNOMEDCT_CORE|Fetal or neonatal effect of transverse lie during labor and delivery|Fetal or neonatal effect of transverse lie during labor and delivery
C0473839|T033|FN|206116006|SNOMEDCT_CORE|Fetal or neonatal effect of transverse lie during labor and delivery|Fetal or neonatal effect of transverse lie during labor and delivery
C0473839|T033|PTGB|206116006|SNOMEDCT_CORE|Fetal or neonatal effect of transverse lie during labour and delivery|Fetal or neonatal effect of transverse lie during labor and delivery
C0473839|T033|OP|206116006|SNOMEDCT_CORE|Fetus or neonate affected by transverse lie during labor and delivery|Fetal or neonatal effect of transverse lie during labor and delivery
C0473839|T033|OF|206116006|SNOMEDCT_CORE|Fetus or neonate affected by transverse lie during labor and delivery|Fetal or neonatal effect of transverse lie during labor and delivery
C0473839|T033|IS|206116006|SNOMEDCT_CORE|Fetus or neonate affected by transverse lie during labour and delivery|Fetal or neonatal effect of transverse lie during labor and delivery
C0473839|T033|SYGB|206116006|SNOMEDCT_CORE|Foetal or neonatal effect of transverse lie during labour and delivery|Fetal or neonatal effect of transverse lie during labor and delivery
C0473839|T033|OP|206116006|SNOMEDCT_CORE|Foetus or neonate affected by transverse lie during labour and delivery|Fetal or neonatal effect of transverse lie during labor and delivery
C0473841|T033|SY|206118007|SNOMEDCT_CORE|Fetal or neonatal effect of cephalopelvic disproportion during labor and delivery|Fetal or neonatal effect of disproportion during labor and delivery
C0473841|T033|IS|206118007|SNOMEDCT_CORE|Fetal or neonatal effect of cephalopelvic disproportion during labour and delivery|Fetal or neonatal effect of disproportion during labor and delivery
C0473841|T033|PT|206118007|SNOMEDCT_CORE|Fetal or neonatal effect of disproportion during labor and delivery|Fetal or neonatal effect of disproportion during labor and delivery
C0473841|T033|FN|206118007|SNOMEDCT_CORE|Fetal or neonatal effect of disproportion during labor and delivery|Fetal or neonatal effect of disproportion during labor and delivery
C0473841|T033|PTGB|206118007|SNOMEDCT_CORE|Fetal or neonatal effect of disproportion during labour and delivery|Fetal or neonatal effect of disproportion during labor and delivery
C0473841|T033|IS|206118007|SNOMEDCT_CORE|Fetus or neonate affected by cephalopelvic disproportion during labor and delivery|Fetal or neonatal effect of disproportion during labor and delivery
C0473841|T033|IS|206118007|SNOMEDCT_CORE|Fetus or neonate affected by cephalopelvic disproportion during labour and delivery|Fetal or neonatal effect of disproportion during labor and delivery
C0473841|T033|OP|206118007|SNOMEDCT_CORE|Fetus or neonate affected by disproportion during labor and delivery|Fetal or neonatal effect of disproportion during labor and delivery
C0473841|T033|OF|206118007|SNOMEDCT_CORE|Fetus or neonate affected by disproportion during labor and delivery|Fetal or neonatal effect of disproportion during labor and delivery
C0473841|T033|IS|206118007|SNOMEDCT_CORE|Fetus or neonate affected by disproportion during labour and delivery|Fetal or neonatal effect of disproportion during labor and delivery
C0473841|T033|SYGB|206118007|SNOMEDCT_CORE|Foetal or neonatal effect of cephalopelvic disproportion during labour and delivery|Fetal or neonatal effect of disproportion during labor and delivery
C0473841|T033|SYGB|206118007|SNOMEDCT_CORE|Foetal or neonatal effect of disproportion during labour and delivery|Fetal or neonatal effect of disproportion during labor and delivery
C0473841|T033|IS|206118007|SNOMEDCT_CORE|Foetus or neonate affected by cephalopelvic disproportion during labour and delivery|Fetal or neonatal effect of disproportion during labor and delivery
C0473841|T033|OP|206118007|SNOMEDCT_CORE|Foetus or neonate affected by disproportion during labour and delivery|Fetal or neonatal effect of disproportion during labor and delivery
C0474298|T033|PTGB|171258008|SNOMEDCT_CORE|Up-to-date with immunisations|Up-to-date with immunizations
C0474298|T033|PT|171258008|SNOMEDCT_CORE|Up-to-date with immunizations|Up-to-date with immunizations
C0474298|T033|FN|171258008|SNOMEDCT_CORE|Up-to-date with immunizations|Up-to-date with immunizations
C0474327|T046|PTGB|246544003|SNOMEDCT_CORE|Partial seizure evolving to secondary generalised seizure|Partial seizure evolving to secondary generalized seizure
C0474327|T046|PT|246544003|SNOMEDCT_CORE|Partial seizure evolving to secondary generalized seizure|Partial seizure evolving to secondary generalized seizure
C0474327|T046|OF|246544003|SNOMEDCT_CORE|Partial seizure evolving to secondary generalized seizure|Partial seizure evolving to secondary generalized seizure
C0474327|T046|FN|246544003|SNOMEDCT_CORE|Partial seizure evolving to secondary generalized seizure|Partial seizure evolving to secondary generalized seizure
C0474413|T048|PT|248036002|SNOMEDCT_CORE|Problematic behavior in children|Problematic behavior in children
C0474413|T048|FN|248036002|SNOMEDCT_CORE|Problematic behavior in children|Problematic behavior in children
C0474413|T048|PTGB|248036002|SNOMEDCT_CORE|Problematic behaviour in children|Problematic behavior in children
C0474481|T033|PT|249166003|SNOMEDCT_CORE|Failure to progress in second stage of labor|Failure to progress in second stage of labor
C0474481|T033|FN|249166003|SNOMEDCT_CORE|Failure to progress in second stage of labor|Failure to progress in second stage of labor
C0474481|T033|PTGB|249166003|SNOMEDCT_CORE|Failure to progress in second stage of labour|Failure to progress in second stage of labor
C0474481|T033|SY|249166003|SNOMEDCT_CORE|No progress in second stage of labor|Failure to progress in second stage of labor
C0474481|T033|SYGB|249166003|SNOMEDCT_CORE|No progress in second stage of labour|Failure to progress in second stage of labor
C0474481|T033|SY|249166003|SNOMEDCT_CORE|No progress with delivery|Failure to progress in second stage of labor
C0474822|T191|PTGB|253032007|SNOMEDCT_CORE|Benign phaeochromocytoma|Benign pheochromocytoma
C0474822|T191|PT|253032007|SNOMEDCT_CORE|Benign pheochromocytoma|Benign pheochromocytoma
C0474822|T191|FN|253032007|SNOMEDCT_CORE|Benign pheochromocytoma|Benign pheochromocytoma
C0475059|T037|OAP|262951009|SNOMEDCT_CORE|Traumatic subdural haematoma|Traumatic subdural haematoma
C0475059|T037|OAP|262951009|SNOMEDCT_CORE|Traumatic subdural hematoma|Traumatic subdural hematoma
C0475059|T037|OAF|262951009|SNOMEDCT_CORE|Traumatic subdural hematoma|Traumatic subdural hematoma
C0475060|T037|SYGB|262952002|SNOMEDCT_CORE|Traumatic cranial subdural haematoma|Traumatic subdural hematoma
C0475060|T037|SY|262952002|SNOMEDCT_CORE|Traumatic cranial subdural hematoma|Traumatic subdural hematoma
C0475060|T037|SYGB|262952002|SNOMEDCT_CORE|Traumatic intracranial subdural haematoma|Traumatic subdural hematoma
C0475060|T037|SY|262952002|SNOMEDCT_CORE|Traumatic intracranial subdural hematoma|Traumatic subdural hematoma
C0475060|T037|FN|262952002|SNOMEDCT_CORE|Traumatic intracranial subdural hematoma|Traumatic subdural hematoma
C0475060|T037|PTGB|262952002|SNOMEDCT_CORE|Traumatic subdural haematoma|Traumatic subdural hematoma
C0475060|T037|PT|262952002|SNOMEDCT_CORE|Traumatic subdural hematoma|Traumatic subdural hematoma
C0475073|T037|PTGB|262955000|SNOMEDCT_CORE|Subarachnoid haemorrhage due to traumatic injury|Subarachnoid hemorrhage due to traumatic injury
C0475073|T037|OAS|262954001|SNOMEDCT_CORE|Subarachnoid haemorrhage following injury|Subarachnoid hemorrhage due to traumatic injury
C0475073|T037|FN|262955000|SNOMEDCT_CORE|Subarachnoid hemorrhage due to traumatic injury|Subarachnoid hemorrhage due to traumatic injury
C0475073|T037|PT|262955000|SNOMEDCT_CORE|Subarachnoid hemorrhage due to traumatic injury|Subarachnoid hemorrhage due to traumatic injury
C0475073|T037|OAS|262954001|SNOMEDCT_CORE|Subarachnoid hemorrhage following injury|Subarachnoid hemorrhage due to traumatic injury
C0475073|T037|SYGB|262955000|SNOMEDCT_CORE|Traumatic cranial subarachnoid haemorrhage|Subarachnoid hemorrhage due to traumatic injury
C0475073|T037|SY|262955000|SNOMEDCT_CORE|Traumatic cranial subarachnoid hemorrhage|Subarachnoid hemorrhage due to traumatic injury
C0475073|T037|SYGB|262955000|SNOMEDCT_CORE|Traumatic haemorrhage into subarachnoid space of neuraxis|Subarachnoid hemorrhage due to traumatic injury
C0475073|T037|SY|262955000|SNOMEDCT_CORE|Traumatic hemorrhage into subarachnoid space of neuraxis|Subarachnoid hemorrhage due to traumatic injury
C0475073|T037|SYGB|262955000|SNOMEDCT_CORE|Traumatic intracranial subarachnoid haemorrhage|Subarachnoid hemorrhage due to traumatic injury
C0475073|T037|SY|262955000|SNOMEDCT_CORE|Traumatic intracranial subarachnoid hemorrhage|Subarachnoid hemorrhage due to traumatic injury
C0475073|T037|OF|262955000|SNOMEDCT_CORE|Traumatic intracranial subarachnoid hemorrhage|Subarachnoid hemorrhage due to traumatic injury
C0475073|T037|OAP|262954001|SNOMEDCT_CORE|Traumatic subarachnoid haemorrhage|Subarachnoid hemorrhage due to traumatic injury
C0475073|T037|OAP|262954001|SNOMEDCT_CORE|Traumatic subarachnoid hemorrhage|Subarachnoid hemorrhage due to traumatic injury
C0475073|T037|OF|262954001|SNOMEDCT_CORE|Traumatic subarachnoid hemorrhage|Subarachnoid hemorrhage due to traumatic injury
C0475073|T037|OAS|262954001|SNOMEDCT_CORE|Traumatic subarachnoid intracranial haemorrhage|Subarachnoid hemorrhage due to traumatic injury
C0475073|T037|OAS|262954001|SNOMEDCT_CORE|Traumatic subarachnoid intracranial hemorrhage|Subarachnoid hemorrhage due to traumatic injury
C0475073|T037|OAF|262954001|SNOMEDCT_CORE|Traumatic subarachnoid intracranial hemorrhage|Subarachnoid hemorrhage due to traumatic injury
C0475172|T033|PTGB|161805006|SNOMEDCT_CORE|H/O: caesarean section|H/O: cesarean section
C0475172|T033|PT|161805006|SNOMEDCT_CORE|H/O: cesarean section|H/O: cesarean section
C0475172|T033|OF|161805006|SNOMEDCT_CORE|History of - cesarean section|H/O: cesarean section
C0475172|T033|IS|161805006|SNOMEDCT_CORE|History of - cesarean section|H/O: cesarean section
C0475172|T033|SYGB|161805006|SNOMEDCT_CORE|History of caesarean section|H/O: cesarean section
C0475172|T033|FN|161805006|SNOMEDCT_CORE|History of cesarean section|H/O: cesarean section
C0475172|T033|SY|161805006|SNOMEDCT_CORE|History of cesarean section|H/O: cesarean section
C0475534|T047|PTGB|191265009|SNOMEDCT_CORE|Anaemia in neoplastic disease|Anemia in neoplastic disease
C0475534|T047|PT|191265009|SNOMEDCT_CORE|Anemia in neoplastic disease|Anemia in neoplastic disease
C0475534|T047|FN|191265009|SNOMEDCT_CORE|Anemia in neoplastic disease|Anemia in neoplastic disease
C0475715|T046|PT|276544005|SNOMEDCT_CORE|Apnea of prematurity|Apnea of prematurity
C0475715|T046|FN|276544005|SNOMEDCT_CORE|Apnea of prematurity|Apnea of prematurity
C0475715|T046|PTGB|276544005|SNOMEDCT_CORE|Apnoea of prematurity|Apnea of prematurity
C0475728|T046|SYGB|276622005|SNOMEDCT_CORE|Epicranial subaponeurotic haemorrhage|Subgaleal hemorrhage
C0475728|T046|SY|276622005|SNOMEDCT_CORE|Epicranial subaponeurotic hemorrhage|Subgaleal hemorrhage
C0475728|T046|FN|276622005|SNOMEDCT_CORE|Epicranial subaponeurotic hemorrhage|Subgaleal hemorrhage
C0475728|T046|IS|276622005|SNOMEDCT_CORE|Subaponeurotic haematoma|Subgaleal hemorrhage
C0475728|T046|SYGB|276622005|SNOMEDCT_CORE|Subaponeurotic haemorrhage|Subgaleal hemorrhage
C0475728|T046|IS|276622005|SNOMEDCT_CORE|Subaponeurotic hematoma|Subgaleal hemorrhage
C0475728|T046|SY|276622005|SNOMEDCT_CORE|Subaponeurotic hemorrhage|Subgaleal hemorrhage
C0475728|T046|IS|276622005|SNOMEDCT_CORE|Subgaleal haematoma|Subgaleal hemorrhage
C0475728|T046|PTGB|276622005|SNOMEDCT_CORE|Subgaleal haemorrhage|Subgaleal hemorrhage
C0475728|T046|IS|276622005|SNOMEDCT_CORE|Subgaleal hematoma|Subgaleal hemorrhage
C0475728|T046|PT|276622005|SNOMEDCT_CORE|Subgaleal hemorrhage|Subgaleal hemorrhage
C0475858|T184|SYGB|276444007|SNOMEDCT_CORE|Generalised itching|Generalized pruritus
C0475858|T184|PTGB|276444007|SNOMEDCT_CORE|Generalised pruritus|Generalized pruritus
C0475858|T184|SY|276444007|SNOMEDCT_CORE|Generalized itching|Generalized pruritus
C0475858|T184|PT|276444007|SNOMEDCT_CORE|Generalized pruritus|Generalized pruritus
C0475858|T184|FN|276444007|SNOMEDCT_CORE|Generalized pruritus|Generalized pruritus
C0476089|T191|IS|254878006|SNOMEDCT_CORE|Endometrial Ca|Endometrial carcinoma
C0476089|T191|PT|254878006|SNOMEDCT_CORE|Endometrial carcinoma|Endometrial carcinoma
C0476089|T191|FN|254878006|SNOMEDCT_CORE|Endometrial carcinoma|Endometrial carcinoma
C0476206|T184|SY|271789005|SNOMEDCT_CORE|Dizziness - giddy|Dizziness and giddiness
C0476206|T184|PT|271789005|SNOMEDCT_CORE|Dizziness and giddiness|Dizziness and giddiness
C0476206|T184|FN|271789005|SNOMEDCT_CORE|Dizziness and giddiness|Dizziness and giddiness
C0476206|T184|IS|271789005|SNOMEDCT_CORE|Giddiness|Dizziness and giddiness
C0476207|T184|IS|399153001|SNOMEDCT_CORE|Vertigo - giddiness|Vertigo - giddiness
C0476241|T033|SY|274625009|SNOMEDCT_CORE|Delayed developmental milestone|Delayed milestone
C0476241|T033|PT|274625009|SNOMEDCT_CORE|Delayed milestone|Delayed milestone
C0476241|T033|FN|274625009|SNOMEDCT_CORE|Delayed milestone|Delayed milestone
C0476250|T184|SY|274751001|SNOMEDCT_CORE|Head and neck mass|Mass in head or neck
C0476250|T184|PT|274751001|SNOMEDCT_CORE|Mass in head or neck|Mass in head or neck
C0476250|T184|FN|274751001|SNOMEDCT_CORE|Mass in head or neck|Mass in head or neck
C0476254|T048|SY|52824009|SNOMEDCT_CORE|Reading disorder|Reading disorder
C0476273|T184|SY|271825005|SNOMEDCT_CORE|Distressed breathing|Respiratory distress
C0476273|T184|PT|271825005|SNOMEDCT_CORE|Respiratory distress|Respiratory distress
C0476273|T184|FN|271825005|SNOMEDCT_CORE|Respiratory distress|Respiratory distress
C0476280|T184|PT|281245003|SNOMEDCT_CORE|Musculoskeletal chest pain|Musculoskeletal chest pain
C0476280|T184|FN|281245003|SNOMEDCT_CORE|Musculoskeletal chest pain|Musculoskeletal chest pain
C0476281|T184|PT|274668005|SNOMEDCT_CORE|Non-cardiac chest pain|Non-cardiac chest pain
C0476281|T184|FN|274668005|SNOMEDCT_CORE|Non-cardiac chest pain|Non-cardiac chest pain
C0476281|T184|SY|274668005|SNOMEDCT_CORE|Noncardiac chest pain|Non-cardiac chest pain
C0476346|T033|PTGB|249625002|SNOMEDCT_CORE|Faeces contents abnormal|Feces contents abnormal
C0476346|T033|PT|249625002|SNOMEDCT_CORE|Feces contents abnormal|Feces contents abnormal
C0476346|T033|FN|249625002|SNOMEDCT_CORE|Feces contents abnormal|Feces contents abnormal
C0476346|T033|SY|249625002|SNOMEDCT_CORE|Stool contents abnormal|Feces contents abnormal
C0476367|T033|PT|274714007|SNOMEDCT_CORE|Shadow of lung|Shadow of lung
C0476367|T033|FN|274714007|SNOMEDCT_CORE|Shadow of lung|Shadow of lung
C0476369|T033|PT|169241000|SNOMEDCT_CORE|Echocardiogram abnormal|Echocardiogram abnormal
C0476369|T033|FN|169241000|SNOMEDCT_CORE|Echocardiogram abnormal|Echocardiogram abnormal
C0476382|T033|PT|441684001|SNOMEDCT_CORE|Lytic lesion of bone on X-ray|Lytic lesion of bone on X-ray
C0476382|T033|FN|441684001|SNOMEDCT_CORE|Lytic lesion of bone on X-ray|Lytic lesion of bone on X-ray
C0476414|T033|PT|312399001|SNOMEDCT_CORE|Thyroid function tests abnormal|Thyroid function tests abnormal
C0476414|T033|FN|312399001|SNOMEDCT_CORE|Thyroid function tests abnormal|Thyroid function tests abnormal
C0476427|T033|FN|439888000|SNOMEDCT_CORE|Abnormal cervical Papanicolaou smear|Abnormal cervical smear
C0476427|T033|PT|439888000|SNOMEDCT_CORE|Abnormal cervical Papanicolaou smear|Abnormal cervical smear
C0476427|T033|PT|309081009|SNOMEDCT_CORE|Abnormal cervical smear|Abnormal cervical smear
C0476427|T033|FN|309081009|SNOMEDCT_CORE|Abnormal cervical smear|Abnormal cervical smear
C0476587|T033|PT|105419003|SNOMEDCT_CORE|Academic underachievement|Academic underachievement
C0476587|T033|FN|105419003|SNOMEDCT_CORE|Academic underachievement|Academic underachievement
C0476587|T033|IS|105419003|SNOMEDCT_CORE|Underachievement in school|Academic underachievement
C0477633|T047|SY|425878001|SNOMEDCT_CORE|Cervical disc disease|Cervical disc disorder
C0477633|T047|PT|425878001|SNOMEDCT_CORE|Cervical disc disorder|Cervical disc disorder
C0477633|T047|FN|425878001|SNOMEDCT_CORE|Cervical disc disorder|Cervical disc disorder
C0478655|T048|SY|5510009|SNOMEDCT_CORE|Paranoid organic state|Paranoid organic state
C0478933|T037|IS|35468003|SNOMEDCT_CORE|Caught, crushed, jammed or pinched in or between objects|Caught, crushed, jammed or pinched in or between objects
C0480203|T037|SY|276853009|SNOMEDCT_CORE|Injury - self-inflicted|Self inflicted injury
C0480203|T037|PT|276853009|SNOMEDCT_CORE|Self inflicted injury|Self inflicted injury
C0480203|T037|OF|276853009|SNOMEDCT_CORE|Self inflicted injury|Self inflicted injury
C0480203|T037|FN|276853009|SNOMEDCT_CORE|Self inflicted injury|Self inflicted injury
C0481354|T037|PT|218247007|SNOMEDCT_CORE|Late effect of motor vehicle accident|Late effect of motor vehicle accident
C0481354|T037|FN|218247007|SNOMEDCT_CORE|Late effect of motor vehicle accident|Late effect of motor vehicle accident
C0481354|T037|IS|218247007|SNOMEDCT_CORE|Late effects of motor vehicle accident|Late effect of motor vehicle accident
C0481354|T037|OF|218247007|SNOMEDCT_CORE|Late effects of motor vehicle accident|Late effect of motor vehicle accident
C0481457|T033|PT|169826009|SNOMEDCT_CORE|Single live birth|Single live birth
C0481457|T033|FN|169826009|SNOMEDCT_CORE|Single live birth|Single live birth
C0489967|T047|PT|9009001|SNOMEDCT_CORE|Low compliance bladder|Low compliance bladder
C0489967|T047|FN|9009001|SNOMEDCT_CORE|Low compliance bladder|Low compliance bladder
C0489985|T046|PT|441630004|SNOMEDCT_CORE|Aphasia as late effect of cerebrovascular disease|Aphasia as late effect of cerebrovascular disease
C0489985|T046|FN|441630004|SNOMEDCT_CORE|Aphasia as late effect of cerebrovascular disease|Aphasia as late effect of cerebrovascular disease
C0490017|T033|PT|430705002|SNOMEDCT_CORE|Family history of malignant neoplasm of ovary|Family history of malignant neoplasm of ovary
C0490017|T033|FN|430705002|SNOMEDCT_CORE|Family history of malignant neoplasm of ovary|Family history of malignant neoplasm of ovary
C0494165|T191|SY|94381002|SNOMEDCT_CORE|Cancer metastatic to liver|Secondary malignant neoplasm of liver
C0494165|T191|SY|94381002|SNOMEDCT_CORE|Hepatic metastasis|Secondary malignant neoplasm of liver
C0494165|T191|SY|94381002|SNOMEDCT_CORE|Liver secondaries|Secondary malignant neoplasm of liver
C0494165|T191|SY|94381002|SNOMEDCT_CORE|Liver secondary cancer|Secondary malignant neoplasm of liver
C0494165|T191|SY|94381002|SNOMEDCT_CORE|Metastasis to liver|Secondary malignant neoplasm of liver
C0494165|T191|SY|94381002|SNOMEDCT_CORE|Metastatic malignant neoplasm to liver|Secondary malignant neoplasm of liver
C0494165|T191|IS|94381002|SNOMEDCT_CORE|Metastatic malignant neoplasm to liver, NOS|Secondary malignant neoplasm of liver
C0494165|T191|SY|94381002|SNOMEDCT_CORE|Secondary malignancy of liver|Secondary malignant neoplasm of liver
C0494165|T191|PT|94381002|SNOMEDCT_CORE|Secondary malignant neoplasm of liver|Secondary malignant neoplasm of liver
C0494165|T191|FN|94381002|SNOMEDCT_CORE|Secondary malignant neoplasm of liver|Secondary malignant neoplasm of liver
C0494165|T191|IS|94381002|SNOMEDCT_CORE|Secondary malignant neoplasm of liver, NOS|Secondary malignant neoplasm of liver
C0494290|T047|IS|313436004|SNOMEDCT_CORE|Non-insulin-dependent diabetes mellitus without complication|Type 2 diabetes mellitus without complication
C0494290|T047|PT|313436004|SNOMEDCT_CORE|Type 2 diabetes mellitus without complication|Type 2 diabetes mellitus without complication
C0494290|T047|FN|313436004|SNOMEDCT_CORE|Type II diabetes mellitus without complication|Type 2 diabetes mellitus without complication
C0494290|T047|SY|313436004|SNOMEDCT_CORE|Type II diabetes mellitus without complication|Type 2 diabetes mellitus without complication
C0494463|T048|IS|66108005|SNOMEDCT_CORE|Alzheimer's disease with late onset|Primary degenerative dementia of the Alzheimer type, senile onset
C0494463|T048|SY|416975007|SNOMEDCT_CORE|Alzheimer's disease with late onset|Primary degenerative dementia of the Alzheimer type, senile onset
C0494463|T048|IS|66108005|SNOMEDCT_CORE|Dementia in Alzheimer's disease - type 1|Primary degenerative dementia of the Alzheimer type, senile onset
C0494463|T048|SY|416975007|SNOMEDCT_CORE|Dementia in Alzheimer's disease - type 1|Primary degenerative dementia of the Alzheimer type, senile onset
C0494463|T048|IS|66108005|SNOMEDCT_CORE|Dementia in Alzheimer's disease with late onset|Primary degenerative dementia of the Alzheimer type, senile onset
C0494463|T048|SY|416975007|SNOMEDCT_CORE|Dementia in Alzheimer's disease with late onset|Primary degenerative dementia of the Alzheimer type, senile onset
C0494463|T048|SY|416975007|SNOMEDCT_CORE|Dementia of the Alzheimers type, late onset|Primary degenerative dementia of the Alzheimer type, senile onset
C0494463|T048|SY|416975007|SNOMEDCT_CORE|Primary degenerative dementia of the Alzheimer type, late onset|Primary degenerative dementia of the Alzheimer type, senile onset
C0494463|T048|PT|416975007|SNOMEDCT_CORE|Primary degenerative dementia of the Alzheimer type, senile onset|Primary degenerative dementia of the Alzheimer type, senile onset
C0494463|T048|FN|416975007|SNOMEDCT_CORE|Primary degenerative dementia of the Alzheimer type, senile onset|Primary degenerative dementia of the Alzheimer type, senile onset
C0494463|T048|IS|66108005|SNOMEDCT_CORE|SDAT - Senile dementia, Alzheimer's type|Primary degenerative dementia of the Alzheimer type, senile onset
C0494463|T048|SY|416975007|SNOMEDCT_CORE|SDAT - Senile dementia, Alzheimer's type|Primary degenerative dementia of the Alzheimer type, senile onset
C0494475|T047|SY|54200006|SNOMEDCT_CORE|Grand mal convulsion|Tonic-clonic seizure
C0494475|T047|SY|54200006|SNOMEDCT_CORE|Grand mal seizure|Tonic-clonic seizure
C0494475|T047|SY|54200006|SNOMEDCT_CORE|Tonic-clonic convulsion|Tonic-clonic seizure
C0494475|T047|PT|54200006|SNOMEDCT_CORE|Tonic-clonic seizure|Tonic-clonic seizure
C0494475|T047|FN|54200006|SNOMEDCT_CORE|Tonic-clonic seizure|Tonic-clonic seizure
C0494475|T047|SY|54200006|SNOMEDCT_CORE|Tonic-clonic seizures|Tonic-clonic seizure
C0494575|T047|PT|194779001|SNOMEDCT_CORE|Hypertensive heart and renal disease with heart failure|Hypertensive heart and renal disease with heart failure
C0494575|T047|FN|194779001|SNOMEDCT_CORE|Hypertensive heart and renal disease with heart failure|Hypertensive heart and renal disease with heart failure
C0494576|T047|PT|194781004|SNOMEDCT_CORE|Hypertensive heart and renal disease with both heart failure and renal failure|Hypertensive heart and renal disease with both heart failure and renal failure
C0494576|T047|FN|194781004|SNOMEDCT_CORE|Hypertensive heart and renal disease with both heart failure and renal failure|Hypertensive heart and renal disease with both heart failure and renal failure
C0494698|T047|SY|371136004|SNOMEDCT_CORE|Abnormal tooth development|Disorder of tooth development
C0494698|T047|PT|371136004|SNOMEDCT_CORE|Disorder of tooth development|Disorder of tooth development
C0494698|T047|FN|371136004|SNOMEDCT_CORE|Disorder of tooth development|Disorder of tooth development
C0494809|T046|PT|235821002|SNOMEDCT_CORE|Postoperative intestinal obstruction|Postoperative intestinal obstruction
C0494809|T046|FN|235821002|SNOMEDCT_CORE|Postoperative intestinal obstruction|Postoperative intestinal obstruction
C0494809|T046|SY|235821002|SNOMEDCT_CORE|Postprocedural intestinal obstruction|Postoperative intestinal obstruction
C0495188|T046|SY|307534009|SNOMEDCT_CORE|Urinary tract infection complicating pregnancy|Urinary tract infection in pregnancy
C0495188|T046|PT|307534009|SNOMEDCT_CORE|Urinary tract infection in pregnancy|Urinary tract infection in pregnancy
C0495188|T046|FN|307534009|SNOMEDCT_CORE|Urinary tract infection in pregnancy|Urinary tract infection in pregnancy
C0495188|T046|SY|307534009|SNOMEDCT_CORE|UTI - urinary tract infection in pregnancy|Urinary tract infection in pregnancy
C0495194|T033|PT|199732004|SNOMEDCT_CORE|Abnormal findings on antenatal screening of mother|Abnormal findings on antenatal screening of mother
C0495194|T033|FN|199732004|SNOMEDCT_CORE|Abnormal findings on antenatal screening of mother|Abnormal findings on antenatal screening of mother
C0495524|T019|PT|275519006|SNOMEDCT_CORE|Peripheral arteriovenous malformation|Peripheral arteriovenous malformation
C0495524|T019|FN|275519006|SNOMEDCT_CORE|Peripheral arteriovenous malformation|Peripheral arteriovenous malformation
C0495676|T033|PT|274719002|SNOMEDCT_CORE|Intra-abdominal and pelvic swelling, mass and lump|Intra-abdominal and pelvic swelling, mass and lump
C0495676|T033|FN|274719002|SNOMEDCT_CORE|Intra-abdominal and pelvic swelling, mass and lump|Intra-abdominal and pelvic swelling, mass and lump
C0495786|T033|PT|274533004|SNOMEDCT_CORE|Abnormal findings on diagnostic imaging of lung|Abnormal findings on diagnostic imaging of lung
C0495786|T033|FN|274533004|SNOMEDCT_CORE|Abnormal findings on diagnostic imaging of lung|Abnormal findings on diagnostic imaging of lung
C0495868|T037|PT|307731004|SNOMEDCT_CORE|Injury of tendon of the rotator cuff of shoulder|Injury of tendon of the rotator cuff of shoulder
C0495868|T037|FN|307731004|SNOMEDCT_CORE|Injury of tendon of the rotator cuff of shoulder|Injury of tendon of the rotator cuff of shoulder
C0495958|T037|PT|125602001|SNOMEDCT_CORE|Injury of lower leg|Injury of lower leg
C0495958|T037|FN|125602001|SNOMEDCT_CORE|Injury of lower leg|Injury of lower leg
C0496779|T191|PT|363411007|SNOMEDCT_CORE|Malignant tumor of appendix|Malignant tumor of appendix
C0496779|T191|FN|363411007|SNOMEDCT_CORE|Malignant tumor of appendix|Malignant tumor of appendix
C0496779|T191|PTGB|363411007|SNOMEDCT_CORE|Malignant tumour of appendix|Malignant tumor of appendix
C0496797|T191|SY|372126009|SNOMEDCT_CORE|Ca skin - trunk|Malignant neoplasm of skin of trunk
C0496797|T191|PT|372126009|SNOMEDCT_CORE|Malignant neoplasm of skin of trunk|Malignant neoplasm of skin of trunk
C0496797|T191|FN|372126009|SNOMEDCT_CORE|Malignant neoplasm of skin of trunk|Malignant neoplasm of skin of trunk
C0496826|T191|SY|188239000|SNOMEDCT_CORE|Malignant neoplasm of trigone of urinary bladder|Malignant tumor of trigone of urinary bladder
C0496826|T191|SY|188239000|SNOMEDCT_CORE|Malignant tumor of trigone of bladder|Malignant tumor of trigone of urinary bladder
C0496826|T191|PT|188239000|SNOMEDCT_CORE|Malignant tumor of trigone of urinary bladder|Malignant tumor of trigone of urinary bladder
C0496826|T191|FN|188239000|SNOMEDCT_CORE|Malignant tumor of trigone of urinary bladder|Malignant tumor of trigone of urinary bladder
C0496826|T191|SYGB|188239000|SNOMEDCT_CORE|Malignant tumour of trigone of bladder|Malignant tumor of trigone of urinary bladder
C0496826|T191|PTGB|188239000|SNOMEDCT_CORE|Malignant tumour of trigone of urinary bladder|Malignant tumor of trigone of urinary bladder
C0496827|T191|SY|188240003|SNOMEDCT_CORE|Malignant neoplasm of dome of urinary bladder|Malignant tumor of vault of bladder
C0496827|T191|SY|188240003|SNOMEDCT_CORE|Malignant neoplasm of vault of bladder|Malignant tumor of vault of bladder
C0496827|T191|SY|188240003|SNOMEDCT_CORE|Malignant tumor of bladder dome|Malignant tumor of vault of bladder
C0496827|T191|PT|188240003|SNOMEDCT_CORE|Malignant tumor of vault of bladder|Malignant tumor of vault of bladder
C0496827|T191|FN|188240003|SNOMEDCT_CORE|Malignant tumor of vault of bladder|Malignant tumor of vault of bladder
C0496827|T191|SYGB|188240003|SNOMEDCT_CORE|Malignant tumour of bladder dome|Malignant tumor of vault of bladder
C0496827|T191|PTGB|188240003|SNOMEDCT_CORE|Malignant tumour of vault of bladder|Malignant tumor of vault of bladder
C0496828|T191|PT|188241004|SNOMEDCT_CORE|Malignant neoplasm of lateral wall of urinary bladder|Malignant neoplasm of lateral wall of urinary bladder
C0496828|T191|FN|188241004|SNOMEDCT_CORE|Malignant neoplasm of lateral wall of urinary bladder|Malignant neoplasm of lateral wall of urinary bladder
C0496899|T191|SY|92030004|SNOMEDCT_CORE|Benign brain tumor|Benign neoplasm of brain
C0496899|T191|SYGB|92030004|SNOMEDCT_CORE|Benign brain tumour|Benign neoplasm of brain
C0496899|T191|PT|92030004|SNOMEDCT_CORE|Benign neoplasm of brain|Benign neoplasm of brain
C0496899|T191|FN|92030004|SNOMEDCT_CORE|Benign neoplasm of brain|Benign neoplasm of brain
C0496899|T191|IS|92030004|SNOMEDCT_CORE|Benign neoplasm of brain, NOS|Benign neoplasm of brain
C0496901|T191|PT|92296004|SNOMEDCT_CORE|Benign neoplasm of pituitary gland|Benign neoplasm of pituitary gland
C0496901|T191|FN|92296004|SNOMEDCT_CORE|Benign neoplasm of pituitary gland|Benign neoplasm of pituitary gland
C0496901|T191|SY|92296004|SNOMEDCT_CORE|Benign tumor of pituitary gland|Benign neoplasm of pituitary gland
C0496901|T191|SYGB|92296004|SNOMEDCT_CORE|Benign tumour of pituitary gland|Benign neoplasm of pituitary gland
C0496927|T191|PT|94889006|SNOMEDCT_CORE|Neoplasm of uncertain behavior of kidney|Neoplasm of uncertain behavior of kidney
C0496927|T191|FN|94889006|SNOMEDCT_CORE|Neoplasm of uncertain behavior of kidney|Neoplasm of uncertain behavior of kidney
C0496927|T191|IS|94889006|SNOMEDCT_CORE|Neoplasm of uncertain behavior of kidney, NOS|Neoplasm of uncertain behavior of kidney
C0496927|T191|PTGB|94889006|SNOMEDCT_CORE|Neoplasm of uncertain behaviour of kidney|Neoplasm of uncertain behavior of kidney
C0496927|T191|SY|94889006|SNOMEDCT_CORE|Renal neoplasm of uncertain behavior|Neoplasm of uncertain behavior of kidney
C0496927|T191|SYGB|94889006|SNOMEDCT_CORE|Renal neoplasm of uncertain behaviour|Neoplasm of uncertain behavior of kidney
C0496930|T191|PT|94754000|SNOMEDCT_CORE|Neoplasm of uncertain behavior of bladder|Neoplasm of uncertain behavior of bladder
C0496930|T191|FN|94754000|SNOMEDCT_CORE|Neoplasm of uncertain behavior of bladder|Neoplasm of uncertain behavior of bladder
C0496930|T191|IS|94754000|SNOMEDCT_CORE|Neoplasm of uncertain behavior of bladder, NOS|Neoplasm of uncertain behavior of bladder
C0496930|T191|PTGB|94754000|SNOMEDCT_CORE|Neoplasm of uncertain behaviour of bladder|Neoplasm of uncertain behavior of bladder
C0496950|T191|PT|94820008|SNOMEDCT_CORE|Neoplasm of uncertain behavior of endocrine gland|Neoplasm of uncertain behavior of endocrine gland
C0496950|T191|FN|94820008|SNOMEDCT_CORE|Neoplasm of uncertain behavior of endocrine gland|Neoplasm of uncertain behavior of endocrine gland
C0496950|T191|IS|94820008|SNOMEDCT_CORE|Neoplasm of uncertain behavior of endocrine gland, NOS|Neoplasm of uncertain behavior of endocrine gland
C0496950|T191|PTGB|94820008|SNOMEDCT_CORE|Neoplasm of uncertain behaviour of endocrine gland|Neoplasm of uncertain behavior of endocrine gland
C0496955|T191|PT|95087004|SNOMEDCT_CORE|Neoplasm of uncertain behavior of skin|Neoplasm of uncertain behavior of skin
C0496955|T191|FN|95087004|SNOMEDCT_CORE|Neoplasm of uncertain behavior of skin|Neoplasm of uncertain behavior of skin
C0496955|T191|IS|95087004|SNOMEDCT_CORE|Neoplasm of uncertain behavior of skin, NOS|Neoplasm of uncertain behavior of skin
C0496955|T191|PTGB|95087004|SNOMEDCT_CORE|Neoplasm of uncertain behaviour of skin|Neoplasm of uncertain behavior of skin
C0497156|T047|IS|30746006|SNOMEDCT_CORE|Enlarged glands|Lymphadenopathy
C0497156|T047|SY|30746006|SNOMEDCT_CORE|Enlargement of lymph nodes|Lymphadenopathy
C0497156|T047|IS|30746006|SNOMEDCT_CORE|Enlargement of lymph nodes, NOS|Lymphadenopathy
C0497156|T047|SY|30746006|SNOMEDCT_CORE|LA - Lymphadenopathy|Lymphadenopathy
C0497156|T047|SY|30746006|SNOMEDCT_CORE|LN - Lymphadenopathy|Lymphadenopathy
C0497156|T047|FN|30746006|SNOMEDCT_CORE|Lymphadenopathy|Lymphadenopathy
C0497156|T047|PT|30746006|SNOMEDCT_CORE|Lymphadenopathy|Lymphadenopathy
C0497156|T047|SY|30746006|SNOMEDCT_CORE|Lymphadenopathy - swelling|Lymphadenopathy
C0497156|T047|IS|30746006|SNOMEDCT_CORE|Lymphadenopathy, NOS|Lymphadenopathy
C0497156|T047|SY|30746006|SNOMEDCT_CORE|Swelling of lymph node|Lymphadenopathy
C0497156|T047|SY|30746006|SNOMEDCT_CORE|Swelling of lymph nodes|Lymphadenopathy
C0497156|T047|IS|30746006|SNOMEDCT_CORE|Swelling of lymph nodes, NOS|Lymphadenopathy
C0497156|T047|IS|30746006|SNOMEDCT_CORE|Swollen glands|Lymphadenopathy
C0497156|T047|SY|30746006|SNOMEDCT_CORE|Swollen lymph glands|Lymphadenopathy
C0497156|T047|SY|30746006|SNOMEDCT_CORE|Swollen lymph nodes|Lymphadenopathy
C0497156|T047|IS|30746006|SNOMEDCT_CORE|Unspecified lymphadenopathy|Lymphadenopathy
C0497247|T033|IS|38341003|SNOMEDCT_CORE|Elevated blood pressure|Elevated blood pressure
C0497247|T033|IS|38341003|SNOMEDCT_CORE|Raised blood pressure|Elevated blood pressure
C0497327|T048|PT|52448006|SNOMEDCT_CORE|Dementia|Dementia
C0497327|T048|FN|52448006|SNOMEDCT_CORE|Dementia|Dementia
C0497327|T048|IS|52448006|SNOMEDCT_CORE|Dementia, NOS|Dementia
C0497327|T048|SY|52448006|SNOMEDCT_CORE|Organic dementia|Dementia
C0497406|T033|PT|238131007|SNOMEDCT_CORE|Overweight|Overweight
C0497406|T033|FN|238131007|SNOMEDCT_CORE|Overweight|Overweight
C0497406|T033|SY|238131007|SNOMEDCT_CORE|Patient overweight|Overweight
C0497481|T184|PT|285375003|SNOMEDCT_CORE|Pain in penis|Pain in penis
C0497481|T184|FN|285375003|SNOMEDCT_CORE|Pain in penis|Pain in penis
C0497481|T184|SY|285375003|SNOMEDCT_CORE|Penile pain|Pain in penis
C0497552|T019|PT|88425004|SNOMEDCT_CORE|Congenital anomaly of nervous system|Congenital anomaly of nervous system
C0497552|T019|FN|88425004|SNOMEDCT_CORE|Congenital anomaly of nervous system|Congenital anomaly of nervous system
C0497552|T019|IS|88425004|SNOMEDCT_CORE|Congenital anomaly of nervous system, NOS|Congenital anomaly of nervous system
C0497552|T019|SY|88425004|SNOMEDCT_CORE|Congenital deformity of nervous system|Congenital anomaly of nervous system
C0497552|T019|IS|88425004|SNOMEDCT_CORE|Congenital deformity of nervous system, NOS|Congenital anomaly of nervous system
C0497552|T019|SY|88425004|SNOMEDCT_CORE|Congenital disease of nervous system|Congenital anomaly of nervous system
C0497552|T019|IS|88425004|SNOMEDCT_CORE|Congenital disease of nervous system, NOS|Congenital anomaly of nervous system
C0497552|T019|SY|88425004|SNOMEDCT_CORE|Congenital lesion of nervous system|Congenital anomaly of nervous system
C0497552|T019|IS|88425004|SNOMEDCT_CORE|Congenital lesion of nervous system, NOS|Congenital anomaly of nervous system
C0497552|T019|SY|88425004|SNOMEDCT_CORE|Congenital malformation of the nervous system|Congenital anomaly of nervous system
C0497556|T191|PT|255166003|SNOMEDCT_CORE|Benign neoplasm of respiratory system|Benign neoplasm of respiratory system
C0497556|T191|FN|255166003|SNOMEDCT_CORE|Benign neoplasm of respiratory system|Benign neoplasm of respiratory system
C0518456|T033|PT|82971005|SNOMEDCT_CORE|Impaired mobility|Impaired mobility
C0518456|T033|FN|82971005|SNOMEDCT_CORE|Impaired mobility|Impaired mobility
C0518456|T033|IS|82971005|SNOMEDCT_CORE|Impaired physical mobility|Impaired mobility
C0518456|T033|SY|82971005|SNOMEDCT_CORE|Physical mobility impairment|Impaired mobility
C0518988|T047|PT|299709002|SNOMEDCT_CORE|Dental abscess|Dental abscess
C0518988|T047|FN|299709002|SNOMEDCT_CORE|Dental abscess|Dental abscess
C0518988|T047|SY|299709002|SNOMEDCT_CORE|Dental sepsis|Dental abscess
C0518988|T047|SY|299709002|SNOMEDCT_CORE|Tooth abscess|Dental abscess
C0519030|T047|SY|64479007|SNOMEDCT_CORE|Pneumonia caused by Klebsiella pneumoniae|Pneumonia due to Klebsiella pneumoniae
C0519030|T047|FN|64479007|SNOMEDCT_CORE|Pneumonia caused by Klebsiella pneumoniae|Pneumonia due to Klebsiella pneumoniae
C0519030|T047|PT|64479007|SNOMEDCT_CORE|Pneumonia due to Klebsiella pneumoniae|Pneumonia due to Klebsiella pneumoniae
C0519030|T047|OF|64479007|SNOMEDCT_CORE|Pneumonia due to Klebsiella pneumoniae|Pneumonia due to Klebsiella pneumoniae
C0520463|T047|SY|197284004|SNOMEDCT_CORE|CAH - Chronic active hepatitis|Chronic active hepatitis
C0520463|T047|SY|197284004|SNOMEDCT_CORE|CAH - Chronic aggressive hepatitis|Chronic active hepatitis
C0520463|T047|PT|197284004|SNOMEDCT_CORE|Chronic active hepatitis|Chronic active hepatitis
C0520463|T047|FN|197284004|SNOMEDCT_CORE|Chronic active hepatitis|Chronic active hepatitis
C0520474|T046|PT|398199007|SNOMEDCT_CORE|Aseptic necrosis of bone|Aseptic necrosis of bone
C0520474|T046|FN|398199007|SNOMEDCT_CORE|Aseptic necrosis of bone|Aseptic necrosis of bone
C0520477|T191|IS|266569009|SNOMEDCT_CORE|Benign adenoma of prostate|Benign adenoma of prostate
C0520482|T048|PTGB|397923000|SNOMEDCT_CORE|Somatisation disorder|Somatization disorder
C0520482|T048|PT|397923000|SNOMEDCT_CORE|Somatization disorder|Somatization disorder
C0520482|T048|FN|397923000|SNOMEDCT_CORE|Somatization disorder|Somatization disorder
C0520556|T190|SY|76545008|SNOMEDCT_CORE|Pilonidal cyst with no abscess|Pilonidal cyst without abscess
C0520556|T190|PT|76545008|SNOMEDCT_CORE|Pilonidal cyst without abscess|Pilonidal cyst without abscess
C0520556|T190|FN|76545008|SNOMEDCT_CORE|Pilonidal cyst without abscess|Pilonidal cyst without abscess
C0520556|T190|IS|76545008|SNOMEDCT_CORE|Pilonidal cyst without mention of abscess|Pilonidal cyst without abscess
C0520556|T190|IS|47639008|SNOMEDCT_CORE|Pilonidal cyst without mention of abscess|Pilonidal cyst without abscess
C0520560|T047|PTGB|60698006|SNOMEDCT_CORE|Haemorrhagic oesophagitis|Hemorrhagic esophagitis
C0520560|T047|PT|60698006|SNOMEDCT_CORE|Hemorrhagic esophagitis|Hemorrhagic esophagitis
C0520560|T047|FN|60698006|SNOMEDCT_CORE|Hemorrhagic esophagitis|Hemorrhagic esophagitis
C0520575|T047|SY|36689008|SNOMEDCT_CORE|Acute kidney infection|Acute pyelonephritis
C0520575|T047|SY|36689008|SNOMEDCT_CORE|Acute PN - pyelonephritis|Acute pyelonephritis
C0520575|T047|PT|36689008|SNOMEDCT_CORE|Acute pyelonephritis|Acute pyelonephritis
C0520575|T047|FN|36689008|SNOMEDCT_CORE|Acute pyelonephritis|Acute pyelonephritis
C0520575|T047|SY|36689008|SNOMEDCT_CORE|APN - Acute pyelonephritis|Acute pyelonephritis
C0520578|T019|SY|21779006|SNOMEDCT_CORE|Pseudocryptorchism|Retractile testis
C0520578|T019|SY|21779006|SNOMEDCT_CORE|Retractible testis|Retractile testis
C0520578|T019|PT|21779006|SNOMEDCT_CORE|Retractile testis|Retractile testis
C0520578|T019|FN|21779006|SNOMEDCT_CORE|Retractile testis|Retractile testis
C0520578|T019|IS|21779006|SNOMEDCT_CORE|Retraction of testis|Retractile testis
C0520578|T019|SY|21779006|SNOMEDCT_CORE|Testicular retraction|Retractile testis
C0520594|T046|PT|44771000|SNOMEDCT_CORE|Microcalcifications of the breast|Microcalcifications of the breast
C0520594|T046|FN|44771000|SNOMEDCT_CORE|Microcalcifications of the breast|Microcalcifications of the breast
C0520602|T047|IS|21584002|SNOMEDCT_CORE|Maternal diabetes mellitus with hypoglycemia affecting fetus or newborn|Maternal diabetes mellitus with hypoglycemia affecting fetus or newborn
C0520627|T048|SY|35481005|SNOMEDCT_CORE|Bipolar I disorder, most recent episode mixed, in remission|Mixed bipolar I disorder in remission
C0520627|T048|IS|35481005|SNOMEDCT_CORE|Mixed bipolar disorder in remission|Mixed bipolar I disorder in remission
C0520627|T048|PT|35481005|SNOMEDCT_CORE|Mixed bipolar I disorder in remission|Mixed bipolar I disorder in remission
C0520627|T048|FN|35481005|SNOMEDCT_CORE|Mixed bipolar I disorder in remission|Mixed bipolar I disorder in remission
C0520676|T048|PT|596004|SNOMEDCT_CORE|Premenstrual dysphoric disorder|Premenstrual dysphoric disorder
C0520676|T048|FN|596004|SNOMEDCT_CORE|Premenstrual dysphoric disorder|Premenstrual dysphoric disorder
C0520679|T047|SY|78275009|SNOMEDCT_CORE|Obstructive sleep apnea|Obstructive sleep apnea syndrome
C0520679|T047|PT|78275009|SNOMEDCT_CORE|Obstructive sleep apnea syndrome|Obstructive sleep apnea syndrome
C0520679|T047|FN|78275009|SNOMEDCT_CORE|Obstructive sleep apnea syndrome|Obstructive sleep apnea syndrome
C0520679|T047|SYGB|78275009|SNOMEDCT_CORE|Obstructive sleep apnoea|Obstructive sleep apnea syndrome
C0520679|T047|PTGB|78275009|SNOMEDCT_CORE|Obstructive sleep apnoea syndrome|Obstructive sleep apnea syndrome
C0520679|T047|SY|78275009|SNOMEDCT_CORE|OSA - Obstructive sleep apnea|Obstructive sleep apnea syndrome
C0520679|T047|SYGB|78275009|SNOMEDCT_CORE|OSA - Obstructive sleep apnoea|Obstructive sleep apnea syndrome
C0520743|T047|PT|52324001|SNOMEDCT_CORE|Mediastinal lymphadenopathy|Mediastinal lymphadenopathy
C0520743|T047|FN|52324001|SNOMEDCT_CORE|Mediastinal lymphadenopathy|Mediastinal lymphadenopathy
C0520753|T033|SY|14448006|SNOMEDCT_CORE|Ingestion of foreign body|Swallowed foreign body
C0520753|T033|IS|33334006|SNOMEDCT_CORE|Swallowed foreign body|Swallowed foreign body
C0520753|T033|PT|14448006|SNOMEDCT_CORE|Swallowed foreign body|Swallowed foreign body
C0520753|T033|FN|14448006|SNOMEDCT_CORE|Swallowed foreign body|Swallowed foreign body
C0520770|T047|PT|6185008|SNOMEDCT_CORE|Helicobacter-associated disease|Helicobacter-associated disease
C0520770|T047|FN|6185008|SNOMEDCT_CORE|Helicobacter-associated disease|Helicobacter-associated disease
C0520770|T047|IS|6185008|SNOMEDCT_CORE|Helicobacter-associated disease, NOS|Helicobacter-associated disease
C0520863|T046|PT|3545003|SNOMEDCT_CORE|Diastolic dysfunction|Diastolic dysfunction
C0520863|T046|FN|3545003|SNOMEDCT_CORE|Diastolic dysfunction|Diastolic dysfunction
C0520955|T033|IS|1855002|SNOMEDCT_CORE|Learning delay|Slow learner
C0520955|T033|IS|1855002|SNOMEDCT_CORE|Slow learner|Slow learner
C0520962|T184|PTGB|112104007|SNOMEDCT_CORE|Localised pain|Localized pain
C0520962|T184|PT|112104007|SNOMEDCT_CORE|Localized pain|Localized pain
C0520962|T184|FN|112104007|SNOMEDCT_CORE|Localized pain|Localized pain
C0520966|T033|SY|302289002|SNOMEDCT_CORE|Abnormal coordination|Coordination problem
C0520966|T033|PT|302289002|SNOMEDCT_CORE|Coordination problem|Coordination problem
C0520966|T033|FN|302289002|SNOMEDCT_CORE|Coordination problem|Coordination problem
C0521168|T037|PT|371128008|SNOMEDCT_CORE|Occupational injury|Occupational injury
C0521168|T037|FN|371128008|SNOMEDCT_CORE|Occupational injury|Occupational injury
C0521169|T046|PT|443395009|SNOMEDCT_CORE|Compression fracture|Compression fracture
C0521169|T046|PT|21947006|SNOMEDCT_CORE|Compression fracture|Compression fracture
C0521169|T046|FN|21947006|SNOMEDCT_CORE|Compression fracture|Compression fracture
C0521169|T046|FN|443395009|SNOMEDCT_CORE|Compression fracture|Compression fracture
C0521170|T047|PT|46675001|SNOMEDCT_CORE|Osteoporotic fracture|Osteoporotic fracture
C0521170|T047|FN|46675001|SNOMEDCT_CORE|Osteoporotic fracture|Osteoporotic fracture
C0521173|T047|PT|443138004|SNOMEDCT_CORE|Granulomatosis|Granulomatosis
C0521173|T047|PT|44328006|SNOMEDCT_CORE|Granulomatosis|Granulomatosis
C0521173|T047|FN|44328006|SNOMEDCT_CORE|Granulomatosis|Granulomatosis
C0521173|T047|FN|443138004|SNOMEDCT_CORE|Granulomatosis|Granulomatosis
C0521173|T047|IS|44328006|SNOMEDCT_CORE|Granulomatosis, NOS|Granulomatosis
C0521208|T037|SY|79573009|SNOMEDCT_CORE|Accident at home|Accident while engaged in household activity
C0521208|T037|IS|79573009|SNOMEDCT_CORE|Accident at home, NOS|Accident while engaged in household activity
C0521208|T037|PT|79573009|SNOMEDCT_CORE|Accident while engaged in household activity|Accident while engaged in household activity
C0521208|T037|OF|79573009|SNOMEDCT_CORE|Accident while engaged in household activity|Accident while engaged in household activity
C0521208|T037|FN|79573009|SNOMEDCT_CORE|Accident while engaged in household activity|Accident while engaged in household activity
C0521208|T037|IS|79573009|SNOMEDCT_CORE|Accident while engaged in household activity, NOS|Accident while engaged in household activity
C0521208|T037|PTGB|79573009|SNOMEDCT_CORE|Accident whilst engaged in household activity|Accident while engaged in household activity
C0521208|T037|SY|79573009|SNOMEDCT_CORE|Household accident|Accident while engaged in household activity
C0521208|T037|IS|79573009|SNOMEDCT_CORE|Household accident, NOS|Accident while engaged in household activity
C0521516|T184|PT|95415006|SNOMEDCT_CORE|Polymyalgia|Polymyalgia
C0521516|T184|FN|95415006|SNOMEDCT_CORE|Polymyalgia|Polymyalgia
C0521516|T184|IS|95415006|SNOMEDCT_CORE|Polymyalgia, NOS|Polymyalgia
C0521518|T046|IS|95418008|SNOMEDCT_CORE|Muscle spasms of head and neck|Muscle spasms of head AND/OR neck
C0521518|T046|PT|95418008|SNOMEDCT_CORE|Muscle spasms of head AND/OR neck|Muscle spasms of head AND/OR neck
C0521518|T046|FN|95418008|SNOMEDCT_CORE|Muscle spasms of head AND/OR neck|Muscle spasms of head AND/OR neck
C0521578|T019|PT|95508001|SNOMEDCT_CORE|Congenital obstruction of lacrimal canal|Congenital obstruction of lacrimal canal
C0521578|T019|FN|95508001|SNOMEDCT_CORE|Congenital obstruction of lacrimal canal|Congenital obstruction of lacrimal canal
C0521595|T046|PTGB|95533003|SNOMEDCT_CORE|Duodenal haemorrhage|Duodenal hemorrhage
C0521595|T046|PT|95533003|SNOMEDCT_CORE|Duodenal hemorrhage|Duodenal hemorrhage
C0521595|T046|FN|95533003|SNOMEDCT_CORE|Duodenal hemorrhage|Duodenal hemorrhage
C0521595|T046|IS|95533003|SNOMEDCT_CORE|Duodenal hemorrhage, NOS|Duodenal hemorrhage
C0521614|T047|PT|95563007|SNOMEDCT_CORE|Gallstone pancreatitis|Gallstone pancreatitis
C0521614|T047|FN|95563007|SNOMEDCT_CORE|Gallstone pancreatitis|Gallstone pancreatitis
C0521618|T190|PT|95574003|SNOMEDCT_CORE|Stenosis of ureter|Stenosis of ureter
C0521618|T190|FN|95574003|SNOMEDCT_CORE|Stenosis of ureter|Stenosis of ureter
C0521618|T190|SY|95574003|SNOMEDCT_CORE|Ureteral stenosis|Stenosis of ureter
C0521618|T190|SY|95574003|SNOMEDCT_CORE|Ureteric stenosis|Stenosis of ureter
C0521619|T046|PT|95575002|SNOMEDCT_CORE|Obstruction of pelviureteric junction|Obstruction of pelviureteric junction
C0521619|T046|FN|95575002|SNOMEDCT_CORE|Obstruction of pelviureteric junction|Obstruction of pelviureteric junction
C0521619|T046|SY|95575002|SNOMEDCT_CORE|Pelviureteric obstruction|Obstruction of pelviureteric junction
C0521619|T046|SY|95575002|SNOMEDCT_CORE|PUJ - Pelviureteric obstruction|Obstruction of pelviureteric junction
C0521619|T046|SY|95575002|SNOMEDCT_CORE|PUO - Pelviureteric obstruction|Obstruction of pelviureteric junction
C0521619|T046|SY|95575002|SNOMEDCT_CORE|UPJ - Ureteropelvic obstruction|Obstruction of pelviureteric junction
C0521619|T046|SY|95575002|SNOMEDCT_CORE|Ureteropelvic obstruction|Obstruction of pelviureteric junction
C0521622|T047|PT|95581005|SNOMEDCT_CORE|Bilateral hydronephrosis|Bilateral hydronephrosis
C0521622|T047|FN|95581005|SNOMEDCT_CORE|Bilateral hydronephrosis|Bilateral hydronephrosis
C0521665|T047|PT|95657009|SNOMEDCT_CORE|Chronic mixed headache syndrome|Chronic mixed headache syndrome
C0521665|T047|FN|95657009|SNOMEDCT_CORE|Chronic mixed headache syndrome|Chronic mixed headache syndrome
C0521687|T047|PTGB|95697007|SNOMEDCT_CORE|Generalised retinal degeneration|Generalized retinal degeneration
C0521687|T047|PT|95697007|SNOMEDCT_CORE|Generalized retinal degeneration|Generalized retinal degeneration
C0521687|T047|FN|95697007|SNOMEDCT_CORE|Generalized retinal degeneration|Generalized retinal degeneration
C0521707|T047|FN|95722004|SNOMEDCT_CORE|Bilateral cataracts|Bilateral cataracts
C0521707|T047|PT|95722004|SNOMEDCT_CORE|Bilateral cataracts|Bilateral cataracts
C0521707|T047|SY|95722004|SNOMEDCT_CORE|Cataracts|Bilateral cataracts
C0521723|T047|IS|373426005|SNOMEDCT_CORE|Anterior membrane corneal dystrophy|Anterior membrane corneal dystrophy
C0521723|T047|IS|373426005|SNOMEDCT_CORE|Basement membrane corneal dystrophy|Anterior membrane corneal dystrophy
C0521723|T047|SY|373426005|SNOMEDCT_CORE|Corneal epithelial and basement membrane dystrophy|Anterior membrane corneal dystrophy
C0521723|T047|OF|373426005|SNOMEDCT_CORE|Corneal epithelial and basement membrane dystrophy|Anterior membrane corneal dystrophy
C0521723|T047|IS|373426005|SNOMEDCT_CORE|Corneal epithelial dystrophy|Anterior membrane corneal dystrophy
C0521723|T047|SY|373426005|SNOMEDCT_CORE|EBMD - Epithelial basement membrane dystrophy|Anterior membrane corneal dystrophy
C0521723|T047|IS|373426005|SNOMEDCT_CORE|Epithelial corneal dystrophy|Anterior membrane corneal dystrophy
C0521730|T047|SY|414521009|SNOMEDCT_CORE|Infected chalazion|Infected cyst of meibomian gland
C0521730|T047|SY|414521009|SNOMEDCT_CORE|Infected cyst of meibomian gland|Infected cyst of meibomian gland
C0521730|T047|SY|414521009|SNOMEDCT_CORE|Infected meibomian cyst|Infected cyst of meibomian gland
C0521730|T047|SY|414521009|SNOMEDCT_CORE|Infection of meibomian gland|Infected cyst of meibomian gland
C0521730|T047|SY|414521009|SNOMEDCT_CORE|Meibomian adenitis|Infected cyst of meibomian gland
C0521770|T047|SY|95800001|SNOMEDCT_CORE|Asteroid hyalitis|Asteroid hyalosis
C0521770|T047|PT|95800001|SNOMEDCT_CORE|Asteroid hyalosis|Asteroid hyalosis
C0521770|T047|FN|95800001|SNOMEDCT_CORE|Asteroid hyalosis|Asteroid hyalosis
C0521770|T047|SY|95800001|SNOMEDCT_CORE|Benson's disease|Asteroid hyalosis
C0521839|T047|SY|95891005|SNOMEDCT_CORE|Flu-like illness|Influenza-like illness
C0521839|T047|SY|95891005|SNOMEDCT_CORE|Influenza like illness|Influenza-like illness
C0521839|T047|PT|95891005|SNOMEDCT_CORE|Influenza-like illness|Influenza-like illness
C0521839|T047|FN|95891005|SNOMEDCT_CORE|Influenza-like illness|Influenza-like illness
C0521861|T033|SY|95919007|SNOMEDCT_CORE|Corticodependence|Dependence on corticoids
C0521861|T033|PT|95919007|SNOMEDCT_CORE|Dependence on corticoids|Dependence on corticoids
C0521861|T033|FN|95919007|SNOMEDCT_CORE|Dependence on corticoids|Dependence on corticoids
C0521861|T033|SY|95919007|SNOMEDCT_CORE|Dependence on corticosteroids|Dependence on corticoids
C0522035|T046|PT|102558002|SNOMEDCT_CORE|Edema of the upper extremity|Edema of the upper extremity
C0522035|T046|FN|102558002|SNOMEDCT_CORE|Edema of the upper extremity|Edema of the upper extremity
C0522035|T046|PTGB|102558002|SNOMEDCT_CORE|Oedema of the upper extremity|Edema of the upper extremity
C0522055|T033|SY|102594003|SNOMEDCT_CORE|Abnormal ECG|Electrocardiogram abnormal
C0522055|T033|OF|102594003|SNOMEDCT_CORE|Abnormal ECG|Electrocardiogram abnormal
C0522055|T033|SY|102594003|SNOMEDCT_CORE|Abnormal EKG finding|Electrocardiogram abnormal
C0522055|T033|PT|102594003|SNOMEDCT_CORE|Electrocardiogram abnormal|Electrocardiogram abnormal
C0522055|T033|FN|102594003|SNOMEDCT_CORE|Electrocardiogram abnormal|Electrocardiogram abnormal
C0522224|T033|SY|44695005|SNOMEDCT_CORE|Palsy|Paralysis
C0522224|T033|PT|44695005|SNOMEDCT_CORE|Paralysis|Paralysis
C0522224|T033|FN|44695005|SNOMEDCT_CORE|Paralysis|Paralysis
C0522224|T033|IS|44695005|SNOMEDCT_CORE|Paralysis, NOS|Paralysis
C0522251|T184|SY|4969004|SNOMEDCT_CORE|Sinus pain|Sinus pain
C0522347|T184|OAS|103280006|SNOMEDCT_CORE|Ear pressure sensation|Ear pressure sensation
C0522347|T184|PT|162403009|SNOMEDCT_CORE|Ear pressure sensation|Ear pressure sensation
C0522347|T184|FN|162403009|SNOMEDCT_CORE|Ear pressure sensation|Ear pressure sensation
C0522347|T184|OAP|103280006|SNOMEDCT_CORE|Sensation of pressure in ear|Ear pressure sensation
C0522347|T184|OAF|103280006|SNOMEDCT_CORE|Sensation of pressure in ear|Ear pressure sensation
C0524385|T033|PT|105530003|SNOMEDCT_CORE|Living in residential institution|Living in residential institution
C0524385|T033|FN|105530003|SNOMEDCT_CORE|Living in residential institution|Living in residential institution
C0524528|T048|PT|35919005|SNOMEDCT_CORE|Autism spectrum disorder|Autism spectrum disorder
C0524528|T048|IS|35919005|SNOMEDCT_CORE|Autistic continuum|Autism spectrum disorder
C0524528|T048|IS|35919005|SNOMEDCT_CORE|Autistic spectrum disorder|Autism spectrum disorder
C0524528|T048|SY|35919005|SNOMEDCT_CORE|Pervasive developmental disorder|Autism spectrum disorder
C0524528|T048|FN|35919005|SNOMEDCT_CORE|Pervasive developmental disorder|Autism spectrum disorder
C0524528|T048|IS|35919005|SNOMEDCT_CORE|Pervasive developmental disorder, NOS|Autism spectrum disorder
C0524528|T048|IS|35919005|SNOMEDCT_CORE|PPD - Pervasive developmental disorder|Autism spectrum disorder
C0524620|T047|SY|237602007|SNOMEDCT_CORE|Dysmetabolic syndrome X|Metabolic syndrome X
C0524620|T047|SY|237602007|SNOMEDCT_CORE|Insulin resistance syndrome|Metabolic syndrome X
C0524620|T047|SY|237602007|SNOMEDCT_CORE|Metabolic syndrome|Metabolic syndrome X
C0524620|T047|PT|237602007|SNOMEDCT_CORE|Metabolic syndrome X|Metabolic syndrome X
C0524620|T047|FN|237602007|SNOMEDCT_CORE|Metabolic syndrome X|Metabolic syndrome X
C0524620|T047|SY|237602007|SNOMEDCT_CORE|Reaven's syndrome|Metabolic syndrome X
C0524662|T048|SY|75544000|SNOMEDCT_CORE|Narcotism|Opioid dependence
C0524662|T048|PT|75544000|SNOMEDCT_CORE|Opioid dependence|Opioid dependence
C0524662|T048|FN|75544000|SNOMEDCT_CORE|Opioid dependence|Opioid dependence
C0524909|T047|PT|61977001|SNOMEDCT_CORE|Chronic type B viral hepatitis|Chronic type B viral hepatitis
C0524909|T047|FN|61977001|SNOMEDCT_CORE|Chronic type B viral hepatitis|Chronic type B viral hepatitis
C0524909|T047|SY|61977001|SNOMEDCT_CORE|Chronic viral hepatitis B|Chronic type B viral hepatitis
C0524910|T047|PT|128302006|SNOMEDCT_CORE|Chronic hepatitis C|Chronic hepatitis C
C0524910|T047|FN|128302006|SNOMEDCT_CORE|Chronic hepatitis C|Chronic hepatitis C
C0524910|T047|SY|128302006|SNOMEDCT_CORE|Chronic type C viral hepatitis|Chronic hepatitis C
C0525045|T048|SY|46206005|SNOMEDCT_CORE|Affective disorder|Mood disorder
C0525045|T048|SY|46206005|SNOMEDCT_CORE|Disorder of affect|Mood disorder
C0525045|T048|PT|46206005|SNOMEDCT_CORE|Mood disorder|Mood disorder
C0525045|T048|FN|46206005|SNOMEDCT_CORE|Mood disorder|Mood disorder
C0525045|T048|IS|46206005|SNOMEDCT_CORE|Mood disorder, NOS|Mood disorder
C0541912|T191|PT|254570009|SNOMEDCT_CORE|Carcinoma of duodenum|Carcinoma of duodenum
C0541912|T191|FN|254570009|SNOMEDCT_CORE|Carcinoma of duodenum|Carcinoma of duodenum
C0541951|T184|PT|290113009|SNOMEDCT_CORE|Bloody nipple discharge|Bloody nipple discharge
C0541951|T184|FN|290113009|SNOMEDCT_CORE|Bloody nipple discharge|Bloody nipple discharge
C0541951|T184|SY|290113009|SNOMEDCT_CORE|Sanguinous nipple discharge|Bloody nipple discharge
C0542322|T047|OAP|410064000|SNOMEDCT_CORE|Non-traumatic subdural haematoma|Non-traumatic subdural haematoma
C0542322|T047|OAP|410064000|SNOMEDCT_CORE|Non-traumatic subdural hematoma|Non-traumatic subdural haematoma
C0542322|T047|OAF|410064000|SNOMEDCT_CORE|Non-traumatic subdural hematoma|Non-traumatic subdural haematoma
C0542322|T047|OAS|410064000|SNOMEDCT_CORE|Nontraumatic subdural haematoma|Non-traumatic subdural haematoma
C0542322|T047|OAS|410064000|SNOMEDCT_CORE|SDH - Non-traumatic subdural haematoma|Non-traumatic subdural haematoma
C0542322|T047|OAS|410064000|SNOMEDCT_CORE|SDH - Non-traumatic subdural hematoma|Non-traumatic subdural haematoma
C0542322|T047|OAS|410064000|SNOMEDCT_CORE|Subdural haematoma - nontraumatic|Non-traumatic subdural haematoma
C0542322|T047|OAS|410064000|SNOMEDCT_CORE|Subdural hematoma - nontraumatic|Non-traumatic subdural haematoma
C0542427|T047|PT|202907005|SNOMEDCT_CORE|Tenosynovitis of ankle|Tenosynovitis of ankle
C0542427|T047|FN|202907005|SNOMEDCT_CORE|Tenosynovitis of ankle|Tenosynovitis of ankle
C0542485|T033|PT|169958000|SNOMEDCT_CORE|Placenta incomplete|Placenta incomplete
C0542485|T033|FN|169958000|SNOMEDCT_CORE|Placenta incomplete|Placenta incomplete
C0542571|T046|PT|445088006|SNOMEDCT_CORE|Edema of face|Edema of face
C0542571|T046|FN|445088006|SNOMEDCT_CORE|Edema of face|Edema of face
C0542571|T046|PTGB|445088006|SNOMEDCT_CORE|Oedema of face|Edema of face
C0543891|T047|SY|38941006|SNOMEDCT_CORE|Neuroleptic induced tardive dyskinesia|Neuroleptic-induced tardive dyskinesia
C0543891|T047|PT|38941006|SNOMEDCT_CORE|Neuroleptic-induced tardive dyskinesia|Neuroleptic-induced tardive dyskinesia
C0543891|T047|FN|38941006|SNOMEDCT_CORE|Neuroleptic-induced tardive dyskinesia|Neuroleptic-induced tardive dyskinesia
C0543947|T048|PT|192041001|SNOMEDCT_CORE|Acute situational disturbance|Acute situational disturbance
C0543947|T048|FN|192041001|SNOMEDCT_CORE|Acute situational disturbance|Acute situational disturbance
C0543947|T048|IS|17226007|SNOMEDCT_CORE|Acute situational disturbance, NOS|Acute situational disturbance
C0544008|T047|PT|392481002|SNOMEDCT_CORE|Chandler syndrome|Chandler syndrome
C0544008|T047|FN|392481002|SNOMEDCT_CORE|Chandler syndrome|Chandler syndrome
C0544008|T047|IS|392481002|SNOMEDCT_CORE|Corneal endothelial dystrophy|Chandler syndrome
C0544008|T047|IS|392481002|SNOMEDCT_CORE|Dystrophy of corneal endothelium|Chandler syndrome
C0544008|T047|IS|392481002|SNOMEDCT_CORE|Endothelial corneal dystrophy|Chandler syndrome
C0544008|T047|OF|392481002|SNOMEDCT_CORE|Endothelial corneal dystrophy|Chandler syndrome
C0544755|T033|OAP|249782009|SNOMEDCT_CORE|Bowing of leg|Bowing of leg
C0544755|T033|OAF|249782009|SNOMEDCT_CORE|Bowing of leg|Bowing of leg
C0546817|T046|SY|21639008|SNOMEDCT_CORE|Fluid excess|Hypervolemia
C0546817|T046|SY|21639008|SNOMEDCT_CORE|Fluid overload|Hypervolemia
C0546817|T046|SY|21639008|SNOMEDCT_CORE|Fluid volume excess|Hypervolemia
C0546817|T046|PTGB|21639008|SNOMEDCT_CORE|Hypervolaemia|Hypervolemia
C0546817|T046|PT|21639008|SNOMEDCT_CORE|Hypervolemia|Hypervolemia
C0546817|T046|FN|21639008|SNOMEDCT_CORE|Hypervolemia|Hypervolemia
C0546817|T046|SY|21639008|SNOMEDCT_CORE|Volume excess|Hypervolemia
C0546826|T047|OAP|266151007|SNOMEDCT_CORE|Dermatophytosis of the body|Dermatophytosis of the body
C0546826|T047|OAF|266151007|SNOMEDCT_CORE|Dermatophytosis of the body|Dermatophytosis of the body
C0546826|T047|SY|84849002|SNOMEDCT_CORE|Dermatophytosis of the trunk|Dermatophytosis of the body
C0546830|T037|PT|217699002|SNOMEDCT_CORE|Bite of nonvenomous snakes and lizards|Bite of nonvenomous snakes and lizards
C0546830|T037|OF|217699002|SNOMEDCT_CORE|Bite of nonvenomous snakes and lizards|Bite of nonvenomous snakes and lizards
C0546830|T037|FN|217699002|SNOMEDCT_CORE|Bite of nonvenomous snakes and lizards|Bite of nonvenomous snakes and lizards
C0546837|T191|SY|363402007|SNOMEDCT_CORE|CA - Cancer of esophagus|Malignant tumor of esophagus
C0546837|T191|SYGB|363402007|SNOMEDCT_CORE|CA - Cancer of oesophagus|Malignant tumor of esophagus
C0546837|T191|SY|363402007|SNOMEDCT_CORE|Cancer of esophagus|Malignant tumor of esophagus
C0546837|T191|SYGB|363402007|SNOMEDCT_CORE|Cancer of oesophagus|Malignant tumor of esophagus
C0546837|T191|SY|363402007|SNOMEDCT_CORE|Esophageal cancer|Malignant tumor of esophagus
C0546837|T191|SY|363402007|SNOMEDCT_CORE|Malignant neoplasm of esophagus|Malignant tumor of esophagus
C0546837|T191|SYGB|363402007|SNOMEDCT_CORE|Malignant neoplasm of oesophagus|Malignant tumor of esophagus
C0546837|T191|PT|363402007|SNOMEDCT_CORE|Malignant tumor of esophagus|Malignant tumor of esophagus
C0546837|T191|FN|363402007|SNOMEDCT_CORE|Malignant tumor of esophagus|Malignant tumor of esophagus
C0546837|T191|PTGB|363402007|SNOMEDCT_CORE|Malignant tumour of oesophagus|Malignant tumor of esophagus
C0546837|T191|SYGB|363402007|SNOMEDCT_CORE|Oesophageal cancer|Malignant tumor of esophagus
C0546884|T033|OAS|28560003|SNOMEDCT_CORE|Depletion of volume of plasma AND/OR extracellular fluid|Hypovolemia
C0546884|T033|IS|28560003|SNOMEDCT_CORE|Depletion of volume of plasma or extracellular fluid|Hypovolemia
C0546884|T033|OAS|28560003|SNOMEDCT_CORE|Fluid depletion|Hypovolemia
C0546884|T033|OAP|37472003|SNOMEDCT_CORE|Fluid volume deficit|Hypovolemia
C0546884|T033|OAS|28560003|SNOMEDCT_CORE|Fluid volume deficit|Hypovolemia
C0546884|T033|OAF|37472003|SNOMEDCT_CORE|Fluid volume deficit|Hypovolemia
C0546884|T033|OAS|28560003|SNOMEDCT_CORE|Fluid volume depletion|Hypovolemia
C0546884|T033|OAP|28560003|SNOMEDCT_CORE|Hypovolaemia|Hypovolemia
C0546884|T033|PTGB|816082000|SNOMEDCT_CORE|Hypovolaemia|Hypovolemia
C0546884|T033|OAP|28560003|SNOMEDCT_CORE|Hypovolemia|Hypovolemia
C0546884|T033|PT|816082000|SNOMEDCT_CORE|Hypovolemia|Hypovolemia
C0546884|T033|FN|816082000|SNOMEDCT_CORE|Hypovolemia|Hypovolemia
C0546884|T033|OAF|28560003|SNOMEDCT_CORE|Hypovolemia|Hypovolemia
C0546884|T033|OAS|28560003|SNOMEDCT_CORE|Sodium and water depletion|Hypovolemia
C0546884|T033|OAS|28560003|SNOMEDCT_CORE|Volume depletion|Hypovolemia
C0546953|T047|IS|27741009|SNOMEDCT_CORE|Subacromial bursitis|Subacromial bursitis
C0546953|T047|PT|40799003|SNOMEDCT_CORE|Subacromial bursitis|Subacromial bursitis
C0546953|T047|FN|40799003|SNOMEDCT_CORE|Subacromial bursitis|Subacromial bursitis
C0546969|T019|SY|204272007|SNOMEDCT_CORE|Congenital preauricular fistula|Preauricular fistula
C0546969|T019|SY|204272007|SNOMEDCT_CORE|Fistula auris congenita|Preauricular fistula
C0546969|T019|PT|204272007|SNOMEDCT_CORE|Preauricular fistula|Preauricular fistula
C0546969|T019|FN|204272007|SNOMEDCT_CORE|Preauricular fistula|Preauricular fistula
C0546969|T019|SY|204272007|SNOMEDCT_CORE|Preauricular sinus|Preauricular fistula
C0546983|T047|SY|40425004|SNOMEDCT_CORE|Nonpsychotic post-traumatic brain syndrome|Postconcussion syndrome
C0546983|T047|SY|40425004|SNOMEDCT_CORE|Post-concussion syndrome|Postconcussion syndrome
C0546983|T047|SY|40425004|SNOMEDCT_CORE|Post-concussional syndrome|Postconcussion syndrome
C0546983|T047|SY|40425004|SNOMEDCT_CORE|Post-contusional encephalopathy|Postconcussion syndrome
C0546983|T047|SY|40425004|SNOMEDCT_CORE|Post-contusional syndrome|Postconcussion syndrome
C0546983|T047|FN|40425004|SNOMEDCT_CORE|Postconcussion syndrome|Postconcussion syndrome
C0546983|T047|PT|40425004|SNOMEDCT_CORE|Postconcussion syndrome|Postconcussion syndrome
C0546983|T047|IS|40425004|SNOMEDCT_CORE|Postconcussion syndrome, NOS|Postconcussion syndrome
C0547030|T033|PT|63102001|SNOMEDCT_CORE|Visual disturbance|Visual disturbance
C0547030|T033|FN|63102001|SNOMEDCT_CORE|Visual disturbance|Visual disturbance
C0547030|T033|IS|63102001|SNOMEDCT_CORE|Visual disturbance, NOS|Visual disturbance
C0547065|T191|IS|22217002|SNOMEDCT_CORE|Mixed oligoastrocytoma|Mixed oligoastrocytoma
C0549106|T033|PT|160932005|SNOMEDCT_CORE|Financial problem|Financial problem
C0549106|T033|FN|160932005|SNOMEDCT_CORE|Financial problem|Financial problem
C0549124|T046|PT|54687002|SNOMEDCT_CORE|Arterial embolism|Arterial embolism
C0549124|T046|FN|54687002|SNOMEDCT_CORE|Arterial embolism|Arterial embolism
C0549124|T046|IS|54687002|SNOMEDCT_CORE|Arterial embolism, NOS, of unspecified artery|Arterial embolism
C0549124|T046|SY|54687002|SNOMEDCT_CORE|Arterial embolus|Arterial embolism
C0549124|T046|SY|54687002|SNOMEDCT_CORE|Embolic arterial occlusion|Arterial embolism
C0549150|T047|FN|399205006|SNOMEDCT_CORE|Pseudofolliculitis barbae|Pseudofolliculitis barbae
C0549150|T047|PT|399205006|SNOMEDCT_CORE|Pseudofolliculitis barbae|Pseudofolliculitis barbae
C0549169|T033|SY|77386006|SNOMEDCT_CORE|Pregnancy confirmed|Pregnancy confirmed
C0549201|T047|OF|201077008|SNOMEDCT_CORE|Asteatotic eczema|Asteatotic eczema
C0549201|T047|PT|201077008|SNOMEDCT_CORE|Asteatotic eczema|Asteatotic eczema
C0549201|T047|FN|201077008|SNOMEDCT_CORE|Asteatotic eczema|Asteatotic eczema
C0549201|T047|IS|201077008|SNOMEDCT_CORE|Eczema craquel|Asteatotic eczema
C0549201|T047|SY|201077008|SNOMEDCT_CORE|Eczema craquele|Asteatotic eczema
C0549206|T033|OP|77386006|SNOMEDCT_CORE|Patient currently pregnant|Pregnant
C0549206|T033|OF|77386006|SNOMEDCT_CORE|Patient currently pregnant|Pregnant
C0549206|T033|SY|77386006|SNOMEDCT_CORE|Pregnancy not delivered|Pregnant
C0549206|T033|PT|77386006|SNOMEDCT_CORE|Pregnant|Pregnant
C0549206|T033|FN|77386006|SNOMEDCT_CORE|Pregnant|Pregnant
C0549315|T191|PT|417044008|SNOMEDCT_CORE|Hydatidiform mole, benign|Hydatidiform mole, benign
C0549315|T191|FN|417044008|SNOMEDCT_CORE|Hydatidiform mole, benign|Hydatidiform mole, benign
C0549374|T047|PT|274137005|SNOMEDCT_CORE|Lumbar disc lesion|Lumbar disc lesion
C0549374|T047|FN|274137005|SNOMEDCT_CORE|Lumbar disc lesion|Lumbar disc lesion
C0549397|T033|PT|126660000|SNOMEDCT_CORE|Deviated nasal septum|Deviated nasal septum
C0549397|T033|FN|126660000|SNOMEDCT_CORE|Deviated nasal septum|Deviated nasal septum
C0549423|T047|PT|230746009|SNOMEDCT_CORE|Obstructive hydrocephalus|Obstructive hydrocephalus
C0549423|T047|FN|230746009|SNOMEDCT_CORE|Obstructive hydrocephalus|Obstructive hydrocephalus
C0549622|T048|PT|56925008|SNOMEDCT_CORE|Abnormal sexual function|Abnormal sexual function
C0549622|T048|FN|56925008|SNOMEDCT_CORE|Abnormal sexual function|Abnormal sexual function
C0549622|T048|SY|56925008|SNOMEDCT_CORE|Sexual dysfunction|Abnormal sexual function
C0549634|T033|PT|166818002|SNOMEDCT_CORE|Lipids abnormal|Lipids abnormal
C0549634|T033|FN|166818002|SNOMEDCT_CORE|Lipids abnormal|Lipids abnormal
C0553570|T047|PT|304930004|SNOMEDCT_CORE|Varicose veins of lower extremity with ulcer|Varicose veins of lower extremity with ulcer
C0553570|T047|FN|304930004|SNOMEDCT_CORE|Varicose veins of lower extremity with ulcer|Varicose veins of lower extremity with ulcer
C0553570|T047|OAP|195445008|SNOMEDCT_CORE|Varicose veins of the leg with ulcer|Varicose veins of lower extremity with ulcer
C0553570|T047|OAF|195445008|SNOMEDCT_CORE|Varicose veins of the leg with ulcer|Varicose veins of lower extremity with ulcer
C0553570|T047|SY|304930004|SNOMEDCT_CORE|Varicose veins with ulcer of lower extremity|Varicose veins of lower extremity with ulcer
C0553587|T047|PT|192999003|SNOMEDCT_CORE|Partial epilepsy with impairment of consciousness|Partial epilepsy with impairment of consciousness
C0553587|T047|FN|192999003|SNOMEDCT_CORE|Partial epilepsy with impairment of consciousness|Partial epilepsy with impairment of consciousness
C0553642|T047|FN|396333008|SNOMEDCT_CORE|Non-articular rheumatism|Non-articular rheumatism
C0553642|T047|PT|396333008|SNOMEDCT_CORE|Non-articular rheumatism|Non-articular rheumatism
C0553656|T047|IS|15033003|SNOMEDCT_CORE|Peritonsillar cellulitis|Peritonsillar cellulitis
C0553686|T190|PT|49453006|SNOMEDCT_CORE|Cerebral herniation|Cerebral herniation
C0553686|T190|FN|49453006|SNOMEDCT_CORE|Cerebral herniation|Cerebral herniation
C0553686|T190|SY|49453006|SNOMEDCT_CORE|Hernia cerebri|Cerebral herniation
C0553690|T047|PT|36179005|SNOMEDCT_CORE|R.I.N.D. syndrome|R.I.N.D. syndrome
C0553690|T047|OF|36179005|SNOMEDCT_CORE|R.I.N.D. syndrome|R.I.N.D. syndrome
C0553690|T047|SYGB|36179005|SNOMEDCT_CORE|Reversible ischaemic neurologic deficit syndrome|R.I.N.D. syndrome
C0553690|T047|SYGB|36179005|SNOMEDCT_CORE|Reversible ischaemic neurological defect|R.I.N.D. syndrome
C0553690|T047|SY|36179005|SNOMEDCT_CORE|Reversible ischemic neurologic deficit syndrome|R.I.N.D. syndrome
C0553690|T047|FN|36179005|SNOMEDCT_CORE|Reversible ischemic neurologic deficit syndrome|R.I.N.D. syndrome
C0553690|T047|SY|36179005|SNOMEDCT_CORE|Reversible ischemic neurological defect|R.I.N.D. syndrome
C0553690|T047|SYGB|36179005|SNOMEDCT_CORE|RIND - Reversible ischaemic neurological defect|R.I.N.D. syndrome
C0553690|T047|SY|36179005|SNOMEDCT_CORE|RIND - Reversible ischemic neurological defect|R.I.N.D. syndrome
C0553718|T047|PT|236488005|SNOMEDCT_CORE|Renal artery occlusion|Renal artery occlusion
C0553718|T047|FN|236488005|SNOMEDCT_CORE|Renal artery occlusion|Renal artery occlusion
C0553723|T191|SY|254651007|SNOMEDCT_CORE|Cutaneous squamous cell carcinoma|Squamous cell carcinoma of skin
C0553723|T191|SY|254651007|SNOMEDCT_CORE|SCC - Cutaneous squamous cell carcinoma|Squamous cell carcinoma of skin
C0553723|T191|SY|254651007|SNOMEDCT_CORE|SCC - Squamous cell carcinoma of skin|Squamous cell carcinoma of skin
C0553723|T191|SY|254651007|SNOMEDCT_CORE|Spinous cell carcinoma|Squamous cell carcinoma of skin
C0553723|T191|PT|254651007|SNOMEDCT_CORE|Squamous cell carcinoma of skin|Squamous cell carcinoma of skin
C0553723|T191|FN|254651007|SNOMEDCT_CORE|Squamous cell carcinoma of skin|Squamous cell carcinoma of skin
C0553727|T033|IS|44695005|SNOMEDCT_CORE|Muscular paralysis|Muscular paralysis
C0553730|T047|SY|239832006|SNOMEDCT_CORE|Calcium pyrophosphate arthritis and periarthritis|Calcium pyrophosphate deposition disease
C0553730|T047|PT|239832006|SNOMEDCT_CORE|Calcium pyrophosphate deposition disease|Calcium pyrophosphate deposition disease
C0553730|T047|FN|239832006|SNOMEDCT_CORE|Calcium pyrophosphate deposition disease|Calcium pyrophosphate deposition disease
C0553730|T047|IS|60782007|SNOMEDCT_CORE|Calcium pyrophosphate deposition disease|Calcium pyrophosphate deposition disease
C0553730|T047|IS|60782007|SNOMEDCT_CORE|Chondrocalcinosis|Calcium pyrophosphate deposition disease
C0553730|T047|OAS|60782007|SNOMEDCT_CORE|Chondrocalcinosis articularis|Calcium pyrophosphate deposition disease
C0553730|T047|OAS|60782007|SNOMEDCT_CORE|Chondrocalcinosis due to pyrophosphate crystals|Calcium pyrophosphate deposition disease
C0553730|T047|PT|201637001|SNOMEDCT_CORE|Chondrocalcinosis due to pyrophosphate crystals|Calcium pyrophosphate deposition disease
C0553730|T047|FN|201637001|SNOMEDCT_CORE|Chondrocalcinosis due to pyrophosphate crystals|Calcium pyrophosphate deposition disease
C0553730|T047|IS|60782007|SNOMEDCT_CORE|CPDD|Calcium pyrophosphate deposition disease
C0553730|T047|SY|239832006|SNOMEDCT_CORE|CPDD - Calcium pyrophosphate deposition disease|Calcium pyrophosphate deposition disease
C0553730|T047|SY|239832006|SNOMEDCT_CORE|CPPD - Calcium pyrophosphate deposition disease|Calcium pyrophosphate deposition disease
C0553730|T047|OAP|60782007|SNOMEDCT_CORE|Pseudogout|Calcium pyrophosphate deposition disease
C0553730|T047|SY|201637001|SNOMEDCT_CORE|Pseudogout|Calcium pyrophosphate deposition disease
C0553757|T047|PT|275462005|SNOMEDCT_CORE|Disorder of smell|Disorder of smell
C0553757|T047|FN|275462005|SNOMEDCT_CORE|Disorder of smell|Disorder of smell
C0553757|T047|OP|275462005|SNOMEDCT_CORE|Disorders of smell|Disorder of smell
C0553757|T047|OF|275462005|SNOMEDCT_CORE|Disorders of smell|Disorder of smell
C0553812|T048|OAP|268641003|SNOMEDCT_CORE|Cannabis type drug dependence|Cannabis type drug dependence
C0553812|T048|OAF|268641003|SNOMEDCT_CORE|Cannabis type drug dependence|Cannabis type drug dependence
C0553968|T047|OAP|275499005|SNOMEDCT_CORE|Acute wheezy bronchitis|Acute wheezy bronchitis
C0553968|T047|OAF|275499005|SNOMEDCT_CORE|Acute wheezy bronchitis|Acute wheezy bronchitis
C0554021|T047|SY|723177002|SNOMEDCT_CORE|Recurrent mouth ulcer|Recurrent ulcer of mouth
C0554021|T047|OAP|281775009|SNOMEDCT_CORE|Recurrent mouth ulcers|Recurrent ulcer of mouth
C0554021|T047|OAF|281775009|SNOMEDCT_CORE|Recurrent mouth ulcers|Recurrent ulcer of mouth
C0554021|T047|OAS|281775009|SNOMEDCT_CORE|Recurrent oral ulceration|Recurrent ulcer of mouth
C0554021|T047|SY|723177002|SNOMEDCT_CORE|Recurrent oral ulceration|Recurrent ulcer of mouth
C0554021|T047|PT|723177002|SNOMEDCT_CORE|Recurrent ulcer of mouth|Recurrent ulcer of mouth
C0554021|T047|FN|723177002|SNOMEDCT_CORE|Recurrent ulcer of mouth|Recurrent ulcer of mouth
C0554021|T047|OAS|281775009|SNOMEDCT_CORE|ROU - Recurrent oral ulceration|Recurrent ulcer of mouth
C0554103|T046|PT|197494007|SNOMEDCT_CORE|Intestinal malabsorption of fat|Intestinal malabsorption of fat
C0554103|T046|FN|197494007|SNOMEDCT_CORE|Intestinal malabsorption of fat|Intestinal malabsorption of fat
C0554122|T020|OAS|18253009|SNOMEDCT_CORE|Unilateral obstructed recurrent inguinal hernia|Unilateral recurrent inguinal hernia with obstruction but no gangrene
C0554122|T020|OAP|18253009|SNOMEDCT_CORE|Unilateral recurrent inguinal hernia with obstruction but no gangrene|Unilateral recurrent inguinal hernia with obstruction but no gangrene
C0554122|T020|OF|18253009|SNOMEDCT_CORE|Unilateral recurrent inguinal hernia with obstruction but no gangrene|Unilateral recurrent inguinal hernia with obstruction but no gangrene
C0554122|T020|OAF|18253009|SNOMEDCT_CORE|Unilateral recurrent inguinal hernia with obstruction but no gangrene|Unilateral recurrent inguinal hernia with obstruction but no gangrene
C0554123|T020|OAP|55993003|SNOMEDCT_CORE|Unilateral inguinal hernia with obstruction but no gangrene|Unilateral inguinal hernia with obstruction but no gangrene
C0554123|T020|OF|55993003|SNOMEDCT_CORE|Unilateral inguinal hernia with obstruction but no gangrene|Unilateral inguinal hernia with obstruction but no gangrene
C0554123|T020|OAF|55993003|SNOMEDCT_CORE|Unilateral inguinal hernia with obstruction but no gangrene|Unilateral inguinal hernia with obstruction but no gangrene
C0554123|T020|OAS|55993003|SNOMEDCT_CORE|Unilateral obstructed inguinal hernia|Unilateral inguinal hernia with obstruction but no gangrene
C0554309|T047|IS|55655006|SNOMEDCT_CORE|Azotaemia|Prerenal uremia syndrome
C0554309|T047|IS|55655006|SNOMEDCT_CORE|Azotemia|Prerenal uremia syndrome
C0554309|T047|OAS|55655006|SNOMEDCT_CORE|Blum's syndrome|Prerenal uremia syndrome
C0554309|T047|OAS|55655006|SNOMEDCT_CORE|Extrarenal uraemia syndrome|Prerenal uremia syndrome
C0554309|T047|OAS|55655006|SNOMEDCT_CORE|Extrarenal uremia syndrome|Prerenal uremia syndrome
C0554309|T047|IS|55655006|SNOMEDCT_CORE|Prerenal azotaemia|Prerenal uremia syndrome
C0554309|T047|IS|55655006|SNOMEDCT_CORE|Prerenal azotemia|Prerenal uremia syndrome
C0554309|T047|OAS|55655006|SNOMEDCT_CORE|Prerenal renal failure|Prerenal uremia syndrome
C0554309|T047|OAS|55655006|SNOMEDCT_CORE|Prerenal uraemia|Prerenal uremia syndrome
C0554309|T047|OAP|55655006|SNOMEDCT_CORE|Prerenal uraemia syndrome|Prerenal uremia syndrome
C0554309|T047|OAS|55655006|SNOMEDCT_CORE|Prerenal uremia|Prerenal uremia syndrome
C0554309|T047|OAP|55655006|SNOMEDCT_CORE|Prerenal uremia syndrome|Prerenal uremia syndrome
C0554309|T047|OAF|55655006|SNOMEDCT_CORE|Prerenal uremia syndrome|Prerenal uremia syndrome
C0554478|T047|PT|275448003|SNOMEDCT_CORE|Perianal dermatitis|Perianal dermatitis
C0554478|T047|FN|275448003|SNOMEDCT_CORE|Perianal dermatitis|Perianal dermatitis
C0554595|T047|PT|202881005|SNOMEDCT_CORE|Tibialis posterior tendinitis|Tibialis posterior tendinitis
C0554595|T047|FN|202881005|SNOMEDCT_CORE|Tibialis posterior tendinitis|Tibialis posterior tendinitis
C0555003|T033|PT|276079004|SNOMEDCT_CORE|Partnership problems|Partnership problems
C0555003|T033|FN|276079004|SNOMEDCT_CORE|Partnership problems|Partnership problems
C0555026|T033|IS|65118005|SNOMEDCT_CORE|Marital problem|Marital problems
C0555026|T033|PT|65118005|SNOMEDCT_CORE|Marital problems|Marital problems
C0555026|T033|FN|65118005|SNOMEDCT_CORE|Marital problems|Marital problems
C0555056|T184|PT|61281005|SNOMEDCT_CORE|Bloodstained sputum|Bloodstained sputum
C0555056|T184|FN|61281005|SNOMEDCT_CORE|Bloodstained sputum|Bloodstained sputum
C0555056|T184|IS|61281005|SNOMEDCT_CORE|Expectoration of blood stained sputum|Bloodstained sputum
C0555056|T184|SY|61281005|SNOMEDCT_CORE|Expectoration of blood tinged sputum|Bloodstained sputum
C0555276|T191|SY|275266006|SNOMEDCT_CORE|Cancer metastatic to digestive organs|Metastasis to digestive organs
C0555276|T191|PT|275266006|SNOMEDCT_CORE|Metastasis to digestive organs|Metastasis to digestive organs
C0555276|T191|FN|275266006|SNOMEDCT_CORE|Metastasis to digestive organs|Metastasis to digestive organs
C0555294|T037|PT|210560004|SNOMEDCT_CORE|Open wound of hand, excluding finger|Open wound of hand, excluding finger
C0555294|T037|FN|210560004|SNOMEDCT_CORE|Open wound of hand, excluding finger|Open wound of hand, excluding finger
C0555295|T037|PT|125653000|SNOMEDCT_CORE|Open wound of finger|Open wound of finger
C0555295|T037|FN|125653000|SNOMEDCT_CORE|Open wound of finger|Open wound of finger
C0555295|T037|SY|125653000|SNOMEDCT_CORE|Open wound, finger|Open wound of finger
C0555297|T037|PT|269183000|SNOMEDCT_CORE|Open wound of foot, excluding toe|Open wound of foot, excluding toe
C0555297|T037|FN|269183000|SNOMEDCT_CORE|Open wound of foot, excluding toe|Open wound of foot, excluding toe
C0555311|T037|PT|275335003|SNOMEDCT_CORE|Ruptured Achilles tendon - traumatic|Ruptured Achilles tendon - traumatic
C0555311|T037|FN|275335003|SNOMEDCT_CORE|Ruptured Achilles tendon - traumatic|Ruptured Achilles tendon - traumatic
C0555315|T037|PT|275334004|SNOMEDCT_CORE|Shoulder strain|Shoulder strain
C0555315|T037|FN|275334004|SNOMEDCT_CORE|Shoulder strain|Shoulder strain
C0555321|T037|PT|275330008|SNOMEDCT_CORE|Current knee cartilage tear|Current knee cartilage tear
C0555321|T037|FN|275330008|SNOMEDCT_CORE|Current knee cartilage tear|Current knee cartilage tear
C0555330|T037|SY|269080004|SNOMEDCT_CORE|Closed fracture of distal end of humerus|Closed fracture of lower end of humerus
C0555330|T037|PT|269080004|SNOMEDCT_CORE|Closed fracture of lower end of humerus|Closed fracture of lower end of humerus
C0555330|T037|SY|269080004|SNOMEDCT_CORE|Closed fracture of the distal humerus|Closed fracture of lower end of humerus
C0555330|T037|FN|269080004|SNOMEDCT_CORE|Closed fracture of the distal humerus|Closed fracture of lower end of humerus
C0555337|T037|PT|274160002|SNOMEDCT_CORE|Fracture of phalanx of thumb|Fracture of phalanx of thumb
C0555337|T037|FN|274160002|SNOMEDCT_CORE|Fracture of phalanx of thumb|Fracture of phalanx of thumb
C0555337|T037|SY|274160002|SNOMEDCT_CORE|Fracture of thumb|Fracture of phalanx of thumb
C0555972|T047|PT|299989006|SNOMEDCT_CORE|Infection of toe|Infection of toe
C0555972|T047|FN|299989006|SNOMEDCT_CORE|Infection of toe|Infection of toe
C0555972|T047|SY|299989006|SNOMEDCT_CORE|Infection toe|Infection of toe
C0555972|T047|OF|299989006|SNOMEDCT_CORE|Infection toe|Infection of toe
C0555977|T037|PT|275453008|SNOMEDCT_CORE|Foreign body - finger|Foreign body - finger
C0555977|T037|FN|275453008|SNOMEDCT_CORE|Foreign body - finger|Foreign body - finger
C0556278|T033|OAS|228142005|SNOMEDCT_CORE|SEN - Special educational needs|Special educational needs
C0556278|T033|OAP|228142005|SNOMEDCT_CORE|Special educational needs|Special educational needs
C0556278|T033|OAF|228142005|SNOMEDCT_CORE|Special educational needs|Special educational needs
C0556279|T033|SY|228146008|SNOMEDCT_CORE|Difficulty with personal care|Personal care impairment
C0556279|T033|PT|228146008|SNOMEDCT_CORE|Personal care impairment|Personal care impairment
C0556279|T033|FN|228146008|SNOMEDCT_CORE|Personal care impairment|Personal care impairment
C0556279|T033|SY|228146008|SNOMEDCT_CORE|Personal condition impairment of self care|Personal care impairment
C0556280|T033|PT|228147004|SNOMEDCT_CORE|Gross motor impairment|Gross motor impairment
C0556280|T033|FN|228147004|SNOMEDCT_CORE|Gross motor impairment|Gross motor impairment
C0556281|T033|PT|228148009|SNOMEDCT_CORE|Fine motor impairment|Fine motor impairment
C0556281|T033|FN|228148009|SNOMEDCT_CORE|Fine motor impairment|Fine motor impairment
C0556338|T033|OAP|228318004|SNOMEDCT_CORE|Regular drinker|Regular drinker
C0556338|T033|OAF|228318004|SNOMEDCT_CORE|Regular drinker|Regular drinker
C0556340|T033|PT|228320001|SNOMEDCT_CORE|Habitual drinker|Habitual drinker
C0556340|T033|FN|228320001|SNOMEDCT_CORE|Habitual drinker|Habitual drinker
C0556389|T033|PT|228371004|SNOMEDCT_CORE|Long-term drug misuser|Long-term drug misuser
C0556389|T033|FN|228371004|SNOMEDCT_CORE|Long-term drug misuser|Long-term drug misuser
C0556390|T033|SY|228372006|SNOMEDCT_CORE|Multi-drug misuser|Poly-drug misuser
C0556390|T033|SY|228372006|SNOMEDCT_CORE|Poly-drug abuser|Poly-drug misuser
C0556390|T033|PT|228372006|SNOMEDCT_CORE|Poly-drug misuser|Poly-drug misuser
C0556390|T033|FN|228372006|SNOMEDCT_CORE|Poly-drug misuser|Poly-drug misuser
C0558116|T048|SY|63384009|SNOMEDCT_CORE|Body image disturbance|Distorted body image
C0558116|T048|PT|63384009|SNOMEDCT_CORE|Distorted body image|Distorted body image
C0558116|T048|FN|63384009|SNOMEDCT_CORE|Distorted body image|Distorted body image
C0558116|T048|SY|63384009|SNOMEDCT_CORE|Disturbed body image|Distorted body image
C0558158|T047|IS|225561003|SNOMEDCT_CORE|Decubitus ulcer of heel|Pressure ulcer of heel
C0558158|T047|SY|225561003|SNOMEDCT_CORE|Pressure sore on heel|Pressure ulcer of heel
C0558158|T047|OF|225561003|SNOMEDCT_CORE|Pressure sore on heel|Pressure ulcer of heel
C0558158|T047|PT|225561003|SNOMEDCT_CORE|Pressure ulcer of heel|Pressure ulcer of heel
C0558158|T047|FN|225561003|SNOMEDCT_CORE|Pressure ulcer of heel|Pressure ulcer of heel
C0558158|T047|SY|225561003|SNOMEDCT_CORE|Pressure ulcer on heel|Pressure ulcer of heel
C0558159|T046|IS|225562005|SNOMEDCT_CORE|Decubitus ulcer of sacrum|Pressure ulcer of sacral region
C0558159|T046|SY|225562005|SNOMEDCT_CORE|Pressure sore on sacrum|Pressure ulcer of sacral region
C0558159|T046|OF|225562005|SNOMEDCT_CORE|Pressure sore on sacrum|Pressure ulcer of sacral region
C0558159|T046|PT|225562005|SNOMEDCT_CORE|Pressure ulcer of sacral region|Pressure ulcer of sacral region
C0558159|T046|FN|225562005|SNOMEDCT_CORE|Pressure ulcer of sacral region|Pressure ulcer of sacral region
C0558159|T046|SY|225562005|SNOMEDCT_CORE|Pressure ulcer on sacrum|Pressure ulcer of sacral region
C0558159|T046|IS|225562005|SNOMEDCT_CORE|Sacral pressure core|Pressure ulcer of sacral region
C0558159|T046|SY|225562005|SNOMEDCT_CORE|Sacral pressure sore|Pressure ulcer of sacral region
C0558160|T047|IS|225563000|SNOMEDCT_CORE|Decubitus ulcer of buttock|Pressure ulcer of buttock
C0558160|T047|SY|225563000|SNOMEDCT_CORE|Pressure sore of buttock|Pressure ulcer of buttock
C0558160|T047|OF|225563000|SNOMEDCT_CORE|Pressure sore of buttock|Pressure ulcer of buttock
C0558160|T047|OP|225563000|SNOMEDCT_CORE|Pressure sore on buttocks|Pressure ulcer of buttock
C0558160|T047|OF|225563000|SNOMEDCT_CORE|Pressure sore on buttocks|Pressure ulcer of buttock
C0558160|T047|PT|225563000|SNOMEDCT_CORE|Pressure ulcer of buttock|Pressure ulcer of buttock
C0558160|T047|FN|225563000|SNOMEDCT_CORE|Pressure ulcer of buttock|Pressure ulcer of buttock
C0558353|T191|PT|269516007|SNOMEDCT_CORE|Tongue carcinoma|Tongue carcinoma
C0558353|T191|FN|269516007|SNOMEDCT_CORE|Tongue carcinoma|Tongue carcinoma
C0558355|T191|PT|274085008|SNOMEDCT_CORE|Tonsil carcinoma|Tonsil carcinoma
C0558355|T191|FN|274085008|SNOMEDCT_CORE|Tonsil carcinoma|Tonsil carcinoma
C0558362|T047|PT|195790000|SNOMEDCT_CORE|Pansinusitis|Pansinusitis
C0558362|T047|FN|195790000|SNOMEDCT_CORE|Pansinusitis|Pansinusitis
C0558368|T033|PT|161816004|SNOMEDCT_CORE|Vaginal irritation|Vaginal irritation
C0558368|T033|FN|161816004|SNOMEDCT_CORE|Vaginal irritation|Vaginal irritation
C0558372|T047|PT|274120003|SNOMEDCT_CORE|Thyroid disease in pregnancy|Thyroid disease in pregnancy
C0558372|T047|FN|274120003|SNOMEDCT_CORE|Thyroid disease in pregnancy|Thyroid disease in pregnancy
C0558382|T047|PT|128276007|SNOMEDCT_CORE|Cellulitis of foot|Cellulitis of foot
C0558382|T047|FN|128276007|SNOMEDCT_CORE|Cellulitis of foot|Cellulitis of foot
C0558385|T047|OF|118939000|SNOMEDCT_CORE|Disease of neck|Disorder of neck
C0558385|T047|IS|118939000|SNOMEDCT_CORE|Disease of neck|Disorder of neck
C0558385|T047|PT|118939000|SNOMEDCT_CORE|Disorder of neck|Disorder of neck
C0558385|T047|FN|118939000|SNOMEDCT_CORE|Disorder of neck|Disorder of neck
C0558399|T037|OAP|269329008|SNOMEDCT_CORE|Arm sprain - upper|Arm sprain - upper
C0558399|T037|OAF|269329008|SNOMEDCT_CORE|Arm sprain - upper|Arm sprain - upper
C0558401|T037|PT|274165007|SNOMEDCT_CORE|Laceration of skin|Laceration of skin
C0558401|T037|FN|274165007|SNOMEDCT_CORE|Laceration of skin|Laceration of skin
C0558407|T037|PT|125652005|SNOMEDCT_CORE|Open wound of hand|Open wound of hand
C0558407|T037|FN|125652005|SNOMEDCT_CORE|Open wound of hand|Open wound of hand
C0558427|T033|PTGB|274203005|SNOMEDCT_CORE|Subungual haematoma of foot|Subungual hematoma of foot
C0558427|T033|OP|274203005|SNOMEDCT_CORE|Subungual haematoma, foot|Subungual hematoma of foot
C0558427|T033|IS|274203005|SNOMEDCT_CORE|Subungual haematoma, foot.|Subungual hematoma of foot
C0558427|T033|PT|274203005|SNOMEDCT_CORE|Subungual hematoma of foot|Subungual hematoma of foot
C0558427|T033|FN|274203005|SNOMEDCT_CORE|Subungual hematoma of foot|Subungual hematoma of foot
C0558427|T033|OP|274203005|SNOMEDCT_CORE|Subungual hematoma, foot|Subungual hematoma of foot
C0558427|T033|OF|274203005|SNOMEDCT_CORE|Subungual hematoma, foot|Subungual hematoma of foot
C0558427|T033|IS|274203005|SNOMEDCT_CORE|Subungual hematoma, foot.|Subungual hematoma of foot
C0558427|T033|OF|274203005|SNOMEDCT_CORE|Subungual hematoma, foot.|Subungual hematoma of foot
C0558441|T037|PT|274227007|SNOMEDCT_CORE|Cut - accidental|Cut - accidental
C0558441|T037|FN|274227007|SNOMEDCT_CORE|Cut - accidental|Cut - accidental
C0558442|T048|PT|274228002|SNOMEDCT_CORE|Drug overdose - suicide|Drug overdose - suicide
C0558442|T048|OF|274228002|SNOMEDCT_CORE|Drug overdose - suicide|Drug overdose - suicide
C0558442|T048|FN|274228002|SNOMEDCT_CORE|Drug overdose - suicide|Drug overdose - suicide
C0558975|T033|IS|275881005|SNOMEDCT_CORE|H/O: sexually trans. disease|History of sexually transmitted disease
C0558975|T033|IS|275881005|SNOMEDCT_CORE|History of - sexually transmitted disease|History of sexually transmitted disease
C0558975|T033|OF|275881005|SNOMEDCT_CORE|History of - sexually transmitted disease|History of sexually transmitted disease
C0558975|T033|PT|275881005|SNOMEDCT_CORE|History of sexually transmitted disease|History of sexually transmitted disease
C0558975|T033|SY|275881005|SNOMEDCT_CORE|History of sexually transmitted disease|History of sexually transmitted disease
C0558975|T033|FN|275881005|SNOMEDCT_CORE|History of sexually transmitted disease|History of sexually transmitted disease
C0558975|T033|SY|275881005|SNOMEDCT_CORE|History of venereal disease|History of sexually transmitted disease
C0558975|T033|IS|275881005|SNOMEDCT_CORE|Sexually transmitted dis H/O|History of sexually transmitted disease
C0558975|T033|OF|275881005|SNOMEDCT_CORE|Sexually transmitted dis H/O|History of sexually transmitted disease
C0558977|T033|PT|275531008|SNOMEDCT_CORE|H/O: pacemaker in situ|H/O: pacemaker in situ
C0558977|T033|OF|275531008|SNOMEDCT_CORE|History of - pacemaker in situ|H/O: pacemaker in situ
C0558977|T033|IS|275531008|SNOMEDCT_CORE|History of - pacemaker in situ|H/O: pacemaker in situ
C0558977|T033|FN|275531008|SNOMEDCT_CORE|History of pacemaker in situ|H/O: pacemaker in situ
C0558977|T033|SY|275531008|SNOMEDCT_CORE|History of pacemaker in situ|H/O: pacemaker in situ
C0559036|T037|PT|111224002|SNOMEDCT_CORE|Derangement of meniscus|Derangement of meniscus
C0559036|T037|FN|111224002|SNOMEDCT_CORE|Derangement of meniscus of knee joint|Derangement of meniscus
C0559036|T037|SY|111224002|SNOMEDCT_CORE|Derangement of meniscus of knee joint|Derangement of meniscus
C0559036|T037|SY|111224002|SNOMEDCT_CORE|Disorder of meniscus of knee|Derangement of meniscus
C0559096|T047|IS|268054009|SNOMEDCT_CORE|Osteoarthritis -multiple joint|Osteoarthritis of multiple joints
C0559096|T047|OF|268054009|SNOMEDCT_CORE|Osteoarthritis -multiple joint|Osteoarthritis of multiple joints
C0559096|T047|FN|268054009|SNOMEDCT_CORE|Osteoarthritis of multiple joints|Osteoarthritis of multiple joints
C0559096|T047|PT|268054009|SNOMEDCT_CORE|Osteoarthritis of multiple joints|Osteoarthritis of multiple joints
C0559112|T033|PT|267004000|SNOMEDCT_CORE|H/O: musculoskeletal disease|H/O: musculoskeletal disease
C0559112|T033|OF|267004000|SNOMEDCT_CORE|History of - musculoskeletal disease|H/O: musculoskeletal disease
C0559112|T033|IS|267004000|SNOMEDCT_CORE|History of - musculoskeletal disease|H/O: musculoskeletal disease
C0559112|T033|FN|267004000|SNOMEDCT_CORE|History of musculoskeletal disease|H/O: musculoskeletal disease
C0559112|T033|SY|267004000|SNOMEDCT_CORE|History of musculoskeletal disease|H/O: musculoskeletal disease
C0559112|T033|SY|267004000|SNOMEDCT_CORE|History of musculoskeletal disorder|H/O: musculoskeletal disease
C0559120|T033|OF|275111003|SNOMEDCT_CORE|Family history: Ovarian carcinoma|FH: Ovarian carcinoma
C0559120|T033|OAF|275111003|SNOMEDCT_CORE|Family history: Ovarian carcinoma|FH: Ovarian carcinoma
C0559120|T033|OAS|275111003|SNOMEDCT_CORE|Family history: Ovarian carcinoma|FH: Ovarian carcinoma
C0559120|T033|OAP|275111003|SNOMEDCT_CORE|FH: Ovarian carcinoma|FH: Ovarian carcinoma
C0559136|T033|OF|275124003|SNOMEDCT_CORE|Family history: Coronary thrombosis|FH: Coronary thrombosis
C0559136|T033|FN|275124003|SNOMEDCT_CORE|Family history: Coronary thrombosis|FH: Coronary thrombosis
C0559136|T033|SY|275124003|SNOMEDCT_CORE|Family history: Coronary thrombosis|FH: Coronary thrombosis
C0559136|T033|PT|275124003|SNOMEDCT_CORE|FH: Coronary thrombosis|FH: Coronary thrombosis
C0559154|T033|OP|275538002|SNOMEDCT_CORE|H/O: anaemia|History of anemia
C0559154|T033|OP|275538002|SNOMEDCT_CORE|H/O: anemia|History of anemia
C0559154|T033|IS|275538002|SNOMEDCT_CORE|History of - anemia|History of anemia
C0559154|T033|OF|275538002|SNOMEDCT_CORE|History of - anemia|History of anemia
C0559154|T033|PTGB|275538002|SNOMEDCT_CORE|History of anaemia|History of anemia
C0559154|T033|PT|275538002|SNOMEDCT_CORE|History of anemia|History of anemia
C0559154|T033|FN|275538002|SNOMEDCT_CORE|History of anemia|History of anemia
C0559157|T033|PT|275544003|SNOMEDCT_CORE|H/O: heart disorder|H/O: heart disorder
C0559157|T033|OF|275544003|SNOMEDCT_CORE|History of - heart disorder|H/O: heart disorder
C0559157|T033|IS|275544003|SNOMEDCT_CORE|History of - heart disorder|H/O: heart disorder
C0559157|T033|FN|275544003|SNOMEDCT_CORE|History of heart disorder|H/O: heart disorder
C0559157|T033|SY|275544003|SNOMEDCT_CORE|History of heart disorder|H/O: heart disorder
C0559159|T033|SY|275526006|SNOMEDCT_CORE|H/O: CVA|History of cerebrovascular accident
C0559159|T033|SY|275526006|SNOMEDCT_CORE|H/O: stroke|History of cerebrovascular accident
C0559159|T033|IS|275526006|SNOMEDCT_CORE|History of - cerebrovascular accident|History of cerebrovascular accident
C0559159|T033|OF|275526006|SNOMEDCT_CORE|History of - cerebrovascular accident|History of cerebrovascular accident
C0559159|T033|OF|275526006|SNOMEDCT_CORE|History of - CVA|History of cerebrovascular accident
C0559159|T033|PT|275526006|SNOMEDCT_CORE|History of cerebrovascular accident|History of cerebrovascular accident
C0559159|T033|FN|275526006|SNOMEDCT_CORE|History of cerebrovascular accident|History of cerebrovascular accident
C0559162|T033|PT|275546001|SNOMEDCT_CORE|H/O: thrombosis|H/O: thrombosis
C0559162|T033|OF|275546001|SNOMEDCT_CORE|History of - thrombosis|H/O: thrombosis
C0559162|T033|IS|275546001|SNOMEDCT_CORE|History of - thrombosis|H/O: thrombosis
C0559162|T033|FN|275546001|SNOMEDCT_CORE|History of thrombosis|H/O: thrombosis
C0559162|T033|SY|275546001|SNOMEDCT_CORE|History of thrombosis|H/O: thrombosis
C0559175|T033|PT|275565009|SNOMEDCT_CORE|H/O: intestinal by-pass|H/O: intestinal by-pass
C0559175|T033|OF|275565009|SNOMEDCT_CORE|History of - intestinal by-pass|H/O: intestinal by-pass
C0559175|T033|IS|275565009|SNOMEDCT_CORE|History of - intestinal by-pass|H/O: intestinal by-pass
C0559175|T033|FN|275565009|SNOMEDCT_CORE|History of intestinal by-pass|H/O: intestinal by-pass
C0559175|T033|SY|275565009|SNOMEDCT_CORE|History of intestinal by-pass|H/O: intestinal by-pass
C0559229|T033|SY|281900007|SNOMEDCT_CORE|NAD - No abnormality detected|No abnormality detected
C0559229|T033|PT|281900007|SNOMEDCT_CORE|No abnormality detected|No abnormality detected
C0559229|T033|FN|281900007|SNOMEDCT_CORE|No abnormality detected|No abnormality detected
C0559258|T047|PT|302935008|SNOMEDCT_CORE|Infective discitis|Infective discitis
C0559258|T047|FN|302935008|SNOMEDCT_CORE|Infective discitis|Infective discitis
C0559260|T019|SY|20944008|SNOMEDCT_CORE|Congenital scoliosis|Congenital scoliosis
C0559260|T019|IS|20944008|SNOMEDCT_CORE|Scoliosis|Congenital scoliosis
C0559444|T037|PT|281544003|SNOMEDCT_CORE|Strain of tendon of foot and ankle|Strain of tendon of foot and ankle
C0559444|T037|FN|281544003|SNOMEDCT_CORE|Strain of tendon of foot and ankle|Strain of tendon of foot and ankle
C0559470|T047|PT|91935009|SNOMEDCT_CORE|Allergy to peanut|Allergy to peanut
C0559470|T047|FN|91935009|SNOMEDCT_CORE|Allergy to peanut|Allergy to peanut
C0559470|T047|SY|91935009|SNOMEDCT_CORE|Allergy to peanuts|Allergy to peanut
C0559470|T047|OF|91935009|SNOMEDCT_CORE|Allergy to peanuts|Allergy to peanut
C0559491|T037|SY|123536004|SNOMEDCT_CORE|Sprain of ligament of upper limb|Sprain of upper extremity
C0559491|T037|SY|123536004|SNOMEDCT_CORE|Sprain of shoulder and upper arm|Sprain of upper extremity
C0559491|T037|PT|123536004|SNOMEDCT_CORE|Sprain of upper extremity|Sprain of upper extremity
C0559491|T037|FN|123536004|SNOMEDCT_CORE|Sprain of upper extremity|Sprain of upper extremity
C0559492|T037|PT|281598004|SNOMEDCT_CORE|Sprain of spinal ligament|Sprain of spinal ligament
C0559492|T037|FN|281598004|SNOMEDCT_CORE|Sprain of spinal ligament|Sprain of spinal ligament
C0559493|T037|PT|281599007|SNOMEDCT_CORE|Sprain of ligament of lower limb|Sprain of ligament of lower limb
C0559493|T037|FN|281599007|SNOMEDCT_CORE|Sprain of ligament of lower limb|Sprain of ligament of lower limb
C0559536|T033|OAP|281638009|SNOMEDCT_CORE|Hepatitis B contact|Hepatitis B contact
C0559536|T033|OAF|281638009|SNOMEDCT_CORE|Hepatitis B contact|Hepatitis B contact
C0559550|T033|PT|281666001|SNOMEDCT_CORE|Family history of disorder|Family history of disorder
C0559550|T033|OF|281666001|SNOMEDCT_CORE|Family history of disorder|Family history of disorder
C0559550|T033|FN|281666001|SNOMEDCT_CORE|Family history of disorder|Family history of disorder
C0559555|T033|SY|266890009|SNOMEDCT_CORE|Alcoholism in family|Family history of alcoholism
C0559555|T033|PT|266890009|SNOMEDCT_CORE|Family history of alcoholism|Family history of alcoholism
C0559555|T033|OF|266890009|SNOMEDCT_CORE|Family history of alcoholism|Family history of alcoholism
C0559555|T033|FN|266890009|SNOMEDCT_CORE|Family history of alcoholism|Family history of alcoholism
C0559555|T033|SY|266890009|SNOMEDCT_CORE|FH - Alcoholism|Family history of alcoholism
C0559567|T037|PT|373600006|SNOMEDCT_CORE|Multiple bruising|Multiple bruising
C0559567|T037|FN|373600006|SNOMEDCT_CORE|Multiple bruising|Multiple bruising
C0559755|T047|PTGB|281864001|SNOMEDCT_CORE|Non-traumatic intracranial subdural haematoma|Non-traumatic intracranial subdural hematoma
C0559755|T047|PT|281864001|SNOMEDCT_CORE|Non-traumatic intracranial subdural hematoma|Non-traumatic intracranial subdural hematoma
C0559755|T047|FN|281864001|SNOMEDCT_CORE|Non-traumatic intracranial subdural hematoma|Non-traumatic intracranial subdural hematoma
C0559893|T047|IS|282028001|SNOMEDCT_CORE|MRSA - Multiple-resistant Staphylococcus aureus infection|Multiple-resistant Staphylococcus aureus infection
C0559893|T047|PT|282028001|SNOMEDCT_CORE|Multiple-resistant Staphylococcus aureus infection|Multiple-resistant Staphylococcus aureus infection
C0559893|T047|FN|282028001|SNOMEDCT_CORE|Multiple-resistant Staphylococcus aureus infection|Multiple-resistant Staphylococcus aureus infection
C0560024|T184|PT|193967004|SNOMEDCT_CORE|Swelling of eyelid|Swelling of eyelid
C0560024|T184|FN|193967004|SNOMEDCT_CORE|Swelling of eyelid|Swelling of eyelid
C0560619|T037|PT|282752000|SNOMEDCT_CORE|Injury of eye region|Injury of eye region
C0560619|T037|FN|282752000|SNOMEDCT_CORE|Injury of eye region|Injury of eye region
C0560619|T037|SY|282752000|SNOMEDCT_CORE|Periocular injury|Injury of eye region
C0560626|T037|PT|282760004|SNOMEDCT_CORE|Clavicle injury|Clavicle injury
C0560626|T037|FN|282760004|SNOMEDCT_CORE|Clavicle injury|Clavicle injury
C0560626|T037|SY|282760004|SNOMEDCT_CORE|Collar bone injury|Clavicle injury
C0560641|T037|PT|282776008|SNOMEDCT_CORE|Injury of toe|Injury of toe
C0560641|T037|FN|282776008|SNOMEDCT_CORE|Injury of toe|Injury of toe
C0560647|T037|PT|282782006|SNOMEDCT_CORE|Injury of scrotum|Injury of scrotum
C0560647|T037|FN|282782006|SNOMEDCT_CORE|Injury of scrotum|Injury of scrotum
C0560960|T037|PT|283062009|SNOMEDCT_CORE|Abrasion of lower limb|Abrasion of lower limb
C0560960|T037|FN|283062009|SNOMEDCT_CORE|Abrasion of lower limb|Abrasion of lower limb
C0560960|T037|SY|283062009|SNOMEDCT_CORE|Graze of leg|Abrasion of lower limb
C0561236|T037|PT|283359004|SNOMEDCT_CORE|Laceration of forehead|Laceration of forehead
C0561236|T037|FN|283359004|SNOMEDCT_CORE|Laceration of forehead|Laceration of forehead
C0561241|T037|PT|283363006|SNOMEDCT_CORE|Laceration of lip|Laceration of lip
C0561241|T037|FN|283363006|SNOMEDCT_CORE|Laceration of lip|Laceration of lip
C0561369|T037|PT|283497000|SNOMEDCT_CORE|Puncture wound of skin|Puncture wound of skin
C0561369|T037|FN|283497000|SNOMEDCT_CORE|Puncture wound of skin|Puncture wound of skin
C0561596|T037|PT|283734005|SNOMEDCT_CORE|Dog bite - wound|Dog bite - wound
C0561596|T037|FN|283734005|SNOMEDCT_CORE|Dog bite - wound|Dog bite - wound
C0561644|T037|PT|283782004|SNOMEDCT_CORE|Cat bite - wound|Cat bite - wound
C0561644|T037|FN|283782004|SNOMEDCT_CORE|Cat bite - wound|Cat bite - wound
C0562083|T037|PT|284220000|SNOMEDCT_CORE|Burn of genitalia|Burn of genitalia
C0562083|T037|FN|284220000|SNOMEDCT_CORE|Burn of genitalia|Burn of genitalia
C0562086|T037|PT|11868005|SNOMEDCT_CORE|Burn of multiple sites of trunk|Burn of multiple sites of trunk
C0562086|T037|FN|11868005|SNOMEDCT_CORE|Burn of multiple sites of trunk|Burn of multiple sites of trunk
C0562086|T037|IS|11868005|SNOMEDCT_CORE|Burn of multiple sites of trunk, NOS|Burn of multiple sites of trunk
C0562086|T037|SY|11868005|SNOMEDCT_CORE|Multiple burns of trunk|Burn of multiple sites of trunk
C0562381|T033|SY|386702006|SNOMEDCT_CORE|Abuse|Victim of abuse
C0562381|T033|IS|386702006|SNOMEDCT_CORE|Abuse, NOS|Victim of abuse
C0562381|T033|SY|386702006|SNOMEDCT_CORE|Abused person|Victim of abuse
C0562381|T033|IS|386702006|SNOMEDCT_CORE|Abused person, NOS|Victim of abuse
C0562381|T033|FN|386702006|SNOMEDCT_CORE|Victim of abuse|Victim of abuse
C0562381|T033|PT|386702006|SNOMEDCT_CORE|Victim of abuse|Victim of abuse
C0562381|T033|IS|386702006|SNOMEDCT_CORE|Victim of abuse, NOS|Victim of abuse
C0562383|T033|PT|225824003|SNOMEDCT_CORE|Victim of physical abuse|Victim of physical abuse
C0562383|T033|FN|225824003|SNOMEDCT_CORE|Victim of physical abuse|Victim of physical abuse
C0562422|T047|OAF|284480000|SNOMEDCT_CORE|Cellulitis of arm|Cellulitis of arm
C0562422|T047|OAP|284480000|SNOMEDCT_CORE|Cellulitis of arm|Cellulitis of arm
C0562512|T037|PT|125664002|SNOMEDCT_CORE|Open wound of toe|Open wound of toe
C0562512|T037|FN|125664002|SNOMEDCT_CORE|Open wound of toe|Open wound of toe
C0562961|T033|PT|285055002|SNOMEDCT_CORE|Does use hearing aid|Does use hearing aid
C0562961|T033|FN|285055002|SNOMEDCT_CORE|Does use hearing aid|Does use hearing aid
C0562961|T033|SY|285055002|SNOMEDCT_CORE|Uses hearing aid|Does use hearing aid
C0563211|T191|PT|285310000|SNOMEDCT_CORE|Carcinoma of anal canal|Carcinoma of anal canal
C0563211|T191|FN|285310000|SNOMEDCT_CORE|Carcinoma of anal canal|Carcinoma of anal canal
C0563242|T037|PT|285348005|SNOMEDCT_CORE|Strain of abdominal muscle|Strain of abdominal muscle
C0563242|T037|FN|285348005|SNOMEDCT_CORE|Strain of abdominal muscle|Strain of abdominal muscle
C0563269|T047|PT|285381006|SNOMEDCT_CORE|Acute infective exacerbation of chronic obstructive airways disease|Acute infective exacerbation of chronic obstructive airways disease
C0563269|T047|FN|285381006|SNOMEDCT_CORE|Acute infective exacerbation of chronic obstructive airways disease|Acute infective exacerbation of chronic obstructive airways disease
C0563273|T033|PT|285384003|SNOMEDCT_CORE|General health deterioration|General health deterioration
C0563273|T033|FN|285384003|SNOMEDCT_CORE|General health deterioration|General health deterioration
C0563276|T184|PT|285387005|SNOMEDCT_CORE|Left sided abdominal pain|Left sided abdominal pain
C0563276|T184|FN|285387005|SNOMEDCT_CORE|Left sided abdominal pain|Left sided abdominal pain
C0564221|T033|SY|286378009|SNOMEDCT_CORE|Difficulty speaking|Difficulty talking
C0564221|T033|PT|286378009|SNOMEDCT_CORE|Difficulty talking|Difficulty talking
C0564221|T033|FN|286378009|SNOMEDCT_CORE|Difficulty talking|Difficulty talking
C0564705|T191|OAP|286892007|SNOMEDCT_CORE|Ca breast - nipple/central|Ca breast - nipple/central
C0564705|T191|OAF|286892007|SNOMEDCT_CORE|Ca breast - nipple/central|Ca breast - nipple/central
C0564708|T191|PT|286895009|SNOMEDCT_CORE|Carcinoma of breast - upper, outer quadrant|Carcinoma of breast - upper, outer quadrant
C0564708|T191|FN|286895009|SNOMEDCT_CORE|Carcinoma of breast - upper, outer quadrant|Carcinoma of breast - upper, outer quadrant
C0564714|T191|OAP|286903005|SNOMEDCT_CORE|Skin - benign mole and naevus|Skin - benign mole and naevus
C0564714|T191|OAP|286903005|SNOMEDCT_CORE|Skin - benign mole and nevus|Skin - benign mole and naevus
C0564714|T191|OAF|286903005|SNOMEDCT_CORE|Skin - benign mole and nevus|Skin - benign mole and naevus
C0564785|T047|PT|287007001|SNOMEDCT_CORE|Rheumatoid arthritis - hand joint|Rheumatoid arthritis - hand joint
C0564785|T047|OF|287007001|SNOMEDCT_CORE|Rheumatoid arthritis - hand joint|Rheumatoid arthritis - hand joint
C0564785|T047|SY|287007001|SNOMEDCT_CORE|Rheumatoid arthritis of hand|Rheumatoid arthritis - hand joint
C0564785|T047|SY|287007001|SNOMEDCT_CORE|Rheumatoid arthritis of hand joint|Rheumatoid arthritis - hand joint
C0564785|T047|FN|287007001|SNOMEDCT_CORE|Rheumatoid arthritis of hand joint|Rheumatoid arthritis - hand joint
C0564794|T047|PT|287018001|SNOMEDCT_CORE|Synovitis/tenosynovitis - elbow|Synovitis/tenosynovitis - elbow
C0564794|T047|FN|287018001|SNOMEDCT_CORE|Synovitis/tenosynovitis - elbow|Synovitis/tenosynovitis - elbow
C0564797|T047|PT|287021004|SNOMEDCT_CORE|Synovitis/tenosynovitis - knee|Synovitis/tenosynovitis - knee
C0564797|T047|FN|287021004|SNOMEDCT_CORE|Synovitis/tenosynovitis - knee|Synovitis/tenosynovitis - knee
C0564837|T046|PT|287065007|SNOMEDCT_CORE|Pathological fracture - upper arm|Pathological fracture - upper arm
C0564837|T046|FN|287065007|SNOMEDCT_CORE|Pathological fracture - upper arm|Pathological fracture - upper arm
C0564837|T046|SY|287065007|SNOMEDCT_CORE|Pathological fracture of humerus|Pathological fracture - upper arm
C0564858|T037|PT|287097007|SNOMEDCT_CORE|Sprained finger/thumb|Sprained finger/thumb
C0564858|T037|FN|287097007|SNOMEDCT_CORE|Sprained finger/thumb|Sprained finger/thumb
C0565822|T047|FN|267727004|SNOMEDCT_CORE|Blind or low vision - both eyes|Blind or low vision - both eyes
C0565822|T047|PT|267727004|SNOMEDCT_CORE|Blind or low vision - both eyes|Blind or low vision - both eyes
C0565848|T037|PT|269795008|SNOMEDCT_CORE|Foreign body accident - orifice|Foreign body accident - orifice
C0565848|T037|OF|269795008|SNOMEDCT_CORE|Foreign body accident - orifice|Foreign body accident - orifice
C0565848|T037|FN|269795008|SNOMEDCT_CORE|Foreign body accident - orifice|Foreign body accident - orifice
C0566602|T047|PT|197441003|SNOMEDCT_CORE|Primary sclerosing cholangitis|Primary sclerosing cholangitis
C0566602|T047|FN|197441003|SNOMEDCT_CORE|Primary sclerosing cholangitis|Primary sclerosing cholangitis
C0566602|T047|SY|197441003|SNOMEDCT_CORE|PSC - Primary sclerosing cholangitis|Primary sclerosing cholangitis
C0566690|T033|FN|289259007|SNOMEDCT_CORE|Vaginal delivery|Vaginal delivery
C0566690|T033|PT|289259007|SNOMEDCT_CORE|Vaginal delivery|Vaginal delivery
C0566871|T033|PT|289439005|SNOMEDCT_CORE|Fetal heart rate absent|Fetal heart rate absent
C0566871|T033|FN|289439005|SNOMEDCT_CORE|Fetal heart rate absent|Fetal heart rate absent
C0566871|T033|SY|289439005|SNOMEDCT_CORE|Foetal heart rate absent|Fetal heart rate absent
C0566908|T033|SY|289477004|SNOMEDCT_CORE|Lump of vulva|Lump of vulva
C0566943|T046|PT|289517005|SNOMEDCT_CORE|Vaginal lesion|Vaginal lesion
C0566943|T046|FN|289517005|SNOMEDCT_CORE|Vaginal lesion|Vaginal lesion
C0566969|T033|SY|271939006|SNOMEDCT_CORE|Observation of vaginal discharge|Observation of vaginal discharge
C0566991|T033|SY|289572007|SNOMEDCT_CORE|No flow of amniotc liquor|No liquor observed vaginally
C0566991|T033|PT|289572007|SNOMEDCT_CORE|No liquor observed vaginally|No liquor observed vaginally
C0566991|T033|FN|289572007|SNOMEDCT_CORE|No liquor observed vaginally|No liquor observed vaginally
C0567312|T033|SY|289903006|SNOMEDCT_CORE|Menopause|Menopause present
C0567312|T033|FN|289903006|SNOMEDCT_CORE|Menopause present|Menopause present
C0567312|T033|PT|289903006|SNOMEDCT_CORE|Menopause present|Menopause present
C0567322|T033|PT|289917002|SNOMEDCT_CORE|History of bladder neoplasm|History of bladder neoplasm
C0567322|T033|OF|289917002|SNOMEDCT_CORE|History of bladder neoplasm|History of bladder neoplasm
C0567322|T033|FN|289917002|SNOMEDCT_CORE|History of bladder neoplasm|History of bladder neoplasm
C0569491|T046|PT|292196008|SNOMEDCT_CORE|Antineoplastic adverse reaction|Antineoplastic adverse reaction
C0569491|T046|FN|292196008|SNOMEDCT_CORE|Antineoplastic adverse reaction|Antineoplastic adverse reaction
C0572025|T037|PT|295124009|SNOMEDCT_CORE|Acetaminophen overdose|Acetaminophen overdose
C0572025|T037|FN|295124009|SNOMEDCT_CORE|Acetaminophen overdose|Acetaminophen overdose
C0572025|T037|PTGB|295124009|SNOMEDCT_CORE|Paracetamol overdose|Acetaminophen overdose
C0572025|T037|OF|295124009|SNOMEDCT_CORE|Paracetamol overdose|Acetaminophen overdose
C0572933|T037|PT|296053004|SNOMEDCT_CORE|Benzodiazepine overdose|Benzodiazepine overdose
C0572933|T037|FN|296053004|SNOMEDCT_CORE|Benzodiazepine overdose|Benzodiazepine overdose
C0573797|T037|PT|47546008|SNOMEDCT_CORE|Warfarin overdosage|Warfarin overdosage
C0573797|T037|FN|47546008|SNOMEDCT_CORE|Warfarin overdosage|Warfarin overdosage
C0573797|T037|SY|47546008|SNOMEDCT_CORE|Warfarin overdose|Warfarin overdosage
C0573993|T191|PT|92380000|SNOMEDCT_CORE|Benign neoplasm of skin of trunk|Benign neoplasm of skin of trunk
C0573993|T191|FN|92380000|SNOMEDCT_CORE|Benign neoplasm of skin of trunk|Benign neoplasm of skin of trunk
C0573993|T191|IS|92380000|SNOMEDCT_CORE|Benign neoplasm of skin of trunk, NOS|Benign neoplasm of skin of trunk
C0574002|T184|FN|102576009|SNOMEDCT_CORE|Edema of foot|Edema of foot
C0574002|T184|PT|102576009|SNOMEDCT_CORE|Edema of foot|Edema of foot
C0574002|T184|SY|102576009|SNOMEDCT_CORE|Foot edema|Edema of foot
C0574002|T184|SYGB|102576009|SNOMEDCT_CORE|Foot oedema|Edema of foot
C0574002|T184|PTGB|102576009|SNOMEDCT_CORE|Oedema of foot|Edema of foot
C0574002|T184|SY|102576009|SNOMEDCT_CORE|Pedal edema|Edema of foot
C0574002|T184|SYGB|102576009|SNOMEDCT_CORE|Pedal oedema|Edema of foot
C0574035|T037|SY|297186008|SNOMEDCT_CORE|Motorbike accident|Motorcycle accident
C0574035|T037|PT|297186008|SNOMEDCT_CORE|Motorcycle accident|Motorcycle accident
C0574035|T037|OF|297186008|SNOMEDCT_CORE|Motorcycle accident|Motorcycle accident
C0574035|T037|FN|297186008|SNOMEDCT_CORE|Motorcycle accident|Motorcycle accident
C0574068|T184|PT|297217002|SNOMEDCT_CORE|Rib pain|Rib pain
C0574068|T184|FN|297217002|SNOMEDCT_CORE|Rib pain|Rib pain
C0574718|T047|PT|297946004|SNOMEDCT_CORE|Lower limb nerve lesion|Lower limb nerve lesion
C0574718|T047|FN|297946004|SNOMEDCT_CORE|Lower limb nerve lesion|Lower limb nerve lesion
C0574785|T184|PT|307541003|SNOMEDCT_CORE|Lower urinary tract symptoms|Lower urinary tract symptoms
C0574785|T184|FN|307541003|SNOMEDCT_CORE|Lower urinary tract symptoms|Lower urinary tract symptoms
C0574785|T184|SY|307541003|SNOMEDCT_CORE|LUTS - Lower urinary tract symptoms|Lower urinary tract symptoms
C0574869|T037|PT|298083004|SNOMEDCT_CORE|Foreign body of skin of finger|Foreign body of skin of finger
C0574869|T037|FN|298083004|SNOMEDCT_CORE|Foreign body of skin of finger|Foreign body of skin of finger
C0574943|T033|IS|298162008|SNOMEDCT_CORE|Shoulder joint active|Shoulder joint inflamed
C0574943|T033|PT|298162008|SNOMEDCT_CORE|Shoulder joint inflamed|Shoulder joint inflamed
C0574943|T033|FN|298162008|SNOMEDCT_CORE|Shoulder joint inflamed|Shoulder joint inflamed
C0574945|T033|IS|298164009|SNOMEDCT_CORE|Wrist joint active|Wrist joint inflamed
C0574945|T033|PT|298164009|SNOMEDCT_CORE|Wrist joint inflamed|Wrist joint inflamed
C0574945|T033|FN|298164009|SNOMEDCT_CORE|Wrist joint inflamed|Wrist joint inflamed
C0574946|T033|IS|298165005|SNOMEDCT_CORE|Hand joint active|Hand joint inflamed
C0574946|T033|PT|298165005|SNOMEDCT_CORE|Hand joint inflamed|Hand joint inflamed
C0574946|T033|FN|298165005|SNOMEDCT_CORE|Hand joint inflamed|Hand joint inflamed
C0574948|T033|IS|298167002|SNOMEDCT_CORE|Finger joint active|Finger joint inflamed
C0574948|T033|PT|298167002|SNOMEDCT_CORE|Finger joint inflamed|Finger joint inflamed
C0574948|T033|FN|298167002|SNOMEDCT_CORE|Finger joint inflamed|Finger joint inflamed
C0574950|T033|IS|298169004|SNOMEDCT_CORE|Hip joint active|Hip joint inflamed
C0574950|T033|PT|298169004|SNOMEDCT_CORE|Hip joint inflamed|Hip joint inflamed
C0574950|T033|FN|298169004|SNOMEDCT_CORE|Hip joint inflamed|Hip joint inflamed
C0574952|T033|IS|298171004|SNOMEDCT_CORE|Ankle joint active|Ankle joint inflamed
C0574952|T033|PT|298171004|SNOMEDCT_CORE|Ankle joint inflamed|Ankle joint inflamed
C0574952|T033|FN|298171004|SNOMEDCT_CORE|Ankle joint inflamed|Ankle joint inflamed
C0574953|T033|IS|298172006|SNOMEDCT_CORE|Foot joint active|Foot joint inflamed
C0574953|T033|PT|298172006|SNOMEDCT_CORE|Foot joint inflamed|Foot joint inflamed
C0574953|T033|FN|298172006|SNOMEDCT_CORE|Foot joint inflamed|Foot joint inflamed
C0574960|T047|PT|55146009|SNOMEDCT_CORE|Inflammation of sacroiliac joint|Inflammation of sacroiliac joint
C0574960|T047|FN|55146009|SNOMEDCT_CORE|Inflammation of sacroiliac joint|Inflammation of sacroiliac joint
C0574960|T047|IS|55146009|SNOMEDCT_CORE|Inflammation of sacroiliac joint, NOS|Inflammation of sacroiliac joint
C0574960|T047|IS|55146009|SNOMEDCT_CORE|Sacroiliac joint active|Inflammation of sacroiliac joint
C0574960|T047|SY|55146009|SNOMEDCT_CORE|Sacroiliac joint inflamed|Inflammation of sacroiliac joint
C0574960|T047|OF|55146009|SNOMEDCT_CORE|Sacroiliac joint inflamed|Inflammation of sacroiliac joint
C0574960|T047|IS|55146009|SNOMEDCT_CORE|Sacroiliitis|Inflammation of sacroiliac joint
C0574960|T047|IS|55146009|SNOMEDCT_CORE|Sacroiliitis, NOS|Inflammation of sacroiliac joint
C0575002|T184|PT|298222004|SNOMEDCT_CORE|Active range of joint movement reduced|Active range of joint movement reduced
C0575002|T184|FN|298222004|SNOMEDCT_CORE|Active range of joint movement reduced|Active range of joint movement reduced
C0575081|T033|PT|22325002|SNOMEDCT_CORE|Abnormal gait|Abnormal gait
C0575081|T033|FN|22325002|SNOMEDCT_CORE|Abnormal gait|Abnormal gait
C0575081|T033|IS|22325002|SNOMEDCT_CORE|Abnormal gait, NOS|Abnormal gait
C0575081|T033|SY|22325002|SNOMEDCT_CORE|Gait abnormality|Abnormal gait
C0575081|T033|IS|22325002|SNOMEDCT_CORE|Gait abnormality, NOS|Abnormal gait
C0575081|T033|SY|22325002|SNOMEDCT_CORE|Gait difficulty|Abnormal gait
C0575081|T033|SY|22325002|SNOMEDCT_CORE|Gait problem|Abnormal gait
C0575081|T033|OF|22325002|SNOMEDCT_CORE|Gait problem|Abnormal gait
C0575152|T033|SY|298375002|SNOMEDCT_CORE|Temporomandibular joint tender|Tenderness of temporomandibular joint
C0575152|T033|OF|298375002|SNOMEDCT_CORE|Temporomandibular joint tender|Tenderness of temporomandibular joint
C0575152|T033|PT|298375002|SNOMEDCT_CORE|Tenderness of temporomandibular joint|Tenderness of temporomandibular joint
C0575152|T033|FN|298375002|SNOMEDCT_CORE|Tenderness of temporomandibular joint|Tenderness of temporomandibular joint
C0575270|T047|SY|298494008|SNOMEDCT_CORE|Scoliosis of dorsal spine|Scoliosis of thoracic spine
C0575270|T047|PT|298494008|SNOMEDCT_CORE|Scoliosis of thoracic spine|Scoliosis of thoracic spine
C0575270|T047|OF|298494008|SNOMEDCT_CORE|Scoliosis of thoracic spine|Scoliosis of thoracic spine
C0575270|T047|FN|298494008|SNOMEDCT_CORE|Scoliosis of thoracic spine|Scoliosis of thoracic spine
C0575367|T033|SY|298591003|SNOMEDCT_CORE|Lumbar spine scoliosis|Scoliosis of lumbar spine
C0575367|T033|OF|298591003|SNOMEDCT_CORE|Lumbar spine scoliosis|Scoliosis of lumbar spine
C0575367|T033|PT|298591003|SNOMEDCT_CORE|Scoliosis of lumbar spine|Scoliosis of lumbar spine
C0575367|T033|FN|298591003|SNOMEDCT_CORE|Scoliosis of lumbar spine|Scoliosis of lumbar spine
C0575503|T033|PT|298731003|SNOMEDCT_CORE|Pain of sternum|Pain of sternum
C0575503|T033|FN|298731003|SNOMEDCT_CORE|Pain of sternum|Pain of sternum
C0575544|T033|PT|298772001|SNOMEDCT_CORE|Shoulder joint deformity|Shoulder joint deformity
C0575544|T033|FN|298772001|SNOMEDCT_CORE|Shoulder joint deformity|Shoulder joint deformity
C0575624|T033|SY|298854003|SNOMEDCT_CORE|Shoulder joint instability|Shoulder joint unstable
C0575624|T033|PT|298854003|SNOMEDCT_CORE|Shoulder joint unstable|Shoulder joint unstable
C0575624|T033|FN|298854003|SNOMEDCT_CORE|Shoulder joint unstable|Shoulder joint unstable
C0575695|T033|SY|298924009|SNOMEDCT_CORE|Elbow joint instability|Elbow joint unstable
C0575695|T033|PT|298924009|SNOMEDCT_CORE|Elbow joint unstable|Elbow joint unstable
C0575695|T033|FN|298924009|SNOMEDCT_CORE|Elbow joint unstable|Elbow joint unstable
C0575805|T033|FN|299037003|SNOMEDCT_CORE|Swelling of hand|Swelling of hand
C0575805|T033|PT|299037003|SNOMEDCT_CORE|Swelling of hand|Swelling of hand
C0575805|T033|SY|299037003|SNOMEDCT_CORE|Swollen hand|Swelling of hand
C0575810|T033|PT|299042006|SNOMEDCT_CORE|Weakness of hand|Weakness of hand
C0575810|T033|FN|299042006|SNOMEDCT_CORE|Weakness of hand|Weakness of hand
C0576091|T190|PT|299328006|SNOMEDCT_CORE|Deformity of knee joint|Deformity of knee joint
C0576091|T190|FN|299328006|SNOMEDCT_CORE|Deformity of knee joint|Deformity of knee joint
C0576404|T033|SY|299647001|SNOMEDCT_CORE|Amputated - transfemoral|Amputated above knee
C0576404|T033|FN|299647001|SNOMEDCT_CORE|Amputated above knee|Amputated above knee
C0576404|T033|PT|299647001|SNOMEDCT_CORE|Amputated above knee|Amputated above knee
C0576456|T033|PT|299698007|SNOMEDCT_CORE|Feeding poor|Feeding poor
C0576456|T033|FN|299698007|SNOMEDCT_CORE|Feeding poor|Feeding poor
C0576456|T033|SY|299698007|SNOMEDCT_CORE|Poor feeding|Feeding poor
C0576825|T033|PT|300092000|SNOMEDCT_CORE|Lesion of external ear|Lesion of external ear
C0576825|T033|FN|300092000|SNOMEDCT_CORE|Lesion of external ear|Lesion of external ear
C0576825|T033|OF|300092000|SNOMEDCT_CORE|Lesion of external ear|Lesion of external ear
C0576971|T033|PT|300246005|SNOMEDCT_CORE|Lesion of tongue|Lesion of tongue
C0576971|T033|FN|300246005|SNOMEDCT_CORE|Lesion of tongue|Lesion of tongue
C0577053|T033|PT|300331000|SNOMEDCT_CORE|Lesion of liver|Lesion of liver
C0577053|T033|FN|300331000|SNOMEDCT_CORE|Lesion of liver|Lesion of liver
C0577180|T033|PT|300457003|SNOMEDCT_CORE|Lesion of bladder|Lesion of bladder
C0577180|T033|FN|300457003|SNOMEDCT_CORE|Lesion of bladder|Lesion of bladder
C0577215|T033|PT|300492006|SNOMEDCT_CORE|Lesion of testis|Lesion of testis
C0577215|T033|FN|300492006|SNOMEDCT_CORE|Lesion of testis|Lesion of testis
C0577559|T033|IS|300848003|SNOMEDCT_CORE|A mass|Mass of body structure
C0577559|T033|SY|300848003|SNOMEDCT_CORE|Lump|Mass of body structure
C0577559|T033|SY|300848003|SNOMEDCT_CORE|Mass|Mass of body structure
C0577559|T033|PT|300848003|SNOMEDCT_CORE|Mass of body structure|Mass of body structure
C0577559|T033|FN|300848003|SNOMEDCT_CORE|Mass of body structure|Mass of body structure
C0577559|T033|SY|300848003|SNOMEDCT_CORE|Observation of a mass|Mass of body structure
C0577598|T046|OAP|300889000|SNOMEDCT_CORE|Swelling of arm|Swelling of upper arm
C0577598|T046|OAF|300889000|SNOMEDCT_CORE|Swelling of arm|Swelling of upper arm
C0577598|T046|PT|449619004|SNOMEDCT_CORE|Swelling of upper arm|Swelling of upper arm
C0577598|T046|FN|449619004|SNOMEDCT_CORE|Swelling of upper arm|Swelling of upper arm
C0577598|T046|OAS|300889000|SNOMEDCT_CORE|Swollen arm|Swelling of upper arm
C0577657|T047|PT|300950007|SNOMEDCT_CORE|Infected hand|Infected hand
C0577657|T047|FN|300950007|SNOMEDCT_CORE|Infected hand|Infected hand
C0577659|T184|SY|300953009|SNOMEDCT_CORE|Axillary pain|Pain in axilla
C0577659|T184|PT|300953009|SNOMEDCT_CORE|Pain in axilla|Pain in axilla
C0577659|T184|FN|300953009|SNOMEDCT_CORE|Pain in axilla|Pain in axilla
C0577688|T020|PT|300984006|SNOMEDCT_CORE|Skin ulcer of calf|Skin ulcer of calf
C0577688|T020|FN|300984006|SNOMEDCT_CORE|Skin ulcer of calf|Skin ulcer of calf
C0577699|T046|PT|300996004|SNOMEDCT_CORE|Controlled atrial fibrillation|Controlled atrial fibrillation
C0577699|T046|FN|300996004|SNOMEDCT_CORE|Controlled atrial fibrillation|Controlled atrial fibrillation
C0577713|T047|OAP|301016007|SNOMEDCT_CORE|Decubitus ulcer of ankle|Pressure ulcer of ankle
C0577713|T047|OAF|301016007|SNOMEDCT_CORE|Decubitus ulcer of ankle|Pressure ulcer of ankle
C0577713|T047|PT|699211004|SNOMEDCT_CORE|Pressure ulcer of ankle|Pressure ulcer of ankle
C0577713|T047|FN|699211004|SNOMEDCT_CORE|Pressure ulcer of ankle|Pressure ulcer of ankle
C0577716|T047|OAP|301019000|SNOMEDCT_CORE|Decubitus ulcer of dorsum of foot|Pressure ulcer of dorsum of foot
C0577716|T047|OAF|301019000|SNOMEDCT_CORE|Decubitus ulcer of dorsum of foot|Pressure ulcer of dorsum of foot
C0577716|T047|PT|699213001|SNOMEDCT_CORE|Pressure ulcer of dorsum of foot|Pressure ulcer of dorsum of foot
C0577716|T047|FN|699213001|SNOMEDCT_CORE|Pressure ulcer of dorsum of foot|Pressure ulcer of dorsum of foot
C0577717|T047|PT|301021005|SNOMEDCT_CORE|Ulcer of toe|Ulcer of toe
C0577717|T047|FN|301021005|SNOMEDCT_CORE|Ulcer of toe|Ulcer of toe
C0577718|T047|PT|301022003|SNOMEDCT_CORE|Ulcer of heel|Ulcer of heel
C0577718|T047|FN|301022003|SNOMEDCT_CORE|Ulcer of heel|Ulcer of heel
C0577719|T047|OAP|301023008|SNOMEDCT_CORE|Ulcer of calf|Ulcer of calf
C0577719|T047|OAF|301023008|SNOMEDCT_CORE|Ulcer of calf|Ulcer of calf
C0577728|T037|PT|301034006|SNOMEDCT_CORE|Fracture of greater trochanter|Fracture of greater trochanter
C0577728|T037|FN|301034006|SNOMEDCT_CORE|Fracture of greater trochanter|Fracture of greater trochanter
C0577730|T033|SY|105485001|SNOMEDCT_CORE|Domestic stress|Family tension
C0577730|T033|IS|105485001|SNOMEDCT_CORE|Family stress|Family tension
C0577730|T033|PT|105485001|SNOMEDCT_CORE|Family tension|Family tension
C0577730|T033|FN|105485001|SNOMEDCT_CORE|Family tension|Family tension
C0577730|T033|SY|105485001|SNOMEDCT_CORE|Stress at home|Family tension
C0577877|T033|PT|301191003|SNOMEDCT_CORE|Lesion of nose|Lesion of nose
C0577877|T033|FN|301191003|SNOMEDCT_CORE|Lesion of nose|Lesion of nose
C0577887|T047|PT|301202006|SNOMEDCT_CORE|Nasal sinus problem|Nasal sinus problem
C0577887|T047|FN|301202006|SNOMEDCT_CORE|Nasal sinus problem|Nasal sinus problem
C0577903|T033|PT|301218000|SNOMEDCT_CORE|Lesion of vocal cord|Lesion of vocal cord
C0577903|T033|FN|301218000|SNOMEDCT_CORE|Lesion of vocal cord|Lesion of vocal cord
C0578026|T033|PT|301336003|SNOMEDCT_CORE|Body weight problem|Body weight problem
C0578026|T033|FN|301336003|SNOMEDCT_CORE|Body weight problem|Body weight problem
C0578040|T033|PT|301350008|SNOMEDCT_CORE|Lesion of lip|Lesion of lip
C0578040|T033|FN|301350008|SNOMEDCT_CORE|Lesion of lip|Lesion of lip
C0578454|T184|PT|301777002|SNOMEDCT_CORE|Neck swelling|Neck swelling
C0578454|T184|FN|301777002|SNOMEDCT_CORE|Neck swelling|Neck swelling
C0578503|T033|PT|301822002|SNOMEDCT_CORE|Abnormal vaginal bleeding|Abnormal vaginal bleeding
C0578503|T033|FN|301822002|SNOMEDCT_CORE|Abnormal vaginal bleeding|Abnormal vaginal bleeding
C0578590|T033|SY|301913002|SNOMEDCT_CORE|Lesion eyelid|Lesion of eyelid
C0578590|T033|PT|301913002|SNOMEDCT_CORE|Lesion of eyelid|Lesion of eyelid
C0578590|T033|FN|301913002|SNOMEDCT_CORE|Lesion of eyelid|Lesion of eyelid
C0578590|T033|SY|301913002|SNOMEDCT_CORE|Lid lesion|Lesion of eyelid
C0578705|T037|PT|81576005|SNOMEDCT_CORE|Closed fracture of phalanx of foot|Closed fracture of phalanx of foot
C0578705|T037|FN|81576005|SNOMEDCT_CORE|Closed fracture of phalanx of foot|Closed fracture of phalanx of foot
C0578705|T037|SY|81576005|SNOMEDCT_CORE|Closed fracture of phalanx of toe|Closed fracture of phalanx of foot
C0578705|T037|SY|81576005|SNOMEDCT_CORE|Closed fracture of toe|Closed fracture of phalanx of foot
C0578706|T037|PT|74395007|SNOMEDCT_CORE|Open fracture of phalanx of foot|Open fracture of phalanx of foot
C0578706|T037|FN|74395007|SNOMEDCT_CORE|Open fracture of phalanx of foot|Open fracture of phalanx of foot
C0578706|T037|SY|74395007|SNOMEDCT_CORE|Open fracture of phalanx of toe|Open fracture of phalanx of foot
C0578706|T037|SY|74395007|SNOMEDCT_CORE|Open fracture of toe|Open fracture of phalanx of foot
C0578735|T046|PT|127189005|SNOMEDCT_CORE|Axillary lymphadenopathy|Axillary lymphadenopathy
C0578735|T046|FN|127189005|SNOMEDCT_CORE|Axillary lymphadenopathy|Axillary lymphadenopathy
C0578736|T047|SY|127199000|SNOMEDCT_CORE|Groin lymphadenopathy|Inguinal lymphadenopathy
C0578736|T047|PT|127199000|SNOMEDCT_CORE|Inguinal lymphadenopathy|Inguinal lymphadenopathy
C0578736|T047|FN|127199000|SNOMEDCT_CORE|Inguinal lymphadenopathy|Inguinal lymphadenopathy
C0578757|T033|PT|102500002|SNOMEDCT_CORE|Good neonatal condition at birth|Good neonatal condition at birth
C0578757|T033|FN|102500002|SNOMEDCT_CORE|Good neonatal condition at birth|Good neonatal condition at birth
C0578757|T033|SY|102500002|SNOMEDCT_CORE|Healthy newborn|Good neonatal condition at birth
C0578757|T033|IS|102500002|SNOMEDCT_CORE|Well newborn|Good neonatal condition at birth
C0578883|T033|PT|271437004|SNOMEDCT_CORE|Problem situation relating to social and personal history|Problem situation relating to social and personal history
C0578883|T033|FN|271437004|SNOMEDCT_CORE|Problem situation relating to social and personal history|Problem situation relating to social and personal history
C0579065|T047|SY|190368000|SNOMEDCT_CORE|Insulin-dependent diabetes mellitus with ulcer|Type 1 diabetes mellitus with ulcer
C0579065|T047|PT|190368000|SNOMEDCT_CORE|Type 1 diabetes mellitus with ulcer|Type 1 diabetes mellitus with ulcer
C0579065|T047|FN|190368000|SNOMEDCT_CORE|Type I diabetes mellitus with ulcer|Type 1 diabetes mellitus with ulcer
C0579065|T047|SY|190368000|SNOMEDCT_CORE|Type I diabetes mellitus with ulcer|Type 1 diabetes mellitus with ulcer
C0579066|T047|IS|190389009|SNOMEDCT_CORE|Non-insulin-dependent diabetes mellitus with ulcer|Type 2 diabetes mellitus with ulcer
C0579066|T047|PT|190389009|SNOMEDCT_CORE|Type 2 diabetes mellitus with ulcer|Type 2 diabetes mellitus with ulcer
C0579066|T047|FN|190389009|SNOMEDCT_CORE|Type II diabetes mellitus with ulcer|Type 2 diabetes mellitus with ulcer
C0579066|T047|SY|190389009|SNOMEDCT_CORE|Type II diabetes mellitus with ulcer|Type 2 diabetes mellitus with ulcer
C0579122|T047|IS|421631007|SNOMEDCT_CORE|Diabetes type 2 with gangrene|Gangrene due to type 2 diabetes mellitus
C0579122|T047|IS|421631007|SNOMEDCT_CORE|Gangrene associated with adult-onside type diabetes mellitus|Gangrene due to type 2 diabetes mellitus
C0579122|T047|IS|421631007|SNOMEDCT_CORE|Gangrene associated with non-insulin dependent diabetes mellitus|Gangrene due to type 2 diabetes mellitus
C0579122|T047|OP|421631007|SNOMEDCT_CORE|Gangrene associated with type 2 diabetes mellitus|Gangrene due to type 2 diabetes mellitus
C0579122|T047|OF|421631007|SNOMEDCT_CORE|Gangrene associated with type II diabetes mellitus|Gangrene due to type 2 diabetes mellitus
C0579122|T047|IS|421631007|SNOMEDCT_CORE|Gangrene associated with type II diabetes mellitus|Gangrene due to type 2 diabetes mellitus
C0579122|T047|PT|421631007|SNOMEDCT_CORE|Gangrene due to type 2 diabetes mellitus|Gangrene due to type 2 diabetes mellitus
C0579122|T047|FN|421631007|SNOMEDCT_CORE|Gangrene due to type 2 diabetes mellitus|Gangrene due to type 2 diabetes mellitus
C0579122|T047|IS|190390000|SNOMEDCT_CORE|Non-insulin-dependent diabetes mellitus with gangrene|Gangrene due to type 2 diabetes mellitus
C0579122|T047|OAP|190390000|SNOMEDCT_CORE|Type 2 diabetes mellitus with gangrene|Gangrene due to type 2 diabetes mellitus
C0579122|T047|OAF|190390000|SNOMEDCT_CORE|Type II diabetes mellitus with gangrene|Gangrene due to type 2 diabetes mellitus
C0579122|T047|OAS|190390000|SNOMEDCT_CORE|Type II diabetes mellitus with gangrene|Gangrene due to type 2 diabetes mellitus
C0579124|T047|OAS|190392008|SNOMEDCT_CORE|Non-insulin-dependent diabetes mellitus - poor control|Type II diabetes mellitus - poor control
C0579124|T047|OAS|190392008|SNOMEDCT_CORE|Type 2 diabetes mellitus - poor control|Type II diabetes mellitus - poor control
C0579124|T047|OAF|190392008|SNOMEDCT_CORE|Type II diabetes mellitus - poor control|Type II diabetes mellitus - poor control
C0579124|T047|OAP|190392008|SNOMEDCT_CORE|Type II diabetes mellitus - poor control|Type II diabetes mellitus - poor control
C0580094|T033|SY|161155000|SNOMEDCT_CORE|School difficulties|School problem
C0580094|T033|FN|161155000|SNOMEDCT_CORE|School problem|School problem
C0580094|T033|PT|161155000|SNOMEDCT_CORE|School problem|School problem
C0580173|T033|SY|303081002|SNOMEDCT_CORE|Intermittent spinal claudication|Neurogenic claudication
C0580173|T033|PT|303081002|SNOMEDCT_CORE|Neurogenic claudication|Neurogenic claudication
C0580173|T033|FN|303081002|SNOMEDCT_CORE|Neurogenic claudication|Neurogenic claudication
C0580173|T033|SY|303081002|SNOMEDCT_CORE|Pseudoclaudication|Neurogenic claudication
C0580173|T033|SY|303081002|SNOMEDCT_CORE|Spinal claudication|Neurogenic claudication
C0580284|T191|PT|303194003|SNOMEDCT_CORE|Metastasis to head and neck lymph node|Metastasis to head and neck lymph node
C0580284|T191|FN|303194003|SNOMEDCT_CORE|Metastasis to head and neck lymph node|Metastasis to head and neck lymph node
C0580467|T033|PT|166584001|SNOMEDCT_CORE|C-reactive protein abnormal|C-reactive protein abnormal
C0580467|T033|FN|166584001|SNOMEDCT_CORE|C-reactive protein abnormal|C-reactive protein abnormal
C0580476|T033|OF|166669000|SNOMEDCT_CORE|Aspartate aminotransferase /serum glutamic oxaloacetic transaminase level raised|Aspartate aminotransferase serum level raised
C0580476|T033|IS|166669000|SNOMEDCT_CORE|Aspartate aminotransferase /serum glutamic oxaloacetic transaminase level raised|Aspartate aminotransferase serum level raised
C0580476|T033|PT|166669000|SNOMEDCT_CORE|Aspartate aminotransferase serum level raised|Aspartate aminotransferase serum level raised
C0580476|T033|FN|166669000|SNOMEDCT_CORE|Aspartate aminotransferase serum level raised|Aspartate aminotransferase serum level raised
C0580476|T033|OF|166669000|SNOMEDCT_CORE|Aspartate aminotransferase/serum glutamic oxaloacetic transaminase level raised|Aspartate aminotransferase serum level raised
C0580476|T033|IS|166669000|SNOMEDCT_CORE|Aspartate aminotransferase/serum glutamic oxaloacetic transaminase level raised|Aspartate aminotransferase serum level raised
C0580476|T033|SY|166669000|SNOMEDCT_CORE|AST serum level raised|Aspartate aminotransferase serum level raised
C0580476|T033|OP|166669000|SNOMEDCT_CORE|AST/SGOT level raised|Aspartate aminotransferase serum level raised
C0580476|T033|OF|166669000|SNOMEDCT_CORE|AST/SGOT level raised|Aspartate aminotransferase serum level raised
C0580476|T033|SY|166669000|SNOMEDCT_CORE|Serum glutamic oxaloacetic transaminase level raised|Aspartate aminotransferase serum level raised
C0580520|T033|OAP|275984001|SNOMEDCT_CORE|Immunisation refused|Immunisation refused
C0580520|T033|OAP|275984001|SNOMEDCT_CORE|Immunization refused|Immunisation refused
C0580520|T033|OAF|275984001|SNOMEDCT_CORE|Immunization refused|Immunisation refused
C0580546|T033|PT|166922008|SNOMEDCT_CORE|Blood glucose abnormal|Blood glucose abnormal
C0580546|T033|FN|166922008|SNOMEDCT_CORE|Blood glucose abnormal|Blood glucose abnormal
C0580555|T033|PT|166160000|SNOMEDCT_CORE|Prostate specific antigen abnormal|Prostate specific antigen abnormal
C0580555|T033|FN|166160000|SNOMEDCT_CORE|Prostate specific antigen abnormal|Prostate specific antigen abnormal
C0580703|T033|PT|183646003|SNOMEDCT_CORE|Postoperative visit|Postoperative visit
C0580703|T033|FN|183646003|SNOMEDCT_CORE|Postoperative visit|Postoperative visit
C0580979|T033|PT|170544002|SNOMEDCT_CORE|Requires a meningitis vaccination|Requires a meningitis vaccination
C0580979|T033|FN|170544002|SNOMEDCT_CORE|Requires a meningitis vaccination|Requires a meningitis vaccination
C0581024|T033|OAP|170536002|SNOMEDCT_CORE|Vaccination required|Vaccination required
C0581024|T033|OAF|170536002|SNOMEDCT_CORE|Vaccination required|Vaccination required
C0581025|T033|IS|170537006|SNOMEDCT_CORE|Requires a booster tetanus|Requires a tetanus booster
C0581025|T033|OF|170537006|SNOMEDCT_CORE|Requires a booster tetanus|Requires a tetanus booster
C0581025|T033|PT|170537006|SNOMEDCT_CORE|Requires a tetanus booster|Requires a tetanus booster
C0581025|T033|FN|170537006|SNOMEDCT_CORE|Requires a tetanus booster|Requires a tetanus booster
C0581027|T033|PT|170539009|SNOMEDCT_CORE|Requires polio vaccination|Requires polio vaccination
C0581027|T033|FN|170539009|SNOMEDCT_CORE|Requires polio vaccination|Requires polio vaccination
C0581077|T033|PT|161626009|SNOMEDCT_CORE|H/O splenectomy|H/O splenectomy
C0581077|T033|OF|161626009|SNOMEDCT_CORE|History of - splenectomy|H/O splenectomy
C0581077|T033|IS|161626009|SNOMEDCT_CORE|History of - splenectomy|H/O splenectomy
C0581077|T033|FN|161626009|SNOMEDCT_CORE|History of splenectomy|H/O splenectomy
C0581077|T033|SY|161626009|SNOMEDCT_CORE|History of splenectomy|H/O splenectomy
C0581118|T033|PT|169255008|SNOMEDCT_CORE|Ultrasound scan abnormal|Ultrasound scan abnormal
C0581118|T033|FN|169255008|SNOMEDCT_CORE|Ultrasound scan abnormal|Ultrasound scan abnormal
C0581275|T047|SY|235774002|SNOMEDCT_CORE|Abscess of colon co-occurrent and due to diverticular disease of colon|Abscess with diverticular disease of colon
C0581275|T047|FN|235774002|SNOMEDCT_CORE|Abscess of colon co-occurrent and due to diverticular disease of colon|Abscess with diverticular disease of colon
C0581275|T047|PT|235774002|SNOMEDCT_CORE|Abscess with diverticular disease of colon|Abscess with diverticular disease of colon
C0581275|T047|SY|235774002|SNOMEDCT_CORE|Colonic diverticular abscess|Abscess with diverticular disease of colon
C0581275|T047|OF|235774002|SNOMEDCT_CORE|Colonic diverticular abscess|Abscess with diverticular disease of colon
C0581275|T047|SY|235774002|SNOMEDCT_CORE|Diverticular abscess|Abscess with diverticular disease of colon
C0581305|T037|PT|211311003|SNOMEDCT_CORE|Foreign body in hand|Foreign body in hand
C0581305|T037|FN|211311003|SNOMEDCT_CORE|Foreign body in hand|Foreign body in hand
C0581351|T033|SY|161882006|SNOMEDCT_CORE|Crick in neck|Crick in neck
C0581352|T047|SY|202805003|SNOMEDCT_CORE|Arthropathy of sacroiliac joint|Sacroiliac disorder
C0581352|T047|PT|202805003|SNOMEDCT_CORE|Sacroiliac disorder|Sacroiliac disorder
C0581352|T047|FN|202805003|SNOMEDCT_CORE|Sacroiliac disorder|Sacroiliac disorder
C0581354|T047|PT|195788001|SNOMEDCT_CORE|Recurrent sinusitis|Recurrent sinusitis
C0581354|T047|FN|195788001|SNOMEDCT_CORE|Recurrent sinusitis|Recurrent sinusitis
C0581360|T047|IS|197092000|SNOMEDCT_CORE|Bleeding diverticulosis|Hemorrhage of large intestine with diverticular disease of large intestine
C0581360|T047|OF|197092000|SNOMEDCT_CORE|Bleeding diverticulosis|Hemorrhage of large intestine with diverticular disease of large intestine
C0581360|T047|SY|197092000|SNOMEDCT_CORE|Bleeding diverticulosis of large intestine|Hemorrhage of large intestine with diverticular disease of large intestine
C0581360|T047|SYGB|197092000|SNOMEDCT_CORE|Haemorrhage of large intestine co-occurrent and due to diverticular disease of large intestine|Hemorrhage of large intestine with diverticular disease of large intestine
C0581360|T047|PTGB|197092000|SNOMEDCT_CORE|Haemorrhage of large intestine with diverticular disease of large intestine|Hemorrhage of large intestine with diverticular disease of large intestine
C0581360|T047|SY|197092000|SNOMEDCT_CORE|Hemorrhage of large intestine co-occurrent and due to diverticular disease of large intestine|Hemorrhage of large intestine with diverticular disease of large intestine
C0581360|T047|FN|197092000|SNOMEDCT_CORE|Hemorrhage of large intestine co-occurrent and due to diverticular disease of large intestine|Hemorrhage of large intestine with diverticular disease of large intestine
C0581360|T047|PT|197092000|SNOMEDCT_CORE|Hemorrhage of large intestine with diverticular disease of large intestine|Hemorrhage of large intestine with diverticular disease of large intestine
C0581362|T184|PT|197232005|SNOMEDCT_CORE|Anorectal pain|Anorectal pain
C0581362|T184|FN|197232005|SNOMEDCT_CORE|Anorectal pain|Anorectal pain
C0581366|T047|PT|197853008|SNOMEDCT_CORE|Recurrent cystitis|Recurrent cystitis
C0581366|T047|FN|197853008|SNOMEDCT_CORE|Recurrent cystitis|Recurrent cystitis
C0581384|T047|PTGB|191268006|SNOMEDCT_CORE|Chronic anaemia|Chronic anemia
C0581384|T047|PT|191268006|SNOMEDCT_CORE|Chronic anemia|Chronic anemia
C0581384|T047|FN|191268006|SNOMEDCT_CORE|Chronic anemia|Chronic anemia
C0581386|T048|PT|191708009|SNOMEDCT_CORE|Chronic anxiety|Chronic anxiety
C0581386|T048|FN|191708009|SNOMEDCT_CORE|Chronic anxiety|Chronic anxiety
C0581394|T046|OAP|275319005|SNOMEDCT_CORE|Swollen legs|Swollen legs
C0581394|T046|OAF|275319005|SNOMEDCT_CORE|Swollen legs|Swollen legs
C0581839|T033|OP|162596006|SNOMEDCT_CORE|Suspected child abuse|Suspected victim of child abuse
C0581839|T033|OF|162596006|SNOMEDCT_CORE|Suspected child abuse|Suspected victim of child abuse
C0581839|T033|PT|162596006|SNOMEDCT_CORE|Suspected victim of child abuse|Suspected victim of child abuse
C0581839|T033|FN|162596006|SNOMEDCT_CORE|Suspected victim of child abuse|Suspected victim of child abuse
C0581869|T184|PT|162042000|SNOMEDCT_CORE|Abdominal wall pain|Abdominal wall pain
C0581869|T184|FN|162042000|SNOMEDCT_CORE|Abdominal wall pain|Abdominal wall pain
C0581896|T033|OAP|160830003|SNOMEDCT_CORE|Child relationship problem|Child relationship problem
C0581896|T033|OAF|160830003|SNOMEDCT_CORE|Child relationship problem|Child relationship problem
C0582114|T033|SY|304253006|SNOMEDCT_CORE|DNAR - Do not attempt resuscitation|Not for resuscitation
C0582114|T033|SY|304253006|SNOMEDCT_CORE|DNR|Not for resuscitation
C0582114|T033|SY|304253006|SNOMEDCT_CORE|Do not resuscitate|Not for resuscitation
C0582114|T033|SY|304253006|SNOMEDCT_CORE|Do not resuscitate status|Not for resuscitation
C0582114|T033|IS|304253006|SNOMEDCT_CORE|Not for attempted cardiopulmonary resuscitation|Not for resuscitation
C0582114|T033|PT|304253006|SNOMEDCT_CORE|Not for resuscitation|Not for resuscitation
C0582114|T033|FN|304253006|SNOMEDCT_CORE|Not for resuscitation|Not for resuscitation
C0582147|T033|PT|78648007|SNOMEDCT_CORE|At risk for infection|At risk for infection
C0582147|T033|FN|78648007|SNOMEDCT_CORE|At risk for infection|At risk for infection
C0582147|T033|IS|78648007|SNOMEDCT_CORE|At risk of infection|At risk for infection
C0582147|T033|OF|78648007|SNOMEDCT_CORE|At risk of infection|At risk for infection
C0582147|T033|SY|78648007|SNOMEDCT_CORE|Potential for infection|At risk for infection
C0582208|T033|PT|304321000|SNOMEDCT_CORE|Decreased range of knee movement|Decreased range of knee movement
C0582208|T033|FN|304321000|SNOMEDCT_CORE|Decreased range of knee movement|Decreased range of knee movement
C0582229|T033|PT|304344002|SNOMEDCT_CORE|Decreased range of cervical spine movement|Decreased range of cervical spine movement
C0582229|T033|FN|304344002|SNOMEDCT_CORE|Decreased range of cervical spine movement|Decreased range of cervical spine movement
C0582415|T047|PT|304527002|SNOMEDCT_CORE|Acute asthma|Acute asthma
C0582415|T047|FN|304527002|SNOMEDCT_CORE|Acute asthma|Acute asthma
C0582730|T037|PTGB|304831001|SNOMEDCT_CORE|Chronic intracranial subdural haematoma|Chronic intracranial subdural hematoma
C0582730|T037|PT|304831001|SNOMEDCT_CORE|Chronic intracranial subdural hematoma|Chronic intracranial subdural hematoma
C0582730|T037|FN|304831001|SNOMEDCT_CORE|Chronic intracranial subdural hematoma|Chronic intracranial subdural hematoma
C0583542|T033|PTGB|305647009|SNOMEDCT_CORE|Seen by paediatrician|Seen by pediatrician
C0583542|T033|PT|305647009|SNOMEDCT_CORE|Seen by pediatrician|Seen by pediatrician
C0583542|T033|FN|305647009|SNOMEDCT_CORE|Seen by pediatrician|Seen by pediatrician
C0584960|T047|SY|307091009|SNOMEDCT_CORE|Factor 5 Leiden mutation|Factor V Leiden mutation
C0584960|T047|PT|307091009|SNOMEDCT_CORE|Factor V Leiden mutation|Factor V Leiden mutation
C0584960|T047|FN|307091009|SNOMEDCT_CORE|Factor V Leiden mutation|Factor V Leiden mutation
C0584983|T047|PT|307115002|SNOMEDCT_CORE|Homozygous Factor V Leiden mutation|Homozygous Factor V Leiden mutation
C0584983|T047|FN|307115002|SNOMEDCT_CORE|Homozygous Factor V Leiden mutation|Homozygous Factor V Leiden mutation
C0584984|T047|PT|307116001|SNOMEDCT_CORE|Heterozygous Factor V Leiden mutation|Heterozygous Factor V Leiden mutation
C0584984|T047|FN|307116001|SNOMEDCT_CORE|Heterozygous Factor V Leiden mutation|Heterozygous Factor V Leiden mutation
C0585008|T047|PT|123608004|SNOMEDCT_CORE|Cholangiectasis|Cholangiectasis
C0585008|T047|FN|123608004|SNOMEDCT_CORE|Cholangiectasis|Cholangiectasis
C0585008|T047|SY|123608004|SNOMEDCT_CORE|Dilation of biliary tract|Cholangiectasis
C0585013|T033|PT|307136000|SNOMEDCT_CORE|Old healed fracture of bone|Old healed fracture of bone
C0585013|T033|OF|307136000|SNOMEDCT_CORE|Old healed fracture of bone|Old healed fracture of bone
C0585013|T033|FN|307136000|SNOMEDCT_CORE|Old healed fracture of bone|Old healed fracture of bone
C0585015|T190|PT|307138004|SNOMEDCT_CORE|Spondylolisthesis L5/S1 level|Spondylolisthesis L5/S1 level
C0585015|T190|FN|307138004|SNOMEDCT_CORE|Spondylolisthesis L5/S1 level|Spondylolisthesis L5/S1 level
C0585017|T047|PT|307140009|SNOMEDCT_CORE|Acute non-Q wave infarction|Acute non-Q wave infarction
C0585017|T047|FN|307140009|SNOMEDCT_CORE|Acute non-Q wave infarction|Acute non-Q wave infarction
C0585104|T047|SY|301000005|SNOMEDCT_CORE|Left basal pneumonia|Left lower zone pneumonia
C0585104|T047|SY|301000005|SNOMEDCT_CORE|Left lower lobe pneumonia|Left lower zone pneumonia
C0585104|T047|PT|301000005|SNOMEDCT_CORE|Left lower zone pneumonia|Left lower zone pneumonia
C0585104|T047|FN|301000005|SNOMEDCT_CORE|Left lower zone pneumonia|Left lower zone pneumonia
C0585104|T047|SY|301000005|SNOMEDCT_CORE|LLL - Left lower lobe pneumonia|Left lower zone pneumonia
C0585104|T047|SY|301000005|SNOMEDCT_CORE|LLZ - Left lower zone pneumonia|Left lower zone pneumonia
C0585104|T047|SY|301000005|SNOMEDCT_CORE|Lobar pneumonia left lower lobe|Left lower zone pneumonia
C0585105|T047|SY|301001009|SNOMEDCT_CORE|Lobar pneumonia right lower lobe|Right lower zone pneumonia
C0585105|T047|SY|301001009|SNOMEDCT_CORE|Right basal pneumonia|Right lower zone pneumonia
C0585105|T047|SY|301001009|SNOMEDCT_CORE|Right lower lobe pneumonia|Right lower zone pneumonia
C0585105|T047|PT|301001009|SNOMEDCT_CORE|Right lower zone pneumonia|Right lower zone pneumonia
C0585105|T047|FN|301001009|SNOMEDCT_CORE|Right lower zone pneumonia|Right lower zone pneumonia
C0585105|T047|SY|301001009|SNOMEDCT_CORE|RLL - Right lower lobe pneumonia|Right lower zone pneumonia
C0585105|T047|SY|301001009|SNOMEDCT_CORE|RLZ - Right lower zone pneumonia|Right lower zone pneumonia
C0585142|T046|PT|307233002|SNOMEDCT_CORE|Bleeding gastric erosion|Bleeding gastric erosion
C0585142|T046|FN|307233002|SNOMEDCT_CORE|Bleeding gastric erosion|Bleeding gastric erosion
C0585362|T191|PT|307502000|SNOMEDCT_CORE|Squamous cell carcinoma of mouth|Squamous cell carcinoma of mouth
C0585362|T191|FN|307502000|SNOMEDCT_CORE|Squamous cell carcinoma of mouth|Squamous cell carcinoma of mouth
C0585442|T191|PT|307576001|SNOMEDCT_CORE|Osteosarcoma of bone|Osteosarcoma of bone
C0585442|T191|FN|307576001|SNOMEDCT_CORE|Osteosarcoma of bone|Osteosarcoma of bone
C0585474|T191|SY|307608006|SNOMEDCT_CORE|Ewing sarcoma of bone|Ewing's sarcoma of bone
C0585474|T191|PT|307608006|SNOMEDCT_CORE|Ewing's sarcoma of bone|Ewing's sarcoma of bone
C0585474|T191|FN|307608006|SNOMEDCT_CORE|Ewing's sarcoma of bone|Ewing's sarcoma of bone
C0585625|T047|PT|307759003|SNOMEDCT_CORE|Helicobacter pylori gastrointestinal tract infection|Helicobacter pylori gastrointestinal tract infection
C0585625|T047|FN|307759003|SNOMEDCT_CORE|Helicobacter pylori gastrointestinal tract infection|Helicobacter pylori gastrointestinal tract infection
C0585894|T033|PTGB|308068007|SNOMEDCT_CORE|H/O: Treatment for ischaemic heart disease|H/O: Treatment for ischemic heart disease
C0585894|T033|PT|308068007|SNOMEDCT_CORE|H/O: Treatment for ischemic heart disease|H/O: Treatment for ischemic heart disease
C0585894|T033|IS|308068007|SNOMEDCT_CORE|History of - Treatment for ischaemic heart disease|H/O: Treatment for ischemic heart disease
C0585894|T033|OF|308068007|SNOMEDCT_CORE|History of - Treatment for ischemic heart disease|H/O: Treatment for ischemic heart disease
C0585894|T033|IS|308068007|SNOMEDCT_CORE|History of - Treatment for ischemic heart disease|H/O: Treatment for ischemic heart disease
C0585894|T033|SYGB|308068007|SNOMEDCT_CORE|History of treatment for ischaemic heart disease|H/O: Treatment for ischemic heart disease
C0585894|T033|FN|308068007|SNOMEDCT_CORE|History of treatment for ischemic heart disease|H/O: Treatment for ischemic heart disease
C0585894|T033|SY|308068007|SNOMEDCT_CORE|History of treatment for ischemic heart disease|H/O: Treatment for ischemic heart disease
C0585952|T047|PT|308129003|SNOMEDCT_CORE|Esophageal varices in cirrhosis of the liver|Esophageal varices in cirrhosis of the liver
C0585952|T047|FN|308129003|SNOMEDCT_CORE|Esophageal varices in cirrhosis of the liver|Esophageal varices in cirrhosis of the liver
C0585952|T047|PTGB|308129003|SNOMEDCT_CORE|Oesophageal varices in cirrhosis of the liver|Esophageal varices in cirrhosis of the liver
C0585965|T037|PT|308153009|SNOMEDCT_CORE|Closed fracture of distal fibula|Closed fracture of distal fibula
C0585965|T037|FN|308153009|SNOMEDCT_CORE|Closed fracture of distal fibula|Closed fracture of distal fibula
C0586285|T033|FN|308684007|SNOMEDCT_CORE|Amputated big toe|Amputated big toe
C0586285|T033|PT|308684007|SNOMEDCT_CORE|Amputated big toe|Amputated big toe
C0586316|T033|OAP|308728002|SNOMEDCT_CORE|Cervical smear biopsy taken|Sampling of cervix for Papanicolaou smear done
C0586316|T033|IS|767357000|SNOMEDCT_CORE|Cervical smear biopsy taken|Sampling of cervix for Papanicolaou smear done
C0586316|T033|OAF|308728002|SNOMEDCT_CORE|Cervical smear biopsy taken|Sampling of cervix for Papanicolaou smear done
C0586316|T033|OAS|308728002|SNOMEDCT_CORE|Cervical smear taken|Sampling of cervix for Papanicolaou smear done
C0586316|T033|OAS|308728002|SNOMEDCT_CORE|Papanicolaou smear taken|Sampling of cervix for Papanicolaou smear done
C0586316|T033|SY|767357000|SNOMEDCT_CORE|Papanicolaou smear taken|Sampling of cervix for Papanicolaou smear done
C0586316|T033|PT|767357000|SNOMEDCT_CORE|Sampling of cervix for Papanicolaou smear done|Sampling of cervix for Papanicolaou smear done
C0586316|T033|FN|767357000|SNOMEDCT_CORE|Sampling of cervix for Papanicolaou smear done|Sampling of cervix for Papanicolaou smear done
C0586316|T033|OAS|308728002|SNOMEDCT_CORE|Smear - cervical:taken|Sampling of cervix for Papanicolaou smear done
C0586384|T046|PTGB|308896002|SNOMEDCT_CORE|Secondary haemorrhage postprocedure|Secondary hemorrhage postprocedure
C0586384|T046|PT|308896002|SNOMEDCT_CORE|Secondary hemorrhage postprocedure|Secondary hemorrhage postprocedure
C0586384|T046|FN|308896002|SNOMEDCT_CORE|Secondary hemorrhage postprocedure|Secondary hemorrhage postprocedure
C0586387|T033|SY|308899009|SNOMEDCT_CORE|Unfavorable living conditions|Unsatisfactory living conditions
C0586387|T033|SYGB|308899009|SNOMEDCT_CORE|Unfavourable living conditions|Unsatisfactory living conditions
C0586387|T033|PT|308899009|SNOMEDCT_CORE|Unsatisfactory living conditions|Unsatisfactory living conditions
C0586387|T033|FN|308899009|SNOMEDCT_CORE|Unsatisfactory living conditions|Unsatisfactory living conditions
C0586553|T033|OAF|131016008|SNOMEDCT_CORE|Increased thyroid stimulating hormone level|Raised TSH level
C0586553|T033|OAP|131016008|SNOMEDCT_CORE|Increased thyroid stimulating hormone level|Raised TSH level
C0586553|T033|FN|309080005|SNOMEDCT_CORE|Raised thyroid stimulating hormone level|Raised TSH level
C0586553|T033|SY|309080005|SNOMEDCT_CORE|Raised thyroid stimulating hormone level|Raised TSH level
C0586553|T033|PT|309080005|SNOMEDCT_CORE|Raised TSH level|Raised TSH level
C0586553|T033|OF|309080005|SNOMEDCT_CORE|Raised TSH level|Raised TSH level
C0586556|T047|PT|309083007|SNOMEDCT_CORE|Abscess of back|Abscess of back
C0586556|T047|FN|309083007|SNOMEDCT_CORE|Abscess of back|Abscess of back
C0586557|T037|SY|17542004|SNOMEDCT_CORE|Accident at work|Accident while engaged in work-related activity
C0586557|T037|IS|17542004|SNOMEDCT_CORE|Accident at work, NOS|Accident while engaged in work-related activity
C0586557|T037|PT|17542004|SNOMEDCT_CORE|Accident while engaged in work-related activity|Accident while engaged in work-related activity
C0586557|T037|OF|17542004|SNOMEDCT_CORE|Accident while engaged in work-related activity|Accident while engaged in work-related activity
C0586557|T037|FN|17542004|SNOMEDCT_CORE|Accident while engaged in work-related activity|Accident while engaged in work-related activity
C0586557|T037|IS|17542004|SNOMEDCT_CORE|Accident while engaged in work-related activity, NOS|Accident while engaged in work-related activity
C0586557|T037|PTGB|17542004|SNOMEDCT_CORE|Accident whilst engaged in work-related activity|Accident while engaged in work-related activity
C0586557|T037|SY|17542004|SNOMEDCT_CORE|Work accident|Accident while engaged in work-related activity
C0586559|T033|PT|309089006|SNOMEDCT_CORE|Prostate mass|Prostate mass
C0586559|T033|FN|309089006|SNOMEDCT_CORE|Prostate mass|Prostate mass
C0586735|T047|SY|309246000|SNOMEDCT_CORE|Degenerative joint disease of foot|Osteoarthritis of foot joint
C0586735|T047|PT|309246000|SNOMEDCT_CORE|Osteoarthritis of foot joint|Osteoarthritis of foot joint
C0586735|T047|FN|309246000|SNOMEDCT_CORE|Osteoarthritis of foot joint|Osteoarthritis of foot joint
C0586979|T033|OF|160297008|SNOMEDCT_CORE|Family history: neoplasm of ovary|FH: neoplasm of ovary
C0586979|T033|FN|160297008|SNOMEDCT_CORE|Family history: neoplasm of ovary|FH: neoplasm of ovary
C0586979|T033|SY|160297008|SNOMEDCT_CORE|Family history: neoplasm of ovary|FH: neoplasm of ovary
C0586979|T033|PT|160297008|SNOMEDCT_CORE|FH: neoplasm of ovary|FH: neoplasm of ovary
C0586989|T047|PT|309465005|SNOMEDCT_CORE|Varicella-zoster virus infection|Varicella-zoster virus infection
C0586989|T047|FN|309465005|SNOMEDCT_CORE|Varicella-zoster virus infection|Varicella-zoster virus infection
C0587046|T033|SY|309523001|SNOMEDCT_CORE|Artificial lens in situ|Artificial lens present
C0587046|T033|PT|309523001|SNOMEDCT_CORE|Artificial lens present|Artificial lens present
C0587046|T033|FN|309523001|SNOMEDCT_CORE|Artificial lens present|Artificial lens present
C0587050|T184|PT|309527000|SNOMEDCT_CORE|Mass of lower limb|Mass of lower limb
C0587050|T184|FN|309527000|SNOMEDCT_CORE|Mass of lower limb|Mass of lower limb
C0587055|T184|PT|309537005|SNOMEDCT_CORE|Numbness of lower limb|Numbness of lower limb
C0587055|T184|FN|309537005|SNOMEDCT_CORE|Numbness of lower limb|Numbness of lower limb
C0587060|T191|PT|269578002|SNOMEDCT_CORE|Malignant melanoma of head and neck|Malignant melanoma of head and neck
C0587060|T191|FN|269578002|SNOMEDCT_CORE|Malignant melanoma of head and neck|Malignant melanoma of head and neck
C0587062|T191|PT|269581007|SNOMEDCT_CORE|Malignant melanoma of lower limb|Malignant melanoma of lower limb
C0587062|T191|FN|269581007|SNOMEDCT_CORE|Malignant melanoma of lower limb|Malignant melanoma of lower limb
C0587094|T033|SY|309587003|SNOMEDCT_CORE|Breast calcification|Calcification of breast
C0587094|T033|PT|309587003|SNOMEDCT_CORE|Calcification of breast|Calcification of breast
C0587094|T033|FN|309587003|SNOMEDCT_CORE|Calcification of breast|Calcification of breast
C0587170|T033|SY|105531004|SNOMEDCT_CORE|Accommodation unsuitable|Housing problem
C0587170|T033|PT|105531004|SNOMEDCT_CORE|Housing problem|Housing problem
C0587170|T033|SY|105531004|SNOMEDCT_CORE|Housing unsatisfactory|Housing problem
C0587170|T033|FN|105531004|SNOMEDCT_CORE|Housing unsatisfactory|Housing problem
C0587170|T033|SY|105531004|SNOMEDCT_CORE|Inadequate housing|Housing problem
C0587170|T033|IS|105531004|SNOMEDCT_CORE|Living in unsatisfactory surroundings|Housing problem
C0587223|T184|PT|309737007|SNOMEDCT_CORE|Abdominal pain in pregnancy|Abdominal pain in pregnancy
C0587223|T184|FN|309737007|SNOMEDCT_CORE|Abdominal pain in pregnancy|Abdominal pain in pregnancy
C0587229|T047|PTGB|309745002|SNOMEDCT_CORE|Osteoporosis localised to spine|Osteoporosis localized to spine
C0587229|T047|PT|309745002|SNOMEDCT_CORE|Osteoporosis localized to spine|Osteoporosis localized to spine
C0587229|T047|FN|309745002|SNOMEDCT_CORE|Osteoporosis localized to spine|Osteoporosis localized to spine
C0587246|T033|IS|309774006|SNOMEDCT_CORE|Loss of power in limb|Muscle weakness of limb
C0587246|T033|SY|713514005|SNOMEDCT_CORE|Loss of power in limb|Muscle weakness of limb
C0587246|T033|PT|713514005|SNOMEDCT_CORE|Muscle weakness of limb|Muscle weakness of limb
C0587246|T033|FN|713514005|SNOMEDCT_CORE|Muscle weakness of limb|Muscle weakness of limb
C0587246|T033|OAP|309774006|SNOMEDCT_CORE|Weakness of limb|Muscle weakness of limb
C0587246|T033|OAF|309774006|SNOMEDCT_CORE|Weakness of limb|Muscle weakness of limb
C0587955|T033|PT|310439007|SNOMEDCT_CORE|Urine cytology abnormal|Urine cytology abnormal
C0587955|T033|FN|310439007|SNOMEDCT_CORE|Urine cytology abnormal|Urine cytology abnormal
C0588006|T048|PT|310495003|SNOMEDCT_CORE|Mild depression|Mild depression
C0588006|T048|FN|310495003|SNOMEDCT_CORE|Mild depression|Mild depression
C0588007|T048|PT|310496002|SNOMEDCT_CORE|Moderate depression|Moderate depression
C0588007|T048|FN|310496002|SNOMEDCT_CORE|Moderate depression|Moderate depression
C0588173|T047|PT|310643001|SNOMEDCT_CORE|Infection of intravenous catheter|Infection of intravenous catheter
C0588173|T047|FN|310643001|SNOMEDCT_CORE|Infection of intravenous catheter|Infection of intravenous catheter
C0588179|T047|PTGB|310647000|SNOMEDCT_CORE|Anaemia secondary to renal failure|Anemia secondary to renal failure
C0588179|T047|PT|310647000|SNOMEDCT_CORE|Anemia secondary to renal failure|Anemia secondary to renal failure
C0588179|T047|FN|310647000|SNOMEDCT_CORE|Anemia secondary to renal failure|Anemia secondary to renal failure
C0589110|T047|PT|213220000|SNOMEDCT_CORE|Postoperative deep vein thrombosis|Postoperative deep vein thrombosis
C0589110|T047|FN|213220000|SNOMEDCT_CORE|Postoperative deep vein thrombosis|Postoperative deep vein thrombosis
C0589379|T020|PT|311806008|SNOMEDCT_CORE|Collapse of cervical vertebra due to osteoporosis|Collapse of cervical vertebra due to osteoporosis
C0589379|T020|FN|311806008|SNOMEDCT_CORE|Collapse of cervical vertebra due to osteoporosis|Collapse of cervical vertebra due to osteoporosis
C0589630|T047|PT|312110005|SNOMEDCT_CORE|Gallbladder and bile duct calculi|Gallbladder and bile duct calculi
C0589630|T047|FN|312110005|SNOMEDCT_CORE|Gallbladder and bile duct calculi|Gallbladder and bile duct calculi
C0589630|T047|SY|312110005|SNOMEDCT_CORE|Gallbladder and bile duct stones|Gallbladder and bile duct calculi
C0595861|T048|OAP|48981002|SNOMEDCT_CORE|Parasuicide|Suicide attempt by inadequate means
C0595861|T048|SY|55554002|SNOMEDCT_CORE|Parasuicide|Suicide attempt by inadequate means
C0595861|T048|OF|48981002|SNOMEDCT_CORE|Parasuicide|Suicide attempt by inadequate means
C0595861|T048|OAF|48981002|SNOMEDCT_CORE|Parasuicide|Suicide attempt by inadequate means
C0595861|T048|PT|55554002|SNOMEDCT_CORE|Suicide attempt by inadequate means|Suicide attempt by inadequate means
C0595861|T048|OF|55554002|SNOMEDCT_CORE|Suicide attempt by inadequate means|Suicide attempt by inadequate means
C0595861|T048|FN|55554002|SNOMEDCT_CORE|Suicide attempt by inadequate means|Suicide attempt by inadequate means
C0595861|T048|SY|55554002|SNOMEDCT_CORE|Suicide gesture|Suicide attempt by inadequate means
C0595861|T048|SY|55554002|SNOMEDCT_CORE|Unsuccessful suicide attempt|Suicide attempt by inadequate means
C0595929|T033|PT|166830008|SNOMEDCT_CORE|Serum cholesterol raised|Serum cholesterol raised
C0595929|T033|FN|166830008|SNOMEDCT_CORE|Serum cholesterol raised|Serum cholesterol raised
C0595948|T047|PT|23374007|SNOMEDCT_CORE|Atypical absence seizure|Atypical absence seizure
C0595948|T047|FN|23374007|SNOMEDCT_CORE|Atypical absence seizure|Atypical absence seizure
C0595948|T047|IS|23374007|SNOMEDCT_CORE|Atypical absence seizures|Atypical absence seizure
C0595989|T191|PT|276975007|SNOMEDCT_CORE|Carcinoma of larynx|Carcinoma of larynx
C0595989|T191|FN|276975007|SNOMEDCT_CORE|Carcinoma of larynx|Carcinoma of larynx
C0595989|T191|SY|276975007|SNOMEDCT_CORE|Laryngeal carcinoma|Carcinoma of larynx
C0595995|T020|PT|203639008|SNOMEDCT_CORE|Idiopathic scoliosis|Idiopathic scoliosis
C0595995|T020|FN|203639008|SNOMEDCT_CORE|Idiopathic scoliosis|Idiopathic scoliosis
C0597984|T190|PT|235921003|SNOMEDCT_CORE|Biliary stricture|Biliary stricture
C0597984|T190|FN|235921003|SNOMEDCT_CORE|Biliary stricture|Biliary stricture
C0598608|T047|PT|419503008|SNOMEDCT_CORE|Hyperhomocysteinemia|Hyperhomocysteinemia
C0598608|T047|FN|419503008|SNOMEDCT_CORE|Hyperhomocysteinemia|Hyperhomocysteinemia
C0598798|T191|PT|414628006|SNOMEDCT_CORE|Lymphoid neoplasm|Lymphoid neoplasm
C0598798|T191|FN|414628006|SNOMEDCT_CORE|Lymphoid neoplasm|Lymphoid neoplasm
C0600040|T047|PT|197834003|SNOMEDCT_CORE|Chronic interstitial cystitis|Chronic interstitial cystitis
C0600040|T047|FN|197834003|SNOMEDCT_CORE|Chronic interstitial cystitis|Chronic interstitial cystitis
C0600040|T047|SY|197834003|SNOMEDCT_CORE|Painful bladder syndrome|Chronic interstitial cystitis
C0600040|T047|SY|197834003|SNOMEDCT_CORE|PBS - Painful bladder syndrome|Chronic interstitial cystitis
C0600106|T037|PT|309464009|SNOMEDCT_CORE|Elbow fracture|Elbow fracture
C0600106|T037|FN|309464009|SNOMEDCT_CORE|Elbow fracture|Elbow fracture
C0600106|T037|SY|309464009|SNOMEDCT_CORE|Fracture of elbow|Elbow fracture
C0600139|T191|SY|254900004|SNOMEDCT_CORE|CA - Carcinoma of prostate|Carcinoma of prostate
C0600139|T191|PT|254900004|SNOMEDCT_CORE|Carcinoma of prostate|Carcinoma of prostate
C0600139|T191|FN|254900004|SNOMEDCT_CORE|Carcinoma of prostate|Carcinoma of prostate
C0600139|T191|SY|254900004|SNOMEDCT_CORE|Prostate cancer|Carcinoma of prostate
C0600139|T191|SY|254900004|SNOMEDCT_CORE|Prostate carcinoma|Carcinoma of prostate
C0600142|T184|SY|198436008|SNOMEDCT_CORE|Hot flashes|Menopausal flushing
C0600142|T184|SY|198436008|SNOMEDCT_CORE|Hot flush|Menopausal flushing
C0600142|T184|SY|198436008|SNOMEDCT_CORE|Hot flushes|Menopausal flushing
C0600142|T184|PT|198436008|SNOMEDCT_CORE|Menopausal flushing|Menopausal flushing
C0600142|T184|FN|198436008|SNOMEDCT_CORE|Menopausal flushing|Menopausal flushing
C0600142|T184|SY|198436008|SNOMEDCT_CORE|Menopausal hot flashes|Menopausal flushing
C0600142|T184|SY|198436008|SNOMEDCT_CORE|Menopausal hot flushes|Menopausal flushing
C0600359|T047|SY|56267009|SNOMEDCT_CORE|Arteriosclerotic dementia|Arteriosclerotic dementia
C0600427|T048|PT|31956009|SNOMEDCT_CORE|Cocaine dependence|Cocaine dependence
C0600427|T048|FN|31956009|SNOMEDCT_CORE|Cocaine dependence|Cocaine dependence
C0677061|T184|PT|267981009|SNOMEDCT_CORE|Pain in thoracic spine|Pain in thoracic spine
C0677061|T184|FN|267981009|SNOMEDCT_CORE|Pain in thoracic spine|Pain in thoracic spine
C0677607|T047|SY|21983002|SNOMEDCT_CORE|Autoimmune lymphocytic chronic thyroiditis|Hashimoto thyroiditis
C0677607|T047|SY|21983002|SNOMEDCT_CORE|Chronic lymphocytic thyroiditis|Hashimoto thyroiditis
C0677607|T047|PT|21983002|SNOMEDCT_CORE|Hashimoto thyroiditis|Hashimoto thyroiditis
C0677607|T047|FN|21983002|SNOMEDCT_CORE|Hashimoto thyroiditis|Hashimoto thyroiditis
C0677607|T047|SY|21983002|SNOMEDCT_CORE|Hashimoto's disease|Hashimoto thyroiditis
C0677607|T047|SY|21983002|SNOMEDCT_CORE|Hashimoto's thyroiditis|Hashimoto thyroiditis
C0677607|T047|SY|21983002|SNOMEDCT_CORE|Lymphocytic thyroiditis|Hashimoto thyroiditis
C0677607|T047|SY|21983002|SNOMEDCT_CORE|Struma lymphomatosa|Hashimoto thyroiditis
C0677607|T047|SY|21983002|SNOMEDCT_CORE|Struma lymphomatosis|Hashimoto thyroiditis
C0677628|T033|SY|247154004|SNOMEDCT_CORE|Drusen of macula|Macular drusen
C0677628|T033|PT|247154004|SNOMEDCT_CORE|Macular drusen|Macular drusen
C0677628|T033|FN|247154004|SNOMEDCT_CORE|Macular drusen|Macular drusen
C0677659|T047|SY|266433003|SNOMEDCT_CORE|Esophageal reflux with esophagitis|Gastro-esophageal reflux disease with esophagitis
C0677659|T047|PT|266433003|SNOMEDCT_CORE|Gastro-esophageal reflux disease with esophagitis|Gastro-esophageal reflux disease with esophagitis
C0677659|T047|PTGB|266433003|SNOMEDCT_CORE|Gastro-oesophageal reflux disease with oesophagitis|Gastro-esophageal reflux disease with esophagitis
C0677659|T047|FN|266433003|SNOMEDCT_CORE|Gastroesophageal reflux disease with esophagitis|Gastro-esophageal reflux disease with esophagitis
C0677659|T047|SY|266433003|SNOMEDCT_CORE|Gastroesophageal reflux disease with esophagitis|Gastro-esophageal reflux disease with esophagitis
C0677659|T047|SYGB|266433003|SNOMEDCT_CORE|Gastroesophageal reflux disease with oesophagitis|Gastro-esophageal reflux disease with esophagitis
C0677659|T047|SYGB|266433003|SNOMEDCT_CORE|Oesophageal reflux with oesophagitis|Gastro-esophageal reflux disease with esophagitis
C0677659|T047|SY|266433003|SNOMEDCT_CORE|Peptic esophagitis|Gastro-esophageal reflux disease with esophagitis
C0677659|T047|SYGB|266433003|SNOMEDCT_CORE|Peptic oesophagitis|Gastro-esophageal reflux disease with esophagitis
C0677659|T047|SY|266433003|SNOMEDCT_CORE|Reflux esophagitis|Gastro-esophageal reflux disease with esophagitis
C0677659|T047|SYGB|266433003|SNOMEDCT_CORE|Reflux oesophagitis|Gastro-esophageal reflux disease with esophagitis
C0677865|T191|PT|444545003|SNOMEDCT_CORE|Glioma of brainstem|Glioma of brainstem
C0677865|T191|FN|444545003|SNOMEDCT_CORE|Glioma of brainstem|Glioma of brainstem
C0678127|T020|SY|201040000|SNOMEDCT_CORE|Tyloma|Tyloma
C0678189|T047|PTGB|267432004|SNOMEDCT_CORE|Pure hypercholesterolaemia|Pure hypercholesterolemia
C0678189|T047|PT|267432004|SNOMEDCT_CORE|Pure hypercholesterolemia|Pure hypercholesterolemia
C0678189|T047|FN|267432004|SNOMEDCT_CORE|Pure hypercholesterolemia|Pure hypercholesterolemia
C0678212|T037|PT|84857004|SNOMEDCT_CORE|Herniation of nucleus pulposus|Herniation of nucleus pulposus
C0678212|T037|FN|84857004|SNOMEDCT_CORE|Herniation of nucleus pulposus|Herniation of nucleus pulposus
C0678212|T037|IS|84857004|SNOMEDCT_CORE|Herniation of nucleus pulposus, NOS|Herniation of nucleus pulposus
C0678222|T191|SY|254838004|SNOMEDCT_CORE|CA - Carcinoma of breast|Carcinoma of breast
C0678222|T191|PT|254838004|SNOMEDCT_CORE|Carcinoma of breast|Carcinoma of breast
C0678222|T191|FN|254838004|SNOMEDCT_CORE|Carcinoma of breast|Carcinoma of breast
C0683369|T033|PT|40917007|SNOMEDCT_CORE|Clouded consciousness|Clouded consciousness
C0683369|T033|FN|40917007|SNOMEDCT_CORE|Clouded consciousness|Clouded consciousness
C0683369|T033|IS|40917007|SNOMEDCT_CORE|Clouding of consciousness|Clouded consciousness
C0683369|T033|SY|40917007|SNOMEDCT_CORE|Confused|Clouded consciousness
C0683369|T033|SY|40917007|SNOMEDCT_CORE|Confusion|Clouded consciousness
C0683369|T033|SY|40917007|SNOMEDCT_CORE|Dazed|Clouded consciousness
C0683369|T033|SY|40917007|SNOMEDCT_CORE|Dazed state|Clouded consciousness
C0683369|T033|SY|40917007|SNOMEDCT_CORE|Dullness of senses|Clouded consciousness
C0683369|T033|SY|40917007|SNOMEDCT_CORE|Foggy mind|Clouded consciousness
C0683369|T033|SY|40917007|SNOMEDCT_CORE|Muddled|Clouded consciousness
C0683369|T033|IS|40917007|SNOMEDCT_CORE|Muzzy headed|Clouded consciousness
C0683369|T033|OP|40917007|SNOMEDCT_CORE|Wooziness|Clouded consciousness
C0683405|T048|SY|425919003|SNOMEDCT_CORE|Chronic organic brain syndrome|Chronic organic mental disorder
C0683405|T048|PT|425919003|SNOMEDCT_CORE|Chronic organic mental disorder|Chronic organic mental disorder
C0683405|T048|FN|425919003|SNOMEDCT_CORE|Chronic organic mental disorder|Chronic organic mental disorder
C0684343|T033|PT|95217000|SNOMEDCT_CORE|Pseudophakia|Pseudophakia
C0684343|T033|FN|95217000|SNOMEDCT_CORE|Pseudophakia|Pseudophakia
C0684364|T191|PT|94022001|SNOMEDCT_CORE|Primary malignant neoplasm of skin of face|Primary malignant neoplasm of skin of face
C0684364|T191|FN|94022001|SNOMEDCT_CORE|Primary malignant neoplasm of skin of face|Primary malignant neoplasm of skin of face
C0684386|T191|IS|94038007|SNOMEDCT_CORE|Malignant neoplasm of skin of scalp|Primary malignant neoplasm of skin of scalp
C0684386|T191|PT|94038007|SNOMEDCT_CORE|Primary malignant neoplasm of skin of scalp|Primary malignant neoplasm of skin of scalp
C0684386|T191|FN|94038007|SNOMEDCT_CORE|Primary malignant neoplasm of skin of scalp|Primary malignant neoplasm of skin of scalp
C0684487|T191|PT|93225001|SNOMEDCT_CORE|Malignant melanoma of skin of face|Malignant melanoma of skin of face
C0684487|T191|FN|93225001|SNOMEDCT_CORE|Malignant melanoma of skin of face|Malignant melanoma of skin of face
C0684487|T191|IS|93225001|SNOMEDCT_CORE|Malignant melanoma of skin of face, NOS|Malignant melanoma of skin of face
C0684498|T191|PT|93651008|SNOMEDCT_CORE|Malignant melanoma of skin of trunk|Malignant melanoma of skin of trunk
C0684498|T191|FN|93651008|SNOMEDCT_CORE|Malignant melanoma of skin of trunk|Malignant melanoma of skin of trunk
C0684498|T191|IS|93651008|SNOMEDCT_CORE|Malignant melanoma of skin of trunk, NOS|Malignant melanoma of skin of trunk
C0684550|T191|SY|94602001|SNOMEDCT_CORE|CA - Secondary cancer of spine|Secondary malignant neoplasm of vertebral column
C0684550|T191|SY|94602001|SNOMEDCT_CORE|Metastasis to spine|Secondary malignant neoplasm of vertebral column
C0684550|T191|SY|94602001|SNOMEDCT_CORE|Metastasis to vertebral column|Secondary malignant neoplasm of vertebral column
C0684550|T191|SY|94602001|SNOMEDCT_CORE|Metastatic malignant neoplasm to spine|Secondary malignant neoplasm of vertebral column
C0684550|T191|IS|94602001|SNOMEDCT_CORE|Metastatic malignant neoplasm to spine, NOS|Secondary malignant neoplasm of vertebral column
C0684550|T191|SY|94602001|SNOMEDCT_CORE|Metastatic malignant neoplasm to vertebral column|Secondary malignant neoplasm of vertebral column
C0684550|T191|IS|94602001|SNOMEDCT_CORE|Metastatic malignant neoplasm to vertebral column, NOS|Secondary malignant neoplasm of vertebral column
C0684550|T191|SY|94602001|SNOMEDCT_CORE|Secondary cancer of spine|Secondary malignant neoplasm of vertebral column
C0684550|T191|SY|94602001|SNOMEDCT_CORE|Secondary malignant neoplasm of spine|Secondary malignant neoplasm of vertebral column
C0684550|T191|IS|94602001|SNOMEDCT_CORE|Secondary malignant neoplasm of spine, NOS|Secondary malignant neoplasm of vertebral column
C0684550|T191|PT|94602001|SNOMEDCT_CORE|Secondary malignant neoplasm of vertebral column|Secondary malignant neoplasm of vertebral column
C0684550|T191|FN|94602001|SNOMEDCT_CORE|Secondary malignant neoplasm of vertebral column|Secondary malignant neoplasm of vertebral column
C0684550|T191|IS|94602001|SNOMEDCT_CORE|Secondary malignant neoplasm of vertebral column, NOS|Secondary malignant neoplasm of vertebral column
C0684550|T191|SY|94602001|SNOMEDCT_CORE|Secondary tumor of spine|Secondary malignant neoplasm of vertebral column
C0684550|T191|SYGB|94602001|SNOMEDCT_CORE|Secondary tumour of spine|Secondary malignant neoplasm of vertebral column
C0684550|T191|SY|94602001|SNOMEDCT_CORE|Spinal metastases|Secondary malignant neoplasm of vertebral column
C0684686|T191|SY|94264008|SNOMEDCT_CORE|Metastasis to soft tissue|Secondary malignant neoplasm of soft tissues
C0684686|T191|SY|94264008|SNOMEDCT_CORE|Metastatic malignant neoplasm to connective and other soft tissues|Secondary malignant neoplasm of soft tissues
C0684686|T191|IS|94264008|SNOMEDCT_CORE|Metastatic malignant neoplasm to connective and other soft tissues, NOS|Secondary malignant neoplasm of soft tissues
C0684686|T191|SY|94264008|SNOMEDCT_CORE|Secondary malignant neoplasm of connective and other soft tissues|Secondary malignant neoplasm of soft tissues
C0684686|T191|IS|94264008|SNOMEDCT_CORE|Secondary malignant neoplasm of connective and other soft tissues, NOS|Secondary malignant neoplasm of soft tissues
C0684686|T191|PT|94264008|SNOMEDCT_CORE|Secondary malignant neoplasm of soft tissues|Secondary malignant neoplasm of soft tissues
C0684686|T191|FN|94264008|SNOMEDCT_CORE|Secondary malignant neoplasm of soft tissues|Secondary malignant neoplasm of soft tissues
C0684699|T191|PT|92401003|SNOMEDCT_CORE|Benign neoplasm of soft tissues of upper limb|Benign neoplasm of soft tissues of upper limb
C0684699|T191|FN|92401003|SNOMEDCT_CORE|Benign neoplasm of soft tissues of upper limb|Benign neoplasm of soft tissues of upper limb
C0684699|T191|SY|92401003|SNOMEDCT_CORE|Benign tumor of soft tissue of upper limb|Benign neoplasm of soft tissues of upper limb
C0684699|T191|SYGB|92401003|SNOMEDCT_CORE|Benign tumour of soft tissue of upper limb|Benign neoplasm of soft tissues of upper limb
C0684706|T191|PT|92394004|SNOMEDCT_CORE|Benign neoplasm of soft tissues of lower limb|Benign neoplasm of soft tissues of lower limb
C0684706|T191|FN|92394004|SNOMEDCT_CORE|Benign neoplasm of soft tissues of lower limb|Benign neoplasm of soft tissues of lower limb
C0684706|T191|SY|92394004|SNOMEDCT_CORE|Benign tumor of soft tissue of leg|Benign neoplasm of soft tissues of lower limb
C0684706|T191|SY|92394004|SNOMEDCT_CORE|Benign tumor of soft tissue of lower limb|Benign neoplasm of soft tissues of lower limb
C0684706|T191|SYGB|92394004|SNOMEDCT_CORE|Benign tumour of soft tissue of leg|Benign neoplasm of soft tissues of lower limb
C0684706|T191|SYGB|92394004|SNOMEDCT_CORE|Benign tumour of soft tissue of lower limb|Benign neoplasm of soft tissues of lower limb
C0684708|T191|IS|94057003|SNOMEDCT_CORE|Malignant neoplasm of soft tissues of lower limb|Primary malignant neoplasm of soft tissues of lower limb
C0684708|T191|PT|94057003|SNOMEDCT_CORE|Primary malignant neoplasm of soft tissues of lower limb|Primary malignant neoplasm of soft tissues of lower limb
C0684708|T191|FN|94057003|SNOMEDCT_CORE|Primary malignant neoplasm of soft tissues of lower limb|Primary malignant neoplasm of soft tissues of lower limb
C0684808|T191|PT|363501002|SNOMEDCT_CORE|Malignant tumor of face|Malignant tumor of face
C0684808|T191|FN|363501002|SNOMEDCT_CORE|Malignant tumor of face|Malignant tumor of face
C0684808|T191|PTGB|363501002|SNOMEDCT_CORE|Malignant tumour of face|Malignant tumor of face
C0684816|T191|PT|94962000|SNOMEDCT_CORE|Neoplasm of uncertain behavior of neck|Neoplasm of uncertain behavior of neck
C0684816|T191|FN|94962000|SNOMEDCT_CORE|Neoplasm of uncertain behavior of neck|Neoplasm of uncertain behavior of neck
C0684816|T191|IS|94962000|SNOMEDCT_CORE|Neoplasm of uncertain behavior of neck, NOS|Neoplasm of uncertain behavior of neck
C0684816|T191|PTGB|94962000|SNOMEDCT_CORE|Neoplasm of uncertain behaviour of neck|Neoplasm of uncertain behavior of neck
C0684830|T191|SY|94180008|SNOMEDCT_CORE|Metastatic malignant neoplasm to axilla|Secondary malignant neoplasm of axilla
C0684830|T191|IS|94180008|SNOMEDCT_CORE|Metastatic malignant neoplasm to axilla, NOS|Secondary malignant neoplasm of axilla
C0684830|T191|PT|94180008|SNOMEDCT_CORE|Secondary malignant neoplasm of axilla|Secondary malignant neoplasm of axilla
C0684830|T191|FN|94180008|SNOMEDCT_CORE|Secondary malignant neoplasm of axilla|Secondary malignant neoplasm of axilla
C0684830|T191|IS|94180008|SNOMEDCT_CORE|Secondary malignant neoplasm of axilla, NOS|Secondary malignant neoplasm of axilla
C0685095|T047|PT|92506005|SNOMEDCT_CORE|Biventricular congestive heart failure|Biventricular congestive heart failure
C0685095|T047|FN|92506005|SNOMEDCT_CORE|Biventricular congestive heart failure|Biventricular congestive heart failure
C0685095|T047|SY|92506005|SNOMEDCT_CORE|Biventricular failure|Biventricular congestive heart failure
C0685707|T019|SY|94706008|SNOMEDCT_CORE|Muscular ventricular septal defect|Muscular ventricular septum defect
C0685707|T019|PT|94706008|SNOMEDCT_CORE|Muscular ventricular septum defect|Muscular ventricular septum defect
C0685707|T019|FN|94706008|SNOMEDCT_CORE|Muscular ventricular septum defect|Muscular ventricular septum defect
C0685925|T047|PT|91945006|SNOMEDCT_CORE|Articular disc disorder of temporomandibular joint|Articular disc disorder of temporomandibular joint
C0685925|T047|FN|91945006|SNOMEDCT_CORE|Articular disc disorder of temporomandibular joint|Articular disc disorder of temporomandibular joint
C0685938|T191|PT|428905002|SNOMEDCT_CORE|Malignant neoplasm of gastrointestinal tract|Malignant neoplasm of gastrointestinal tract
C0685938|T191|FN|428905002|SNOMEDCT_CORE|Malignant neoplasm of gastrointestinal tract|Malignant neoplasm of gastrointestinal tract
C0686055|T191|SY|94286009|SNOMEDCT_CORE|Cancer metastatic to esophagus|Secondary malignant neoplasm of esophagus
C0686055|T191|SY|94286009|SNOMEDCT_CORE|Metastatic malignant neoplasm to esophagus|Secondary malignant neoplasm of esophagus
C0686055|T191|IS|94286009|SNOMEDCT_CORE|Metastatic malignant neoplasm to esophagus, NOS|Secondary malignant neoplasm of esophagus
C0686055|T191|SYGB|94286009|SNOMEDCT_CORE|Metastatic malignant neoplasm to oesophagus|Secondary malignant neoplasm of esophagus
C0686055|T191|PT|94286009|SNOMEDCT_CORE|Secondary malignant neoplasm of esophagus|Secondary malignant neoplasm of esophagus
C0686055|T191|FN|94286009|SNOMEDCT_CORE|Secondary malignant neoplasm of esophagus|Secondary malignant neoplasm of esophagus
C0686055|T191|IS|94286009|SNOMEDCT_CORE|Secondary malignant neoplasm of esophagus, NOS|Secondary malignant neoplasm of esophagus
C0686055|T191|PTGB|94286009|SNOMEDCT_CORE|Secondary malignant neoplasm of oesophagus|Secondary malignant neoplasm of esophagus
C0686241|T191|SY|94281004|SNOMEDCT_CORE|Metastatic malignant neoplasm to endometrium|Secondary malignant neoplasm of endometrium
C0686241|T191|PT|94281004|SNOMEDCT_CORE|Secondary malignant neoplasm of endometrium|Secondary malignant neoplasm of endometrium
C0686241|T191|FN|94281004|SNOMEDCT_CORE|Secondary malignant neoplasm of endometrium|Secondary malignant neoplasm of endometrium
C0686344|T184|PT|91957002|SNOMEDCT_CORE|Back pain complicating pregnancy|Back pain complicating pregnancy
C0686344|T184|FN|91957002|SNOMEDCT_CORE|Back pain complicating pregnancy|Back pain complicating pregnancy
C0686347|T047|IS|38941006|SNOMEDCT_CORE|Tardive dyskinesia|Tardive dyskinesia
C0686366|T047|SY|41446000|SNOMEDCT_CORE|Inflammation of lid margin|Marginal blepharitis
C0686366|T047|SY|41446000|SNOMEDCT_CORE|Marginal blepharitis|Marginal blepharitis
C0686377|T191|SY|94243009|SNOMEDCT_CORE|Cancer metastatic to CNS|Secondary malignant neoplasm of central nervous system
C0686377|T191|SY|94243009|SNOMEDCT_CORE|Metastatic malignant neoplasm to central nervous system|Secondary malignant neoplasm of central nervous system
C0686377|T191|IS|94243009|SNOMEDCT_CORE|Metastatic malignant neoplasm to central nervous system, NOS|Secondary malignant neoplasm of central nervous system
C0686377|T191|PT|94243009|SNOMEDCT_CORE|Secondary malignant neoplasm of central nervous system|Secondary malignant neoplasm of central nervous system
C0686377|T191|FN|94243009|SNOMEDCT_CORE|Secondary malignant neoplasm of central nervous system|Secondary malignant neoplasm of central nervous system
C0686377|T191|IS|94243009|SNOMEDCT_CORE|Secondary malignant neoplasm of central nervous system, NOS|Secondary malignant neoplasm of central nervous system
C0686557|T191|PT|93199007|SNOMEDCT_CORE|Malignant lymphoma of extranodal AND/OR solid organ site|Malignant lymphoma of extranodal AND/OR solid organ site
C0686557|T191|FN|93199007|SNOMEDCT_CORE|Malignant lymphoma of extranodal AND/OR solid organ site|Malignant lymphoma of extranodal AND/OR solid organ site
C0686557|T191|IS|93199007|SNOMEDCT_CORE|Malignant lymphoma, NOS of unspecified, extranodal or solid organ site|Malignant lymphoma of extranodal AND/OR solid organ site
C0686587|T191|IS|91855006|SNOMEDCT_CORE|Acute leukemia, NOS, without mention of remission|Acute leukemia, NOS, without mention of remission
C0686588|T191|IS|92812005|SNOMEDCT_CORE|Chronic leukemia, NOS, without mention of remission|Chronic leukemia, NOS, without mention of remission
C0686619|T191|SY|94392001|SNOMEDCT_CORE|Cancer metastatic to lymph nodes|Secondary malignant neoplasm of lymph node
C0686619|T191|SY|94392001|SNOMEDCT_CORE|Metastatic malignant neoplasm to lymph node|Secondary malignant neoplasm of lymph node
C0686619|T191|IS|94392001|SNOMEDCT_CORE|Metastatic malignant neoplasm to lymph node, NOS|Secondary malignant neoplasm of lymph node
C0686619|T191|SY|94392001|SNOMEDCT_CORE|Secondary lymph node cancer|Secondary malignant neoplasm of lymph node
C0686619|T191|PT|94392001|SNOMEDCT_CORE|Secondary malignant neoplasm of lymph node|Secondary malignant neoplasm of lymph node
C0686619|T191|FN|94392001|SNOMEDCT_CORE|Secondary malignant neoplasm of lymph node|Secondary malignant neoplasm of lymph node
C0686619|T191|IS|94392001|SNOMEDCT_CORE|Secondary malignant neoplasm of lymph node, NOS|Secondary malignant neoplasm of lymph node
C0686623|T191|SY|94393006|SNOMEDCT_CORE|Cancer metastatic to lymph nodes of face|Secondary malignant neoplasm of lymph nodes of face
C0686623|T191|SY|94393006|SNOMEDCT_CORE|Metastatic malignant neoplasm to lymph nodes of face|Secondary malignant neoplasm of lymph nodes of face
C0686623|T191|IS|94393006|SNOMEDCT_CORE|Metastatic malignant neoplasm to lymph nodes of face, NOS|Secondary malignant neoplasm of lymph nodes of face
C0686623|T191|PT|94393006|SNOMEDCT_CORE|Secondary malignant neoplasm of lymph nodes of face|Secondary malignant neoplasm of lymph nodes of face
C0686623|T191|FN|94393006|SNOMEDCT_CORE|Secondary malignant neoplasm of lymph nodes of face|Secondary malignant neoplasm of lymph nodes of face
C0686623|T191|IS|94393006|SNOMEDCT_CORE|Secondary malignant neoplasm of lymph nodes of face, NOS|Secondary malignant neoplasm of lymph nodes of face
C0686625|T191|SY|94397007|SNOMEDCT_CORE|Cancer metastatic to neck lymph nodes|Secondary malignant neoplasm of lymph nodes of neck
C0686625|T191|SY|94397007|SNOMEDCT_CORE|Metastasis to cervical lymph nodes|Secondary malignant neoplasm of lymph nodes of neck
C0686625|T191|SY|94397007|SNOMEDCT_CORE|Metastatic malignant neoplasm to lymph nodes of neck|Secondary malignant neoplasm of lymph nodes of neck
C0686625|T191|IS|94397007|SNOMEDCT_CORE|Metastatic malignant neoplasm to lymph nodes of neck, NOS|Secondary malignant neoplasm of lymph nodes of neck
C0686625|T191|PT|94397007|SNOMEDCT_CORE|Secondary malignant neoplasm of lymph nodes of neck|Secondary malignant neoplasm of lymph nodes of neck
C0686625|T191|FN|94397007|SNOMEDCT_CORE|Secondary malignant neoplasm of lymph nodes of neck|Secondary malignant neoplasm of lymph nodes of neck
C0686625|T191|IS|94397007|SNOMEDCT_CORE|Secondary malignant neoplasm of lymph nodes of neck, NOS|Secondary malignant neoplasm of lymph nodes of neck
C0686645|T191|SY|94351005|SNOMEDCT_CORE|Cancer metastatic to intrathoracic lymph nodes|Secondary malignant neoplasm of intrathoracic lymph nodes
C0686645|T191|SY|94351005|SNOMEDCT_CORE|Metastatic malignant neoplasm to intrathoracic lymph nodes|Secondary malignant neoplasm of intrathoracic lymph nodes
C0686645|T191|IS|94351005|SNOMEDCT_CORE|Metastatic malignant neoplasm to intrathoracic lymph nodes, NOS|Secondary malignant neoplasm of intrathoracic lymph nodes
C0686645|T191|PT|94351005|SNOMEDCT_CORE|Secondary malignant neoplasm of intrathoracic lymph nodes|Secondary malignant neoplasm of intrathoracic lymph nodes
C0686645|T191|FN|94351005|SNOMEDCT_CORE|Secondary malignant neoplasm of intrathoracic lymph nodes|Secondary malignant neoplasm of intrathoracic lymph nodes
C0686645|T191|IS|94351005|SNOMEDCT_CORE|Secondary malignant neoplasm of intrathoracic lymph nodes, NOS|Secondary malignant neoplasm of intrathoracic lymph nodes
C0686655|T191|SY|94347008|SNOMEDCT_CORE|Cancer metastatic to intra-abdominal lymph nodes|Secondary malignant neoplasm of intra-abdominal lymph nodes
C0686655|T191|SY|94347008|SNOMEDCT_CORE|Metastatic malignant neoplasm to intra-abdominal lymph nodes|Secondary malignant neoplasm of intra-abdominal lymph nodes
C0686655|T191|IS|94347008|SNOMEDCT_CORE|Metastatic malignant neoplasm to intra-abdominal lymph nodes, NOS|Secondary malignant neoplasm of intra-abdominal lymph nodes
C0686655|T191|PT|94347008|SNOMEDCT_CORE|Secondary malignant neoplasm of intra-abdominal lymph nodes|Secondary malignant neoplasm of intra-abdominal lymph nodes
C0686655|T191|FN|94347008|SNOMEDCT_CORE|Secondary malignant neoplasm of intra-abdominal lymph nodes|Secondary malignant neoplasm of intra-abdominal lymph nodes
C0686655|T191|IS|94347008|SNOMEDCT_CORE|Secondary malignant neoplasm of intra-abdominal lymph nodes, NOS|Secondary malignant neoplasm of intra-abdominal lymph nodes
C0686689|T191|SY|94350006|SNOMEDCT_CORE|Cancer metastatic to intrapelvic lymph nodes|Secondary malignant neoplasm of intrapelvic lymph nodes
C0686689|T191|SY|94350006|SNOMEDCT_CORE|Metastatic malignant neoplasm to intrapelvic lymph nodes|Secondary malignant neoplasm of intrapelvic lymph nodes
C0686689|T191|IS|94350006|SNOMEDCT_CORE|Metastatic malignant neoplasm to intrapelvic lymph nodes, NOS|Secondary malignant neoplasm of intrapelvic lymph nodes
C0686689|T191|PT|94350006|SNOMEDCT_CORE|Secondary malignant neoplasm of intrapelvic lymph nodes|Secondary malignant neoplasm of intrapelvic lymph nodes
C0686689|T191|FN|94350006|SNOMEDCT_CORE|Secondary malignant neoplasm of intrapelvic lymph nodes|Secondary malignant neoplasm of intrapelvic lymph nodes
C0686689|T191|IS|94350006|SNOMEDCT_CORE|Secondary malignant neoplasm of intrapelvic lymph nodes, NOS|Secondary malignant neoplasm of intrapelvic lymph nodes
C0686724|T033|FN|95317002|SNOMEDCT_CORE|Victim of terrorism|Victim of terrorism
C0686724|T033|PT|95317002|SNOMEDCT_CORE|Victim of terrorism|Victim of terrorism
C0687140|T191|PTGB|93471006|SNOMEDCT_CORE|Haemangioma of skin|Hemangioma of skin
C0687140|T191|PT|93471006|SNOMEDCT_CORE|Hemangioma of skin|Hemangioma of skin
C0687140|T191|FN|93471006|SNOMEDCT_CORE|Hemangioma of skin|Hemangioma of skin
C0687707|T047|PT|426867001|SNOMEDCT_CORE|Anorectal disorder|Anorectal disorder
C0687707|T047|FN|426867001|SNOMEDCT_CORE|Anorectal disorder|Anorectal disorder
C0687720|T047|SY|45369008|SNOMEDCT_CORE|Central diabetes insipidus|Neurohypophyseal diabetes insipidus
C0687720|T047|IS|15771004|SNOMEDCT_CORE|Cranial diabetes insipidus|Neurohypophyseal diabetes insipidus
C0687720|T047|SY|45369008|SNOMEDCT_CORE|Cranial diabetes insipidus|Neurohypophyseal diabetes insipidus
C0687720|T047|SY|45369008|SNOMEDCT_CORE|Diabetes insipidus - pituitary|Neurohypophyseal diabetes insipidus
C0687720|T047|SY|45369008|SNOMEDCT_CORE|Diabetes insipidus secondary to vasopressin deficiency|Neurohypophyseal diabetes insipidus
C0687720|T047|IS|15771004|SNOMEDCT_CORE|Neurogenic diabetes insipidus|Neurohypophyseal diabetes insipidus
C0687720|T047|SY|45369008|SNOMEDCT_CORE|Neurogenic diabetes insipidus|Neurohypophyseal diabetes insipidus
C0687720|T047|PT|45369008|SNOMEDCT_CORE|Neurohypophyseal diabetes insipidus|Neurohypophyseal diabetes insipidus
C0687720|T047|FN|45369008|SNOMEDCT_CORE|Neurohypophyseal diabetes insipidus|Neurohypophyseal diabetes insipidus
C0687720|T047|IS|15771004|SNOMEDCT_CORE|Neurohypophyseal diabetes insipidus, NOS|Neurohypophyseal diabetes insipidus
C0687720|T047|IS|45369008|SNOMEDCT_CORE|Neurohypophyseal diabetes insipidus, NOS|Neurohypophyseal diabetes insipidus
C0687720|T047|IS|15771004|SNOMEDCT_CORE|Pituitary diabetes insipidus|Neurohypophyseal diabetes insipidus
C0687720|T047|SY|45369008|SNOMEDCT_CORE|Pituitary diabetes insipidus|Neurohypophyseal diabetes insipidus
C0687720|T047|IS|15771004|SNOMEDCT_CORE|Primary central diabetes insipidus|Neurohypophyseal diabetes insipidus
C0687720|T047|SY|45369008|SNOMEDCT_CORE|Primary central diabetes insipidus|Neurohypophyseal diabetes insipidus
C0687720|T047|SY|45369008|SNOMEDCT_CORE|Vasopressin deficiency|Neurohypophyseal diabetes insipidus
C0687720|T047|IS|15771004|SNOMEDCT_CORE|Vasopressin deficiency syndrome|Neurohypophyseal diabetes insipidus
C0687720|T047|SY|45369008|SNOMEDCT_CORE|Vasopressin deficiency syndrome|Neurohypophyseal diabetes insipidus
C0687754|T047|SYGB|276549000|SNOMEDCT_CORE|Transient neonatal hyperbilirubinaemia|Transient neonatal hyperbilirubinemia
C0687754|T047|SY|276549000|SNOMEDCT_CORE|Transient neonatal hyperbilirubinemia|Transient neonatal hyperbilirubinemia
C0694499|T047|IS|195029002|SNOMEDCT_CORE|Cardiomyopathy in disease EC|Cardiomyopathy in disease EC
C0694499|T047|OF|195029002|SNOMEDCT_CORE|Cardiomyopathy in disease EC|Cardiomyopathy in disease EC
C0694536|T033|SY|441668002|SNOMEDCT_CORE|Drug seeking|Drug seeking behavior
C0694536|T033|PT|441668002|SNOMEDCT_CORE|Drug seeking behavior|Drug seeking behavior
C0694536|T033|FN|441668002|SNOMEDCT_CORE|Drug seeking behavior|Drug seeking behavior
C0694536|T033|PTGB|441668002|SNOMEDCT_CORE|Drug seeking behaviour|Drug seeking behavior
C0694539|T047|PT|426749004|SNOMEDCT_CORE|Chronic atrial fibrillation|Chronic atrial fibrillation
C0694539|T047|FN|426749004|SNOMEDCT_CORE|Chronic atrial fibrillation|Chronic atrial fibrillation
C0694541|T047|SY|64715009|SNOMEDCT_CORE|Hypertensive cardiomegaly|Hypertensive cardiomegaly
C0694548|T047|PT|409663006|SNOMEDCT_CORE|Cough variant asthma|Cough variant asthma
C0694548|T047|FN|409663006|SNOMEDCT_CORE|Cough variant asthma|Cough variant asthma
C0694549|T047|PT|385093006|SNOMEDCT_CORE|Community acquired pneumonia|Community acquired pneumonia
C0694549|T047|FN|385093006|SNOMEDCT_CORE|Community acquired pneumonia|Community acquired pneumonia
C0694551|T184|PT|301754002|SNOMEDCT_CORE|Right lower quadrant pain|Right lower quadrant pain
C0694551|T184|FN|301754002|SNOMEDCT_CORE|Right lower quadrant pain|Right lower quadrant pain
C0695242|T047|PT|425671009|SNOMEDCT_CORE|Neurogenic bowel|Neurogenic bowel
C0695242|T047|FN|425671009|SNOMEDCT_CORE|Neurogenic bowel|Neurogenic bowel
C0699757|T048|SY|25702006|SNOMEDCT_CORE|Acute alcoholism|Acute alcoholism
C0699790|T191|PT|269533000|SNOMEDCT_CORE|Carcinoma of colon|Carcinoma of colon
C0699790|T191|FN|269533000|SNOMEDCT_CORE|Carcinoma of colon|Carcinoma of colon
C0699791|T191|PT|372143007|SNOMEDCT_CORE|Carcinoma of stomach|Carcinoma of stomach
C0699791|T191|FN|372143007|SNOMEDCT_CORE|Carcinoma of stomach|Carcinoma of stomach
C0699791|T191|SY|372143007|SNOMEDCT_CORE|Gastric carcinoma|Carcinoma of stomach
C0699815|T033|PT|274540003|SNOMEDCT_CORE|Feeding difficulties and mismanagement|Feeding difficulties and mismanagement
C0699815|T033|FN|274540003|SNOMEDCT_CORE|Feeding difficulties and mismanagement|Feeding difficulties and mismanagement
C0699885|T191|PT|255108000|SNOMEDCT_CORE|Carcinoma of bladder|Carcinoma of bladder
C0699885|T191|FN|255108000|SNOMEDCT_CORE|Carcinoma of bladder|Carcinoma of bladder
C0700031|T048|PT|300895004|SNOMEDCT_CORE|Anxiety attack|Anxiety attack
C0700031|T048|FN|300895004|SNOMEDCT_CORE|Anxiety attack|Anxiety attack
C0700101|T191|SY|363459007|SNOMEDCT_CORE|CA - Cancer of urethra|CA - Cancer of urethra
C0700101|T191|SY|363459007|SNOMEDCT_CORE|Urethral Ca|CA - Cancer of urethra
C0700184|T184|IS|405737000|SNOMEDCT_CORE|Irritation of the throat|Irritation of the throat
C0700198|T046|SY|68052005|SNOMEDCT_CORE|Aspiration|Pulmonary aspiration
C0700198|T046|IS|68052005|SNOMEDCT_CORE|Aspiration, NOS|Pulmonary aspiration
C0700198|T046|PT|68052005|SNOMEDCT_CORE|Pulmonary aspiration|Pulmonary aspiration
C0700198|T046|FN|68052005|SNOMEDCT_CORE|Pulmonary aspiration|Pulmonary aspiration
C0700198|T046|IS|68052005|SNOMEDCT_CORE|Pulmonary aspiration, NOS|Pulmonary aspiration
C0700200|T184|PT|427461000|SNOMEDCT_CORE|Near syncope|Near syncope
C0700200|T184|FN|427461000|SNOMEDCT_CORE|Near syncope|Near syncope
C0700200|T184|SY|427461000|SNOMEDCT_CORE|Presyncope|Near syncope
C0700201|T048|PT|44186003|SNOMEDCT_CORE|Dyssomnia|Dyssomnia
C0700201|T048|FN|44186003|SNOMEDCT_CORE|Dyssomnia|Dyssomnia
C0700201|T048|IS|44186003|SNOMEDCT_CORE|Dyssomnia, NOS|Dyssomnia
C0700201|T048|SY|44186003|SNOMEDCT_CORE|Sleep disturbance|Dyssomnia
C0700201|T048|SY|44186003|SNOMEDCT_CORE|Sleep problem|Dyssomnia
C0700208|T020|PT|111266001|SNOMEDCT_CORE|Acquired scoliosis|Acquired scoliosis
C0700208|T020|FN|111266001|SNOMEDCT_CORE|Acquired scoliosis|Acquired scoliosis
C0700208|T020|IS|111266001|SNOMEDCT_CORE|Scoliosis|Acquired scoliosis
C0700211|T047|IS|66071002|SNOMEDCT_CORE|Viral hepatitis B without mention of hepatic coma|Viral hepatitis B without mention of hepatic coma
C0700225|T033|PT|166717003|SNOMEDCT_CORE|Serum creatinine raised|Serum creatinine raised
C0700225|T033|FN|166717003|SNOMEDCT_CORE|Serum creatinine raised|Serum creatinine raised
C0700226|T047|PT|373435003|SNOMEDCT_CORE|Battey disease|Battey disease
C0700226|T047|FN|373435003|SNOMEDCT_CORE|Battey disease|Battey disease
C0700226|T047|IS|373435003|SNOMEDCT_CORE|Pulmonary mycobacterium avium-intracellulare infection|Battey disease
C0700226|T047|SY|373435003|SNOMEDCT_CORE|Pulmonary mycobacterium intracellulare infection|Battey disease
C0700251|T047|SY|3548001|SNOMEDCT_CORE|BPN - Brachial plexus neuropathy|Brachial plexus disorder
C0700251|T047|PT|3548001|SNOMEDCT_CORE|Brachial plexus disorder|Brachial plexus disorder
C0700251|T047|FN|3548001|SNOMEDCT_CORE|Brachial plexus disorder|Brachial plexus disorder
C0700251|T047|SY|3548001|SNOMEDCT_CORE|Brachial plexus neuropathy|Brachial plexus disorder
C0700251|T047|IS|3548001|SNOMEDCT_CORE|Brachial plexus neuropathy, NOS|Brachial plexus disorder
C0700292|T033|SYGB|389087006|SNOMEDCT_CORE|Arterial hypoxaemia|Hypoxemia
C0700292|T033|SY|389087006|SNOMEDCT_CORE|Arterial hypoxemia|Hypoxemia
C0700292|T033|PTGB|389087006|SNOMEDCT_CORE|Hypoxaemia|Hypoxemia
C0700292|T033|PT|389087006|SNOMEDCT_CORE|Hypoxemia|Hypoxemia
C0700292|T033|FN|389087006|SNOMEDCT_CORE|Hypoxemia|Hypoxemia
C0700318|T047|SY|89155008|SNOMEDCT_CORE|Thibierge-Weissenbach syndrome|Thibierge-Weissenbach syndrome
C0700345|T047|PT|72605008|SNOMEDCT_CORE|Candidal vulvovaginitis|Candidal vulvovaginitis
C0700345|T047|FN|72605008|SNOMEDCT_CORE|Candidal vulvovaginitis|Candidal vulvovaginitis
C0700345|T047|SY|72605008|SNOMEDCT_CORE|Monilial vulvovaginitis|Candidal vulvovaginitis
C0700345|T047|SY|72605008|SNOMEDCT_CORE|Vulvovaginal thrush|Candidal vulvovaginitis
C0700440|T033|PT|274710003|SNOMEDCT_CORE|Lung field abnormal|Lung field abnormal
C0700440|T033|FN|274710003|SNOMEDCT_CORE|Lung field abnormal|Lung field abnormal
C0700501|T019|PT|64635004|SNOMEDCT_CORE|Congenital nystagmus|Congenital nystagmus
C0700501|T019|FN|64635004|SNOMEDCT_CORE|Congenital nystagmus|Congenital nystagmus
C0700502|T047|PT|111566002|SNOMEDCT_CORE|Acquired hypothyroidism|Acquired hypothyroidism
C0700502|T047|FN|111566002|SNOMEDCT_CORE|Acquired hypothyroidism|Acquired hypothyroidism
C0700502|T047|IS|111566002|SNOMEDCT_CORE|Acquired hypothyroidism, NOS|Acquired hypothyroidism
C0700502|T047|SY|111566002|SNOMEDCT_CORE|Primary hypothyroidism|Acquired hypothyroidism
C0700509|T047|PT|128287004|SNOMEDCT_CORE|Chronic peptic ulcer|Chronic peptic ulcer
C0700509|T047|FN|128287004|SNOMEDCT_CORE|Chronic peptic ulcer|Chronic peptic ulcer
C0700590|T033|SY|52613005|SNOMEDCT_CORE|Diaphoresis|Excessive sweating
C0700590|T033|PT|52613005|SNOMEDCT_CORE|Excessive sweating|Excessive sweating
C0700590|T033|FN|52613005|SNOMEDCT_CORE|Excessive sweating|Excessive sweating
C0700590|T033|IS|52613005|SNOMEDCT_CORE|Increased sweating|Excessive sweating
C0700590|T033|SY|52613005|SNOMEDCT_CORE|Profuse sweating|Excessive sweating
C0700590|T033|SY|52613005|SNOMEDCT_CORE|Sweating profusely|Excessive sweating
C0700594|T047|SY|72274001|SNOMEDCT_CORE|Radiculopathy|Radiculopathy
C0700594|T047|IS|72274001|SNOMEDCT_CORE|Radiculopathy, NOS|Radiculopathy
C0700613|T048|IS|207363009|SNOMEDCT_CORE|Anxiety state|Anxiety state
C0700613|T048|PT|198288003|SNOMEDCT_CORE|Anxiety state|Anxiety state
C0700613|T048|FN|198288003|SNOMEDCT_CORE|Anxiety state|Anxiety state
C0701807|T047|SY|4927003|SNOMEDCT_CORE|AAU - acute anterior uveitis|Acute anterior uveitis
C0701807|T047|PT|4927003|SNOMEDCT_CORE|Acute anterior uveitis|Acute anterior uveitis
C0701807|T047|FN|4927003|SNOMEDCT_CORE|Acute anterior uveitis|Acute anterior uveitis
C0701811|T048|PT|247592009|SNOMEDCT_CORE|Poor short-term memory|Poor short-term memory
C0701811|T048|FN|247592009|SNOMEDCT_CORE|Poor short-term memory|Poor short-term memory
C0701811|T048|SY|247592009|SNOMEDCT_CORE|Short term memory loss|Poor short-term memory
C0701811|T048|SY|247592009|SNOMEDCT_CORE|Short-term memory loss|Poor short-term memory
C0701847|T047|SY|16607004|SNOMEDCT_CORE|Fetal death before 22 weeks with retention of dead fetus|Fetal death before 22 weeks with retention of dead fetus
C0702157|T047|PTGB|19442009|SNOMEDCT_CORE|Heterozygous thalassaemia|Heterozygous thalassemia
C0702157|T047|PT|19442009|SNOMEDCT_CORE|Heterozygous thalassemia|Heterozygous thalassemia
C0702157|T047|FN|19442009|SNOMEDCT_CORE|Heterozygous thalassemia|Heterozygous thalassemia
C0702157|T047|IS|19442009|SNOMEDCT_CORE|Heterozygous thalassemia, NOS|Heterozygous thalassemia
C0702157|T047|SYGB|19442009|SNOMEDCT_CORE|Thalassaemia trait|Heterozygous thalassemia
C0702157|T047|SY|19442009|SNOMEDCT_CORE|Thalassemia trait|Heterozygous thalassemia
C0702157|T047|IS|19442009|SNOMEDCT_CORE|Thalassemia trait, NOS|Heterozygous thalassemia
C0702166|T047|PT|11381005|SNOMEDCT_CORE|Acne|Acne
C0702166|T047|OF|11381005|SNOMEDCT_CORE|Acne|Acne
C0702166|T047|SY|11381005|SNOMEDCT_CORE|Acne vulgaris|Acne
C0702166|T047|FN|11381005|SNOMEDCT_CORE|Acne vulgaris|Acne
C0702166|T047|IS|11381005|SNOMEDCT_CORE|Acne, NOS|Acne
C0702166|T047|SY|11381005|SNOMEDCT_CORE|Common acne|Acne
C0702176|T047|FN|6284004|SNOMEDCT_CORE|Abscess of neck|Cervical abscess
C0702176|T047|SY|6284004|SNOMEDCT_CORE|Cervical abscess|Cervical abscess
C0728711|T033|SY|429011007|SNOMEDCT_CORE|Family history of lung cancer|Family history of malignant neoplasm of lung
C0728711|T033|PT|429011007|SNOMEDCT_CORE|Family history of malignant neoplasm of lung|Family history of malignant neoplasm of lung
C0728711|T033|FN|429011007|SNOMEDCT_CORE|Family history of malignant neoplasm of lung|Family history of malignant neoplasm of lung
C0728731|T033|OAS|44247006|SNOMEDCT_CORE|Prematurity|Prematurity of fetus
C0728731|T033|OAP|44247006|SNOMEDCT_CORE|Prematurity of fetus|Prematurity of fetus
C0728731|T033|OAF|44247006|SNOMEDCT_CORE|Prematurity of fetus|Prematurity of fetus
C0728731|T033|IS|44247006|SNOMEDCT_CORE|Prematurity of fetus, NOS|Prematurity of fetus
C0728731|T033|OAS|44247006|SNOMEDCT_CORE|Prematurity of foetus|Prematurity of fetus
C0728731|T033|IS|44247006|SNOMEDCT_CORE|Prematurity, NOS|Prematurity of fetus
C0728731|T033|OAS|44247006|SNOMEDCT_CORE|Preterm infant|Prematurity of fetus
C0728731|T033|IS|44247006|SNOMEDCT_CORE|Preterm infant, NOS|Prematurity of fetus
C0728864|T191|SY|363422006|SNOMEDCT_CORE|Malignant neoplasm of nasal cavities|Malignant tumor of nasal cavity
C0728864|T191|PT|363422006|SNOMEDCT_CORE|Malignant tumor of nasal cavity|Malignant tumor of nasal cavity
C0728864|T191|FN|363422006|SNOMEDCT_CORE|Malignant tumor of nasal cavity|Malignant tumor of nasal cavity
C0728864|T191|PTGB|363422006|SNOMEDCT_CORE|Malignant tumour of nasal cavity|Malignant tumor of nasal cavity
C0728936|T047|SY|49601007|SNOMEDCT_CORE|Disorder of circulatory system|Disorder of circulatory system
C0728936|T047|IS|49601007|SNOMEDCT_CORE|Disorder of circulatory system, NOS|Disorder of circulatory system
C0728936|T047|SY|49601007|SNOMEDCT_CORE|Disorder of the circulatory system|Disorder of circulatory system
C0729245|T047|FN|196682000|SNOMEDCT_CORE|Acute peptic ulcer|Acute peptic ulcer
C0729245|T047|PT|196682000|SNOMEDCT_CORE|Acute peptic ulcer|Acute peptic ulcer
C0729248|T033|OAP|267129008|SNOMEDCT_CORE|Inadequate housing|Inadequate housing
C0729248|T033|OAF|267129008|SNOMEDCT_CORE|Inadequate housing|Inadequate housing
C0729262|T033|SY|35298007|SNOMEDCT_CORE|Colonic constipation|Slow transit constipation
C0729262|T033|SY|35298007|SNOMEDCT_CORE|Constipation by delayed colonic transit|Slow transit constipation
C0729262|T033|PT|35298007|SNOMEDCT_CORE|Slow transit constipation|Slow transit constipation
C0729262|T033|FN|35298007|SNOMEDCT_CORE|Slow transit constipation|Slow transit constipation
C0729264|T046|SY|312974005|SNOMEDCT_CORE|PPROM - Preterm premature rupture of membranes|Preterm premature rupture of membranes
C0729264|T046|FN|312974005|SNOMEDCT_CORE|Preterm premature rupture of membranes|Preterm premature rupture of membranes
C0729264|T046|PT|312974005|SNOMEDCT_CORE|Preterm premature rupture of membranes|Preterm premature rupture of membranes
C0729728|T190|PT|312373008|SNOMEDCT_CORE|Femoral false aneurysm|Femoral false aneurysm
C0729728|T190|FN|312373008|SNOMEDCT_CORE|Femoral false aneurysm|Femoral false aneurysm
C0729728|T190|SY|312373008|SNOMEDCT_CORE|Pseudoaneurysm of femoral artery|Femoral false aneurysm
C0729733|T047|PT|233956002|SNOMEDCT_CORE|Aortoiliac atherosclerosis|Aortoiliac atherosclerosis
C0729733|T047|FN|233956002|SNOMEDCT_CORE|Aortoiliac atherosclerosis|Aortoiliac atherosclerosis
C0729733|T047|SY|233956002|SNOMEDCT_CORE|Aortoiliac disease|Aortoiliac atherosclerosis
C0729790|T033|PT|312442005|SNOMEDCT_CORE|H/O: atrial fibrillation|H/O: atrial fibrillation
C0729790|T033|OF|312442005|SNOMEDCT_CORE|History of - atrial fibrillation|H/O: atrial fibrillation
C0729790|T033|IS|312442005|SNOMEDCT_CORE|History of - atrial fibrillation|H/O: atrial fibrillation
C0729790|T033|FN|312442005|SNOMEDCT_CORE|History of atrial fibrillation|H/O: atrial fibrillation
C0729790|T033|SY|312442005|SNOMEDCT_CORE|History of atrial fibrillation|H/O: atrial fibrillation
C0729949|T046|SY|90958004|SNOMEDCT_CORE|Lower limb arterial thrombosis|Thrombosis of arteries of lower extremity
C0729949|T046|PT|90958004|SNOMEDCT_CORE|Thrombosis of arteries of lower extremity|Thrombosis of arteries of lower extremity
C0729949|T046|FN|90958004|SNOMEDCT_CORE|Thrombosis of arteries of lower extremity|Thrombosis of arteries of lower extremity
C0730194|T047|PT|123798002|SNOMEDCT_CORE|Lumbosacral spondylosis|Lumbosacral spondylosis
C0730194|T047|FN|123798002|SNOMEDCT_CORE|Lumbosacral spondylosis|Lumbosacral spondylosis
C0730200|T033|PT|312824007|SNOMEDCT_CORE|Family history of cancer of colon|Family history of cancer of colon
C0730200|T033|OF|312824007|SNOMEDCT_CORE|Family history of cancer of colon|Family history of cancer of colon
C0730200|T033|FN|312824007|SNOMEDCT_CORE|Family history of cancer of colon|Family history of cancer of colon
C0730226|T033|PT|312850006|SNOMEDCT_CORE|H/O: Disorder|H/O: Disorder
C0730226|T033|OF|312850006|SNOMEDCT_CORE|History of - disorder|H/O: Disorder
C0730226|T033|IS|312850006|SNOMEDCT_CORE|History of - disorder|H/O: Disorder
C0730226|T033|FN|312850006|SNOMEDCT_CORE|History of disorder|H/O: Disorder
C0730226|T033|SY|312850006|SNOMEDCT_CORE|History of disorder|H/O: Disorder
C0730276|T047|IS|312903003|SNOMEDCT_CORE|Mild non proliferative diabetic retinopathy|Mild nonproliferative retinopathy due to diabetes mellitus
C0730276|T047|OF|312903003|SNOMEDCT_CORE|Mild non proliferative diabetic retinopathy|Mild nonproliferative retinopathy due to diabetes mellitus
C0730276|T047|SY|312903003|SNOMEDCT_CORE|Mild non proliferative retinopathy|Mild nonproliferative retinopathy due to diabetes mellitus
C0730276|T047|SY|312903003|SNOMEDCT_CORE|Mild non-proliferative diabetic retinopathy|Mild nonproliferative retinopathy due to diabetes mellitus
C0730276|T047|OF|312903003|SNOMEDCT_CORE|Mild non-proliferative diabetic retinopathy|Mild nonproliferative retinopathy due to diabetes mellitus
C0730276|T047|SY|312903003|SNOMEDCT_CORE|Mild nonproliferative diabetic retinopathy|Mild nonproliferative retinopathy due to diabetes mellitus
C0730276|T047|SY|312903003|SNOMEDCT_CORE|Mild nonproliferative retinopathy|Mild nonproliferative retinopathy due to diabetes mellitus
C0730276|T047|OF|312903003|SNOMEDCT_CORE|Mild nonproliferative retinopathy co-occurrent and due to diabetes mellitus|Mild nonproliferative retinopathy due to diabetes mellitus
C0730276|T047|IS|312903003|SNOMEDCT_CORE|Mild nonproliferative retinopathy co-occurrent and due to diabetes mellitus|Mild nonproliferative retinopathy due to diabetes mellitus
C0730276|T047|PT|312903003|SNOMEDCT_CORE|Mild nonproliferative retinopathy due to diabetes mellitus|Mild nonproliferative retinopathy due to diabetes mellitus
C0730276|T047|FN|312903003|SNOMEDCT_CORE|Mild nonproliferative retinopathy due to diabetes mellitus|Mild nonproliferative retinopathy due to diabetes mellitus
C0730277|T047|OF|312904009|SNOMEDCT_CORE|Moderate non proliferative diabetic retinopathy|Moderate nonproliferative retinopathy due to diabetes mellitus
C0730277|T047|IS|312904009|SNOMEDCT_CORE|Moderate non proliferative diabetic retinopathy|Moderate nonproliferative retinopathy due to diabetes mellitus
C0730277|T047|SY|312904009|SNOMEDCT_CORE|Moderate non-proliferative diabetic retinopathy|Moderate nonproliferative retinopathy due to diabetes mellitus
C0730277|T047|OF|312904009|SNOMEDCT_CORE|Moderate nonproliferative diabetic retinopathy|Moderate nonproliferative retinopathy due to diabetes mellitus
C0730277|T047|SY|312904009|SNOMEDCT_CORE|Moderate nonproliferative diabetic retinopathy|Moderate nonproliferative retinopathy due to diabetes mellitus
C0730277|T047|SY|312904009|SNOMEDCT_CORE|Moderate nonproliferative retinopathy|Moderate nonproliferative retinopathy due to diabetes mellitus
C0730277|T047|OF|312904009|SNOMEDCT_CORE|Moderate nonproliferative retinopathy co-occurrent and due to diabetes mellitus|Moderate nonproliferative retinopathy due to diabetes mellitus
C0730277|T047|IS|312904009|SNOMEDCT_CORE|Moderate nonproliferative retinopathy co-occurrent and due to diabetes mellitus|Moderate nonproliferative retinopathy due to diabetes mellitus
C0730277|T047|PT|312904009|SNOMEDCT_CORE|Moderate nonproliferative retinopathy due to diabetes mellitus|Moderate nonproliferative retinopathy due to diabetes mellitus
C0730277|T047|FN|312904009|SNOMEDCT_CORE|Moderate nonproliferative retinopathy due to diabetes mellitus|Moderate nonproliferative retinopathy due to diabetes mellitus
C0730278|T047|OF|312905005|SNOMEDCT_CORE|Severe non proliferative diabetic retinopathy|Severe nonproliferative retinopathy due to diabetes mellitus
C0730278|T047|IS|312905005|SNOMEDCT_CORE|Severe non proliferative diabetic retinopathy|Severe nonproliferative retinopathy due to diabetes mellitus
C0730278|T047|SY|312905005|SNOMEDCT_CORE|Severe nonproliferative diabetic retinopathy|Severe nonproliferative retinopathy due to diabetes mellitus
C0730278|T047|OF|312905005|SNOMEDCT_CORE|Severe nonproliferative diabetic retinopathy|Severe nonproliferative retinopathy due to diabetes mellitus
C0730278|T047|SY|312905005|SNOMEDCT_CORE|Severe nonproliferative retinopathy|Severe nonproliferative retinopathy due to diabetes mellitus
C0730278|T047|OF|312905005|SNOMEDCT_CORE|Severe nonproliferative retinopathy co-occurrent and due to diabetes mellitus|Severe nonproliferative retinopathy due to diabetes mellitus
C0730278|T047|IS|312905005|SNOMEDCT_CORE|Severe nonproliferative retinopathy co-occurrent and due to diabetes mellitus|Severe nonproliferative retinopathy due to diabetes mellitus
C0730278|T047|FN|312905005|SNOMEDCT_CORE|Severe nonproliferative retinopathy due to diabetes mellitus|Severe nonproliferative retinopathy due to diabetes mellitus
C0730278|T047|PT|312905005|SNOMEDCT_CORE|Severe nonproliferative retinopathy due to diabetes mellitus|Severe nonproliferative retinopathy due to diabetes mellitus
C0730278|T047|SY|312905005|SNOMEDCT_CORE|Severe NPDR|Severe nonproliferative retinopathy due to diabetes mellitus
C0730278|T047|IS|312905005|SNOMEDCT_CORE|Severe NPDR|Severe nonproliferative retinopathy due to diabetes mellitus
C0730285|T047|SY|312912001|SNOMEDCT_CORE|Diabetic macular edema|Macular edema due to diabetes mellitus
C0730285|T047|OF|312912001|SNOMEDCT_CORE|Diabetic macular edema|Macular edema due to diabetes mellitus
C0730285|T047|SYGB|312912001|SNOMEDCT_CORE|Diabetic macular oedema|Macular edema due to diabetes mellitus
C0730285|T047|IS|312912001|SNOMEDCT_CORE|Macular edema co-occurrent and due to diabetes mellitus|Macular edema due to diabetes mellitus
C0730285|T047|OF|312912001|SNOMEDCT_CORE|Macular edema co-occurrent and due to diabetes mellitus|Macular edema due to diabetes mellitus
C0730285|T047|PT|312912001|SNOMEDCT_CORE|Macular edema due to diabetes mellitus|Macular edema due to diabetes mellitus
C0730285|T047|FN|312912001|SNOMEDCT_CORE|Macular edema due to diabetes mellitus|Macular edema due to diabetes mellitus
C0730285|T047|IS|312912001|SNOMEDCT_CORE|Macular oedema co-occurrent and due to diabetes mellitus|Macular edema due to diabetes mellitus
C0730285|T047|OP|312912001|SNOMEDCT_CORE|Macular oedema due to diabetes mallitus|Macular edema due to diabetes mellitus
C0730285|T047|PTGB|312912001|SNOMEDCT_CORE|Macular oedema due to diabetes mellitus|Macular edema due to diabetes mellitus
C0730328|T047|PT|312956001|SNOMEDCT_CORE|Central serous chorioretinopathy|Central serous chorioretinopathy
C0730328|T047|FN|312956001|SNOMEDCT_CORE|Central serous chorioretinopathy|Central serous chorioretinopathy
C0730328|T047|SY|312956001|SNOMEDCT_CORE|Central serous choroidopathy|Central serous chorioretinopathy
C0730328|T047|SY|312956001|SNOMEDCT_CORE|Central serous retinopathy|Central serous chorioretinopathy
C0730328|T047|IS|312956001|SNOMEDCT_CORE|central serous retinopathy|Central serous chorioretinopathy
C0730328|T047|SY|312956001|SNOMEDCT_CORE|CSC - Central serous choroidopathy|Central serous chorioretinopathy
C0730328|T047|SY|312956001|SNOMEDCT_CORE|CSR - central serous retinopathy|Central serous chorioretinopathy
C0730345|T033|PT|312975006|SNOMEDCT_CORE|Microalbuminuria|Microalbuminuria
C0730345|T033|FN|312975006|SNOMEDCT_CORE|Microalbuminuria|Microalbuminuria
C0730345|T033|SY|312975006|SNOMEDCT_CORE|Moderately increased albuminuria|Microalbuminuria
C0730504|T047|PT|313157004|SNOMEDCT_CORE|Pseudostrabismus|Pseudostrabismus
C0730504|T047|FN|313157004|SNOMEDCT_CORE|Pseudostrabismus|Pseudostrabismus
C0730525|T048|PT|313182004|SNOMEDCT_CORE|Chronic post-traumatic stress disorder|Chronic post-traumatic stress disorder
C0730525|T048|FN|313182004|SNOMEDCT_CORE|Chronic post-traumatic stress disorder|Chronic post-traumatic stress disorder
C0730576|T047|PTGB|313259008|SNOMEDCT_CORE|Localised, primary osteoarthritis of elbow|Localized, primary osteoarthritis of elbow
C0730576|T047|PT|313259008|SNOMEDCT_CORE|Localized, primary osteoarthritis of elbow|Localized, primary osteoarthritis of elbow
C0730576|T047|FN|313259008|SNOMEDCT_CORE|Localized, primary osteoarthritis of elbow|Localized, primary osteoarthritis of elbow
C0730604|T047|PT|313296004|SNOMEDCT_CORE|Mild chronic obstructive pulmonary disease|Mild chronic obstructive pulmonary disease
C0730604|T047|FN|313296004|SNOMEDCT_CORE|Mild chronic obstructive pulmonary disease|Mild chronic obstructive pulmonary disease
C0730605|T047|PT|313297008|SNOMEDCT_CORE|Moderate chronic obstructive pulmonary disease|Moderate chronic obstructive pulmonary disease
C0730605|T047|FN|313297008|SNOMEDCT_CORE|Moderate chronic obstructive pulmonary disease|Moderate chronic obstructive pulmonary disease
C0730607|T047|PT|313299006|SNOMEDCT_CORE|Severe chronic obstructive pulmonary disease|Severe chronic obstructive pulmonary disease
C0730607|T047|FN|313299006|SNOMEDCT_CORE|Severe chronic obstructive pulmonary disease|Severe chronic obstructive pulmonary disease
C0740083|T191|PT|372103002|SNOMEDCT_CORE|Carcinoma of glottis|Carcinoma of glottis
C0740083|T191|FN|372103002|SNOMEDCT_CORE|Carcinoma of glottis|Carcinoma of glottis
C0740394|T047|PTGB|35885006|SNOMEDCT_CORE|Hyperuricaemia|Hyperuricemia
C0740394|T047|PT|35885006|SNOMEDCT_CORE|Hyperuricemia|Hyperuricemia
C0740394|T047|FN|35885006|SNOMEDCT_CORE|Hyperuricemia|Hyperuricemia
C0740394|T047|IS|35885006|SNOMEDCT_CORE|Hyperuricemia, NOS|Hyperuricemia
C0740394|T047|SYGB|35885006|SNOMEDCT_CORE|Uricacidaemia|Hyperuricemia
C0740394|T047|SY|35885006|SNOMEDCT_CORE|Uricacidemia|Hyperuricemia
C0740394|T047|IS|35885006|SNOMEDCT_CORE|Uricacidemia, NOS|Hyperuricemia
C0740418|T184|PT|134407002|SNOMEDCT_CORE|Chronic back pain|Chronic back pain
C0740418|T184|OF|134407002|SNOMEDCT_CORE|Chronic back pain|Chronic back pain
C0740418|T184|FN|134407002|SNOMEDCT_CORE|Chronic back pain|Chronic back pain
C0740421|T047|PT|371036001|SNOMEDCT_CORE|Postsurgical menopause|Postsurgical menopause
C0740421|T047|FN|371036001|SNOMEDCT_CORE|Postsurgical menopause|Postsurgical menopause
C0740421|T047|SY|371036001|SNOMEDCT_CORE|Surgical menopause|Postsurgical menopause
C0740447|T047|PT|424736006|SNOMEDCT_CORE|Diabetic peripheral neuropathy|Diabetic peripheral neuropathy
C0740447|T047|OF|424736006|SNOMEDCT_CORE|Diabetic peripheral neuropathy|Diabetic peripheral neuropathy
C0740447|T047|OF|424736006|SNOMEDCT_CORE|Peripheral neuropathy co-occurrent and due to diabetes mellitus|Diabetic peripheral neuropathy
C0740447|T047|IS|424736006|SNOMEDCT_CORE|Peripheral neuropathy co-occurrent and due to diabetes mellitus|Diabetic peripheral neuropathy
C0740447|T047|FN|424736006|SNOMEDCT_CORE|Peripheral neuropathy due to diabetes mellitus|Diabetic peripheral neuropathy
C0740447|T047|SY|424736006|SNOMEDCT_CORE|Peripheral neuropathy due to diabetes mellitus|Diabetic peripheral neuropathy
C0740457|T191|SY|363518003|SNOMEDCT_CORE|CA - Cancer of kidney|Malignant tumor of kidney
C0740457|T191|SY|363518003|SNOMEDCT_CORE|CA - Renal cancer|Malignant tumor of kidney
C0740457|T191|PT|363518003|SNOMEDCT_CORE|Malignant tumor of kidney|Malignant tumor of kidney
C0740457|T191|FN|363518003|SNOMEDCT_CORE|Malignant tumor of kidney|Malignant tumor of kidney
C0740457|T191|PTGB|363518003|SNOMEDCT_CORE|Malignant tumour of kidney|Malignant tumor of kidney
C0740457|T191|SY|363518003|SNOMEDCT_CORE|Renal cancer|Malignant tumor of kidney
C0740457|T191|SY|363518003|SNOMEDCT_CORE|Renal malignant tumor|Malignant tumor of kidney
C0740457|T191|SYGB|363518003|SNOMEDCT_CORE|Renal malignant tumour|Malignant tumor of kidney
C0740577|T184|IS|9991008|SNOMEDCT_CORE|Acute abdominal pain|Acute abdominal pain
C0740858|T048|SY|66214007|SNOMEDCT_CORE|Harmful substance use|Substance abuse
C0740858|T048|SY|66214007|SNOMEDCT_CORE|Nondependent abuse of substance|Substance abuse
C0740858|T048|PT|66214007|SNOMEDCT_CORE|Substance abuse|Substance abuse
C0740858|T048|FN|66214007|SNOMEDCT_CORE|Substance abuse|Substance abuse
C0741085|T047|PT|419193008|SNOMEDCT_CORE|Ankle ulcer|Ankle ulcer
C0741085|T047|FN|419193008|SNOMEDCT_CORE|Ankle ulcer|Ankle ulcer
C0741151|T047|PT|444569004|SNOMEDCT_CORE|Aneurysm of infrarenal abdominal aorta|Aneurysm of infrarenal abdominal aorta
C0741151|T047|FN|444569004|SNOMEDCT_CORE|Aneurysm of infrarenal abdominal aorta|Aneurysm of infrarenal abdominal aorta
C0741292|T046|PT|427665004|SNOMEDCT_CORE|Paroxysmal atrial flutter|Paroxysmal atrial flutter
C0741292|T046|FN|427665004|SNOMEDCT_CORE|Paroxysmal atrial flutter|Paroxysmal atrial flutter
C0741521|T037|PT|403149008|SNOMEDCT_CORE|Spider bite wound|Spider bite wound
C0741521|T037|FN|403149008|SNOMEDCT_CORE|Spider bite wound|Spider bite wound
C0741521|T037|OF|403149008|SNOMEDCT_CORE|Spider bite wound|Spider bite wound
C0742078|T047|SY|422840005|SNOMEDCT_CORE|Brain mass|Mass lesion of brain
C0742078|T047|PT|422840005|SNOMEDCT_CORE|Mass lesion of brain|Mass lesion of brain
C0742078|T047|FN|422840005|SNOMEDCT_CORE|Mass lesion of brain|Mass lesion of brain
C0742078|T047|SY|422840005|SNOMEDCT_CORE|Space-occupying lesion of brain|Mass lesion of brain
C0742186|T047|PT|54404000|SNOMEDCT_CORE|Cervical radiculopathy|Cervical radiculopathy
C0742186|T047|FN|54404000|SNOMEDCT_CORE|Cervical radiculopathy|Cervical radiculopathy
C0742186|T047|SY|54404000|SNOMEDCT_CORE|Cervical root lesion|Cervical radiculopathy
C0742186|T047|IS|54404000|SNOMEDCT_CORE|Cervical root lesion, NOS|Cervical radiculopathy
C0742186|T047|SY|54404000|SNOMEDCT_CORE|Cervical root neuropathy|Cervical radiculopathy
C0742352|T033|PT|441124000|SNOMEDCT_CORE|Mass of chest wall|Mass of chest wall
C0742352|T033|FN|441124000|SNOMEDCT_CORE|Mass of chest wall|Mass of chest wall
C0742724|T033|PT|116224001|SNOMEDCT_CORE|Complication of procedure|Complication of procedure
C0742724|T033|FN|116224001|SNOMEDCT_CORE|Complication of procedure|Complication of procedure
C0743841|T047|PTGB|416113008|SNOMEDCT_CORE|Disorder characterised by fever|Disorder characterized by fever
C0743841|T047|PT|416113008|SNOMEDCT_CORE|Disorder characterized by fever|Disorder characterized by fever
C0743841|T047|SY|416113008|SNOMEDCT_CORE|Febrile disorder|Disorder characterized by fever
C0743841|T047|FN|416113008|SNOMEDCT_CORE|Febrile disorder|Disorder characterized by fever
C0743841|T047|SY|416113008|SNOMEDCT_CORE|Febrile illness|Disorder characterized by fever
C0743841|T047|SY|416113008|SNOMEDCT_CORE|Febrile syndrome|Disorder characterized by fever
C0743988|T037|PT|447395005|SNOMEDCT_CORE|Closed fracture of fibula|Closed fracture of fibula
C0743988|T037|FN|447395005|SNOMEDCT_CORE|Closed fracture of fibula|Closed fracture of fibula
C0744595|T047|PT|423778009|SNOMEDCT_CORE|Tenosynovitis of hand|Tenosynovitis of hand
C0744595|T047|FN|423778009|SNOMEDCT_CORE|Tenosynovitis of hand|Tenosynovitis of hand
C0745138|T047|PT|443482000|SNOMEDCT_CORE|Hypertensive urgency|Hypertensive urgency
C0745138|T047|FN|443482000|SNOMEDCT_CORE|Hypertensive urgency|Hypertensive urgency
C0745890|T047|OAP|408662006|SNOMEDCT_CORE|Reflex sympathetic dystrophy of lower extremity|Reflex sympathetic dystrophy of lower extremity
C0745890|T047|OAF|408662006|SNOMEDCT_CORE|Reflex sympathetic dystrophy of lower extremity|Reflex sympathetic dystrophy of lower extremity
C0745961|T047|PT|449711005|SNOMEDCT_CORE|Cellulitis of lower leg|Cellulitis of lower leg
C0745961|T047|FN|449711005|SNOMEDCT_CORE|Cellulitis of lower leg|Cellulitis of lower leg
C0745966|T046|PT|449707004|SNOMEDCT_CORE|Edema of lower leg|Edema of lower leg
C0745966|T046|FN|449707004|SNOMEDCT_CORE|Edema of lower leg|Edema of lower leg
C0745966|T046|PTGB|449707004|SNOMEDCT_CORE|Oedema of lower leg|Edema of lower leg
C0746011|T037|PT|426646004|SNOMEDCT_CORE|Compression fracture of lumbar spine|Compression fracture of lumbar spine
C0746011|T037|FN|426646004|SNOMEDCT_CORE|Compression fracture of lumbar spine|Compression fracture of lumbar spine
C0746102|T047|PT|413839001|SNOMEDCT_CORE|Chronic lung disease|Chronic lung disease
C0746102|T047|FN|413839001|SNOMEDCT_CORE|Chronic lung disease|Chronic lung disease
C0746787|T191|PT|363489000|SNOMEDCT_CORE|Malignant tumor of neck|Malignant tumor of neck
C0746787|T191|FN|363489000|SNOMEDCT_CORE|Malignant tumor of neck|Malignant tumor of neck
C0746787|T191|PTGB|363489000|SNOMEDCT_CORE|Malignant tumour of neck|Malignant tumor of neck
C0746883|T047|PT|409089005|SNOMEDCT_CORE|Febrile neutropenia|Febrile neutropenia
C0746883|T047|FN|409089005|SNOMEDCT_CORE|Febrile neutropenia|Febrile neutropenia
C0746883|T047|SYGB|409089005|SNOMEDCT_CORE|Neutropaenic fever|Febrile neutropenia
C0746883|T047|SY|409089005|SNOMEDCT_CORE|Neutropenic fever|Febrile neutropenia
C0746935|T033|PT|129834002|SNOMEDCT_CORE|Noncompliance with medication regimen|Noncompliance with medication regimen
C0746935|T033|FN|129834002|SNOMEDCT_CORE|Noncompliance with medication regimen|Noncompliance with medication regimen
C0746935|T033|SY|129834002|SNOMEDCT_CORE|Noncompliance: medication regimen|Noncompliance with medication regimen
C0747102|T047|PT|111550004|SNOMEDCT_CORE|Ovarian failure|Ovarian failure
C0747102|T047|FN|111550004|SNOMEDCT_CORE|Ovarian failure|Ovarian failure
C0747273|T191|SY|363379000|SNOMEDCT_CORE|CA - Cancer of parotid gland|Malignant tumor of parotid gland
C0747273|T191|SY|363379000|SNOMEDCT_CORE|Cancer of parotid gland|Malignant tumor of parotid gland
C0747273|T191|PT|363379000|SNOMEDCT_CORE|Malignant tumor of parotid gland|Malignant tumor of parotid gland
C0747273|T191|FN|363379000|SNOMEDCT_CORE|Malignant tumor of parotid gland|Malignant tumor of parotid gland
C0747273|T191|PTGB|363379000|SNOMEDCT_CORE|Malignant tumour of parotid gland|Malignant tumor of parotid gland
C0747635|T047|PT|425802001|SNOMEDCT_CORE|Bilateral pleural effusion|Bilateral pleural effusion
C0747635|T047|FN|425802001|SNOMEDCT_CORE|Bilateral pleural effusion|Bilateral pleural effusion
C0747752|T048|PT|445273005|SNOMEDCT_CORE|Polysubstance abuse|Polysubstance abuse
C0747752|T048|FN|445273005|SNOMEDCT_CORE|Polysubstance abuse|Polysubstance abuse
C0748164|T033|PT|445249002|SNOMEDCT_CORE|Multiple nodules of lung|Multiple nodules of lung
C0748164|T033|FN|445249002|SNOMEDCT_CORE|Multiple nodules of lung|Multiple nodules of lung
C0748164|T033|SY|445249002|SNOMEDCT_CORE|Multiple pulmonary nodules|Multiple nodules of lung
C0748226|T047|PT|16644004|SNOMEDCT_CORE|Radial neuropathy|Radial neuropathy
C0748226|T047|FN|16644004|SNOMEDCT_CORE|Radial neuropathy|Radial neuropathy
C0748226|T047|OF|16644004|SNOMEDCT_CORE|Radial neuropathy|Radial neuropathy
C0748315|T047|PT|425369003|SNOMEDCT_CORE|Chronic progressive renal failure|Chronic progressive renal failure
C0748315|T047|FN|425369003|SNOMEDCT_CORE|Chronic progressive renal failure|Chronic progressive renal failure
C0748315|T047|SY|425369003|SNOMEDCT_CORE|Chronic progressive renal insufficiency|Chronic progressive renal failure
C0748390|T046|PT|127154008|SNOMEDCT_CORE|Retroperitoneal lymphadenopathy|Retroperitoneal lymphadenopathy
C0748390|T046|FN|127154008|SNOMEDCT_CORE|Retroperitoneal lymphadenopathy|Retroperitoneal lymphadenopathy
C0748505|T191|PT|443144000|SNOMEDCT_CORE|Metastatic sarcoma|Sarcoma, metastatic
C0748505|T191|FN|443144000|SNOMEDCT_CORE|Metastatic sarcoma|Sarcoma, metastatic
C0748505|T191|PT|372152003|SNOMEDCT_CORE|Sarcoma, metastatic|Sarcoma, metastatic
C0748505|T191|FN|372152003|SNOMEDCT_CORE|Sarcoma, metastatic|Sarcoma, metastatic
C0748712|T046|PT|444605001|SNOMEDCT_CORE|Symptomatic sinus bradycardia|Symptomatic sinus bradycardia
C0748712|T046|FN|444605001|SNOMEDCT_CORE|Symptomatic sinus bradycardia|Symptomatic sinus bradycardia
C0748731|T047|PT|444814009|SNOMEDCT_CORE|Viral sinusitis|Viral sinusitis
C0748731|T047|FN|444814009|SNOMEDCT_CORE|Viral sinusitis|Viral sinusitis
C0749225|T046|PT|371037005|SNOMEDCT_CORE|Systolic dysfunction|Systolic dysfunction
C0749225|T046|FN|371037005|SNOMEDCT_CORE|Systolic dysfunction|Systolic dysfunction
C0750175|T020|FN|414474001|SNOMEDCT_CORE|Incisional hernia of anterior abdominal wall|Ventral incisional hernia
C0750175|T020|SY|414474001|SNOMEDCT_CORE|Incisional hernia of anterior abdominal wall|Ventral incisional hernia
C0750175|T020|PT|414474001|SNOMEDCT_CORE|Ventral incisional hernia|Ventral incisional hernia
C0750197|T047|PT|426525004|SNOMEDCT_CORE|Sustained ventricular tachycardia|Sustained ventricular tachycardia
C0750197|T047|FN|426525004|SNOMEDCT_CORE|Sustained ventricular tachycardia|Sustained ventricular tachycardia
C0750461|T047|PT|423810002|SNOMEDCT_CORE|Tendinitis of wrist|Tendinitis of wrist
C0750461|T047|FN|423810002|SNOMEDCT_CORE|Tendinitis of wrist|Tendinitis of wrist
C0750461|T047|SY|423810002|SNOMEDCT_CORE|Tendonitis of wrist|Tendinitis of wrist
C0750876|T047|SY|2477008|SNOMEDCT_CORE|Superficial phlebitis|Superficial phlebitis
C0750903|T047|PT|35600002|SNOMEDCT_CORE|Strabismic amblyopia|Strabismic amblyopia
C0750903|T047|FN|35600002|SNOMEDCT_CORE|Strabismic amblyopia|Strabismic amblyopia
C0750903|T047|SY|35600002|SNOMEDCT_CORE|Suppression amblyopia|Strabismic amblyopia
C0750929|T019|SY|253185002|SNOMEDCT_CORE|Arnold Chiari type 1|Chiari malformation type I
C0750929|T019|PT|253185002|SNOMEDCT_CORE|Chiari malformation type I|Chiari malformation type I
C0750929|T019|FN|253185002|SNOMEDCT_CORE|Chiari malformation type I|Chiari malformation type I
C0750944|T047|PT|128123007|SNOMEDCT_CORE|Disorder of peripheral autonomic nervous system|Disorder of peripheral autonomic nervous system
C0750944|T047|FN|128123007|SNOMEDCT_CORE|Disorder of peripheral autonomic nervous system|Disorder of peripheral autonomic nervous system
C0750944|T047|IS|15241006|SNOMEDCT_CORE|Disorder of peripheral autonomic nervous system, NOS|Disorder of peripheral autonomic nervous system
C0750955|T047|PT|425596001|SNOMEDCT_CORE|Spastic neurogenic bladder|Spastic neurogenic bladder
C0750955|T047|FN|425596001|SNOMEDCT_CORE|Spastic neurogenic bladder|Spastic neurogenic bladder
C0750955|T047|SY|425596001|SNOMEDCT_CORE|Spastic neuropathic bladder|Spastic neurogenic bladder
C0751186|T184|PT|445511002|SNOMEDCT_CORE|Orthostatic headache|Orthostatic headache
C0751186|T184|FN|445511002|SNOMEDCT_CORE|Orthostatic headache|Orthostatic headache
C0751188|T184|IS|398987004|SNOMEDCT_CORE|PDPH - Post dural puncture headache|PDPH - Post dural puncture headache
C0751188|T184|IS|398987004|SNOMEDCT_CORE|Post dural puncture headache|PDPH - Post dural puncture headache
C0751203|T047|PT|721537005|SNOMEDCT_CORE|Acquired Horner syndrome|Acquired Horner syndrome
C0751203|T047|FN|721537005|SNOMEDCT_CORE|Acquired Horner syndrome|Acquired Horner syndrome
C0751265|T048|SY|1855002|SNOMEDCT_CORE|General learning disability|General learning disability
C0751265|T048|SY|1855002|SNOMEDCT_CORE|Learning disability|General learning disability
C0751340|T047|PT|230684008|SNOMEDCT_CORE|Ocular myasthenia|Ocular myasthenia
C0751340|T047|FN|230684008|SNOMEDCT_CORE|Ocular myasthenia|Ocular myasthenia
C0751362|T047|PT|193042000|SNOMEDCT_CORE|Cataplexy and narcolepsy|Cataplexy and narcolepsy
C0751362|T047|FN|193042000|SNOMEDCT_CORE|Cataplexy and narcolepsy|Cataplexy and narcolepsy
C0751373|T184|SY|16269008|SNOMEDCT_CORE|Paroxysmal nerve pain|Paroxysmal nerve pain
C0751396|T191|PT|443936004|SNOMEDCT_CORE|Oligodendroglioma|Oligodendroglioma
C0751396|T191|FN|443936004|SNOMEDCT_CORE|Oligodendroglioma|Oligodendroglioma
C0751409|T184|PT|249944006|SNOMEDCT_CORE|Monoparesis - arm|Monoparesis - arm
C0751409|T184|FN|249944006|SNOMEDCT_CORE|Monoparesis - arm|Monoparesis - arm
C0751409|T184|SY|249944006|SNOMEDCT_CORE|Weakness of arm|Monoparesis - arm
C0751410|T184|SY|102568007|SNOMEDCT_CORE|Muscle weakness of lower extremity|Paresis of lower extremity
C0751410|T184|PT|102568007|SNOMEDCT_CORE|Paresis of lower extremity|Paresis of lower extremity
C0751410|T184|FN|102568007|SNOMEDCT_CORE|Paresis of lower extremity|Paresis of lower extremity
C0751434|T047|PT|7573000|SNOMEDCT_CORE|Classical phenylketonuria|Classical phenylketonuria
C0751434|T047|FN|7573000|SNOMEDCT_CORE|Classical phenylketonuria|Classical phenylketonuria
C0751434|T047|SY|7573000|SNOMEDCT_CORE|Folling's syndrome|Classical phenylketonuria
C0751434|T047|SYGB|7573000|SNOMEDCT_CORE|Hyperphenylalaninaemia, type I|Classical phenylketonuria
C0751434|T047|SY|7573000|SNOMEDCT_CORE|Hyperphenylalaninemia, type I|Classical phenylketonuria
C0751434|T047|SY|7573000|SNOMEDCT_CORE|Imbecilitus phenylpyruvica|Classical phenylketonuria
C0751434|T047|SY|7573000|SNOMEDCT_CORE|Oligophrenia phenylpyruvica|Classical phenylketonuria
C0751434|T047|SY|7573000|SNOMEDCT_CORE|PAH - Phenylalanine hydroxylase deficiency|Classical phenylketonuria
C0751434|T047|SY|7573000|SNOMEDCT_CORE|PAH deficiency|Classical phenylketonuria
C0751434|T047|SY|7573000|SNOMEDCT_CORE|Phenylalanine hydroxylase deficiency|Classical phenylketonuria
C0751434|T047|SY|7573000|SNOMEDCT_CORE|Phenylketonuria|Classical phenylketonuria
C0751434|T047|IS|7573000|SNOMEDCT_CORE|Phenylketonuria, NOS|Classical phenylketonuria
C0751434|T047|SY|7573000|SNOMEDCT_CORE|Phenylpyruvic oligophrenia|Classical phenylketonuria
C0751434|T047|SY|7573000|SNOMEDCT_CORE|PKU|Classical phenylketonuria
C0751434|T047|SY|7573000|SNOMEDCT_CORE|PKU - Phenylketonuria|Classical phenylketonuria
C0751434|T047|SY|7573000|SNOMEDCT_CORE|PKU1 - Phenylketonuria|Classical phenylketonuria
C0751434|T047|SY|7573000|SNOMEDCT_CORE|Severe phenylalanine hydroxylase deficiency|Classical phenylketonuria
C0751437|T047|SY|51742006|SNOMEDCT_CORE|Anterior pituitary disease|Disorder of anterior pituitary
C0751437|T047|IS|51742006|SNOMEDCT_CORE|Disease of anterior pituitary|Disorder of anterior pituitary
C0751437|T047|OF|51742006|SNOMEDCT_CORE|Disease of anterior pituitary|Disorder of anterior pituitary
C0751437|T047|IS|51742006|SNOMEDCT_CORE|Disease of anterior pituitary, NOS|Disorder of anterior pituitary
C0751437|T047|SY|51742006|SNOMEDCT_CORE|Disorder of adenohypophysis|Disorder of anterior pituitary
C0751437|T047|PT|51742006|SNOMEDCT_CORE|Disorder of anterior pituitary|Disorder of anterior pituitary
C0751437|T047|FN|51742006|SNOMEDCT_CORE|Disorder of anterior pituitary|Disorder of anterior pituitary
C0751437|T047|IS|51742006|SNOMEDCT_CORE|Disorder of anterior pituitary, NOS|Disorder of anterior pituitary
C0751449|T047|SY|42345000|SNOMEDCT_CORE|Acquired polyneuropathy|Acquired polyneuropathy
C0751449|T047|IS|42345000|SNOMEDCT_CORE|Acquired polyneuropathy, NOS|Acquired polyneuropathy
C0751495|T047|SY|29753000|SNOMEDCT_CORE|Focal seizure|Partial seizure
C0751495|T047|SY|29753000|SNOMEDCT_CORE|Local convulsion|Partial seizure
C0751495|T047|SY|29753000|SNOMEDCT_CORE|Local seizure|Partial seizure
C0751495|T047|PT|29753000|SNOMEDCT_CORE|Partial seizure|Partial seizure
C0751495|T047|FN|29753000|SNOMEDCT_CORE|Partial seizure|Partial seizure
C0751495|T047|SY|29753000|SNOMEDCT_CORE|Partial seizures|Partial seizure
C0751495|T047|IS|29753000|SNOMEDCT_CORE|Partial seizures, NOS|Partial seizure
C0751498|T191|PT|285312008|SNOMEDCT_CORE|Carcinoma of sigmoid colon|Carcinoma of sigmoid colon
C0751498|T191|FN|285312008|SNOMEDCT_CORE|Carcinoma of sigmoid colon|Carcinoma of sigmoid colon
C0751540|T047|IS|111496009|SNOMEDCT_CORE|Morvan's disease|Morvan's disease
C0751544|T047|SYGB|15346004|SNOMEDCT_CORE|A - alphalipoproteinaemia neuropathy|Alphalipoproteinemia neuropathy
C0751544|T047|SY|15346004|SNOMEDCT_CORE|A - alphalipoproteinemia neuropathy|Alphalipoproteinemia neuropathy
C0751544|T047|SYGB|15346004|SNOMEDCT_CORE|Alphalipoproteinaemia neuropathy|Alphalipoproteinemia neuropathy
C0751544|T047|SY|15346004|SNOMEDCT_CORE|Alphalipoproteinemia neuropathy|Alphalipoproteinemia neuropathy
C0751560|T191|SY|363393007|SNOMEDCT_CORE|CA - Cancer of tonsil|Malignant tumor of tonsil
C0751560|T191|SY|363393007|SNOMEDCT_CORE|Cancer of tonsil|Malignant tumor of tonsil
C0751560|T191|SY|363393007|SNOMEDCT_CORE|Malignant neoplasm of faucial tonsil|Malignant tumor of tonsil
C0751560|T191|SY|363393007|SNOMEDCT_CORE|Malignant neoplasm of palatine tonsil|Malignant tumor of tonsil
C0751560|T191|SY|363393007|SNOMEDCT_CORE|Malignant tumor of faucial tonsil|Malignant tumor of tonsil
C0751560|T191|SY|363393007|SNOMEDCT_CORE|Malignant tumor of palatine tonsil|Malignant tumor of tonsil
C0751560|T191|PT|363393007|SNOMEDCT_CORE|Malignant tumor of tonsil|Malignant tumor of tonsil
C0751560|T191|FN|363393007|SNOMEDCT_CORE|Malignant tumor of tonsil|Malignant tumor of tonsil
C0751560|T191|SYGB|363393007|SNOMEDCT_CORE|Malignant tumour of faucial tonsil|Malignant tumor of tonsil
C0751560|T191|SYGB|363393007|SNOMEDCT_CORE|Malignant tumour of palatine tonsil|Malignant tumor of tonsil
C0751560|T191|PTGB|363393007|SNOMEDCT_CORE|Malignant tumour of tonsil|Malignant tumor of tonsil
C0751571|T191|SY|363517008|SNOMEDCT_CORE|Malignant tumor of urinary tract|Malignant tumor of urinary tract proper
C0751571|T191|OF|363517008|SNOMEDCT_CORE|Malignant tumor of urinary tract|Malignant tumor of urinary tract proper
C0751571|T191|PT|363517008|SNOMEDCT_CORE|Malignant tumor of urinary tract proper|Malignant tumor of urinary tract proper
C0751571|T191|FN|363517008|SNOMEDCT_CORE|Malignant tumor of urinary tract proper|Malignant tumor of urinary tract proper
C0751571|T191|SYGB|363517008|SNOMEDCT_CORE|Malignant tumour of urinary tract|Malignant tumor of urinary tract proper
C0751571|T191|PTGB|363517008|SNOMEDCT_CORE|Malignant tumour of urinary tract proper|Malignant tumor of urinary tract proper
C0751576|T047|IS|302912005|SNOMEDCT_CORE|Vocal cord paresis|Vocal cord paresis
C0751658|T047|PT|277188003|SNOMEDCT_CORE|Ulnar nerve entrapment|Ulnar nerve entrapment
C0751658|T047|FN|277188003|SNOMEDCT_CORE|Ulnar nerve entrapment|Ulnar nerve entrapment
C0751772|T048|SY|415238003|SNOMEDCT_CORE|Rapid eye movement sleep behavior disorder|REM sleep behavior disorder
C0751772|T048|FN|415238003|SNOMEDCT_CORE|Rapid eye movement sleep behavior disorder|REM sleep behavior disorder
C0751772|T048|SYGB|415238003|SNOMEDCT_CORE|Rapid eye movement sleep behaviour disorder|REM sleep behavior disorder
C0751772|T048|PT|415238003|SNOMEDCT_CORE|REM sleep behavior disorder|REM sleep behavior disorder
C0751772|T048|PTGB|415238003|SNOMEDCT_CORE|REM sleep behaviour disorder|REM sleep behavior disorder
C0751772|T048|SY|415238003|SNOMEDCT_CORE|REM sleep disorder|REM sleep behavior disorder
C0751774|T047|PT|418763003|SNOMEDCT_CORE|Periodic limb movement disorder|Periodic limb movement disorder
C0751774|T047|FN|418763003|SNOMEDCT_CORE|Periodic limb movement disorder|Periodic limb movement disorder
C0751815|T047|PT|705066004|SNOMEDCT_CORE|Dissection of internal carotid artery|Dissection of internal carotid artery
C0751815|T047|FN|705066004|SNOMEDCT_CORE|Dissection of internal carotid artery|Dissection of internal carotid artery
C0751815|T047|OP|705066004|SNOMEDCT_CORE|Internal carotid artery dissection|Dissection of internal carotid artery
C0751815|T047|OF|705066004|SNOMEDCT_CORE|Internal carotid artery dissection|Dissection of internal carotid artery
C0751908|T047|SY|186738001|SNOMEDCT_CORE|Acute epidemic vertigo|Epidemic vertigo
C0751908|T047|SY|186738001|SNOMEDCT_CORE|Acute vestibular neuronitis|Epidemic vertigo
C0751908|T047|SY|186738001|SNOMEDCT_CORE|Epidemic neurolabyrinthitis|Epidemic vertigo
C0751908|T047|PT|186738001|SNOMEDCT_CORE|Epidemic vertigo|Epidemic vertigo
C0751908|T047|FN|186738001|SNOMEDCT_CORE|Epidemic vertigo|Epidemic vertigo
C0751908|T047|SY|186738001|SNOMEDCT_CORE|Vestibular neuritis|Epidemic vertigo
C0751908|T047|SY|186738001|SNOMEDCT_CORE|Vestibular neuronitis|Epidemic vertigo
C0751908|T047|SY|186738001|SNOMEDCT_CORE|Vestibular neuropathy|Epidemic vertigo
C0751922|T047|SY|397828008|SNOMEDCT_CORE|Median nerve palsy|Median neuropathy
C0751922|T047|PT|397828008|SNOMEDCT_CORE|Median neuropathy|Median neuropathy
C0751922|T047|FN|397828008|SNOMEDCT_CORE|Median neuropathy|Median neuropathy
C0751922|T047|OF|397828008|SNOMEDCT_CORE|Median neuropathy|Median neuropathy
C0751925|T047|PT|247390002|SNOMEDCT_CORE|Sciatic nerve palsy|Sciatic nerve palsy
C0751925|T047|FN|247390002|SNOMEDCT_CORE|Sciatic nerve palsy|Sciatic nerve palsy
C0751926|T047|PT|399081005|SNOMEDCT_CORE|Common peroneal neuropathy|Common peroneal neuropathy
C0751926|T047|FN|399081005|SNOMEDCT_CORE|Common peroneal neuropathy|Common peroneal neuropathy
C0751926|T047|SY|399081005|SNOMEDCT_CORE|Lateral popliteal neuropathy|Common peroneal neuropathy
C0751965|T047|SY|425500002|SNOMEDCT_CORE|Multiple sclerosis secondary progressive|Secondary progressive multiple sclerosis
C0751965|T047|PT|425500002|SNOMEDCT_CORE|Secondary progressive multiple sclerosis|Secondary progressive multiple sclerosis
C0751965|T047|FN|425500002|SNOMEDCT_CORE|Secondary progressive multiple sclerosis|Secondary progressive multiple sclerosis
C0751967|T047|SY|426373005|SNOMEDCT_CORE|Multiple sclerosis relapsing remitting|Relapsing remitting multiple sclerosis
C0751967|T047|PT|426373005|SNOMEDCT_CORE|Relapsing remitting multiple sclerosis|Relapsing remitting multiple sclerosis
C0751967|T047|FN|426373005|SNOMEDCT_CORE|Relapsing remitting multiple sclerosis|Relapsing remitting multiple sclerosis
C0752235|T047|IS|23502006|SNOMEDCT_CORE|Bannwarth syndrome|Bannwarth syndrome
C0752235|T047|IS|23502006|SNOMEDCT_CORE|Bannworth's syndrome|Bannwarth syndrome
C0752242|T020|IS|6654000|SNOMEDCT_CORE|Hallux limitus|Hallux limitus
C0752347|T047|SY|80098002|SNOMEDCT_CORE|CLBD - Cortical Lewy body disease|Diffuse Lewy body disease
C0752347|T047|SY|80098002|SNOMEDCT_CORE|Cortical Lewy body disease|Diffuse Lewy body disease
C0752347|T047|SY|80098002|SNOMEDCT_CORE|Dementia of the Lewy body type|Diffuse Lewy body disease
C0752347|T047|PT|80098002|SNOMEDCT_CORE|Diffuse Lewy body disease|Diffuse Lewy body disease
C0752347|T047|FN|80098002|SNOMEDCT_CORE|Diffuse Lewy body disease|Diffuse Lewy body disease
C0752347|T047|SY|80098002|SNOMEDCT_CORE|DLBD - Diffuse Lewy body disease|Diffuse Lewy body disease
C0752347|T047|SY|80098002|SNOMEDCT_CORE|LBD - Lewy body disease|Diffuse Lewy body disease
C0752347|T047|SY|312991009|SNOMEDCT_CORE|Lewy body dementia|Diffuse Lewy body disease
C0752347|T047|SY|80098002|SNOMEDCT_CORE|Lewy body variant of Alzheimer's disease|Diffuse Lewy body disease
C0752347|T047|SY|312991009|SNOMEDCT_CORE|SDLT - senile dementia of Lewy body type|Diffuse Lewy body disease
C0752347|T047|IS|80098002|SNOMEDCT_CORE|SDLT - Senile dementia of the Lewy body type|Diffuse Lewy body disease
C0752347|T047|PT|312991009|SNOMEDCT_CORE|Senile dementia of the Lewy body type|Diffuse Lewy body disease
C0752347|T047|FN|312991009|SNOMEDCT_CORE|Senile dementia of the Lewy body type|Diffuse Lewy body disease
C0795687|T047|SY|71444005|SNOMEDCT_CORE|Cerebral arterial thrombosis|Cerebral thrombosis
C0795687|T047|FN|71444005|SNOMEDCT_CORE|Cerebral arterial thrombosis|Cerebral thrombosis
C0795687|T047|PT|71444005|SNOMEDCT_CORE|Cerebral thrombosis|Cerebral thrombosis
C0795687|T047|SY|71444005|SNOMEDCT_CORE|CT - Cerebral thrombosis|Cerebral thrombosis
C0795687|T047|SY|71444005|SNOMEDCT_CORE|Thrombosis of cerebral arteries|Cerebral thrombosis
C0795690|T019|SY|18735004|SNOMEDCT_CORE|Amniocele|Congenital omphalocele
C0795690|T019|PT|18735004|SNOMEDCT_CORE|Congenital omphalocele|Congenital omphalocele
C0795690|T019|FN|18735004|SNOMEDCT_CORE|Congenital omphalocele|Congenital omphalocele
C0795690|T019|SY|18735004|SNOMEDCT_CORE|Omphalocele|Congenital omphalocele
C0812413|T191|PT|254645002|SNOMEDCT_CORE|Malignant mesothelioma of pleura|Malignant mesothelioma of pleura
C0812413|T191|FN|254645002|SNOMEDCT_CORE|Malignant mesothelioma of pleura|Malignant mesothelioma of pleura
C0812413|T191|SY|254645002|SNOMEDCT_CORE|Malignant pleural mesothelioma|Malignant mesothelioma of pleura
C0812454|T047|IS|359837005|SNOMEDCT_CORE|Ulnar nerve palsy|Ulnar nerve palsy
C0812470|T046|OAS|16863000|SNOMEDCT_CORE|Incomplete abortion|Incomplete abortion
C0812470|T046|OAF|16863000|SNOMEDCT_CORE|Incomplete abortion|Incomplete abortion
C0812470|T046|OF|156072005|SNOMEDCT_CORE|Incomplete miscarriage|Incomplete miscarriage
C0813142|T047|SY|271794005|SNOMEDCT_CORE|Circadian dysregulation|Circadian dysregulation
C0813178|T184|SY|40917007|SNOMEDCT_CORE|Bewilderment|Bewilderment
C0815316|T047|SYGB|49472006|SNOMEDCT_CORE|Megaloblastic anaemia due to cobalamin deficiency|Megaloblastic anemia due to vitamin B>12< deficiency
C0815316|T047|MTH_PTGB|49472006|SNOMEDCT_CORE|Megaloblastic anaemia due to vitamin B<sub>12</sub> deficiency|Megaloblastic anemia due to vitamin B>12< deficiency
C0815316|T047|PTGB|49472006|SNOMEDCT_CORE|Megaloblastic anaemia due to vitamin B>12< deficiency|Megaloblastic anemia due to vitamin B>12< deficiency
C0815316|T047|MTH_PTGB|49472006|SNOMEDCT_CORE|Megaloblastic anaemia due to vitamin B12 deficiency|Megaloblastic anemia due to vitamin B>12< deficiency
C0815316|T047|SY|49472006|SNOMEDCT_CORE|Megaloblastic anemia due to cobalamin deficiency|Megaloblastic anemia due to vitamin B>12< deficiency
C0815316|T047|MTH_FN|49472006|SNOMEDCT_CORE|Megaloblastic anemia due to vitamin B<sub>12</sub> deficiency|Megaloblastic anemia due to vitamin B>12< deficiency
C0815316|T047|MTH_PT|49472006|SNOMEDCT_CORE|Megaloblastic anemia due to vitamin B<sub>12</sub> deficiency|Megaloblastic anemia due to vitamin B>12< deficiency
C0815316|T047|PT|49472006|SNOMEDCT_CORE|Megaloblastic anemia due to vitamin B>12< deficiency|Megaloblastic anemia due to vitamin B>12< deficiency
C0815316|T047|FN|49472006|SNOMEDCT_CORE|Megaloblastic anemia due to vitamin B>12< deficiency|Megaloblastic anemia due to vitamin B>12< deficiency
C0815316|T047|MTH_FN|49472006|SNOMEDCT_CORE|Megaloblastic anemia due to vitamin B12 deficiency|Megaloblastic anemia due to vitamin B>12< deficiency
C0815316|T047|MTH_PT|49472006|SNOMEDCT_CORE|Megaloblastic anemia due to vitamin B12 deficiency|Megaloblastic anemia due to vitamin B>12< deficiency
C0815316|T047|SYGB|49472006|SNOMEDCT_CORE|Vitamin B12-deficient megaloblastic anaemia|Megaloblastic anemia due to vitamin B>12< deficiency
C0815316|T047|SY|49472006|SNOMEDCT_CORE|Vitamin B12-deficient megaloblastic anemia|Megaloblastic anemia due to vitamin B>12< deficiency
C0836911|T033|OAP|37757003|SNOMEDCT_CORE|Communicable disease contact|Communicable disease contact
C0836911|T033|OAF|37757003|SNOMEDCT_CORE|Communicable disease contact|Communicable disease contact
C0836911|T033|OAS|37757003|SNOMEDCT_CORE|Contact - infectious disease|Communicable disease contact
C0836911|T033|IS|37757003|SNOMEDCT_CORE|Contact state, infectious agent|Communicable disease contact
C0836924|T047|SYGB|6631009|SNOMEDCT_CORE|Thrombocythaemia|Thrombocytosis
C0836924|T047|SY|6631009|SNOMEDCT_CORE|Thrombocythemia|Thrombocytosis
C0836924|T047|PT|6631009|SNOMEDCT_CORE|Thrombocytosis|Thrombocytosis
C0836924|T047|FN|6631009|SNOMEDCT_CORE|Thrombocytosis|Thrombocytosis
C0837144|T047|PT|713029000|SNOMEDCT_CORE|Dissection of thoracoabdominal aorta|Dissection of thoracoabdominal aorta
C0837144|T047|FN|713029000|SNOMEDCT_CORE|Dissection of thoracoabdominal aorta|Dissection of thoracoabdominal aorta
C0848377|T037|SY|128069005|SNOMEDCT_CORE|Abdominal injury|Injury of abdomen
C0848377|T037|FN|128069005|SNOMEDCT_CORE|Injury of abdomen|Injury of abdomen
C0848377|T037|PT|128069005|SNOMEDCT_CORE|Injury of abdomen|Injury of abdomen
C0848548|T047|SY|38481006|SNOMEDCT_CORE|Hypertensive nephropathy|Hypertensive renal disease
C0848548|T047|IS|38481006|SNOMEDCT_CORE|Hypertensive nephropathy, NOS|Hypertensive renal disease
C0848548|T047|PT|38481006|SNOMEDCT_CORE|Hypertensive renal disease|Hypertensive renal disease
C0848548|T047|FN|38481006|SNOMEDCT_CORE|Hypertensive renal disease|Hypertensive renal disease
C0848548|T047|IS|38481006|SNOMEDCT_CORE|Hypertensive renal disease, NOS|Hypertensive renal disease
C0848548|T047|SY|38481006|SNOMEDCT_CORE|Renal disease due to hypertension|Hypertensive renal disease
C0848558|T019|PT|416010008|SNOMEDCT_CORE|Hypospadias|Hypospadias
C0848558|T019|FN|416010008|SNOMEDCT_CORE|Hypospadias|Hypospadias
C0849970|T033|SY|224960004|SNOMEDCT_CORE|Feeling tired|Tired
C0849970|T033|PT|224960004|SNOMEDCT_CORE|Tired|Tired
C0849970|T033|FN|224960004|SNOMEDCT_CORE|Tired|Tired
C0849993|T184|PT|444951002|SNOMEDCT_CORE|Fussy infant|Fussy infant
C0849993|T184|FN|444951002|SNOMEDCT_CORE|Fussy infant|Fussy infant
C0849993|T184|SY|444951002|SNOMEDCT_CORE|Unsettled infant|Fussy infant
C0850572|T191|PT|428054006|SNOMEDCT_CORE|Adenomatous polyp of colon|Adenomatous polyp of colon
C0850572|T191|FN|428054006|SNOMEDCT_CORE|Adenomatous polyp of colon|Adenomatous polyp of colon
C0851043|T033|PT|124042003|SNOMEDCT_CORE|Increased lipid|Increased lipid
C0851043|T033|FN|124042003|SNOMEDCT_CORE|Increased lipid|Increased lipid
C0851140|T191|SY|92564006|SNOMEDCT_CORE|Carcinoma in situ of cervix uteri|Carcinoma in situ of uterine cervix
C0851140|T191|PT|92564006|SNOMEDCT_CORE|Carcinoma in situ of uterine cervix|Carcinoma in situ of uterine cervix
C0851140|T191|FN|92564006|SNOMEDCT_CORE|Carcinoma in situ of uterine cervix|Carcinoma in situ of uterine cervix
C0851140|T191|PT|252991009|SNOMEDCT_CORE|Cervical intraepithelial neoplasia grade III with severe dysplasia|Carcinoma in situ of uterine cervix
C0851140|T191|FN|252991009|SNOMEDCT_CORE|Cervical intraepithelial neoplasia grade III with severe dysplasia|Carcinoma in situ of uterine cervix
C0851140|T191|SY|92564006|SNOMEDCT_CORE|CIN 3 - Cervical intraepithelial neoplasia grade 3|Carcinoma in situ of uterine cervix
C0851140|T191|SY|252991009|SNOMEDCT_CORE|CIN III - Cervical intraepithelial neoplasia grade III with severe dysplasia|Carcinoma in situ of uterine cervix
C0851140|T191|SY|92564006|SNOMEDCT_CORE|CIS - Carcinoma in situ of cervix|Carcinoma in situ of uterine cervix
C0851207|T047|PT|609564002|SNOMEDCT_CORE|Pre-existing type 1 diabetes mellitus in pregnancy|Pre-existing type 1 diabetes mellitus in pregnancy
C0851207|T047|FN|609564002|SNOMEDCT_CORE|Pre-existing type 1 diabetes mellitus in pregnancy|Pre-existing type 1 diabetes mellitus in pregnancy
C0851258|T047|SY|17059001|SNOMEDCT_CORE|Beat knee|Prepatellar bursitis
C0851258|T047|PT|17059001|SNOMEDCT_CORE|Prepatellar bursitis|Prepatellar bursitis
C0851258|T047|FN|17059001|SNOMEDCT_CORE|Prepatellar bursitis|Prepatellar bursitis
C0851578|T048|PT|39898005|SNOMEDCT_CORE|Sleep disorder|Sleep disorder
C0851578|T048|FN|39898005|SNOMEDCT_CORE|Sleep disorder|Sleep disorder
C0851578|T048|IS|39898005|SNOMEDCT_CORE|Sleep disorder, NOS|Sleep disorder
C0852036|T047|SY|48194001|SNOMEDCT_CORE|Gestational hypertension|Pregnancy-induced hypertension
C0852036|T047|SY|48194001|SNOMEDCT_CORE|GH - Gestational hypertension|Pregnancy-induced hypertension
C0852036|T047|SY|48194001|SNOMEDCT_CORE|Hypertension induced by pregnancy|Pregnancy-induced hypertension
C0852036|T047|SY|48194001|SNOMEDCT_CORE|PIH - Pregnancy-induced hypertension|Pregnancy-induced hypertension
C0852036|T047|PT|48194001|SNOMEDCT_CORE|Pregnancy-induced hypertension|Pregnancy-induced hypertension
C0852036|T047|FN|48194001|SNOMEDCT_CORE|Pregnancy-induced hypertension|Pregnancy-induced hypertension
C0852036|T047|IS|48194001|SNOMEDCT_CORE|Pregnancy-induced hypertension, NOS|Pregnancy-induced hypertension
C0852949|T047|SY|359557001|SNOMEDCT_CORE|Arterial disease|Disorder of artery
C0852949|T047|SY|39823006|SNOMEDCT_CORE|Arteriopath|Disorder of artery
C0852949|T047|SY|39823006|SNOMEDCT_CORE|Arteriopathy|Disorder of artery
C0852949|T047|IS|359557001|SNOMEDCT_CORE|Disease of artery|Disorder of artery
C0852949|T047|OF|359557001|SNOMEDCT_CORE|Disease of artery|Disorder of artery
C0852949|T047|PT|359557001|SNOMEDCT_CORE|Disorder of artery|Disorder of artery
C0852949|T047|FN|359557001|SNOMEDCT_CORE|Disorder of artery|Disorder of artery
C0853193|T048|SY|371596008|SNOMEDCT_CORE|Bipolar 1 disorder|Bipolar I disorder
C0853193|T048|PT|371596008|SNOMEDCT_CORE|Bipolar I disorder|Bipolar I disorder
C0853193|T048|FN|371596008|SNOMEDCT_CORE|Bipolar I disorder|Bipolar I disorder
C0853225|T033|PT|313341008|SNOMEDCT_CORE|INR raised|INR raised
C0853225|T033|OF|313341008|SNOMEDCT_CORE|INR raised|INR raised
C0853225|T033|SYGB|313341008|SNOMEDCT_CORE|International Normalised Ratio raised|INR raised
C0853225|T033|FN|313341008|SNOMEDCT_CORE|International Normalized Ratio raised|INR raised
C0853225|T033|SY|313341008|SNOMEDCT_CORE|International Normalized Ratio raised|INR raised
C0853225|T033|OF|313341008|SNOMEDCT_CORE|International Normalized Ratio raised|INR raised
C0853697|T033|PT|165517008|SNOMEDCT_CORE|Neutropenia|Neutropenia
C0853697|T033|FN|165517008|SNOMEDCT_CORE|Neutropenia|Neutropenia
C0853697|T033|SY|165517008|SNOMEDCT_CORE|Neutrophil count below reference range|Neutropenia
C0854165|T047|PT|416878008|SNOMEDCT_CORE|Papillary conjunctivitis|Papillary conjunctivitis
C0854165|T047|FN|416878008|SNOMEDCT_CORE|Papillary conjunctivitis|Papillary conjunctivitis
C0854248|T047|SY|430395005|SNOMEDCT_CORE|Gram negative pneumonia|Pneumonia due to Gram negative bacteria
C0854248|T047|SY|430395005|SNOMEDCT_CORE|Pneumonia caused by Gram negative bacteria|Pneumonia due to Gram negative bacteria
C0854248|T047|FN|430395005|SNOMEDCT_CORE|Pneumonia caused by Gram negative bacteria|Pneumonia due to Gram negative bacteria
C0854248|T047|SY|430395005|SNOMEDCT_CORE|Pneumonia caused by Gram-negative bacteria|Pneumonia due to Gram negative bacteria
C0854248|T047|PT|430395005|SNOMEDCT_CORE|Pneumonia due to Gram negative bacteria|Pneumonia due to Gram negative bacteria
C0854248|T047|OF|430395005|SNOMEDCT_CORE|Pneumonia due to Gram negative bacteria|Pneumonia due to Gram negative bacteria
C0854248|T047|SY|430395005|SNOMEDCT_CORE|Pneumonia due to Gram-negative bacteria|Pneumonia due to Gram negative bacteria
C0856169|T047|SY|233845001|SNOMEDCT_CORE|Endothelial dysfunction|Endothelial dysfunction
C0856695|T047|IS|195951007|SNOMEDCT_CORE|Acute exacerbation of chronic bronchitis|Acute exacerbation of chronic bronchitis
C0856747|T047|PT|425963007|SNOMEDCT_CORE|Aneurysm of ascending aorta|Aneurysm of ascending aorta
C0856747|T047|FN|425963007|SNOMEDCT_CORE|Aneurysm of ascending aorta|Aneurysm of ascending aorta
C0857460|T033|SY|6631009|SNOMEDCT_CORE|Increased platelets|Increased platelets
C0858617|T047|PT|315353005|SNOMEDCT_CORE|Posterior subcapsular cataract|Posterior subcapsular cataract
C0858617|T047|FN|315353005|SNOMEDCT_CORE|Posterior subcapsular cataract|Posterior subcapsular cataract
C0858617|T047|SY|315353005|SNOMEDCT_CORE|PSC - posterior subcapsular cataract|Posterior subcapsular cataract
C0859897|T033|PT|134290008|SNOMEDCT_CORE|Vocal cord dysfunction|Vocal cord dysfunction
C0859897|T033|FN|134290008|SNOMEDCT_CORE|Vocal cord dysfunction|Vocal cord dysfunction
C0860096|T033|SY|127364007|SNOMEDCT_CORE|First pregnancy|Primigravida
C0860096|T033|SY|127364007|SNOMEDCT_CORE|Gravida 1|Primigravida
C0860096|T033|FN|127364007|SNOMEDCT_CORE|Primigravida|Primigravida
C0860096|T033|PT|127364007|SNOMEDCT_CORE|Primigravida|Primigravida
C0860096|T033|SY|127364007|SNOMEDCT_CORE|Primip|Primigravida
C0860207|T047|SY|427399008|SNOMEDCT_CORE|Drug induced hepatotoxicity|Drug-induced disorder of liver
C0860207|T047|FN|427399008|SNOMEDCT_CORE|Drug-induced disorder of liver|Drug-induced disorder of liver
C0860207|T047|PT|427399008|SNOMEDCT_CORE|Drug-induced disorder of liver|Drug-induced disorder of liver
C0860594|T191|PT|372158004|SNOMEDCT_CORE|Malignant melanoma, metastatic|Malignant melanoma, metastatic
C0860594|T191|FN|372158004|SNOMEDCT_CORE|Malignant melanoma, metastatic|Malignant melanoma, metastatic
C0860594|T191|PT|443493003|SNOMEDCT_CORE|Metastatic malignant melanoma|Malignant melanoma, metastatic
C0860594|T191|FN|443493003|SNOMEDCT_CORE|Metastatic malignant melanoma|Malignant melanoma, metastatic
C0865424|T048|SY|444613000|SNOMEDCT_CORE|Adult attention deficit disorder|Adult attention deficit hyperactivity disorder
C0865424|T048|PT|444613000|SNOMEDCT_CORE|Adult attention deficit hyperactivity disorder|Adult attention deficit hyperactivity disorder
C0865424|T048|FN|444613000|SNOMEDCT_CORE|Adult attention deficit hyperactivity disorder|Adult attention deficit hyperactivity disorder
C0866713|T020|IS|52012001|SNOMEDCT_CORE|Acquired deformity of the knee|Acquired deformity of the knee
C0869256|T184|SY|413343005|SNOMEDCT_CORE|Mixed incontinence|Mixed urinary incontinence
C0869256|T184|FN|413343005|SNOMEDCT_CORE|Mixed incontinence|Mixed urinary incontinence
C0869256|T184|PT|413343005|SNOMEDCT_CORE|Mixed urinary incontinence|Mixed urinary incontinence
C0870082|T047|OAS|396228006|SNOMEDCT_CORE|HK - Hyperkeratosis|Hyperkeratosis
C0870082|T047|OAP|396228006|SNOMEDCT_CORE|Hyperkeratosis|Hyperkeratosis
C0870082|T047|OAF|396228006|SNOMEDCT_CORE|Hyperkeratosis|Hyperkeratosis
C0870082|T047|OAS|396228006|SNOMEDCT_CORE|Hyperkeratosis of skin|Hyperkeratosis
C0876926|T037|PT|127295002|SNOMEDCT_CORE|Traumatic brain injury|Traumatic brain injury
C0876926|T037|FN|127295002|SNOMEDCT_CORE|Traumatic brain injury|Traumatic brain injury
C0877377|T037|SY|428220001|SNOMEDCT_CORE|Skin tear|Tear of skin
C0877377|T037|PT|428220001|SNOMEDCT_CORE|Tear of skin|Tear of skin
C0877377|T037|FN|428220001|SNOMEDCT_CORE|Traumatic tear of skin|Tear of skin
C0877377|T037|SY|428220001|SNOMEDCT_CORE|Traumatic tear of skin|Tear of skin
C0877425|T033|PT|425810000|SNOMEDCT_CORE|Mass of pancreas|Mass of pancreas
C0877425|T033|FN|425810000|SNOMEDCT_CORE|Mass of pancreas|Mass of pancreas
C0877425|T033|SY|425810000|SNOMEDCT_CORE|Pancreatic mass|Mass of pancreas
C0877792|T046|SY|271794005|SNOMEDCT_CORE|Circadian rhythm sleep-wake disorder|Disorder of sleep-wake cycle
C0877792|T046|PT|271794005|SNOMEDCT_CORE|Disorder of sleep-wake cycle|Disorder of sleep-wake cycle
C0877792|T046|FN|271794005|SNOMEDCT_CORE|Disorder of sleep-wake cycle|Disorder of sleep-wake cycle
C0877792|T046|IS|271794005|SNOMEDCT_CORE|Disorder of sleep-wake schedule|Disorder of sleep-wake cycle
C0877792|T046|IS|271794005|SNOMEDCT_CORE|Disorders of the sleep-wake schedule|Disorder of sleep-wake cycle
C0877792|T046|SY|271794005|SNOMEDCT_CORE|Disturbed nyctohemeral rhythm|Disorder of sleep-wake cycle
C0878521|T047|PTGB|269175006|SNOMEDCT_CORE|Beta thalassaemia trait|Beta thalassemia trait
C0878521|T047|PT|269175006|SNOMEDCT_CORE|Beta thalassemia trait|Beta thalassemia trait
C0878521|T047|FN|269175006|SNOMEDCT_CORE|Beta thalassemia trait|Beta thalassemia trait
C0878544|T047|PT|85898001|SNOMEDCT_CORE|Cardiomyopathy|Cardiomyopathy
C0878544|T047|FN|85898001|SNOMEDCT_CORE|Cardiomyopathy|Cardiomyopathy
C0878544|T047|IS|85898001|SNOMEDCT_CORE|Cardiomyopathy, NOS|Cardiomyopathy
C0878544|T047|SY|85898001|SNOMEDCT_CORE|Myocardiopathy|Cardiomyopathy
C0878544|T047|IS|85898001|SNOMEDCT_CORE|Myocardiopathy, NOS|Cardiomyopathy
C0878697|T047|PTGB|444808002|SNOMEDCT_CORE|Benign localised hyperplasia of prostate|Benign localized hyperplasia of prostate
C0878697|T047|PT|444808002|SNOMEDCT_CORE|Benign localized hyperplasia of prostate|Benign localized hyperplasia of prostate
C0878697|T047|FN|444808002|SNOMEDCT_CORE|Benign localized hyperplasia of prostate|Benign localized hyperplasia of prostate
C0878697|T047|SYGB|444808002|SNOMEDCT_CORE|Localised BPH|Benign localized hyperplasia of prostate
C0878697|T047|SY|444808002|SNOMEDCT_CORE|Localized BPH|Benign localized hyperplasia of prostate
C0878773|T047|SY|786457000|SNOMEDCT_CORE|Bladder instability|Overactive bladder
C0878773|T047|OAS|236633002|SNOMEDCT_CORE|Hyperactive bladder|Overactive bladder
C0878773|T047|SY|786457000|SNOMEDCT_CORE|Hyperactive bladder|Overactive bladder
C0878773|T047|SY|9009001|SNOMEDCT_CORE|Hypertonic bladder|Overactive bladder
C0878773|T047|IS|9009001|SNOMEDCT_CORE|Hypertonicity of bladder|Overactive bladder
C0878773|T047|SY|786457000|SNOMEDCT_CORE|Instability of bladder|Overactive bladder
C0878773|T047|OAS|236633002|SNOMEDCT_CORE|Overactive bladder|Overactive bladder
C0878773|T047|PT|786457000|SNOMEDCT_CORE|Overactive bladder|Overactive bladder
C0878773|T047|FN|786457000|SNOMEDCT_CORE|Overactive bladder|Overactive bladder
C0917799|T047|SY|77692006|SNOMEDCT_CORE|Excessive sleep|Hypersomnia
C0917799|T047|SY|77692006|SNOMEDCT_CORE|Excessive sleepiness|Hypersomnia
C0917799|T047|PT|77692006|SNOMEDCT_CORE|Hypersomnia|Hypersomnia
C0917799|T047|FN|77692006|SNOMEDCT_CORE|Hypersomnia|Hypersomnia
C0917799|T047|SY|77692006|SNOMEDCT_CORE|Hypersomnia|Hypersomnia
C0917799|T047|IS|77692006|SNOMEDCT_CORE|Hypersomnia, NOS|Hypersomnia
C0917799|T047|SY|77692006|SNOMEDCT_CORE|Sleeps too much|Hypersomnia
C0917801|T184|PT|193462001|SNOMEDCT_CORE|Insomnia|Insomnia
C0917801|T184|FN|193462001|SNOMEDCT_CORE|Insomnia|Insomnia
C0917801|T184|SY|193462001|SNOMEDCT_CORE|Sleeplessness|Insomnia
C0917804|T019|SY|234142008|SNOMEDCT_CORE|AVM - Cerebral arteriovenous malformation|Cerebral arteriovenous malformation
C0917804|T019|PT|234142008|SNOMEDCT_CORE|Cerebral arteriovenous malformation|Cerebral arteriovenous malformation
C0917804|T019|FN|234142008|SNOMEDCT_CORE|Cerebral arteriovenous malformation|Cerebral arteriovenous malformation
C0917804|T019|SY|234142008|SNOMEDCT_CORE|Congenital cerebral arteriovenous malformation|Cerebral arteriovenous malformation
C0917996|T047|IS|128609009|SNOMEDCT_CORE|Cerebral aneurysm|Cerebral aneurysm
C0919267|T191|PT|123843001|SNOMEDCT_CORE|Neoplasm of ovary|Neoplasm of ovary
C0919267|T191|FN|123843001|SNOMEDCT_CORE|Neoplasm of ovary|Neoplasm of ovary
C0919267|T191|SY|123843001|SNOMEDCT_CORE|Ovarian tumor|Neoplasm of ovary
C0919267|T191|SYGB|123843001|SNOMEDCT_CORE|Ovarian tumour|Neoplasm of ovary
C0919267|T191|SY|123843001|SNOMEDCT_CORE|Tumor of ovary|Neoplasm of ovary
C0919267|T191|SYGB|123843001|SNOMEDCT_CORE|Tumour of ovary|Neoplasm of ovary
C0920296|T048|PT|52824009|SNOMEDCT_CORE|Developmental reading disorder|Developmental reading disorder
C0920296|T048|FN|52824009|SNOMEDCT_CORE|Developmental reading disorder|Developmental reading disorder
C0920350|T047|IS|21983002|SNOMEDCT_CORE|Autoimmune thyroiditis|Autoimmune thyroiditis
C0920350|T047|PT|66944004|SNOMEDCT_CORE|Autoimmune thyroiditis|Autoimmune thyroiditis
C0920350|T047|FN|66944004|SNOMEDCT_CORE|Autoimmune thyroiditis|Autoimmune thyroiditis
C0920350|T047|IS|66944004|SNOMEDCT_CORE|Autoimmune thyroiditis, NOS|Autoimmune thyroiditis
C0936227|T033|SY|267024001|SNOMEDCT_CORE|Abnormal decrease in weight|Abnormal weight loss
C0936227|T033|FN|267024001|SNOMEDCT_CORE|Abnormal weight loss|Abnormal weight loss
C0936227|T033|PT|267024001|SNOMEDCT_CORE|Abnormal weight loss|Abnormal weight loss
C0947622|T047|SY|235919008|SNOMEDCT_CORE|Cholecystolithiasis|Gallstone
C0947622|T047|SY|235919008|SNOMEDCT_CORE|Gallbladder calculus|Gallstone
C0947622|T047|FN|235919008|SNOMEDCT_CORE|Gallbladder calculus|Gallstone
C0947622|T047|SY|235919008|SNOMEDCT_CORE|Gallbladder stones|Gallstone
C0947622|T047|PT|235919008|SNOMEDCT_CORE|Gallstone|Gallstone
C0947622|T047|SY|235919008|SNOMEDCT_CORE|Gallstones|Gallstone
C0947622|T047|SY|235919008|SNOMEDCT_CORE|GS - Gallstone|Gallstone
C0948008|T047|PTGB|422504002|SNOMEDCT_CORE|Ischaemic stroke|Ischemic stroke
C0948008|T047|PT|422504002|SNOMEDCT_CORE|Ischemic stroke|Ischemic stroke
C0948008|T047|FN|422504002|SNOMEDCT_CORE|Ischemic stroke|Ischemic stroke
C0948089|T047|SY|394659003|SNOMEDCT_CORE|ACS - Acute coronary syndrome|Acute coronary syndrome
C0948089|T047|PT|394659003|SNOMEDCT_CORE|Acute coronary syndrome|Acute coronary syndrome
C0948089|T047|FN|394659003|SNOMEDCT_CORE|Acute coronary syndrome|Acute coronary syndrome
C0948187|T047|PT|95434006|SNOMEDCT_CORE|Tracheomalacia|Tracheomalacia
C0948187|T047|FN|95434006|SNOMEDCT_CORE|Tracheomalacia|Tracheomalacia
C0948657|T033|SY|432519008|SNOMEDCT_CORE|Elevated cancer antigen 125|Increased cancer antigen 125
C0948657|T033|PT|432519008|SNOMEDCT_CORE|Increased cancer antigen 125|Increased cancer antigen 125
C0948657|T033|FN|432519008|SNOMEDCT_CORE|Increased cancer antigen 125|Increased cancer antigen 125
C0948657|T033|SY|432519008|SNOMEDCT_CORE|Raised cancer antigen 125|Increased cancer antigen 125
C0948672|T047|SYGB|402843003|SNOMEDCT_CORE|Acquired venous haemangioma|Venous lake
C0948672|T047|SY|402843003|SNOMEDCT_CORE|Acquired venous hemangioma|Venous lake
C0948672|T047|PT|402843003|SNOMEDCT_CORE|Venous lake|Venous lake
C0948672|T047|FN|402843003|SNOMEDCT_CORE|Venous lake|Venous lake
C0948824|T047|PTGB|413532003|SNOMEDCT_CORE|Anaemia due to blood loss|Anemia due to blood loss
C0948824|T047|PT|413532003|SNOMEDCT_CORE|Anemia due to blood loss|Anemia due to blood loss
C0948824|T047|FN|413532003|SNOMEDCT_CORE|Anemia due to blood loss|Anemia due to blood loss
C0948968|T191|SY|307651005|SNOMEDCT_CORE|Osteomyelofibrosis|Osteomyelofibrosis
C0949690|T047|PT|371082009|SNOMEDCT_CORE|Arthritis of spine|Arthritis of spine
C0949690|T047|FN|371082009|SNOMEDCT_CORE|Arthritis of spine|Arthritis of spine
C0949690|T047|SY|371082009|SNOMEDCT_CORE|Inflammatory spondylopathy|Arthritis of spine
C0949690|T047|IS|371082009|SNOMEDCT_CORE|Spondylarthritis|Arthritis of spine
C0949690|T047|IS|371082009|SNOMEDCT_CORE|Spondyloarthritis|Arthritis of spine
C0949691|T047|FN|372109003|SNOMEDCT_CORE|Disorder of joint of spine|Disorder of joint of spine
C0949691|T047|PT|372109003|SNOMEDCT_CORE|Disorder of joint of spine|Disorder of joint of spine
C0949691|T047|SY|8847002|SNOMEDCT_CORE|Spondarthropathy|Disorder of joint of spine
C0949691|T047|SY|8847002|SNOMEDCT_CORE|Spondylarthrosis|Disorder of joint of spine
C0949691|T047|IS|8847002|SNOMEDCT_CORE|Spondylarthrosis, NOS|Disorder of joint of spine
C0949691|T047|IS|372109003|SNOMEDCT_CORE|Spondyloarthropathy|Disorder of joint of spine
C0949691|T047|SY|372109003|SNOMEDCT_CORE|Spondyloarthropathy|Disorder of joint of spine
C0973461|T047|PT|20301004|SNOMEDCT_CORE|Dysphasia|Dysphasia
C0973461|T047|FN|20301004|SNOMEDCT_CORE|Dysphasia|Dysphasia
C1096063|T047|SY|445355009|SNOMEDCT_CORE|Intractable epilepsy|Refractory epilepsy
C1096063|T047|PT|445355009|SNOMEDCT_CORE|Refractory epilepsy|Refractory epilepsy
C1096063|T047|FN|445355009|SNOMEDCT_CORE|Refractory epilepsy|Refractory epilepsy
C1096519|T037|PT|444356002|SNOMEDCT_CORE|Exposure to Human immunodeficiency virus|Exposure to Human immunodeficiency virus
C1096519|T037|FN|444356002|SNOMEDCT_CORE|Exposure to Human immunodeficiency virus|Exposure to Human immunodeficiency virus
C1096624|T033|SY|443503005|SNOMEDCT_CORE|Periumbilical abdominal pain|Periumbilical pain
C1096624|T033|PT|443503005|SNOMEDCT_CORE|Periumbilical pain|Periumbilical pain
C1096624|T033|FN|443503005|SNOMEDCT_CORE|Periumbilical pain|Periumbilical pain
C1112213|T047|PT|433237003|SNOMEDCT_CORE|Cholestasis in newborn|Cholestasis in newborn
C1112213|T047|FN|433237003|SNOMEDCT_CORE|Cholestasis in newborn|Cholestasis in newborn
C1112213|T047|SY|433237003|SNOMEDCT_CORE|Neonatal cholestasis|Cholestasis in newborn
C1134719|T191|FN|408643008|SNOMEDCT_CORE|Infiltrating duct carcinoma of breast|Infiltrating duct carcinoma of breast
C1134719|T191|PT|408643008|SNOMEDCT_CORE|Infiltrating duct carcinoma of breast|Infiltrating duct carcinoma of breast
C1134719|T191|SY|408643008|SNOMEDCT_CORE|Infiltrating ductal carcinoma of breast|Infiltrating duct carcinoma of breast
C1134719|T191|SY|408643008|SNOMEDCT_CORE|Invasive duct carcinoma of breast|Infiltrating duct carcinoma of breast
C1134719|T191|SY|408643008|SNOMEDCT_CORE|Invasive ductal carcinoma of breast|Infiltrating duct carcinoma of breast
C1135191|T047|PT|417996009|SNOMEDCT_CORE|Systolic heart failure|Systolic heart failure
C1135191|T047|FN|417996009|SNOMEDCT_CORE|Systolic heart failure|Systolic heart failure
C1135194|T047|PT|441481004|SNOMEDCT_CORE|Chronic systolic heart failure|Chronic systolic heart failure
C1135194|T047|FN|441481004|SNOMEDCT_CORE|Chronic systolic heart failure|Chronic systolic heart failure
C1135196|T047|PT|418304008|SNOMEDCT_CORE|Diastolic heart failure|Diastolic heart failure
C1135196|T047|FN|418304008|SNOMEDCT_CORE|Diastolic heart failure|Diastolic heart failure
C1135812|T037|SY|263029007|SNOMEDCT_CORE|Dislocated patella|Dislocation of patellofemoral joint
C1135812|T037|PT|263029007|SNOMEDCT_CORE|Dislocation of patellofemoral joint|Dislocation of patellofemoral joint
C1135812|T037|FN|263029007|SNOMEDCT_CORE|Dislocation of patellofemoral joint|Dislocation of patellofemoral joint
C1136085|T191|SY|109983007|SNOMEDCT_CORE|Monoclonal gammopathy|Monoclonal gammopathy
C1136085|T191|PT|109983007|SNOMEDCT_CORE|Monoclonal gammopathy|Monoclonal gammopathy
C1136085|T191|FN|109983007|SNOMEDCT_CORE|Monoclonal gammopathy|Monoclonal gammopathy
C1136085|T191|SYGB|109983007|SNOMEDCT_CORE|Monoclonal paraproteinaemia|Monoclonal gammopathy
C1136085|T191|SY|109983007|SNOMEDCT_CORE|Monoclonal paraproteinemia|Monoclonal gammopathy
C1136179|T190|PT|122481008|SNOMEDCT_CORE|Hammer toe|Hammer toe
C1136179|T190|FN|122481008|SNOMEDCT_CORE|Hammer toe|Hammer toe
C1140680|T191|SY|363443007|SNOMEDCT_CORE|CA - Cancer of ovary|Malignant tumor of ovary
C1140680|T191|SY|363443007|SNOMEDCT_CORE|Cancer of ovary|Malignant tumor of ovary
C1140680|T191|IS|93934004|SNOMEDCT_CORE|Malignant neoplasm of ovary|Malignant tumor of ovary
C1140680|T191|PT|363443007|SNOMEDCT_CORE|Malignant tumor of ovary|Malignant tumor of ovary
C1140680|T191|FN|363443007|SNOMEDCT_CORE|Malignant tumor of ovary|Malignant tumor of ovary
C1140680|T191|PTGB|363443007|SNOMEDCT_CORE|Malignant tumour of ovary|Malignant tumor of ovary
C1140680|T191|IS|363443007|SNOMEDCT_CORE|Ovarian Ca|Malignant tumor of ovary
C1140680|T191|SY|363443007|SNOMEDCT_CORE|Ovarian cancer|Malignant tumor of ovary
C1140716|T046|PT|126944002|SNOMEDCT_CORE|Brain damage due to hypoxia|Brain damage due to hypoxia
C1140716|T046|FN|126944002|SNOMEDCT_CORE|Brain disorder resulting from a period of impaired oxygen delivery to the brain|Brain damage due to hypoxia
C1140716|T046|SY|126944002|SNOMEDCT_CORE|Brain disorder resulting from a period of impaired oxygen delivery to the brain|Brain damage due to hypoxia
C1140716|T046|SY|126944002|SNOMEDCT_CORE|Hypoxic brain damage|Brain damage due to hypoxia
C1140716|T046|IS|126944002|SNOMEDCT_CORE|Hypoxic-ischaemic brain injury|Brain damage due to hypoxia
C1140716|T046|IS|126944002|SNOMEDCT_CORE|Hypoxic-ischemic brain injury|Brain damage due to hypoxia
C1142430|T048|SY|191714002|SNOMEDCT_CORE|Psychogenic seizures|Psychogenic seizures
C1142491|T191|PT|314515006|SNOMEDCT_CORE|Papilloma of eyelid|Papilloma of eyelid
C1142491|T191|FN|314515006|SNOMEDCT_CORE|Papilloma of eyelid|Papilloma of eyelid
C1145628|T047|PT|15241006|SNOMEDCT_CORE|Disorder of autonomic nervous system|Disorder of autonomic nervous system
C1145628|T047|FN|15241006|SNOMEDCT_CORE|Disorder of autonomic nervous system|Disorder of autonomic nervous system
C1145628|T047|IS|15241006|SNOMEDCT_CORE|Disorder of autonomic nervous system, NOS|Disorder of autonomic nervous system
C1145628|T047|SY|15241006|SNOMEDCT_CORE|Disorder of vegetative system|Disorder of autonomic nervous system
C1145628|T047|IS|15241006|SNOMEDCT_CORE|Disorder of vegetative system, NOS|Disorder of autonomic nervous system
C1145628|T047|SY|15241006|SNOMEDCT_CORE|Disorders of autonomic nervous system|Disorder of autonomic nervous system
C1145670|T047|PT|409622000|SNOMEDCT_CORE|Respiratory failure|Respiratory failure
C1145670|T047|FN|409622000|SNOMEDCT_CORE|Respiratory failure|Respiratory failure
C1153706|T191|PT|123845008|SNOMEDCT_CORE|Adenocarcinoma of endometrium|Adenocarcinoma of endometrium
C1153706|T191|FN|123845008|SNOMEDCT_CORE|Adenocarcinoma of endometrium|Adenocarcinoma of endometrium
C1153706|T191|SY|123845008|SNOMEDCT_CORE|Endometrial adenocarcinoma|Adenocarcinoma of endometrium
C1168250|T047|PT|414581006|SNOMEDCT_CORE|Laryngopharyngeal reflux|Laryngopharyngeal reflux
C1168250|T047|FN|414581006|SNOMEDCT_CORE|Laryngopharyngeal reflux|Laryngopharyngeal reflux
C1253936|T046|SY|387637008|SNOMEDCT_CORE|Effusion into joint|Effusion of joint
C1253936|T046|PT|387637008|SNOMEDCT_CORE|Effusion of joint|Effusion of joint
C1253936|T046|FN|387637008|SNOMEDCT_CORE|Effusion of joint|Effusion of joint
C1253936|T046|SY|387637008|SNOMEDCT_CORE|Hydrarthrosis|Effusion of joint
C1253936|T046|SY|387637008|SNOMEDCT_CORE|Joint effusion|Effusion of joint
C1257843|T047|OAS|397683000|SNOMEDCT_CORE|PMC - Pseudomembranous colitis|PMC - Pseudomembranous colitis
C1257843|T047|OAS|397683000|SNOMEDCT_CORE|Pseudomembranous colitis|PMC - Pseudomembranous colitis
C1258215|T047|IS|81060008|SNOMEDCT_CORE|Ileus|Ileus
C1258215|T047|IS|81060008|SNOMEDCT_CORE|Ileus, NOS|Ileus
C1258666|T047|SY|71307009|SNOMEDCT_CORE|Benign cystic mucinous tumor|Ganglion cyst
C1258666|T047|IS|71307009|SNOMEDCT_CORE|Benign cystic mucinous tumor, NOS|Ganglion cyst
C1258666|T047|SYGB|71307009|SNOMEDCT_CORE|Benign cystic mucinous tumour|Ganglion cyst
C1258666|T047|SY|71307009|SNOMEDCT_CORE|Ganglion|Ganglion cyst
C1258666|T047|PT|445008009|SNOMEDCT_CORE|Ganglion cyst|Ganglion cyst
C1258666|T047|PT|71307009|SNOMEDCT_CORE|Ganglion cyst|Ganglion cyst
C1258666|T047|FN|71307009|SNOMEDCT_CORE|Ganglion cyst|Ganglion cyst
C1258666|T047|FN|445008009|SNOMEDCT_CORE|Ganglion cyst|Ganglion cyst
C1258666|T047|IS|71307009|SNOMEDCT_CORE|Ganglion, NOS|Ganglion cyst
C1258666|T047|SY|78435003|SNOMEDCT_CORE|Mucous cyst of skin|Ganglion cyst
C1258666|T047|SY|71307009|SNOMEDCT_CORE|Myxoid cyst|Ganglion cyst
C1260873|T047|SY|8722008|SNOMEDCT_CORE|Aortic valve disease|Aortic valve disorder
C1260873|T047|PT|8722008|SNOMEDCT_CORE|Aortic valve disorder|Aortic valve disorder
C1260873|T047|FN|8722008|SNOMEDCT_CORE|Aortic valve disorder|Aortic valve disorder
C1260873|T047|IS|8722008|SNOMEDCT_CORE|Aortic valve disorder, NOS|Aortic valve disorder
C1260873|T047|SY|8722008|SNOMEDCT_CORE|AVD - Aortic valve disease|Aortic valve disorder
C1260880|T184|SY|64531003|SNOMEDCT_CORE|Discharge from nose|Nasal discharge
C1260880|T184|SY|64531003|SNOMEDCT_CORE|Nasal catarrh|Nasal discharge
C1260880|T184|PT|64531003|SNOMEDCT_CORE|Nasal discharge|Nasal discharge
C1260880|T184|FN|64531003|SNOMEDCT_CORE|Nasal discharge|Nasal discharge
C1260880|T184|OF|64531003|SNOMEDCT_CORE|Nasal discharge|Nasal discharge
C1260880|T184|SY|64531003|SNOMEDCT_CORE|Rhinorrhea|Nasal discharge
C1260880|T184|SYGB|64531003|SNOMEDCT_CORE|Rhinorrhoea|Nasal discharge
C1260883|T047|SY|91335003|SNOMEDCT_CORE|Endocardial thrombosis|Mural thrombus of heart
C1260883|T047|SY|91335003|SNOMEDCT_CORE|Mural thrombosis|Mural thrombus of heart
C1260883|T047|PT|91335003|SNOMEDCT_CORE|Mural thrombus of heart|Mural thrombus of heart
C1260883|T047|FN|91335003|SNOMEDCT_CORE|Mural thrombus of heart|Mural thrombus of heart
C1260915|T047|PT|186903006|SNOMEDCT_CORE|Late latent syphilis|Late latent syphilis
C1260915|T047|FN|186903006|SNOMEDCT_CORE|Late latent syphilis|Late latent syphilis
C1261120|T047|SY|195957006|SNOMEDCT_CORE|Bullous emphysema|Chronic bullous emphysema
C1261120|T047|PT|195957006|SNOMEDCT_CORE|Chronic bullous emphysema|Chronic bullous emphysema
C1261120|T047|FN|195957006|SNOMEDCT_CORE|Chronic bullous emphysema|Chronic bullous emphysema
C1261262|T047|IS|48194001|SNOMEDCT_CORE|Hypertension complicating pregnancy, childbirth AND/OR puerperium|Hypertension complicating pregnancy, childbirth AND/OR puerperium
C1261262|T047|IS|48194001|SNOMEDCT_CORE|Unspecified hypertension complicating pregnancy, childbirth or puerperium|Hypertension complicating pregnancy, childbirth AND/OR puerperium
C1261276|T019|SY|268242003|SNOMEDCT_CORE|Congenital subluxation of hip, unilateral|Congenital unilateral subluxation of hip
C1261276|T019|OF|268242003|SNOMEDCT_CORE|Congenital subluxation of hip, unilateral|Congenital unilateral subluxation of hip
C1261276|T019|PT|268242003|SNOMEDCT_CORE|Congenital unilateral subluxation of hip|Congenital unilateral subluxation of hip
C1261276|T019|FN|268242003|SNOMEDCT_CORE|Congenital unilateral subluxation of hip|Congenital unilateral subluxation of hip
C1261281|T046|SY|58797008|SNOMEDCT_CORE|Complication of transplanted kidney|Disorder of transplanted kidney
C1261281|T046|FN|58797008|SNOMEDCT_CORE|Complication of transplanted kidney|Disorder of transplanted kidney
C1261281|T046|PT|58797008|SNOMEDCT_CORE|Disorder of transplanted kidney|Disorder of transplanted kidney
C1261282|T046|PT|33167004|SNOMEDCT_CORE|Complication of transplanted liver|Complication of transplanted liver
C1261282|T046|FN|33167004|SNOMEDCT_CORE|Complication of transplanted liver|Complication of transplanted liver
C1261325|T033|PT|429740004|SNOMEDCT_CORE|Family history of breast cancer|Family history of breast cancer
C1261325|T033|SY|429740004|SNOMEDCT_CORE|Family history of malignant neoplasm of breast|Family history of breast cancer
C1261325|T033|FN|429740004|SNOMEDCT_CORE|Family history of malignant neoplasm of breast|Family history of breast cancer
C1261327|T033|PT|160377001|SNOMEDCT_CORE|Family history of asthma|Family history of asthma
C1261327|T033|SY|160377001|SNOMEDCT_CORE|Family history: Asthma|Family history of asthma
C1261327|T033|OF|160377001|SNOMEDCT_CORE|Family history: Asthma|Family history of asthma
C1261327|T033|FN|160377001|SNOMEDCT_CORE|Family history: Asthma|Family history of asthma
C1261327|T033|SY|160377001|SNOMEDCT_CORE|FH: Asthma|Family history of asthma
C1261329|T033|SY|160417009|SNOMEDCT_CORE|Family history: Congenital anomaly|FH: Congenital anomaly
C1261329|T033|OF|160417009|SNOMEDCT_CORE|Family history: Congenital anomaly|FH: Congenital anomaly
C1261329|T033|FN|160417009|SNOMEDCT_CORE|Family history: Congenital anomaly|FH: Congenital anomaly
C1261329|T033|PT|160417009|SNOMEDCT_CORE|FH: Congenital anomaly|FH: Congenital anomaly
C1261331|T047|PT|267612009|SNOMEDCT_CORE|Degeneration of macula due to cyst, hole or pseudohole|Degeneration of macula due to cyst, hole or pseudohole
C1261331|T047|FN|267612009|SNOMEDCT_CORE|Degeneration of macula due to cyst, hole or pseudohole|Degeneration of macula due to cyst, hole or pseudohole
C1261367|T033|SY|275104002|SNOMEDCT_CORE|Family history of CVA|Family history of stroke
C1261367|T033|PT|275104002|SNOMEDCT_CORE|Family history of stroke|Family history of stroke
C1261367|T033|OF|275104002|SNOMEDCT_CORE|Family history of stroke|Family history of stroke
C1261367|T033|FN|275104002|SNOMEDCT_CORE|Family history of stroke|Family history of stroke
C1261367|T033|SY|275104002|SNOMEDCT_CORE|FH: CVA|Family history of stroke
C1261367|T033|SY|275104002|SNOMEDCT_CORE|FH: Stroke|Family history of stroke
C1261368|T033|SY|275134007|SNOMEDCT_CORE|Family history: Arthritis|FH: Arthritis
C1261368|T033|OF|275134007|SNOMEDCT_CORE|Family history: Arthritis|FH: Arthritis
C1261368|T033|FN|275134007|SNOMEDCT_CORE|Family history: Arthritis|FH: Arthritis
C1261368|T033|PT|275134007|SNOMEDCT_CORE|FH: Arthritis|FH: Arthritis
C1261473|T191|PT|424413001|SNOMEDCT_CORE|Sarcoma|Sarcoma
C1261473|T191|FN|424413001|SNOMEDCT_CORE|Sarcoma|Sarcoma
C1261562|T047|OAS|61033006|SNOMEDCT_CORE|Detrusor dyssynergia|Idiopathic detrusor overactivity
C1261562|T047|SY|786496006|SNOMEDCT_CORE|Detrusor dyssynergia|Idiopathic detrusor overactivity
C1261562|T047|OAS|61033006|SNOMEDCT_CORE|Detrusor instability|Idiopathic detrusor overactivity
C1261562|T047|SY|786496006|SNOMEDCT_CORE|Detrusor instability|Idiopathic detrusor overactivity
C1261562|T047|OAP|61033006|SNOMEDCT_CORE|Detrusor instability of bladder|Idiopathic detrusor overactivity
C1261562|T047|SY|786496006|SNOMEDCT_CORE|Detrusor instability of bladder|Idiopathic detrusor overactivity
C1261562|T047|OAF|61033006|SNOMEDCT_CORE|Detrusor instability of bladder|Idiopathic detrusor overactivity
C1261562|T047|SY|786496006|SNOMEDCT_CORE|DI - detrusor instability|Idiopathic detrusor overactivity
C1261562|T047|OAS|61033006|SNOMEDCT_CORE|DI - Detrusor instability|Idiopathic detrusor overactivity
C1261562|T047|PT|786496006|SNOMEDCT_CORE|Idiopathic detrusor overactivity|Idiopathic detrusor overactivity
C1261562|T047|FN|786496006|SNOMEDCT_CORE|Idiopathic detrusor overactivity|Idiopathic detrusor overactivity
C1262206|T047|PT|423849004|SNOMEDCT_CORE|Iliotibial band friction syndrome|Iliotibial band friction syndrome
C1262206|T047|FN|423849004|SNOMEDCT_CORE|Iliotibial band friction syndrome|Iliotibial band friction syndrome
C1262206|T047|SY|423849004|SNOMEDCT_CORE|Iliotibial band syndrome|Iliotibial band friction syndrome
C1262477|T033|PT|262285001|SNOMEDCT_CORE|Weight decreased|Weight decreased
C1262477|T033|OF|262285001|SNOMEDCT_CORE|Weight decreased|Weight decreased
C1262477|T033|FN|262285001|SNOMEDCT_CORE|Weight decreased|Weight decreased
C1263682|T191|PT|126789008|SNOMEDCT_CORE|Neoplasm of submaxillary gland|Neoplasm of submaxillary gland
C1263682|T191|FN|126789008|SNOMEDCT_CORE|Neoplasm of submaxillary gland|Neoplasm of submaxillary gland
C1263682|T191|SY|126789008|SNOMEDCT_CORE|Tumor of submandibular gland|Neoplasm of submaxillary gland
C1263682|T191|SYGB|126789008|SNOMEDCT_CORE|Tumour of submandibular gland|Neoplasm of submaxillary gland
C1263764|T047|PT|106002000|SNOMEDCT_CORE|Disorder associated with menstruation AND/OR menopause|Disorder associated with menstruation AND/OR menopause
C1263764|T047|FN|106002000|SNOMEDCT_CORE|Disorder associated with menstruation AND/OR menopause|Disorder associated with menstruation AND/OR menopause
C1263820|T046|PT|106008001|SNOMEDCT_CORE|Delivery AND/OR maternal condition affecting management|Delivery AND/OR maternal condition affecting management
C1263820|T046|FN|106008001|SNOMEDCT_CORE|Delivery AND/OR maternal condition affecting management|Delivery AND/OR maternal condition affecting management
C1263821|T047|OAP|111443000|SNOMEDCT_CORE|Congenital OR acquired abnormality of cervix affecting pregnancy|Congenital OR acquired abnormality of cervix affecting pregnancy
C1263821|T047|OAF|111443000|SNOMEDCT_CORE|Congenital OR acquired abnormality of cervix affecting pregnancy|Congenital OR acquired abnormality of cervix affecting pregnancy
C1263846|T048|SY|406506008|SNOMEDCT_CORE|ADHD - Attention deficit disorder with hyperactivity|Attention deficit hyperactivity disorder
C1263846|T048|PT|406506008|SNOMEDCT_CORE|Attention deficit hyperactivity disorder|Attention deficit hyperactivity disorder
C1263846|T048|FN|406506008|SNOMEDCT_CORE|Attention deficit hyperactivity disorder|Attention deficit hyperactivity disorder
C1263846|T048|SY|406506008|SNOMEDCT_CORE|Attention deficit hyperkinetic disorder|Attention deficit hyperactivity disorder
C1263846|T048|SY|406506008|SNOMEDCT_CORE|Hyperkinetic disorder|Attention deficit hyperactivity disorder
C1263846|T048|SY|406506008|SNOMEDCT_CORE|Hyperkinetic syndrome|Attention deficit hyperactivity disorder
C1263846|T048|SY|406506008|SNOMEDCT_CORE|Overactive child syndrome|Attention deficit hyperactivity disorder
C1263853|T047|PT|116288000|SNOMEDCT_CORE|Paralytic stroke|Paralytic stroke
C1263853|T047|FN|116288000|SNOMEDCT_CORE|Paralytic stroke|Paralytic stroke
C1263855|T047|PT|128196005|SNOMEDCT_CORE|Lumbar radiculopathy|Lumbar radiculopathy
C1263855|T047|FN|128196005|SNOMEDCT_CORE|Lumbar radiculopathy|Lumbar radiculopathy
C1263855|T047|IS|2415007|SNOMEDCT_CORE|Lumbar radiculopathy, NOS|Lumbar radiculopathy
C1263878|T033|PT|126946000|SNOMEDCT_CORE|Excessive cerumen in ear canal|Excessive cerumen in ear canal
C1263878|T033|FN|126946000|SNOMEDCT_CORE|Excessive cerumen in ear canal|Excessive cerumen in ear canal
C1264038|T037|PT|109957002|SNOMEDCT_CORE|Drug-induced purpura|Drug-induced purpura
C1264038|T037|FN|109957002|SNOMEDCT_CORE|Drug-induced purpura|Drug-induced purpura
C1264190|T191|SY|109972003|SNOMEDCT_CORE|Follicular lymphoma grade 3|Follicular non-Hodgkin's lymphoma, large cell
C1264190|T191|SY|109972003|SNOMEDCT_CORE|Follicular non-Hodgkin lymphoma, large cell|Follicular non-Hodgkin's lymphoma, large cell
C1264190|T191|OAS|277641001|SNOMEDCT_CORE|Follicular non-Hodgkin's large cell lymphoma|Follicular non-Hodgkin's lymphoma, large cell
C1264190|T191|SY|109972003|SNOMEDCT_CORE|Follicular non-Hodgkin's lymphoma, large cell|Follicular non-Hodgkin's lymphoma, large cell
C1264190|T191|PT|109972003|SNOMEDCT_CORE|Follicular non-Hodgkin's lymphoma, large cell|Follicular non-Hodgkin's lymphoma, large cell
C1264190|T191|FN|109972003|SNOMEDCT_CORE|Follicular non-Hodgkin's lymphoma, large cell|Follicular non-Hodgkin's lymphoma, large cell
C1264240|T037|PTGB|111593004|SNOMEDCT_CORE|Closed fracture of vault of skull with intracranial haemorrhage|Closed fracture of vault of skull with intracranial hemorrhage
C1264240|T037|PT|111593004|SNOMEDCT_CORE|Closed fracture of vault of skull with intracranial hemorrhage|Closed fracture of vault of skull with intracranial hemorrhage
C1264240|T037|OF|111593004|SNOMEDCT_CORE|Closed fracture of vault of skull with intracranial hemorrhage|Closed fracture of vault of skull with intracranial hemorrhage
C1264240|T037|SY|111593004|SNOMEDCT_CORE|Intracranial hemorrhage co-occurrent and due to closed fracture of vault of skull|Closed fracture of vault of skull with intracranial hemorrhage
C1264240|T037|FN|111593004|SNOMEDCT_CORE|Intracranial hemorrhage co-occurrent and due to closed fracture of vault of skull|Closed fracture of vault of skull with intracranial hemorrhage
C1264284|T037|PT|111653006|SNOMEDCT_CORE|Sprain of sacroiliac region|Sprain of sacroiliac region
C1264284|T037|FN|111653006|SNOMEDCT_CORE|Sprain of sacroiliac region|Sprain of sacroiliac region
C1264517|T046|PT|269406001|SNOMEDCT_CORE|Post-traumatic wound infection|Post-traumatic wound infection
C1264517|T046|FN|269406001|SNOMEDCT_CORE|Post-traumatic wound infection|Post-traumatic wound infection
C1264620|T047|PT|111853008|SNOMEDCT_CORE|Herpes simplex without complication|Herpes simplex without complication
C1264620|T047|FN|111853008|SNOMEDCT_CORE|Herpes simplex without complication|Herpes simplex without complication
C1264622|T047|PT|111859007|SNOMEDCT_CORE|Herpes zoster without complication|Herpes zoster without complication
C1264622|T047|FN|111859007|SNOMEDCT_CORE|Herpes zoster without complication|Herpes zoster without complication
C1266194|T191|SY|118607005|SNOMEDCT_CORE|Hodgkin lymphoma, lymphocyte-rich|Lymphocyte-rich classical Hodgkin lymphoma
C1266194|T191|FN|118607005|SNOMEDCT_CORE|Hodgkin lymphoma, lymphocyte-rich|Lymphocyte-rich classical Hodgkin lymphoma
C1266194|T191|IS|118607005|SNOMEDCT_CORE|Hodgkin's disease, lymphocytic predominance|Lymphocyte-rich classical Hodgkin lymphoma
C1266194|T191|IS|118607005|SNOMEDCT_CORE|Hodgkin's disease, lymphocytic-histiocytic predominance|Lymphocyte-rich classical Hodgkin lymphoma
C1266194|T191|PT|118607005|SNOMEDCT_CORE|Lymphocyte-rich classical Hodgkin lymphoma|Lymphocyte-rich classical Hodgkin lymphoma
C1268712|T033|PT|129788004|SNOMEDCT_CORE|Mammographic breast mass|Mammographic breast mass
C1268712|T033|FN|129788004|SNOMEDCT_CORE|Mammographic breast mass finding|Mammographic breast mass
C1268712|T033|SY|129788004|SNOMEDCT_CORE|Mammographic breast mass finding|Mammographic breast mass
C1268740|T033|PT|129839007|SNOMEDCT_CORE|At risk for falls|At risk for falls
C1268740|T033|FN|129839007|SNOMEDCT_CORE|At risk for falls|At risk for falls
C1268740|T033|SY|129839007|SNOMEDCT_CORE|At risk of falls|At risk for falls
C1268740|T033|SY|129839007|SNOMEDCT_CORE|Fall risk|At risk for falls
C1268942|T047|PTGB|371132002|SNOMEDCT_CORE|Gastro-oesophageal reflux disease with hiatal hernia|Gastroesophageal reflux disease with hiatal hernia
C1268942|T047|PT|371132002|SNOMEDCT_CORE|Gastroesophageal reflux disease with hiatal hernia|Gastroesophageal reflux disease with hiatal hernia
C1268942|T047|SYGB|371132002|SNOMEDCT_CORE|Hiatal hernia with gastro-oesophageal reflux disease|Gastroesophageal reflux disease with hiatal hernia
C1268942|T047|SY|371132002|SNOMEDCT_CORE|Hiatal hernia with gastroesophageal reflux disease|Gastroesophageal reflux disease with hiatal hernia
C1268942|T047|FN|371132002|SNOMEDCT_CORE|Hiatal hernia with gastroesophageal reflux disease|Gastroesophageal reflux disease with hiatal hernia
C1269683|T048|IS|35489007|SNOMEDCT_CORE|Major depression|Major depressive disorder
C1269683|T048|SY|370143000|SNOMEDCT_CORE|Major depression|Major depressive disorder
C1269683|T048|IS|35489007|SNOMEDCT_CORE|Major depression, NOS|Major depressive disorder
C1269683|T048|IS|35489007|SNOMEDCT_CORE|Major depressive disorder|Major depressive disorder
C1269683|T048|PT|370143000|SNOMEDCT_CORE|Major depressive disorder|Major depressive disorder
C1269683|T048|FN|370143000|SNOMEDCT_CORE|Major depressive disorder|Major depressive disorder
C1269683|T048|IS|35489007|SNOMEDCT_CORE|Major depressive disorder, NOS|Major depressive disorder
C1269757|T047|OAS|371095004|SNOMEDCT_CORE|Infection due to penicillin-resistant organism|Infection due to penicillin-resistant organism
C1269757|T047|OAP|371095004|SNOMEDCT_CORE|Infection resistant to penicillin|Infection due to penicillin-resistant organism
C1269757|T047|OAF|371095004|SNOMEDCT_CORE|Infection resistant to penicillin|Infection due to penicillin-resistant organism
C1269831|T047|OAS|372292006|SNOMEDCT_CORE|Infection caused by resistant organism|Infection due to resistant organism
C1269831|T047|OAF|372292006|SNOMEDCT_CORE|Infection caused by resistant organism|Infection due to resistant organism
C1269831|T047|OF|372292006|SNOMEDCT_CORE|Infection due to resistant organism|Infection due to resistant organism
C1269831|T047|OAP|372292006|SNOMEDCT_CORE|Infection due to resistant organism|Infection due to resistant organism
C1269831|T047|OAS|372292006|SNOMEDCT_CORE|Resistant infection|Infection due to resistant organism
C1269832|T033|PT|373108000|SNOMEDCT_CORE|Post percutaneous transluminal coronary angioplasty|Post percutaneous transluminal coronary angioplasty
C1269832|T033|FN|373108000|SNOMEDCT_CORE|Post percutaneous transluminal coronary angioplasty|Post percutaneous transluminal coronary angioplasty
C1269832|T033|SY|373108000|SNOMEDCT_CORE|Post PTCA|Post percutaneous transluminal coronary angioplasty
C1270972|T048|PT|386805003|SNOMEDCT_CORE|Mild cognitive disorder|Mild cognitive disorder
C1270972|T048|FN|386805003|SNOMEDCT_CORE|Mild cognitive disorder|Mild cognitive disorder
C1270972|T048|SY|386805003|SNOMEDCT_CORE|Mild cognitive impairment|Mild cognitive disorder
C1271045|T033|SY|394877006|SNOMEDCT_CORE|Family history of Alzheimers|FH: Alzheimer's disease
C1271045|T033|SY|394877006|SNOMEDCT_CORE|Family history: Alzheimer disease|FH: Alzheimer's disease
C1271045|T033|SY|394877006|SNOMEDCT_CORE|Family history: Alzheimer's disease|FH: Alzheimer's disease
C1271045|T033|FN|394877006|SNOMEDCT_CORE|Family history: Alzheimer's disease|FH: Alzheimer's disease
C1271045|T033|PT|394877006|SNOMEDCT_CORE|FH: Alzheimer's disease|FH: Alzheimer's disease
C1271045|T033|OF|394877006|SNOMEDCT_CORE|FH: Alzheimer's disease|FH: Alzheimer's disease
C1271398|T047|FN|392133001|SNOMEDCT_CORE|Pigment dispersion syndrome|Pigment dispersion syndrome
C1271398|T047|PT|392133001|SNOMEDCT_CORE|Pigment dispersion syndrome|Pigment dispersion syndrome
C1272060|T033|PT|391083006|SNOMEDCT_CORE|H/O: bilateral oophorectomy|H/O: bilateral oophorectomy
C1272060|T033|OF|391083006|SNOMEDCT_CORE|H/O: bilateral oophorectomy|H/O: bilateral oophorectomy
C1272060|T033|OF|391083006|SNOMEDCT_CORE|History of - bilateral oophorectomy|H/O: bilateral oophorectomy
C1272060|T033|IS|391083006|SNOMEDCT_CORE|History of - bilateral oophorectomy|H/O: bilateral oophorectomy
C1272060|T033|FN|391083006|SNOMEDCT_CORE|History of bilateral oophorectomy|H/O: bilateral oophorectomy
C1272060|T033|SY|391083006|SNOMEDCT_CORE|History of bilateral oophorectomy|H/O: bilateral oophorectomy
C1272092|T033|SY|390951007|SNOMEDCT_CORE|Impaired fasting glucose|Impaired fasting glycemia
C1272092|T033|PTGB|390951007|SNOMEDCT_CORE|Impaired fasting glycaemia|Impaired fasting glycemia
C1272092|T033|OF|390951007|SNOMEDCT_CORE|Impaired fasting glycaemia|Impaired fasting glycemia
C1272092|T033|PT|390951007|SNOMEDCT_CORE|Impaired fasting glycemia|Impaired fasting glycemia
C1272092|T033|FN|390951007|SNOMEDCT_CORE|Impaired fasting glycemia|Impaired fasting glycemia
C1272097|T033|PT|390943009|SNOMEDCT_CORE|Serum ferritin high|Serum ferritin high
C1272097|T033|FN|390943009|SNOMEDCT_CORE|Serum ferritin high|Serum ferritin high
C1272167|T047|FN|390833005|SNOMEDCT_CORE|Osteoporosis caused by corticosteroid|Osteoporosis due to corticosteroid
C1272167|T047|SY|390833005|SNOMEDCT_CORE|Osteoporosis caused by corticosteroid|Osteoporosis due to corticosteroid
C1272167|T047|PT|390833005|SNOMEDCT_CORE|Osteoporosis due to corticosteroid|Osteoporosis due to corticosteroid
C1272167|T047|OP|390833005|SNOMEDCT_CORE|Osteoporosis due to corticosteroids|Osteoporosis due to corticosteroid
C1272167|T047|OF|390833005|SNOMEDCT_CORE|Osteoporosis due to corticosteroids|Osteoporosis due to corticosteroid
C1272176|T033|OAP|390845001|SNOMEDCT_CORE|Breast screening declined|Breast screening declined
C1272176|T033|OAF|390845001|SNOMEDCT_CORE|Breast screening declined|Breast screening declined
C1272587|T033|PT|386138005|SNOMEDCT_CORE|Stented coronary artery|Stented coronary artery
C1272587|T033|FN|386138005|SNOMEDCT_CORE|Stented coronary artery|Stented coronary artery
C1273070|T047|PT|395704004|SNOMEDCT_CORE|Left ventricular diastolic dysfunction|Left ventricular diastolic dysfunction
C1273070|T047|FN|395704004|SNOMEDCT_CORE|Left ventricular diastolic dysfunction|Left ventricular diastolic dysfunction
C1273099|T191|PTGB|395692003|SNOMEDCT_CORE|Benign paraproteinaemia|Benign paraproteinemia
C1273099|T191|OF|395692003|SNOMEDCT_CORE|Benign paraproteinaemia|Benign paraproteinemia
C1273099|T191|PT|395692003|SNOMEDCT_CORE|Benign paraproteinemia|Benign paraproteinemia
C1273099|T191|FN|395692003|SNOMEDCT_CORE|Benign paraproteinemia|Benign paraproteinemia
C1273344|T047|PT|395204000|SNOMEDCT_CORE|Hyperosmolar non-ketotic state due to type 2 diabetes mellitus|Hyperosmolar non-ketotic state due to type 2 diabetes mellitus
C1273344|T047|FN|395204000|SNOMEDCT_CORE|Hyperosmolar non-ketotic state due to type 2 diabetes mellitus|Hyperosmolar non-ketotic state due to type 2 diabetes mellitus
C1273344|T047|OF|395204000|SNOMEDCT_CORE|Hyperosmolar non-ketotic state in type 2 diabetes mellitus|Hyperosmolar non-ketotic state due to type 2 diabetes mellitus
C1273344|T047|SY|395204000|SNOMEDCT_CORE|Hyperosmolar non-ketotic state in type 2 diabetes mellitus|Hyperosmolar non-ketotic state due to type 2 diabetes mellitus
C1273544|T033|PT|394888000|SNOMEDCT_CORE|Hormone replacement therapy requested|Hormone replacement therapy requested
C1273544|T033|OF|394888000|SNOMEDCT_CORE|Hormone replacement therapy requested|Hormone replacement therapy requested
C1273544|T033|FN|394888000|SNOMEDCT_CORE|Hormone replacement therapy requested|Hormone replacement therapy requested
C1274148|T047|PT|402698005|SNOMEDCT_CORE|Dermatitis of external ear|Dermatitis of external ear
C1274148|T047|FN|402698005|SNOMEDCT_CORE|Dermatitis of external ear|Dermatitis of external ear
C1274258|T191|PT|402818009|SNOMEDCT_CORE|Basal cell carcinoma of nose|Basal cell carcinoma of nose
C1274258|T191|FN|402818009|SNOMEDCT_CORE|Basal cell carcinoma of nose|Basal cell carcinoma of nose
C1274258|T191|SY|402818009|SNOMEDCT_CORE|Cancer of nose, basal cell|Basal cell carcinoma of nose
C1274260|T191|PT|402820007|SNOMEDCT_CORE|Basal cell carcinoma of ear|Basal cell carcinoma of ear
C1274260|T191|FN|402820007|SNOMEDCT_CORE|Basal cell carcinoma of ear|Basal cell carcinoma of ear
C1274260|T191|SY|402820007|SNOMEDCT_CORE|Cancer of skin of ear, basal cell|Basal cell carcinoma of ear
C1274323|T047|PT|402894005|SNOMEDCT_CORE|Recurrent genital herpes simplex|Recurrent genital herpes simplex
C1274323|T047|FN|402894005|SNOMEDCT_CORE|Recurrent genital herpes simplex|Recurrent genital herpes simplex
C1274323|T047|SY|402894005|SNOMEDCT_CORE|Recurrent herpes genitalis|Recurrent genital herpes simplex
C1274361|T047|PT|402944008|SNOMEDCT_CORE|Condylomata lata of perianal skin|Condylomata lata of perianal skin
C1274361|T047|FN|402944008|SNOMEDCT_CORE|Condylomata lata of perianal skin|Condylomata lata of perianal skin
C1274392|T047|OF|402981007|SNOMEDCT_CORE|Mycobacterium chelonae infection of skin|Mycobacteroides chelonae infection of skin
C1274392|T047|SY|402981007|SNOMEDCT_CORE|Mycobacterium chelonae infection of skin|Mycobacteroides chelonae infection of skin
C1274392|T047|PT|402981007|SNOMEDCT_CORE|Mycobacteroides chelonae infection of skin|Mycobacteroides chelonae infection of skin
C1274392|T047|FN|402981007|SNOMEDCT_CORE|Mycobacteroides chelonae infection of skin|Mycobacteroides chelonae infection of skin
C1274581|T033|PT|403180003|SNOMEDCT_CORE|Decorative tattoo|Decorative tattoo
C1274581|T033|OF|403180003|SNOMEDCT_CORE|Decorative tattoo|Decorative tattoo
C1274581|T033|FN|403180003|SNOMEDCT_CORE|Decorative tattoo of skin|Decorative tattoo
C1274581|T033|SY|403180003|SNOMEDCT_CORE|Decorative tattoo of skin|Decorative tattoo
C1275179|T191|SY|403891008|SNOMEDCT_CORE|Cancer of the scalp, squamous cell|Squamous cell carcinoma of scalp
C1275179|T191|PT|403891008|SNOMEDCT_CORE|Squamous cell carcinoma of scalp|Squamous cell carcinoma of scalp
C1275179|T191|FN|403891008|SNOMEDCT_CORE|Squamous cell carcinoma of scalp|Squamous cell carcinoma of scalp
C1275180|T191|SY|403892001|SNOMEDCT_CORE|Squamous cell cancer of skin of face|Squamous cell carcinoma of skin of face
C1275180|T191|PT|403892001|SNOMEDCT_CORE|Squamous cell carcinoma of skin of face|Squamous cell carcinoma of skin of face
C1275180|T191|FN|403892001|SNOMEDCT_CORE|Squamous cell carcinoma of skin of face|Squamous cell carcinoma of skin of face
C1275184|T191|PT|403896003|SNOMEDCT_CORE|Squamous cell carcinoma of hand|Squamous cell carcinoma of hand
C1275184|T191|FN|403896003|SNOMEDCT_CORE|Squamous cell carcinoma of hand|Squamous cell carcinoma of hand
C1275186|T191|SY|403898002|SNOMEDCT_CORE|Squamous cell cancer of skin of lower limb|Squamous cell carcinoma of skin of lower extremity
C1275186|T191|PT|403898002|SNOMEDCT_CORE|Squamous cell carcinoma of skin of lower extremity|Squamous cell carcinoma of skin of lower extremity
C1275186|T191|FN|403898002|SNOMEDCT_CORE|Squamous cell carcinoma of skin of lower extremity|Squamous cell carcinoma of skin of lower extremity
C1275187|T191|PT|403899005|SNOMEDCT_CORE|Squamous cell carcinoma of skin of trunk|Squamous cell carcinoma of skin of trunk
C1275187|T191|FN|403899005|SNOMEDCT_CORE|Squamous cell carcinoma of skin of trunk|Squamous cell carcinoma of skin of trunk
C1275194|T191|PT|403915004|SNOMEDCT_CORE|Basal cell carcinoma of scalp|Basal cell carcinoma of scalp
C1275194|T191|FN|403915004|SNOMEDCT_CORE|Basal cell carcinoma of scalp|Basal cell carcinoma of scalp
C1275194|T191|SY|403915004|SNOMEDCT_CORE|Cancer of scalp, basal cell|Basal cell carcinoma of scalp
C1275289|T190|PT|404098005|SNOMEDCT_CORE|Digital mucous cyst|Digital mucous cyst
C1275289|T190|FN|404098005|SNOMEDCT_CORE|Digital mucous cyst|Digital mucous cyst
C1275289|T190|SY|404098005|SNOMEDCT_CORE|Digital myxoid cyst|Digital mucous cyst
C1275289|T190|SY|404098005|SNOMEDCT_CORE|Digital synovial cyst|Digital mucous cyst
C1275668|T191|SY|83217000|SNOMEDCT_CORE|Melanotic medulloblastoma|Melanotic medulloblastoma
C1275684|T047|PT|397549002|SNOMEDCT_CORE|Meibomian gland dysfunction|Meibomian gland dysfunction
C1275684|T047|FN|397549002|SNOMEDCT_CORE|Meibomian gland dysfunction|Meibomian gland dysfunction
C1275684|T047|SY|397549002|SNOMEDCT_CORE|MGD-Meibomian gland dysfunction|Meibomian gland dysfunction
C1275684|T047|SY|397549002|SNOMEDCT_CORE|Posterior blepharitis|Meibomian gland dysfunction
C1275835|T033|OP|399211009|SNOMEDCT_CORE|History of - myocardial infarction|History of myocardial infarction
C1275835|T033|OF|399211009|SNOMEDCT_CORE|History of - myocardial infarction|History of myocardial infarction
C1275835|T033|PT|399211009|SNOMEDCT_CORE|History of myocardial infarction|History of myocardial infarction
C1275835|T033|FN|399211009|SNOMEDCT_CORE|History of myocardial infarction|History of myocardial infarction
C1275835|T033|SY|399211009|SNOMEDCT_CORE|Past history of myocardial infarction|History of myocardial infarction
C1275842|T033|OP|399261000|SNOMEDCT_CORE|History of - coronary artery bypass grafting|History of coronary artery bypass grafting
C1275842|T033|OF|399261000|SNOMEDCT_CORE|History of - coronary artery bypass grafting|History of coronary artery bypass grafting
C1275842|T033|PT|399261000|SNOMEDCT_CORE|History of coronary artery bypass grafting|History of coronary artery bypass grafting
C1275842|T033|FN|399261000|SNOMEDCT_CORE|History of coronary artery bypass grafting|History of coronary artery bypass grafting
C1275842|T033|SY|399261000|SNOMEDCT_CORE|Past history of coronary artery bypass grafting|History of coronary artery bypass grafting
C1275854|T033|SY|399374009|SNOMEDCT_CORE|Regional lymph node involvement present|Regional lymph node metastasis present
C1275854|T033|PT|399374009|SNOMEDCT_CORE|Regional lymph node metastasis present|Regional lymph node metastasis present
C1275854|T033|FN|399374009|SNOMEDCT_CORE|Regional lymph node metastasis present|Regional lymph node metastasis present
C1275952|T047|OF|399872003|SNOMEDCT_CORE|Severe nonproliferative diabetic retinopathy with clinically significant macular edema|Severe nonproliferative diabetic retinopathy with clinically significant macular edema
C1275952|T047|SY|399872003|SNOMEDCT_CORE|Severe nonproliferative diabetic retinopathy with clinically significant macular edema|Severe nonproliferative diabetic retinopathy with clinically significant macular edema
C1275952|T047|SYGB|399872003|SNOMEDCT_CORE|Severe nonproliferative diabetic retinopathy with clinically significant macular oedema|Severe nonproliferative diabetic retinopathy with clinically significant macular edema
C1275952|T047|IS|399872003|SNOMEDCT_CORE|Severe NPDR with CSME|Severe nonproliferative diabetic retinopathy with clinically significant macular edema
C1276053|T033|PT|401206008|SNOMEDCT_CORE|At risk for deliberate self harm|At risk for deliberate self harm
C1276053|T033|FN|401206008|SNOMEDCT_CORE|At risk for deliberate self harm|At risk for deliberate self harm
C1276053|T033|SY|401206008|SNOMEDCT_CORE|At risk of DSH - deliberate self harm|At risk for deliberate self harm
C1276061|T047|FN|401314000|SNOMEDCT_CORE|Acute non-ST segment elevation myocardial infarction|Acute non-ST segment elevation myocardial infarction
C1276061|T047|PT|401314000|SNOMEDCT_CORE|Acute non-ST segment elevation myocardial infarction|Acute non-ST segment elevation myocardial infarction
C1276061|T047|SY|401314000|SNOMEDCT_CORE|NSTEMI - Non-ST segment elevation MI|Acute non-ST segment elevation myocardial infarction
C1276131|T191|SY|402555001|SNOMEDCT_CORE|Moles multiple benign|Multiple benign melanocytic nevi
C1276131|T191|PTGB|402555001|SNOMEDCT_CORE|Multiple benign melanocytic naevi|Multiple benign melanocytic nevi
C1276131|T191|PT|402555001|SNOMEDCT_CORE|Multiple benign melanocytic nevi|Multiple benign melanocytic nevi
C1276131|T191|FN|402555001|SNOMEDCT_CORE|Multiple benign melanocytic nevi|Multiple benign melanocytic nevi
C1277595|T033|PT|314938000|SNOMEDCT_CORE|Poor sleep pattern|Poor sleep pattern
C1277595|T033|FN|314938000|SNOMEDCT_CORE|Poor sleep pattern|Poor sleep pattern
C1277629|T033|PT|315284009|SNOMEDCT_CORE|Mass of parotid gland|Mass of parotid gland
C1277629|T033|FN|315284009|SNOMEDCT_CORE|Mass of parotid gland|Mass of parotid gland
C1277629|T033|SY|315284009|SNOMEDCT_CORE|Parotid lump|Mass of parotid gland
C1277644|T033|PT|315249005|SNOMEDCT_CORE|Persistent breast nodularity|Persistent breast nodularity
C1277644|T033|FN|315249005|SNOMEDCT_CORE|Persistent breast nodularity|Persistent breast nodularity
C1277644|T033|SY|315249005|SNOMEDCT_CORE|Persistent nodularity|Persistent breast nodularity
C1278395|T033|PT|314956000|SNOMEDCT_CORE|Borderline blood pressure|Borderline blood pressure
C1278395|T033|FN|314956000|SNOMEDCT_CORE|Borderline blood pressure|Borderline blood pressure
C1278535|T047|PT|314116003|SNOMEDCT_CORE|Post infarct angina|Post infarct angina
C1278535|T047|FN|314116003|SNOMEDCT_CORE|Post infarct angina|Post infarct angina
C1278558|T037|SY|35468003|SNOMEDCT_CORE|Caught, crushed, jammed or pinched in or between objects|Crushed in between objects
C1278558|T037|PT|35468003|SNOMEDCT_CORE|Crushed in between objects|Crushed in between objects
C1278558|T037|OF|35468003|SNOMEDCT_CORE|Crushed in between objects|Crushed in between objects
C1278558|T037|FN|35468003|SNOMEDCT_CORE|Crushed in between objects|Crushed in between objects
C1278558|T037|IS|35468003|SNOMEDCT_CORE|Crushed in between objects, NOS|Crushed in between objects
C1279224|T047|OAP|186156007|SNOMEDCT_CORE|Infectious colitis, enteritis and gastroenteritis|Infectious colitis, enteritis and gastroenteritis
C1279224|T047|OAF|186156007|SNOMEDCT_CORE|Infectious colitis, enteritis and gastroenteritis|Infectious colitis, enteritis and gastroenteritis
C1279258|T191|PT|188189001|SNOMEDCT_CORE|Malignant neoplasm of corpus uteri, excluding isthmus|Malignant neoplasm of corpus uteri, excluding isthmus
C1279258|T191|FN|188189001|SNOMEDCT_CORE|Malignant neoplasm of corpus uteri, excluding isthmus|Malignant neoplasm of corpus uteri, excluding isthmus
C1279296|T191|PTGB|92812005|SNOMEDCT_CORE|Chronic leukaemia|Chronic leukemia
C1279296|T191|SYGB|92812005|SNOMEDCT_CORE|Chronic leukaemia, disease|Chronic leukemia
C1279296|T191|PT|92812005|SNOMEDCT_CORE|Chronic leukemia|Chronic leukemia
C1279296|T191|FN|92812005|SNOMEDCT_CORE|Chronic leukemia, disease|Chronic leukemia
C1279296|T191|SY|92812005|SNOMEDCT_CORE|Chronic leukemia, disease|Chronic leukemia
C1279315|T047|IS|314904008|SNOMEDCT_CORE|Non-insulin dependent diabetes mellitus with neuropathic arthropathy|Type 2 diabetes mellitus with neuropathic arthropathy
C1279315|T047|PT|314904008|SNOMEDCT_CORE|Type 2 diabetes mellitus with neuropathic arthropathy|Type 2 diabetes mellitus with neuropathic arthropathy
C1279315|T047|FN|314904008|SNOMEDCT_CORE|Type II diabetes mellitus with neuropathic arthropathy|Type 2 diabetes mellitus with neuropathic arthropathy
C1279315|T047|SY|314904008|SNOMEDCT_CORE|Type II diabetes mellitus with neuropathic arthropathy|Type 2 diabetes mellitus with neuropathic arthropathy
C1279369|T047|PT|315348000|SNOMEDCT_CORE|Asymptomatic coronary heart disease|Asymptomatic coronary heart disease
C1279369|T047|FN|315348000|SNOMEDCT_CORE|Asymptomatic coronary heart disease|Asymptomatic coronary heart disease
C1279386|T047|PT|314978007|SNOMEDCT_CORE|Postoperative pneumonia|Postoperative pneumonia
C1279386|T047|FN|314978007|SNOMEDCT_CORE|Postoperative pneumonia|Postoperative pneumonia
C1279420|T048|FN|207363009|SNOMEDCT_CORE|Anxiety neurosis|Anxiety neurosis
C1279420|T048|PT|207363009|SNOMEDCT_CORE|Anxiety neurosis|Anxiety neurosis
C1279702|T047|IS|415530009|SNOMEDCT_CORE|Calorie overload|Calorie overload
C1279945|T047|IS|45157009|SNOMEDCT_CORE|Idiopathic fibrosing alveolitis, acute fatal form|Idiopathic fibrosing alveolitis, acute fatal form
C1280798|T047|SY|128105004|SNOMEDCT_CORE|von Willebrand disease, platelet type|von Willebrand disease, platelet type
C1281429|T033|SY|415530009|SNOMEDCT_CORE|Alimentary obesity|Exogenous obesity
C1281429|T033|SY|415530009|SNOMEDCT_CORE|Exogenous obesity|Exogenous obesity
C1281489|T047|PT|297713002|SNOMEDCT_CORE|Varicose veins of lower extremity without ulcer AND without inflammation|Varicose veins of lower extremity without ulcer AND without inflammation
C1281489|T047|FN|297713002|SNOMEDCT_CORE|Varicose veins of lower extremity without ulcer AND without inflammation|Varicose veins of lower extremity without ulcer AND without inflammation
C1281551|T033|PT|302109006|SNOMEDCT_CORE|Gastrostomy present|Gastrostomy present
C1281551|T033|FN|302109006|SNOMEDCT_CORE|Gastrostomy present|Gastrostomy present
C1281553|T033|FN|302111002|SNOMEDCT_CORE|Ileostomy present|Ileostomy present
C1281553|T033|PT|302111002|SNOMEDCT_CORE|Ileostomy present|Ileostomy present
C1281553|T033|SY|302111002|SNOMEDCT_CORE|Ileostomy, has currently|Ileostomy present
C1281554|T033|PT|302112009|SNOMEDCT_CORE|Colostomy present|Colostomy present
C1281554|T033|FN|302112009|SNOMEDCT_CORE|Colostomy present|Colostomy present
C1281729|T037|PT|307945003|SNOMEDCT_CORE|Current tear of medial cartilage AND/OR meniscus of knee|Current tear of medial cartilage AND/OR meniscus of knee
C1281729|T037|FN|307945003|SNOMEDCT_CORE|Current tear of medial cartilage AND/OR meniscus of knee|Current tear of medial cartilage AND/OR meniscus of knee
C1281794|T037|PT|308849005|SNOMEDCT_CORE|Current tear of lateral cartilage AND/OR meniscus of knee|Current tear of lateral cartilage AND/OR meniscus of knee
C1281794|T037|FN|308849005|SNOMEDCT_CORE|Current tear of lateral cartilage AND/OR meniscus of knee|Current tear of lateral cartilage AND/OR meniscus of knee
C1281931|T033|OF|314022009|SNOMEDCT_CORE|Nasolacrimal duct obstructed|Obstruction of nasolacrimal duct
C1281931|T033|SY|314022009|SNOMEDCT_CORE|Nasolacrimal duct obstructed|Obstruction of nasolacrimal duct
C1281931|T033|OAP|417162001|SNOMEDCT_CORE|Nasolacrimal duct obstruction|Obstruction of nasolacrimal duct
C1281931|T033|SY|231841004|SNOMEDCT_CORE|Nasolacrimal duct obstruction|Obstruction of nasolacrimal duct
C1281931|T033|OAF|417162001|SNOMEDCT_CORE|Nasolacrimal duct obstruction|Obstruction of nasolacrimal duct
C1281931|T033|OAS|417162001|SNOMEDCT_CORE|NLDO - nasolacrimal duct obstruction|Obstruction of nasolacrimal duct
C1281931|T033|PT|314022009|SNOMEDCT_CORE|Obstruction of nasolacrimal duct|Obstruction of nasolacrimal duct
C1281931|T033|FN|314022009|SNOMEDCT_CORE|Obstruction of nasolacrimal duct|Obstruction of nasolacrimal duct
C1281995|T037|PT|314201008|SNOMEDCT_CORE|Dislocation of hip joint prosthesis|Dislocation of hip joint prosthesis
C1281995|T037|FN|314201008|SNOMEDCT_CORE|Dislocation of hip joint prosthesis|Dislocation of hip joint prosthesis
C1281999|T047|PT|314208002|SNOMEDCT_CORE|Rapid atrial fibrillation|Rapid atrial fibrillation
C1281999|T047|FN|314208002|SNOMEDCT_CORE|Rapid atrial fibrillation|Rapid atrial fibrillation
C1282208|T047|PT|314516007|SNOMEDCT_CORE|Preseptal cellulitis|Preseptal cellulitis
C1282208|T047|FN|314516007|SNOMEDCT_CORE|Preseptal cellulitis|Preseptal cellulitis
C1282376|T047|PT|314788004|SNOMEDCT_CORE|Divergence insufficiency|Divergence insufficiency
C1282376|T047|FN|314788004|SNOMEDCT_CORE|Divergence insufficiency|Divergence insufficiency
C1282471|T191|PT|314955001|SNOMEDCT_CORE|Local recurrence of malignant tumor of breast|Local recurrence of malignant tumor of breast
C1282471|T191|FN|314955001|SNOMEDCT_CORE|Local recurrence of malignant tumor of breast|Local recurrence of malignant tumor of breast
C1282471|T191|PTGB|314955001|SNOMEDCT_CORE|Local recurrence of malignant tumour of breast|Local recurrence of malignant tumor of breast
C1282478|T191|PT|314965007|SNOMEDCT_CORE|Local recurrence of malignant tumor of colon|Local recurrence of malignant tumor of colon
C1282478|T191|FN|314965007|SNOMEDCT_CORE|Local recurrence of malignant tumor of colon|Local recurrence of malignant tumor of colon
C1282478|T191|PTGB|314965007|SNOMEDCT_CORE|Local recurrence of malignant tumour of colon|Local recurrence of malignant tumor of colon
C1282479|T191|PT|314966008|SNOMEDCT_CORE|Local recurrence of malignant tumor of rectum|Local recurrence of malignant tumor of rectum
C1282479|T191|FN|314966008|SNOMEDCT_CORE|Local recurrence of malignant tumor of rectum|Local recurrence of malignant tumor of rectum
C1282479|T191|PTGB|314966008|SNOMEDCT_CORE|Local recurrence of malignant tumour of rectum|Local recurrence of malignant tumor of rectum
C1282492|T191|PT|314990009|SNOMEDCT_CORE|Metastasis from malignant tumor of bone|Metastasis from malignant tumor of bone
C1282492|T191|FN|314990009|SNOMEDCT_CORE|Metastasis from malignant tumor of bone|Metastasis from malignant tumor of bone
C1282492|T191|PTGB|314990009|SNOMEDCT_CORE|Metastasis from malignant tumour of bone|Metastasis from malignant tumor of bone
C1282512|T033|SY|315016007|SNOMEDCT_CORE|At risk of CHD|At risk of coronary heart disease
C1282512|T033|PT|315016007|SNOMEDCT_CORE|At risk of coronary heart disease|At risk of coronary heart disease
C1282512|T033|FN|315016007|SNOMEDCT_CORE|At risk of coronary heart disease|At risk of coronary heart disease
C1282926|T047|PT|359532006|SNOMEDCT_CORE|Rotator cuff impingement syndrome|Rotator cuff impingement syndrome
C1282926|T047|FN|359532006|SNOMEDCT_CORE|Rotator cuff impingement syndrome|Rotator cuff impingement syndrome
C1285577|T033|SY|2776000|SNOMEDCT_CORE|Acute confusional state|Acute confusional state
C1288279|T047|PT|367475009|SNOMEDCT_CORE|Lesion of ulnar nerve|Lesion of ulnar nerve
C1288279|T047|FN|367475009|SNOMEDCT_CORE|Lesion of ulnar nerve|Lesion of ulnar nerve
C1290118|T191|PTGB|109269004|SNOMEDCT_CORE|Melanocytic naevus of face|Melanocytic nevus of face
C1290118|T191|PT|109269004|SNOMEDCT_CORE|Melanocytic nevus of face|Melanocytic nevus of face
C1290118|T191|FN|109269004|SNOMEDCT_CORE|Melanocytic nevus of face|Melanocytic nevus of face
C1290139|T047|IS|48245008|SNOMEDCT_CORE|Arthropathy associated with bacterial disease|Arthropathy associated with bacterial disease
C1290145|T047|PT|128049000|SNOMEDCT_CORE|Disorder of cervical spine|Disorder of cervical spine
C1290145|T047|FN|128049000|SNOMEDCT_CORE|Disorder of cervical spine|Disorder of cervical spine
C1290147|T047|PT|129139009|SNOMEDCT_CORE|Disorder of lumbar spine|Disorder of lumbar spine
C1290147|T047|FN|129139009|SNOMEDCT_CORE|Disorder of lumbar spine|Disorder of lumbar spine
C1290398|T047|PT|128608001|SNOMEDCT_CORE|Cerebral arterial aneurysm|Cerebral arterial aneurysm
C1290398|T047|IS|42994005|SNOMEDCT_CORE|Cerebral arterial aneurysm|Cerebral arterial aneurysm
C1290398|T047|FN|128608001|SNOMEDCT_CORE|Cerebral arterial aneurysm|Cerebral arterial aneurysm
C1290398|T047|IS|128608001|SNOMEDCT_CORE|Intracranial arterial aneurysm|Cerebral arterial aneurysm
C1290603|T019|OAP|111333002|SNOMEDCT_CORE|Congenital anomaly of genital system|Congenital anomaly of genital system
C1290603|T019|OAF|111333002|SNOMEDCT_CORE|Congenital anomaly of genital system|Congenital anomaly of genital system
C1290739|T033|SY|109728009|SNOMEDCT_CORE|Abnormal tooth restoration|Defective dental restoration
C1290739|T033|PT|109728009|SNOMEDCT_CORE|Defective dental restoration|Defective dental restoration
C1290739|T033|FN|109728009|SNOMEDCT_CORE|Defective dental restoration|Defective dental restoration
C1290739|T033|SY|109728009|SNOMEDCT_CORE|Defective restoration of teeth|Defective dental restoration
C1290807|T047|IS|43240000|SNOMEDCT_CORE|Diarrheal disease, NOS|Diarrheal disease, NOS
C1290807|T047|IS|43240000|SNOMEDCT_CORE|Diarrhoeal disease, NOS|Diarrhoeal disease, NOS
C1290810|T047|IS|40468003|SNOMEDCT_CORE|Viral hepatitis A without mention of hepatic coma|Viral hepatitis A without mention of hepatic coma
C1290859|T047|OF|118944007|SNOMEDCT_CORE|Disease of shoulder|Disorder of shoulder
C1290859|T047|IS|118944007|SNOMEDCT_CORE|Disease of shoulder|Disorder of shoulder
C1290859|T047|PT|118944007|SNOMEDCT_CORE|Disorder of shoulder|Disorder of shoulder
C1290859|T047|FN|118944007|SNOMEDCT_CORE|Disorder of shoulder region|Disorder of shoulder
C1290859|T047|SY|118944007|SNOMEDCT_CORE|Disorder of shoulder region|Disorder of shoulder
C1290875|T047|OF|128133004|SNOMEDCT_CORE|Disease of elbow|Disorder of elbow
C1290875|T047|IS|128133004|SNOMEDCT_CORE|Disease of elbow|Disorder of elbow
C1290875|T047|PT|128133004|SNOMEDCT_CORE|Disorder of elbow|Disorder of elbow
C1290875|T047|FN|128133004|SNOMEDCT_CORE|Disorder of elbow|Disorder of elbow
C1290876|T047|OF|118937003|SNOMEDCT_CORE|Disease of lower extremity|Disorder of lower extremity
C1290876|T047|IS|118937003|SNOMEDCT_CORE|Disease of lower extremity|Disorder of lower extremity
C1290876|T047|PT|118937003|SNOMEDCT_CORE|Disorder of lower extremity|Disorder of lower extremity
C1290876|T047|FN|118937003|SNOMEDCT_CORE|Disorder of lower extremity|Disorder of lower extremity
C1290879|T047|OF|128136007|SNOMEDCT_CORE|Disease of knee|Disorder of knee
C1290879|T047|IS|128136007|SNOMEDCT_CORE|Disease of knee|Disorder of knee
C1290879|T047|PT|128136007|SNOMEDCT_CORE|Disorder of knee|Disorder of knee
C1290879|T047|FN|128136007|SNOMEDCT_CORE|Disorder of knee|Disorder of knee
C1291077|T184|IS|116289008|SNOMEDCT_CORE|Abdomen feels bloated|Abdominal bloating
C1291077|T184|PT|116289008|SNOMEDCT_CORE|Abdominal bloating|Abdominal bloating
C1291077|T184|FN|116289008|SNOMEDCT_CORE|Abdominal bloating|Abdominal bloating
C1291077|T184|SY|60728008|SNOMEDCT_CORE|Bloat|Abdominal bloating
C1291077|T184|SY|60728008|SNOMEDCT_CORE|Bloated abdomen|Abdominal bloating
C1291077|T184|SY|60728008|SNOMEDCT_CORE|Bloating|Abdominal bloating
C1291077|T184|IS|60728008|SNOMEDCT_CORE|Gassiness|Abdominal bloating
C1291077|T184|SY|60728008|SNOMEDCT_CORE|Meteorism|Abdominal bloating
C1291077|T184|IS|60728008|SNOMEDCT_CORE|Tympanites|Abdominal bloating
C1291748|T033|PT|110368006|SNOMEDCT_CORE|Decreased estrogen level|Decreased estrogen level
C1291748|T033|FN|110368006|SNOMEDCT_CORE|Decreased estrogen level|Decreased estrogen level
C1291748|T033|PTGB|110368006|SNOMEDCT_CORE|Decreased oestrogen level|Decreased estrogen level
C1292769|T191|PT|277571004|SNOMEDCT_CORE|B-cell acute lymphoblastic leukemia|B-cell acute lymphoblastic leukemia
C1292769|T191|FN|277571004|SNOMEDCT_CORE|B-cell acute lymphoblastic leukemia|B-cell acute lymphoblastic leukemia
C1292769|T191|SYGB|277571004|SNOMEDCT_CORE|Mature B-cell leukaemia Burkitt type|B-cell acute lymphoblastic leukemia
C1292769|T191|SY|277571004|SNOMEDCT_CORE|Mature B-cell leukemia Burkitt type|B-cell acute lymphoblastic leukemia
C1295654|T033|PT|131078003|SNOMEDCT_CORE|Decreased testosterone level|Decreased testosterone level
C1295654|T033|FN|131078003|SNOMEDCT_CORE|Decreased testosterone level|Decreased testosterone level
C1295654|T033|SY|131078003|SNOMEDCT_CORE|Low testosterone|Decreased testosterone level
C1297929|T046|PT|369462000|SNOMEDCT_CORE|Atypical hyperplasia of breast|Atypical hyperplasia of breast
C1297929|T046|FN|369462000|SNOMEDCT_CORE|Atypical hyperplasia of breast|Atypical hyperplasia of breast
C1298685|T047|PT|373621006|SNOMEDCT_CORE|Chronic pain syndrome|Chronic pain syndrome
C1298685|T047|FN|373621006|SNOMEDCT_CORE|Chronic pain syndrome|Chronic pain syndrome
C1298714|T019|PT|373584008|SNOMEDCT_CORE|Congenital pelviureteric junction obstruction|Congenital pelviureteric junction obstruction
C1298714|T019|FN|373584008|SNOMEDCT_CORE|Congenital pelviureteric junction obstruction|Congenital pelviureteric junction obstruction
C1299237|T191|FN|372098004|SNOMEDCT_CORE|Carcinoma of endocervix|Carcinoma of endocervix
C1299237|T191|PT|372098004|SNOMEDCT_CORE|Carcinoma of endocervix|Carcinoma of endocervix
C1299238|T191|FN|372100004|SNOMEDCT_CORE|Carcinoma of exocervix|Carcinoma of exocervix
C1299238|T191|PT|372100004|SNOMEDCT_CORE|Carcinoma of exocervix|Carcinoma of exocervix
C1299242|T191|PT|372111007|SNOMEDCT_CORE|Carcinoma of lower lobe, bronchus or lung|Carcinoma of lower lobe, bronchus or lung
C1299242|T191|FN|372111007|SNOMEDCT_CORE|Carcinoma of lower lobe, bronchus or lung|Carcinoma of lower lobe, bronchus or lung
C1299244|T191|PT|372113005|SNOMEDCT_CORE|Carcinoma of middle lobe, bronchus or lung|Carcinoma of middle lobe, bronchus or lung
C1299244|T191|FN|372113005|SNOMEDCT_CORE|Carcinoma of middle lobe, bronchus or lung|Carcinoma of middle lobe, bronchus or lung
C1299250|T191|PT|372120003|SNOMEDCT_CORE|Carcinoma of main bronchus|Carcinoma of main bronchus
C1299250|T191|FN|372120003|SNOMEDCT_CORE|Carcinoma of main bronchus|Carcinoma of main bronchus
C1299257|T191|PT|372136001|SNOMEDCT_CORE|Carcinoma of upper lobe, bronchus or lung|Carcinoma of upper lobe, bronchus or lung
C1299257|T191|FN|372136001|SNOMEDCT_CORE|Carcinoma of upper lobe, bronchus or lung|Carcinoma of upper lobe, bronchus or lung
C1299297|T191|PT|372003004|SNOMEDCT_CORE|Primary malignant neoplasm of pancreas|Primary malignant neoplasm of pancreas
C1299297|T191|FN|372003004|SNOMEDCT_CORE|Primary malignant neoplasm of pancreas|Primary malignant neoplasm of pancreas
C1299302|T191|PT|372010005|SNOMEDCT_CORE|Primary malignant neoplasm of soft tissues|Primary malignant neoplasm of soft tissues
C1299302|T191|FN|372010005|SNOMEDCT_CORE|Primary malignant neoplasm of soft tissues|Primary malignant neoplasm of soft tissues
C1299307|T191|PT|372016004|SNOMEDCT_CORE|Primary malignant neoplasm of the peritoneum|Primary malignant neoplasm of the peritoneum
C1299307|T191|FN|372016004|SNOMEDCT_CORE|Primary malignant neoplasm of the peritoneum|Primary malignant neoplasm of the peritoneum
C1299435|T047|OP|371806006|SNOMEDCT_CORE|Progressive Angina|Progressive angina
C1299435|T047|PT|371806006|SNOMEDCT_CORE|Progressive angina|Progressive angina
C1299435|T047|FN|371806006|SNOMEDCT_CORE|Progressive angina|Progressive angina
C1299435|T047|OF|371806006|SNOMEDCT_CORE|Progressive Angina|Progressive angina
C1299471|T047|SY|371686006|SNOMEDCT_CORE|Infection caused by Mycobacterium avium complex|Infection due to Mycobacterium avium-intracellulare group
C1299471|T047|SY|371686006|SNOMEDCT_CORE|Infection caused by Mycobacterium avium-intracellulare group|Infection due to Mycobacterium avium-intracellulare group
C1299471|T047|FN|371686006|SNOMEDCT_CORE|Infection caused by Mycobacterium avium-intracellulare group|Infection due to Mycobacterium avium-intracellulare group
C1299471|T047|SY|371686006|SNOMEDCT_CORE|Infection due to Mycobacterium avium complex|Infection due to Mycobacterium avium-intracellulare group
C1299471|T047|PT|371686006|SNOMEDCT_CORE|Infection due to Mycobacterium avium-intracellulare group|Infection due to Mycobacterium avium-intracellulare group
C1299471|T047|OF|371686006|SNOMEDCT_CORE|Infection due to Mycobacterium avium-intracellulare group|Infection due to Mycobacterium avium-intracellulare group
C1299544|T033|SY|371435006|SNOMEDCT_CORE|H/O: drug abuse|History of drug abuse
C1299544|T033|OF|371435006|SNOMEDCT_CORE|History of drug abuse|History of drug abuse
C1299544|T033|PT|371435006|SNOMEDCT_CORE|History of drug abuse|History of drug abuse
C1299544|T033|FN|371435006|SNOMEDCT_CORE|History of drug abuse|History of drug abuse
C1299615|T046|PT|371060002|SNOMEDCT_CORE|Visual loss after cataract extraction|Visual loss after cataract extraction
C1299615|T046|FN|371060002|SNOMEDCT_CORE|Visual loss after cataract extraction|Visual loss after cataract extraction
C1299624|T047|PT|371073003|SNOMEDCT_CORE|Postural orthostatic tachycardia syndrome|Postural orthostatic tachycardia syndrome
C1299624|T047|FN|371073003|SNOMEDCT_CORE|Postural orthostatic tachycardia syndrome|Postural orthostatic tachycardia syndrome
C1299631|T020|PT|371084005|SNOMEDCT_CORE|Partially edentulous mandible|Partially edentulous mandible
C1299631|T020|FN|371084005|SNOMEDCT_CORE|Partially edentulous mandible|Partially edentulous mandible
C1299633|T047|PT|371088008|SNOMEDCT_CORE|Reactive airways dysfunction syndrome|Reactive airways dysfunction syndrome
C1299633|T047|FN|371088008|SNOMEDCT_CORE|Reactive airways dysfunction syndrome|Reactive airways dysfunction syndrome
C1299634|T047|PT|371090009|SNOMEDCT_CORE|Cholestasis of parenteral nutrition|Cholestasis of parenteral nutrition
C1299634|T047|FN|371090009|SNOMEDCT_CORE|Cholestasis of parenteral nutrition|Cholestasis of parenteral nutrition
C1299881|T020|PT|370471003|SNOMEDCT_CORE|Lumbosacral stenosis|Lumbosacral stenosis
C1299881|T020|FN|370471003|SNOMEDCT_CORE|Lumbosacral stenosis|Lumbosacral stenosis
C1299881|T020|OAF|428513007|SNOMEDCT_CORE|Stenosis of lumbosacral spine|Lumbosacral stenosis
C1299881|T020|OAP|428513007|SNOMEDCT_CORE|Stenosis of lumbosacral spine|Lumbosacral stenosis
C1299932|T033|PT|370532003|SNOMEDCT_CORE|Head tilt|Head tilt
C1299932|T033|FN|370532003|SNOMEDCT_CORE|Head tilt|Head tilt
C1299938|T046|FN|370540009|SNOMEDCT_CORE|Adverse reaction caused by food|Adverse reaction to food
C1299938|T046|SY|370540009|SNOMEDCT_CORE|Adverse reaction caused by food|Adverse reaction to food
C1299938|T046|PT|370540009|SNOMEDCT_CORE|Adverse reaction to food|Adverse reaction to food
C1299938|T046|OF|370540009|SNOMEDCT_CORE|Adverse reaction to food|Adverse reaction to food
C1299975|T037|PT|370240005|SNOMEDCT_CORE|Superficial laceration of foot|Superficial laceration of foot
C1299975|T037|FN|370240005|SNOMEDCT_CORE|Superficial laceration of foot|Superficial laceration of foot
C1299978|T037|IS|274172008|SNOMEDCT_CORE|Superficial laceration of finger|Superficial laceration of finger
C1299979|T037|IS|284549007|SNOMEDCT_CORE|Superficial laceration of hand|Superficial laceration of hand
C1299979|T037|PT|370244001|SNOMEDCT_CORE|Superficial laceration of hand|Superficial laceration of hand
C1299979|T037|FN|370244001|SNOMEDCT_CORE|Superficial laceration of hand|Superficial laceration of hand
C1299982|T037|PT|370247008|SNOMEDCT_CORE|Facial laceration|Facial laceration
C1299982|T037|FN|370247008|SNOMEDCT_CORE|Facial laceration|Facial laceration
C1301626|T047|IS|46764007|SNOMEDCT_CORE|Hypertension with albuminuria|Hypertension with albuminuria
C1302248|T047|PTGB|399194009|SNOMEDCT_CORE|Disorder characterised by back pain|Disorder characterized by back pain
C1302248|T047|PT|399194009|SNOMEDCT_CORE|Disorder characterized by back pain|Disorder characterized by back pain
C1302248|T047|FN|399194009|SNOMEDCT_CORE|Disorder characterized by back pain|Disorder characterized by back pain
C1302652|T191|PT|399730005|SNOMEDCT_CORE|Adenoma of rectum|Adenoma of rectum
C1302652|T191|FN|399730005|SNOMEDCT_CORE|Adenoma of rectum|Adenoma of rectum
C1302709|T047|PT|399901005|SNOMEDCT_CORE|Acquired plantar keratoderma|Acquired plantar keratoderma
C1302709|T047|FN|399901005|SNOMEDCT_CORE|Acquired plantar keratoderma|Acquired plantar keratoderma
C1302713|T037|PT|399907009|SNOMEDCT_CORE|Animal bite wound|Animal bite wound
C1302713|T037|FN|399907009|SNOMEDCT_CORE|Animal bite wound|Animal bite wound
C1302713|T037|SY|399907009|SNOMEDCT_CORE|Injury caused by animal bite|Animal bite wound
C1302752|T037|PT|399963005|SNOMEDCT_CORE|Abrasion|Abrasion
C1302752|T037|FN|399963005|SNOMEDCT_CORE|Abrasion|Abrasion
C1302752|T037|SY|399963005|SNOMEDCT_CORE|Graze|Abrasion
C1302752|T037|SY|399963005|SNOMEDCT_CORE|Superficial abrasion|Abrasion
C1302790|T047|PT|400038003|SNOMEDCT_CORE|Congenital malformation syndrome|Congenital malformation syndrome
C1302790|T047|FN|400038003|SNOMEDCT_CORE|Congenital malformation syndrome|Congenital malformation syndrome
C1302790|T047|SY|400038003|SNOMEDCT_CORE|Multiple congenital anomalies|Congenital malformation syndrome
C1302790|T047|SY|400038003|SNOMEDCT_CORE|Multiple congenital malformations|Congenital malformation syndrome
C1302856|T191|PT|443250000|SNOMEDCT_CORE|Malignant fibromatous neoplasm|Malignant fibromatous neoplasm
C1302856|T191|FN|443250000|SNOMEDCT_CORE|Malignant fibromatous neoplasm|Malignant fibromatous neoplasm
C1303112|T047|OAP|401110002|SNOMEDCT_CORE|Type 1 diabetes mellitus with persistent microalbuminuria|Type 1 diabetes mellitus with persistent microalbuminuria
C1303112|T047|OAF|401110002|SNOMEDCT_CORE|Type 1 diabetes mellitus with persistent microalbuminuria|Type 1 diabetes mellitus with persistent microalbuminuria
C1303147|T033|PT|401169009|SNOMEDCT_CORE|Not yet walking|Not yet walking
C1303147|T033|FN|401169009|SNOMEDCT_CORE|Not yet walking|Not yet walking
C1303258|T047|FN|401303003|SNOMEDCT_CORE|Acute ST segment elevation myocardial infarction|Acute ST segment elevation myocardial infarction
C1303258|T047|PT|401303003|SNOMEDCT_CORE|Acute ST segment elevation myocardial infarction|Acute ST segment elevation myocardial infarction
C1303258|T047|SY|401303003|SNOMEDCT_CORE|STEMI - ST elevation myocardial infarction|Acute ST segment elevation myocardial infarction
C1304281|T191|PT|402509003|SNOMEDCT_CORE|Basal cell carcinoma of neck|Basal cell carcinoma of neck
C1304281|T191|FN|402509003|SNOMEDCT_CORE|Basal cell carcinoma of neck|Basal cell carcinoma of neck
C1304281|T191|SY|402509003|SNOMEDCT_CORE|Cancer of skin of neck, basal cell|Basal cell carcinoma of neck
C1304291|T191|PT|402519009|SNOMEDCT_CORE|Basal cell carcinoma of face|Basal cell carcinoma of face
C1304291|T191|FN|402519009|SNOMEDCT_CORE|Basal cell carcinoma of face|Basal cell carcinoma of face
C1304291|T191|SY|402519009|SNOMEDCT_CORE|Cancer of skin of face, basal cell|Basal cell carcinoma of face
C1304293|T191|PT|402522006|SNOMEDCT_CORE|Basal cell carcinoma of lower extremity|Basal cell carcinoma of lower extremity
C1304293|T191|FN|402522006|SNOMEDCT_CORE|Basal cell carcinoma of lower extremity|Basal cell carcinoma of lower extremity
C1304293|T191|SY|402522006|SNOMEDCT_CORE|Cancer of skin of lower limb, basal cell|Basal cell carcinoma of lower extremity
C1304294|T191|PT|402523001|SNOMEDCT_CORE|Basal cell carcinoma of truncal skin|Basal cell carcinoma of truncal skin
C1304294|T191|FN|402523001|SNOMEDCT_CORE|Basal cell carcinoma of truncal skin|Basal cell carcinoma of truncal skin
C1304294|T191|SY|402523001|SNOMEDCT_CORE|Cancer of skin of trunk, basal cell|Basal cell carcinoma of truncal skin
C1305267|T191|SY|14990007|SNOMEDCT_CORE|Fibrochondrosarcoma|Fibrochondrosarcoma
C1305875|T047|SY|23260002|SNOMEDCT_CORE|Fibroadenosis breast|Fibroadenosis of breast
C1305875|T047|PT|23260002|SNOMEDCT_CORE|Fibroadenosis of breast|Fibroadenosis of breast
C1305875|T047|FN|23260002|SNOMEDCT_CORE|Fibroadenosis of breast|Fibroadenosis of breast
C1305875|T047|IS|23260002|SNOMEDCT_CORE|Fibroadenosis of breast, NOS|Fibroadenosis of breast
C1305887|T191|PT|269579005|SNOMEDCT_CORE|Malignant melanoma of trunk|Malignant melanoma of trunk
C1305887|T191|FN|269579005|SNOMEDCT_CORE|Malignant melanoma of trunk|Malignant melanoma of trunk
C1305936|T047|SY|70759006|SNOMEDCT_CORE|Pustuloderma|Pustuloderma
C1305951|T047|SY|86279000|SNOMEDCT_CORE|Acute suppurative otitis media with discharge|Acute suppurative otitis media with discharge
C1305953|T033|SY|195957006|SNOMEDCT_CORE|Emphysematous bulla|Emphysematous bulla
C1306041|T046|OF|156073000|SNOMEDCT_CORE|Complete miscarriage|Complete miscarriage
C1306041|T046|PT|156073000|SNOMEDCT_CORE|Complete miscarriage|Complete miscarriage
C1306041|T046|FN|156073000|SNOMEDCT_CORE|Complete miscarriage|Complete miscarriage
C1306041|T046|OAS|69124005|SNOMEDCT_CORE|Complete spontaneous abortion|Complete miscarriage
C1306041|T046|SY|156073000|SNOMEDCT_CORE|Complete spontaneous abortion|Complete miscarriage
C1306063|T047|IS|85232009|SNOMEDCT_CORE|Acute edema of lung with heart disease|Acute edema of lung with heart disease
C1306063|T047|IS|85232009|SNOMEDCT_CORE|Acute pulmonary edema with heart disease|Acute edema of lung with heart disease
C1306068|T047|SY|766834007|SNOMEDCT_CORE|After-cataract|Secondary cataract
C1306068|T047|OAP|47337003|SNOMEDCT_CORE|After-cataract|Secondary cataract
C1306068|T047|OF|47337003|SNOMEDCT_CORE|After-cataract|Secondary cataract
C1306068|T047|IS|47337003|SNOMEDCT_CORE|After-cataract, NOS|Secondary cataract
C1306068|T047|OAS|47337003|SNOMEDCT_CORE|Capsular fibrosis|Secondary cataract
C1306068|T047|OAS|47337003|SNOMEDCT_CORE|Cloudy posterior capsule|Secondary cataract
C1306068|T047|OAS|47337003|SNOMEDCT_CORE|PCF - Posterior capsular fibrosis|Secondary cataract
C1306068|T047|OAS|47337003|SNOMEDCT_CORE|PCO - Posterior capsule opacification|Secondary cataract
C1306068|T047|OAF|47337003|SNOMEDCT_CORE|Posterior capsular opacification|Secondary cataract
C1306068|T047|OAS|47337003|SNOMEDCT_CORE|Posterior capsular opacification|Secondary cataract
C1306068|T047|SY|766834007|SNOMEDCT_CORE|Posterior capsular opacification|Secondary cataract
C1306068|T047|IS|47337003|SNOMEDCT_CORE|Secondary cataract|Secondary cataract
C1306068|T047|PT|766834007|SNOMEDCT_CORE|Secondary cataract|Secondary cataract
C1306068|T047|FN|766834007|SNOMEDCT_CORE|Secondary cataract|Secondary cataract
C1306265|T020|PT|62730001|SNOMEDCT_CORE|Female proctocele without uterine prolapse|Female proctocele without uterine prolapse
C1306265|T020|FN|62730001|SNOMEDCT_CORE|Female proctocele without uterine prolapse|Female proctocele without uterine prolapse
C1306265|T020|SY|62730001|SNOMEDCT_CORE|Female rectocele without uterine prolapse|Female proctocele without uterine prolapse
C1306274|T048|SY|89765005|SNOMEDCT_CORE|Tabagism|Tabagism
C1306310|T191|PT|94098005|SNOMEDCT_CORE|Primary malignant neoplasm of thyroid gland|Primary malignant neoplasm of thyroid gland
C1306310|T191|FN|94098005|SNOMEDCT_CORE|Primary malignant neoplasm of thyroid gland|Primary malignant neoplasm of thyroid gland
C1306339|T048|IS|91138005|SNOMEDCT_CORE|Mental retardation, severity unspecified|Mental retardation, severity unspecified
C1306341|T048|IS|1855002|SNOMEDCT_CORE|Mental disability|Mental handicap
C1306341|T048|IS|1855002|SNOMEDCT_CORE|Mental handicap|Mental handicap
C1306341|T048|IS|1855002|SNOMEDCT_CORE|Mental impairment|Mental handicap
C1306341|T048|IS|1855002|SNOMEDCT_CORE|Mental subnormality|Mental handicap
C1306341|T048|IS|1855002|SNOMEDCT_CORE|MH - Mental handicap|Mental handicap
C1306460|T191|SY|93880001|SNOMEDCT_CORE|Lung cancer|Primary malignant neoplasm of lung
C1306460|T191|PT|93880001|SNOMEDCT_CORE|Primary malignant neoplasm of lung|Primary malignant neoplasm of lung
C1306460|T191|FN|93880001|SNOMEDCT_CORE|Primary malignant neoplasm of lung|Primary malignant neoplasm of lung
C1306468|T191|PT|93934004|SNOMEDCT_CORE|Primary malignant neoplasm of ovary|Primary malignant neoplasm of ovary
C1306468|T191|FN|93934004|SNOMEDCT_CORE|Primary malignant neoplasm of ovary|Primary malignant neoplasm of ovary
C1306503|T019|OAP|5867007|SNOMEDCT_CORE|Congenital exomphalos|Congenital exomphalos
C1306503|T019|OAF|5867007|SNOMEDCT_CORE|Congenital exomphalos|Congenital exomphalos
C1306503|T019|SY|396347007|SNOMEDCT_CORE|Exomphalos|Congenital exomphalos
C1306503|T019|SY|396347007|SNOMEDCT_CORE|Exumbilication|Congenital exomphalos
C1306557|T047|SY|20696009|SNOMEDCT_CORE|Chronic venous insufficiency|Chronic venous insufficiency
C1306557|T047|IS|20696009|SNOMEDCT_CORE|Chronic venous insufficiency, NOS|Chronic venous insufficiency
C1306571|T046|SY|59927004|SNOMEDCT_CORE|Hepatic insufficiency|Hepatic insufficiency
C1306571|T046|IS|59927004|SNOMEDCT_CORE|Hepatic insufficiency, NOS|Hepatic insufficiency
C1306578|T047|SY|23560001|SNOMEDCT_CORE|Schizoid disorder of childhood|Schizoid disorder of childhood
C1306587|T047|IS|2776000|SNOMEDCT_CORE|Acute encephalopathy|Acute encephalopathy
C1306587|T047|IS|2776000|SNOMEDCT_CORE|Acute encephalopathy, NOS|Acute encephalopathy
C1306588|T048|SY|2776000|SNOMEDCT_CORE|Acute organic reaction|Acute psycho-organic syndrome
C1306588|T048|SY|2776000|SNOMEDCT_CORE|Acute psycho-organic syndrome|Acute psycho-organic syndrome
C1306600|T047|IS|16644004|SNOMEDCT_CORE|Radial nerve palsy|Radial nerve palsy
C1306601|T047|SY|398114001|SNOMEDCT_CORE|Dermatorrhexis with dermatochalasis AND arthrochalasis|Dermatorrhexis with dermatochalasis AND arthrochalasis
C1306835|T047|SY|399114005|SNOMEDCT_CORE|Periarthritis of shoulder|Periarthritis of shoulder
C1306838|T047|SY|69896004|SNOMEDCT_CORE|Proliferative arthritis|Proliferative arthritis
C1306848|T047|IS|36989005|SNOMEDCT_CORE|Mumps without mention of complication|Mumps without mention of complication
C1306869|T191|SY|266569009|SNOMEDCT_CORE|Benign fibroma of prostate|Benign fibroma of prostate
C1306871|T191|SY|266569009|SNOMEDCT_CORE|Benign myoma of prostate|Benign myoma of prostate
C1306879|T037|SY|127287001|SNOMEDCT_CORE|Extracapsular fracture of neck of femur|Trochanteric fracture of neck of femur
C1306879|T037|SY|127287001|SNOMEDCT_CORE|Trochanteric fracture of neck of femur|Trochanteric fracture of neck of femur
C1306889|T047|SY|399957001|SNOMEDCT_CORE|PAD - Peripheral arterial disease|Peripheral arterial occlusive disease
C1306889|T047|SY|399957001|SNOMEDCT_CORE|PAOD - Peripheral arterial occlusive disease|Peripheral arterial occlusive disease
C1306889|T047|PT|399957001|SNOMEDCT_CORE|Peripheral arterial occlusive disease|Peripheral arterial occlusive disease
C1306889|T047|FN|399957001|SNOMEDCT_CORE|Peripheral arterial occlusive disease|Peripheral arterial occlusive disease
C1306889|T047|SY|399957001|SNOMEDCT_CORE|Peripheral artery occlusive disease|Peripheral arterial occlusive disease
C1313876|T033|PT|189445003|SNOMEDCT_CORE|Light-for-dates without fetal malnutrition|Light-for-dates without fetal malnutrition
C1313876|T033|FN|189445003|SNOMEDCT_CORE|Light-for-dates without fetal malnutrition|Light-for-dates without fetal malnutrition
C1313876|T033|SY|189445003|SNOMEDCT_CORE|Light-for-dates without foetal malnutrition|Light-for-dates without fetal malnutrition
C1313876|T033|IS|189445003|SNOMEDCT_CORE|Light-for-dates without mention of fetal malnutrition|Light-for-dates without fetal malnutrition
C1313937|T033|PT|160303001|SNOMEDCT_CORE|Family history of diabetes mellitus|Family history of diabetes mellitus
C1313937|T033|FN|160303001|SNOMEDCT_CORE|Family history of diabetes mellitus|Family history of diabetes mellitus
C1313937|T033|SY|160303001|SNOMEDCT_CORE|Family history: Diabetes mellitus|Family history of diabetes mellitus
C1313937|T033|OF|160303001|SNOMEDCT_CORE|Family history: Diabetes mellitus|Family history of diabetes mellitus
C1313937|T033|SY|160303001|SNOMEDCT_CORE|FH: Diabetes mellitus|Family history of diabetes mellitus
C1313946|T047|SY|91487003|SNOMEDCT_CORE|Urine-induced contact dermatitis|Urine-induced contact dermatitis
C1313967|T033|PTGB|185903001|SNOMEDCT_CORE|Needs influenza immunisation|Needs influenza immunization
C1313967|T033|PT|185903001|SNOMEDCT_CORE|Needs influenza immunization|Needs influenza immunization
C1313967|T033|FN|185903001|SNOMEDCT_CORE|Needs influenza immunization|Needs influenza immunization
C1313980|T033|PTGB|297242006|SNOMEDCT_CORE|Family history of ischaemic heart disease|Family history of ischemic heart disease
C1313980|T033|PT|297242006|SNOMEDCT_CORE|Family history of ischemic heart disease|Family history of ischemic heart disease
C1313980|T033|OF|297242006|SNOMEDCT_CORE|Family history of ischemic heart disease|Family history of ischemic heart disease
C1313980|T033|FN|297242006|SNOMEDCT_CORE|Family history of ischemic heart disease|Family history of ischemic heart disease
C1313980|T033|SYGB|297242006|SNOMEDCT_CORE|FH: Ischaemic heart disease|Family history of ischemic heart disease
C1313980|T033|SY|297242006|SNOMEDCT_CORE|FH: Ischemic heart disease|Family history of ischemic heart disease
C1313983|T047|OAP|240066005|SNOMEDCT_CORE|Acute contagious conjunctivitis|Acute contagious conjunctivitis
C1313983|T047|OAF|240066005|SNOMEDCT_CORE|Acute contagious conjunctivitis|Acute contagious conjunctivitis
C1313984|T033|SY|266997008|SNOMEDCT_CORE|H/O: intestinal disease|H/O: intestinal disease
C1314667|T191|PT|93980002|SNOMEDCT_CORE|Primary malignant neoplasm of rectosigmoid junction|Primary malignant neoplasm of rectosigmoid junction
C1314667|T191|FN|93980002|SNOMEDCT_CORE|Primary malignant neoplasm of rectosigmoid junction|Primary malignant neoplasm of rectosigmoid junction
C1314696|T191|SY|254622008|SNOMEDCT_CORE|SCC - Squamous cell carcinoma of bronchus|Squamous cell carcinoma of bronchus
C1314696|T191|PT|254622008|SNOMEDCT_CORE|Squamous cell carcinoma of bronchus|Squamous cell carcinoma of bronchus
C1314696|T191|FN|254622008|SNOMEDCT_CORE|Squamous cell carcinoma of bronchus|Squamous cell carcinoma of bronchus
C1314741|T191|IS|419603000|SNOMEDCT_CORE|Steatoma|Steatoma
C1314752|T047|IS|48194001|SNOMEDCT_CORE|Hypertension complicating childbirth|Hypertension complicating childbirth
C1314753|T046|IS|48194001|SNOMEDCT_CORE|Hypertension complicating pregnancy|Hypertension complicating pregnancy
C1314769|T047|IS|39629007|SNOMEDCT_CORE|Septic granuloma of skin|Septic granuloma of skin
C1318500|T047|PT|190236006|SNOMEDCT_CORE|Non-toxic nodular goiter|Non-toxic nodular goiter
C1318500|T047|FN|190236006|SNOMEDCT_CORE|Non-toxic nodular goiter|Non-toxic nodular goiter
C1318500|T047|PTGB|190236006|SNOMEDCT_CORE|Non-toxic nodular goitre|Non-toxic nodular goiter
C1318500|T047|SY|190236006|SNOMEDCT_CORE|Nontoxic nodular thyroid goiter|Non-toxic nodular goiter
C1318500|T047|SYGB|190236006|SNOMEDCT_CORE|Nontoxic nodular thyroid goitre|Non-toxic nodular goiter
C1318518|T019|SY|367489004|SNOMEDCT_CORE|Autosomal recessive lethal osteopetrosis|Infantile malignant osteopetrosis
C1318518|T019|SY|367489004|SNOMEDCT_CORE|Autosomal recessive malignant osteopetrosis|Infantile malignant osteopetrosis
C1318518|T019|PT|367489004|SNOMEDCT_CORE|Infantile malignant osteopetrosis|Infantile malignant osteopetrosis
C1318518|T019|FN|367489004|SNOMEDCT_CORE|Infantile malignant osteopetrosis|Infantile malignant osteopetrosis
C1318518|T019|IS|367489004|SNOMEDCT_CORE|Osteopetrosis - precocious type|Infantile malignant osteopetrosis
C1318518|T019|IS|367489004|SNOMEDCT_CORE|Severe osteopetrosis|Infantile malignant osteopetrosis
C1318520|T047|PTGB|11791001|SNOMEDCT_CORE|Necrotising vasculitis|Necrotizing vasculitis
C1318520|T047|PT|11791001|SNOMEDCT_CORE|Necrotizing vasculitis|Necrotizing vasculitis
C1318520|T047|FN|11791001|SNOMEDCT_CORE|Necrotizing vasculitis|Necrotizing vasculitis
C1318520|T047|IS|11791001|SNOMEDCT_CORE|Necrotizing vasculitis, NOS|Necrotizing vasculitis
C1318533|T047|SYGB|44865000|SNOMEDCT_CORE|Acquired polycythaemia|Secondary polycythemia
C1318533|T047|IS|44865000|SNOMEDCT_CORE|Acquired polycythaemia, NOS|Secondary polycythemia
C1318533|T047|SY|44865000|SNOMEDCT_CORE|Acquired polycythemia|Secondary polycythemia
C1318533|T047|IS|44865000|SNOMEDCT_CORE|Acquired polycythemia, NOS|Secondary polycythemia
C1318533|T047|SY|44865000|SNOMEDCT_CORE|Secondary erythrocytosis|Secondary polycythemia
C1318533|T047|IS|44865000|SNOMEDCT_CORE|Secondary erythrocytosis, NOS|Secondary polycythemia
C1318533|T047|PTGB|44865000|SNOMEDCT_CORE|Secondary polycythaemia|Secondary polycythemia
C1318533|T047|IS|44865000|SNOMEDCT_CORE|Secondary polycythaemia, NOS|Secondary polycythemia
C1318533|T047|PT|44865000|SNOMEDCT_CORE|Secondary polycythemia|Secondary polycythemia
C1318533|T047|FN|44865000|SNOMEDCT_CORE|Secondary polycythemia|Secondary polycythemia
C1318533|T047|IS|44865000|SNOMEDCT_CORE|Secondary polycythemia, NOS|Secondary polycythemia
C1318543|T191|PT|310605004|SNOMEDCT_CORE|Fibrous histiocytoma of tendon sheath|Fibrous histiocytoma of tendon sheath
C1318543|T191|FN|310605004|SNOMEDCT_CORE|Fibrous histiocytoma of tendon sheath|Fibrous histiocytoma of tendon sheath
C1318558|T191|SYGB|398696001|SNOMEDCT_CORE|Congenital melanocytic naevus|Congenital pigmented melanocytic nevus
C1318558|T191|SY|398696001|SNOMEDCT_CORE|Congenital melanocytic nevus|Congenital pigmented melanocytic nevus
C1318558|T191|PTGB|398696001|SNOMEDCT_CORE|Congenital pigmented melanocytic naevus|Congenital pigmented melanocytic nevus
C1318558|T191|FN|398696001|SNOMEDCT_CORE|Congenital pigmented melanocytic nevus|Congenital pigmented melanocytic nevus
C1318558|T191|PT|398696001|SNOMEDCT_CORE|Congenital pigmented melanocytic nevus|Congenital pigmented melanocytic nevus
C1318558|T191|SYGB|398696001|SNOMEDCT_CORE|Congenital pigmented naevus|Congenital pigmented melanocytic nevus
C1318558|T191|SY|398696001|SNOMEDCT_CORE|Congenital pigmented nevus|Congenital pigmented melanocytic nevus
C1318710|T047|SY|407450002|SNOMEDCT_CORE|Herpes simplex 2|Herpes simplex type 2 infection
C1318710|T047|SY|407450002|SNOMEDCT_CORE|Herpes simplex 2 infection|Herpes simplex type 2 infection
C1318710|T047|PT|407450002|SNOMEDCT_CORE|Herpes simplex type 2 infection|Herpes simplex type 2 infection
C1318710|T047|FN|407450002|SNOMEDCT_CORE|Herpes simplex type 2 infection|Herpes simplex type 2 infection
C1318710|T047|IS|407450002|SNOMEDCT_CORE|Herpex simplex 2|Herpes simplex type 2 infection
C1318711|T047|SY|407451003|SNOMEDCT_CORE|Herpes simplex 1|Herpes simplex type 1 infection
C1318711|T047|SY|407451003|SNOMEDCT_CORE|Herpes simplex 1 infection|Herpes simplex type 1 infection
C1318711|T047|PT|407451003|SNOMEDCT_CORE|Herpes simplex type 1 infection|Herpes simplex type 1 infection
C1318711|T047|FN|407451003|SNOMEDCT_CORE|Herpes simplex type 1 infection|Herpes simplex type 1 infection
C1319000|T047|SY|405633009|SNOMEDCT_CORE|Infantile group B strep infection|Streptococcus group B infection of the infant
C1319000|T047|PT|405633009|SNOMEDCT_CORE|Streptococcus group B infection of the infant|Streptococcus group B infection of the infant
C1319000|T047|FN|405633009|SNOMEDCT_CORE|Streptococcus group B infection of the infant|Streptococcus group B infection of the infant
C1319018|T047|PT|405944004|SNOMEDCT_CORE|Asthmatic bronchitis|Asthmatic bronchitis
C1319018|T047|FN|405944004|SNOMEDCT_CORE|Asthmatic bronchitis|Asthmatic bronchitis
C1319018|T047|IS|405944004|SNOMEDCT_CORE|Wheezy bronchitis|Asthmatic bronchitis
C1319314|T191|PT|408642003|SNOMEDCT_CORE|Transitional cell carcinoma of kidney|Transitional cell carcinoma of kidney
C1319314|T191|FN|408642003|SNOMEDCT_CORE|Transitional cell carcinoma of kidney|Transitional cell carcinoma of kidney
C1319315|T191|PT|408645001|SNOMEDCT_CORE|Adenocarcinoma of large intestine|Adenocarcinoma of large intestine
C1319315|T191|FN|408645001|SNOMEDCT_CORE|Adenocarcinoma of large intestine|Adenocarcinoma of large intestine
C1319321|T033|PT|408546009|SNOMEDCT_CORE|Coronary artery bypass graft occlusion|Coronary artery bypass graft occlusion
C1319321|T033|FN|408546009|SNOMEDCT_CORE|Coronary artery bypass graft occlusion|Coronary artery bypass graft occlusion
C1319384|T047|PT|408418009|SNOMEDCT_CORE|Upper airway resistance syndrome|Upper airway resistance syndrome
C1319384|T047|FN|408418009|SNOMEDCT_CORE|Upper airway resistance syndrome|Upper airway resistance syndrome
C1319441|T033|SY|408512008|SNOMEDCT_CORE|Body mass index 40+ - morbidly obese|Body mass index 40+ - severely obese
C1319441|T033|PT|408512008|SNOMEDCT_CORE|Body mass index 40+ - severely obese|Body mass index 40+ - severely obese
C1319441|T033|FN|408512008|SNOMEDCT_CORE|Body mass index 40+ - severely obese|Body mass index 40+ - severely obese
C1319441|T033|SY|408512008|SNOMEDCT_CORE|Obese class III|Body mass index 40+ - severely obese
C1319851|T033|FN|407669000|SNOMEDCT_CORE|Magnetic resonance imaging of brain abnormal|Magnetic resonance imaging of brain abnormal
C1319851|T033|PT|407669000|SNOMEDCT_CORE|Magnetic resonance imaging of brain abnormal|Magnetic resonance imaging of brain abnormal
C1319898|T033|PT|407560009|SNOMEDCT_CORE|At risk of sexually transmitted infection|At risk of sexually transmitted infection
C1319898|T033|FN|407560009|SNOMEDCT_CORE|At risk of sexually transmitted infection|At risk of sexually transmitted infection
C1320640|T047|OAF|405721006|SNOMEDCT_CORE|Peripheral degeneration of retina|Peripheral retinal degeneration
C1320640|T047|OAP|405721006|SNOMEDCT_CORE|Peripheral degeneration of retina|Peripheral retinal degeneration
C1320640|T047|SY|61536007|SNOMEDCT_CORE|Peripheral degeneration of retina|Peripheral retinal degeneration
C1320640|T047|PT|61536007|SNOMEDCT_CORE|Peripheral retinal degeneration|Peripheral retinal degeneration
C1320640|T047|FN|61536007|SNOMEDCT_CORE|Peripheral retinal degeneration|Peripheral retinal degeneration
C1320640|T047|IS|61536007|SNOMEDCT_CORE|Peripheral retinal degeneration, NOS|Peripheral retinal degeneration
C1320654|T033|PT|405748007|SNOMEDCT_CORE|Already on aspirin|Already on aspirin
C1320654|T033|FN|405748007|SNOMEDCT_CORE|Already on aspirin|Already on aspirin
C1320835|T046|SY|405543000|SNOMEDCT_CORE|Drug fever|Drug-induced hyperpyrexia
C1320835|T046|PT|405543000|SNOMEDCT_CORE|Drug-induced hyperpyrexia|Drug-induced hyperpyrexia
C1320835|T046|FN|405543000|SNOMEDCT_CORE|Drug-induced hyperpyrexia|Drug-induced hyperpyrexia
C1320845|T047|PT|405557003|SNOMEDCT_CORE|Occlusion of lower limb artery|Occlusion of lower limb artery
C1320845|T047|FN|405557003|SNOMEDCT_CORE|Occlusion of lower limb artery|Occlusion of lower limb artery
C1321321|T047|PT|404670008|SNOMEDCT_CORE|Cholesterol retinal embolus|Cholesterol retinal embolus
C1321321|T047|FN|404670008|SNOMEDCT_CORE|Cholesterol retinal embolus|Cholesterol retinal embolus
C1321321|T047|SY|404670008|SNOMEDCT_CORE|Hollenhorst plaque|Cholesterol retinal embolus
C1321782|T047|IS|46764007|SNOMEDCT_CORE|Gestosis|Gestosis
C1321896|T037|IS|25604001|SNOMEDCT_CORE|Injury of peroneal nerve|Peroneal nerve injury
C1321896|T037|SY|212317001|SNOMEDCT_CORE|Injury of peroneal nerve|Peroneal nerve injury
C1321896|T037|FN|212317001|SNOMEDCT_CORE|Injury of peroneal nerve|Peroneal nerve injury
C1321896|T037|PT|212317001|SNOMEDCT_CORE|Peroneal nerve injury|Peroneal nerve injury
C1321896|T037|OF|212317001|SNOMEDCT_CORE|Peroneal nerve injury|Peroneal nerve injury
C1321898|T184|IS|2901004|SNOMEDCT_CORE|Blood in stool|Blood in stool
C1321905|T048|SY|406506008|SNOMEDCT_CORE|MBD - Minimal brain dysfunction|MBD - Minimal brain dysfunction
C1321905|T048|SY|406506008|SNOMEDCT_CORE|Minimal brain dysfunction|MBD - Minimal brain dysfunction
C1328248|T047|SY|196341005|SNOMEDCT_CORE|Alveolar abscess|Alveolar abscess
C1328479|T191|PT|254612002|SNOMEDCT_CORE|Carcinoma of endocrine pancreas|Carcinoma of endocrine pancreas
C1328479|T191|FN|254612002|SNOMEDCT_CORE|Carcinoma of endocrine pancreas|Carcinoma of endocrine pancreas
C1328479|T191|SY|254612002|SNOMEDCT_CORE|Endocrine pancreatic carcinoma|Carcinoma of endocrine pancreas
C1328971|T047|IS|70218004|SNOMEDCT_CORE|Discogenic syndrome, NOS|Displacement of intervertebral disc without myelopathy
C1328971|T047|PT|70218004|SNOMEDCT_CORE|Displacement of intervertebral disc without myelopathy|Displacement of intervertebral disc without myelopathy
C1328971|T047|FN|70218004|SNOMEDCT_CORE|Displacement of intervertebral disc without myelopathy|Displacement of intervertebral disc without myelopathy
C1328971|T047|IS|70218004|SNOMEDCT_CORE|Displacement of intervertebral disc, site unspecified without myelopathy|Displacement of intervertebral disc without myelopathy
C1330959|T191|PT|93974005|SNOMEDCT_CORE|Primary malignant neoplasm of prostate|Primary malignant neoplasm of prostate
C1330959|T191|FN|93974005|SNOMEDCT_CORE|Primary malignant neoplasm of prostate|Primary malignant neoplasm of prostate
C1330966|T033|PT|1855002|SNOMEDCT_CORE|Developmental academic disorder|Developmental academic disorder
C1330966|T033|FN|1855002|SNOMEDCT_CORE|Developmental academic disorder|Developmental academic disorder
C1330966|T033|IS|1855002|SNOMEDCT_CORE|Developmental academic disorder, NOS|Developmental academic disorder
C1330966|T033|SY|1855002|SNOMEDCT_CORE|Developmental disorder of scholastic skill|Developmental academic disorder
C1331537|T047|SY|67754003|SNOMEDCT_CORE|Aortic sclerosis|Aortic sclerosis
C1331543|T047|PT|237348005|SNOMEDCT_CORE|Puerperal pyrexia|Puerperal pyrexia
C1331543|T047|FN|237348005|SNOMEDCT_CORE|Puerperal pyrexia|Puerperal pyrexia
C1331979|T046|SY|81642009|SNOMEDCT_CORE|Sequelae of injury of spinal cord|Sequelae of injury of spinal cord
C1331981|T046|SY|110270004|SNOMEDCT_CORE|Sequelae of poliomyelitis|Sequelae of poliomyelitis
C1333990|T191|SY|315058005|SNOMEDCT_CORE|Hereditary nonpolyposis colon cancer|HNPCC - hereditary nonpolyposis colon cancer
C1333990|T191|FN|315058005|SNOMEDCT_CORE|Hereditary nonpolyposis colon cancer|HNPCC - hereditary nonpolyposis colon cancer
C1333990|T191|PT|315058005|SNOMEDCT_CORE|HNPCC - hereditary nonpolyposis colon cancer|HNPCC - hereditary nonpolyposis colon cancer
C1333990|T191|SY|315058005|SNOMEDCT_CORE|HNPCC - hereditary nonpolyposis colorectal cancer|HNPCC - hereditary nonpolyposis colon cancer
C1334177|T191|SY|423973006|SNOMEDCT_CORE|Cancer of uterine cervix, invasive|Carcinoma of uterine cervix, invasive
C1334177|T191|FN|423973006|SNOMEDCT_CORE|Carcinoma of uterine cervix, invasive|Carcinoma of uterine cervix, invasive
C1334177|T191|PT|423973006|SNOMEDCT_CORE|Carcinoma of uterine cervix, invasive|Carcinoma of uterine cervix, invasive
C1334177|T191|SY|423973006|SNOMEDCT_CORE|Invasive cervical cancer|Carcinoma of uterine cervix, invasive
C1334237|T191|PTGB|445513004|SNOMEDCT_CORE|Intracranial cavernous haemangioma|Intracranial cavernous hemangioma
C1334237|T191|PT|445513004|SNOMEDCT_CORE|Intracranial cavernous hemangioma|Intracranial cavernous hemangioma
C1334237|T191|FN|445513004|SNOMEDCT_CORE|Intracranial cavernous hemangioma|Intracranial cavernous hemangioma
C1337102|T033|SY|214264003|SNOMEDCT_CORE|Lack of vitality|Lack of vitality
C1363843|T047|SY|57534004|SNOMEDCT_CORE|Changes in retinal vascular appearance|Changes in retinal vascular appearance
C1367166|T037|SYGB|209987007|SNOMEDCT_CORE|Subdural haemorrhage following injury|Traumatic subdural hemorrhage
C1367166|T037|SY|209987007|SNOMEDCT_CORE|Subdural hemorrhage following injury|Traumatic subdural hemorrhage
C1367166|T037|PTGB|209987007|SNOMEDCT_CORE|Traumatic subdural haemorrhage|Traumatic subdural hemorrhage
C1367166|T037|PT|209987007|SNOMEDCT_CORE|Traumatic subdural hemorrhage|Traumatic subdural hemorrhage
C1367166|T037|OF|209987007|SNOMEDCT_CORE|Traumatic subdural hemorrhage|Traumatic subdural hemorrhage
C1367166|T037|SYGB|209987007|SNOMEDCT_CORE|Traumatic subdural intracranial haemorrhage|Traumatic subdural hemorrhage
C1367166|T037|SY|209987007|SNOMEDCT_CORE|Traumatic subdural intracranial hemorrhage|Traumatic subdural hemorrhage
C1367166|T037|FN|209987007|SNOMEDCT_CORE|Traumatic subdural intracranial hemorrhage|Traumatic subdural hemorrhage
C1367974|T047|IS|34250006|SNOMEDCT_CORE|Benign mucous membrane pemphigoid without ocular involvement|Benign mucous membrane pemphigoid without ocular involvement
C1368020|T047|SY|67782005|SNOMEDCT_CORE|Post-traumatic pulmonary insufficiency|Pulmonary insufficiency following trauma
C1368020|T047|IS|67782005|SNOMEDCT_CORE|Pulmonary insufficiency following trauma|Pulmonary insufficiency following trauma
C1368020|T047|SY|67782005|SNOMEDCT_CORE|Traumatic wet lung|Pulmonary insufficiency following trauma
C1368021|T047|IS|67782005|SNOMEDCT_CORE|Pulmonary insufficiency following shock|Pulmonary insufficiency following shock
C1368022|T046|IS|67782005|SNOMEDCT_CORE|Pulmonary insufficiency following surgery|Pulmonary insufficiency following surgery
C1370500|T191|IS|57706008|SNOMEDCT_CORE|Tanycytic ependymoma|Tanycytic ependymoma
C1370867|T037|PT|17383000|SNOMEDCT_CORE|Toxic effect of carbon monoxide|Toxic effect of carbon monoxide
C1370867|T037|FN|17383000|SNOMEDCT_CORE|Toxic effect of carbon monoxide|Toxic effect of carbon monoxide
C1378703|T191|IS|254915003|SNOMEDCT_CORE|Carcinoma of kidney|Carcinoma of kidney
C1383860|T046|IS|8186001|SNOMEDCT_CORE|Cardiac hypertrophy|Cardiac hypertrophy
C1384403|T191|IS|57706008|SNOMEDCT_CORE|Cellular ependymoma|Clear cell ependymoma
C1384403|T191|IS|57706008|SNOMEDCT_CORE|Clear cell ependymoma|Clear cell ependymoma
C1384457|T020|PT|240244006|SNOMEDCT_CORE|Acquired deformity of joint of foot|Acquired deformity of joint of foot
C1384457|T020|FN|240244006|SNOMEDCT_CORE|Acquired deformity of joint of foot|Acquired deformity of joint of foot
C1384485|T033|PT|48782003|SNOMEDCT_CORE|Delivery normal|Delivery normal
C1384485|T033|OF|48782003|SNOMEDCT_CORE|Delivery normal|Delivery normal
C1384485|T033|FN|48782003|SNOMEDCT_CORE|Delivery normal|Delivery normal
C1384485|T033|IS|48782003|SNOMEDCT_CORE|Delivery of fetus, completely normal case|Delivery normal
C1384485|T033|SY|48782003|SNOMEDCT_CORE|FTND - Full term normal delivery|Delivery normal
C1384485|T033|SY|48782003|SNOMEDCT_CORE|Normal delivery|Delivery normal
C1384485|T033|SY|48782003|SNOMEDCT_CORE|Spontaneous vaginal delivery|Delivery normal
C1384485|T033|SY|48782003|SNOMEDCT_CORE|SVD - Spontaneous vaginal delivery|Delivery normal
C1384498|T047|PT|235651006|SNOMEDCT_CORE|Gastric erosion|Gastric erosion
C1384498|T047|FN|235651006|SNOMEDCT_CORE|Gastric erosion|Gastric erosion
C1384514|T047|SY|190507007|SNOMEDCT_CORE|Conn syndrome|Primary aldosteronism
C1384514|T047|SY|190507007|SNOMEDCT_CORE|Conn's syndrome|Primary aldosteronism
C1384514|T047|PT|190507007|SNOMEDCT_CORE|Primary aldosteronism|Primary aldosteronism
C1384514|T047|SY|190507007|SNOMEDCT_CORE|Primary hyperaldosteronism|Primary aldosteronism
C1384514|T047|FN|190507007|SNOMEDCT_CORE|Primary hyperaldosteronism|Primary aldosteronism
C1384582|T047|SY|370997001|SNOMEDCT_CORE|Primary failure of the testes|Primary testicular failure
C1384582|T047|SY|48723006|SNOMEDCT_CORE|Primary gonadal failure|Primary testicular failure
C1384582|T047|SY|48723006|SNOMEDCT_CORE|Primary male hypogonadism|Primary testicular failure
C1384582|T047|IS|48723006|SNOMEDCT_CORE|Primary testicular failure|Primary testicular failure
C1384582|T047|PT|370997001|SNOMEDCT_CORE|Primary testicular failure|Primary testicular failure
C1384582|T047|FN|370997001|SNOMEDCT_CORE|Primary testicular failure|Primary testicular failure
C1384584|T047|PT|201819000|SNOMEDCT_CORE|Degenerative joint disease involving multiple joints|Degenerative joint disease involving multiple joints
C1384584|T047|SYGB|201819000|SNOMEDCT_CORE|Generalised osteoarthritis|Degenerative joint disease involving multiple joints
C1384584|T047|SYGB|201819000|SNOMEDCT_CORE|Generalised osteoarthrosis|Degenerative joint disease involving multiple joints
C1384584|T047|SY|201819000|SNOMEDCT_CORE|Generalized osteoarthritis|Degenerative joint disease involving multiple joints
C1384584|T047|FN|201819000|SNOMEDCT_CORE|Generalized osteoarthritis|Degenerative joint disease involving multiple joints
C1384584|T047|SY|201819000|SNOMEDCT_CORE|Generalized osteoarthrosis|Degenerative joint disease involving multiple joints
C1384584|T047|SYGB|201819000|SNOMEDCT_CORE|GOA - Generalised osteoarthritis|Degenerative joint disease involving multiple joints
C1384584|T047|SY|201819000|SNOMEDCT_CORE|GOA - Generalized osteoarthritis|Degenerative joint disease involving multiple joints
C1384584|T047|SY|201819000|SNOMEDCT_CORE|Polyarticular osteoarthritis|Degenerative joint disease involving multiple joints
C1384589|T047|PT|399029005|SNOMEDCT_CORE|Tinea cruris|Tinea cruris
C1384589|T047|FN|399029005|SNOMEDCT_CORE|Tinea cruris|Tinea cruris
C1384600|T047|SY|201796004|SNOMEDCT_CORE|Juvenile arthritis with systemic onset|Systemic onset juvenile chronic arthritis
C1384600|T047|SY|201796004|SNOMEDCT_CORE|Systemic juvenile idiopathic arthritis|Systemic onset juvenile chronic arthritis
C1384600|T047|PT|201796004|SNOMEDCT_CORE|Systemic onset juvenile chronic arthritis|Systemic onset juvenile chronic arthritis
C1384600|T047|FN|201796004|SNOMEDCT_CORE|Systemic onset juvenile chronic arthritis|Systemic onset juvenile chronic arthritis
C1384600|T047|SY|201796004|SNOMEDCT_CORE|Systemic onset juvenile rheumatoid arthritis|Systemic onset juvenile chronic arthritis
C1384641|T047|PT|387800004|SNOMEDCT_CORE|Cervical spondylosis|Cervical spondylosis
C1384641|T047|FN|387800004|SNOMEDCT_CORE|Cervical spondylosis|Cervical spondylosis
C1384641|T047|SY|387800004|SNOMEDCT_CORE|CS - Cervical spondylosis|Cervical spondylosis
C1384666|T047|PT|103276001|SNOMEDCT_CORE|Decreased hearing|Hearing loss
C1384666|T047|FN|103276001|SNOMEDCT_CORE|Decreased hearing|Hearing loss
C1384666|T047|SY|15188001|SNOMEDCT_CORE|Difficulty hearing|Hearing loss
C1384666|T047|SY|15188001|SNOMEDCT_CORE|Hard of hearing|Hearing loss
C1384666|T047|SY|15188001|SNOMEDCT_CORE|Hearing impaired|Hearing loss
C1384666|T047|SY|15188001|SNOMEDCT_CORE|Hearing impairment|Hearing loss
C1384666|T047|PT|15188001|SNOMEDCT_CORE|Hearing loss|Hearing loss
C1384666|T047|OF|15188001|SNOMEDCT_CORE|Hearing loss|Hearing loss
C1384666|T047|FN|15188001|SNOMEDCT_CORE|Hearing loss|Hearing loss
C1384666|T047|IS|15188001|SNOMEDCT_CORE|Hearing loss, NOS|Hearing loss
C1384666|T047|SY|15188001|SNOMEDCT_CORE|HI - Hearing impairment|Hearing loss
C1384666|T047|SY|15188001|SNOMEDCT_CORE|HL - Hearing loss|Hearing loss
C1384666|T047|SY|15188001|SNOMEDCT_CORE|HOH - Hard of hearing|Hearing loss
C1384666|T047|SY|15188001|SNOMEDCT_CORE|Hypoacusis|Hearing loss
C1384666|T047|SY|15188001|SNOMEDCT_CORE|Impaired hearing|Hearing loss
C1384670|T019|SY|204470001|SNOMEDCT_CORE|Congenital absence of umbilical artery|Single umbilical artery
C1384670|T019|PT|204470001|SNOMEDCT_CORE|Single umbilical artery|Single umbilical artery
C1384670|T019|FN|204470001|SNOMEDCT_CORE|Single umbilical artery|Single umbilical artery
C1384674|T033|SYGB|200144004|SNOMEDCT_CORE|Caesarean delivery|Deliveries by cesarean
C1384674|T033|SY|200144004|SNOMEDCT_CORE|Cesarean delivery|Deliveries by cesarean
C1384674|T033|PTGB|200144004|SNOMEDCT_CORE|Deliveries by caesarean|Deliveries by cesarean
C1384674|T033|PT|200144004|SNOMEDCT_CORE|Deliveries by cesarean|Deliveries by cesarean
C1384674|T033|FN|200144004|SNOMEDCT_CORE|Deliveries by cesarean|Deliveries by cesarean
C1387400|T033|SY|415077006|SNOMEDCT_CORE|H/O: malignant neoplasm of bronchus|History of malignant neoplasm of bronchus
C1387400|T033|PT|415077006|SNOMEDCT_CORE|History of malignant neoplasm of bronchus|History of malignant neoplasm of bronchus
C1387400|T033|OF|415077006|SNOMEDCT_CORE|Personal history of primary malignant neoplasm of bronchus|History of malignant neoplasm of bronchus
C1387400|T033|SY|415077006|SNOMEDCT_CORE|Personal history of primary malignant neoplasm of bronchus|History of malignant neoplasm of bronchus
C1387400|T033|FN|415077006|SNOMEDCT_CORE|Personal history of primary malignant neoplasm of bronchus|History of malignant neoplasm of bronchus
C1387403|T033|OAS|415084003|SNOMEDCT_CORE|H/O: malignant neoplasm of skin|History of malignant neoplasm of skin
C1387403|T033|OAS|415084003|SNOMEDCT_CORE|H/O: primary malignant neoplasm of skin|History of malignant neoplasm of skin
C1387403|T033|OAP|415084003|SNOMEDCT_CORE|History of malignant neoplasm of skin|History of malignant neoplasm of skin
C1387403|T033|OAS|415084003|SNOMEDCT_CORE|Personal history of primary malignant neoplasm of skin|History of malignant neoplasm of skin
C1387403|T033|OF|415084003|SNOMEDCT_CORE|Personal history of primary malignant neoplasm of skin|History of malignant neoplasm of skin
C1387403|T033|OAF|415084003|SNOMEDCT_CORE|Personal history of primary malignant neoplasm of skin|History of malignant neoplasm of skin
C1387404|T033|SY|415082004|SNOMEDCT_CORE|H/O: malignant neoplasm of lung|History of malignant neoplasm of lung
C1387404|T033|PT|415082004|SNOMEDCT_CORE|History of malignant neoplasm of lung|History of malignant neoplasm of lung
C1387404|T033|OF|415082004|SNOMEDCT_CORE|Personal history of primary malignant neoplasm of lung|History of malignant neoplasm of lung
C1387404|T033|SY|415082004|SNOMEDCT_CORE|Personal history of primary malignant neoplasm of lung|History of malignant neoplasm of lung
C1387404|T033|FN|415082004|SNOMEDCT_CORE|Personal history of primary malignant neoplasm of lung|History of malignant neoplasm of lung
C1387407|T033|IS|415076002|SNOMEDCT_CORE|H/O: malignant neoplasm of breast|Personal history of primary malignant neoplasm of breast
C1387407|T033|IS|415076002|SNOMEDCT_CORE|History of malignant neoplasm of breast|Personal history of primary malignant neoplasm of breast
C1387407|T033|PT|415076002|SNOMEDCT_CORE|Personal history of primary malignant neoplasm of breast|Personal history of primary malignant neoplasm of breast
C1387407|T033|OF|415076002|SNOMEDCT_CORE|Personal history of primary malignant neoplasm of breast|Personal history of primary malignant neoplasm of breast
C1387407|T033|FN|415076002|SNOMEDCT_CORE|Personal history of primary malignant neoplasm of breast|Personal history of primary malignant neoplasm of breast
C1387408|T033|SY|415081006|SNOMEDCT_CORE|H/O: malignant neoplasm of kidney|History of malignant neoplasm of kidney
C1387408|T033|PT|415081006|SNOMEDCT_CORE|History of malignant neoplasm of kidney|History of malignant neoplasm of kidney
C1387408|T033|OF|415081006|SNOMEDCT_CORE|Personal history of primary malignant neoplasm of kidney|History of malignant neoplasm of kidney
C1387408|T033|SY|415081006|SNOMEDCT_CORE|Personal history of primary malignant neoplasm of kidney|History of malignant neoplasm of kidney
C1387408|T033|FN|415081006|SNOMEDCT_CORE|Personal history of primary malignant neoplasm of kidney|History of malignant neoplasm of kidney
C1389527|T047|PT|444599008|SNOMEDCT_CORE|Relaxation of pelvic floor|Relaxation of pelvic floor
C1389527|T047|FN|444599008|SNOMEDCT_CORE|Relaxation of pelvic floor|Relaxation of pelvic floor
C1389941|T047|PT|427482006|SNOMEDCT_CORE|Flaccid neurogenic bladder|Flaccid neurogenic bladder
C1389941|T047|FN|427482006|SNOMEDCT_CORE|Flaccid neurogenic bladder|Flaccid neurogenic bladder
C1389941|T047|SY|427482006|SNOMEDCT_CORE|Flaccid neuropathic bladder|Flaccid neurogenic bladder
C1394494|T047|SY|252005008|SNOMEDCT_CORE|Bladder cystocele|Cystocele
C1394494|T047|PT|252005008|SNOMEDCT_CORE|Cystocele|Cystocele
C1394494|T047|OF|252005008|SNOMEDCT_CORE|Cystocele|Cystocele
C1394494|T047|SY|252005008|SNOMEDCT_CORE|Female cystocele|Cystocele
C1394494|T047|FN|252005008|SNOMEDCT_CORE|Female cystocele|Cystocele
C1394494|T047|SY|252005008|SNOMEDCT_CORE|Vaginal cystocele|Cystocele
C1395852|T019|SY|205135003|SNOMEDCT_CORE|Accessory thumb|Accessory thumb
C1399226|T047|SY|33413000|SNOMEDCT_CORE|Ectopic rhythm abnormality|Ectopic rhythm abnormality
C1399226|T047|IS|33413000|SNOMEDCT_CORE|Ectopic rhythm disorder|Ectopic rhythm abnormality
C1399729|T033|PT|432525007|SNOMEDCT_CORE|Mass of head|Mass of head
C1399729|T033|FN|432525007|SNOMEDCT_CORE|Mass of head|Mass of head
C1400137|T047|SY|418103007|SNOMEDCT_CORE|Enlarged lingual tonsil|Hypertrophy of lingual tonsil
C1400137|T047|PT|418103007|SNOMEDCT_CORE|Hypertrophy of lingual tonsil|Hypertrophy of lingual tonsil
C1400137|T047|FN|418103007|SNOMEDCT_CORE|Hypertrophy of lingual tonsil|Hypertrophy of lingual tonsil
C1402450|T046|SY|429656004|SNOMEDCT_CORE|Late effect of brain injury|Late effect of traumatic injury to brain
C1402450|T046|PT|429656004|SNOMEDCT_CORE|Late effect of traumatic injury to brain|Late effect of traumatic injury to brain
C1402450|T046|FN|429656004|SNOMEDCT_CORE|Late effect of traumatic injury to brain|Late effect of traumatic injury to brain
C1410927|T047|SY|419422001|SNOMEDCT_CORE|Angle narrow|Narrow angle
C1410927|T047|PT|419422001|SNOMEDCT_CORE|Narrow angle|Narrow angle
C1410927|T047|FN|419422001|SNOMEDCT_CORE|Narrow angle|Narrow angle
C1410927|T047|SY|419422001|SNOMEDCT_CORE|Narrow angle anterior chamber|Narrow angle
C1412002|T047|PT|233606009|SNOMEDCT_CORE|Atypical pneumonia|Atypical pneumonia
C1412002|T047|FN|233606009|SNOMEDCT_CORE|Atypical pneumonia|Atypical pneumonia
C1442826|T047|OF|206525008|SNOMEDCT_CORE|Neonatal necrotising enterocolitis|Neonatal necrotizing enterocolitis
C1442826|T047|PTGB|206525008|SNOMEDCT_CORE|Neonatal necrotising enterocolitis|Neonatal necrotizing enterocolitis
C1442826|T047|PT|206525008|SNOMEDCT_CORE|Neonatal necrotizing enterocolitis|Neonatal necrotizing enterocolitis
C1442826|T047|FN|206525008|SNOMEDCT_CORE|Neonatal necrotizing enterocolitis|Neonatal necrotizing enterocolitis
C1442826|T047|SYGB|206525008|SNOMEDCT_CORE|NNE - Neonatal necrotising enterocolitis|Neonatal necrotizing enterocolitis
C1442826|T047|SY|206525008|SNOMEDCT_CORE|NNE - Neonatal necrotizing enterocolitis|Neonatal necrotizing enterocolitis
C1442826|T047|SYGB|206525008|SNOMEDCT_CORE|NNEC - Neonatal necrotising enterocolitis|Neonatal necrotizing enterocolitis
C1442826|T047|SY|206525008|SNOMEDCT_CORE|NNEC - Neonatal necrotizing enterocolitis|Neonatal necrotizing enterocolitis
C1442835|T047|OAS|23346002|SNOMEDCT_CORE|Solar dermatitis|Solar dermatitis
C1442861|T033|SY|367423000|SNOMEDCT_CORE|Black eye|Black eye
C1442861|T033|IS|367423000|SNOMEDCT_CORE|Black eye, NOS|Black eye
C1442867|T047|IS|48210000|SNOMEDCT_CORE|Lumbar and sacral osteoarthritis|Lumbar and sacral osteoarthritis
C1442867|T047|IS|48210000|SNOMEDCT_CORE|Lumbar AND/OR sacral osteoarthritis|Lumbar and sacral osteoarthritis
C1442868|T047|SY|387800004|SNOMEDCT_CORE|Cervical spine degeneration|Cervical spine degeneration
C1442869|T047|SY|239880009|SNOMEDCT_CORE|Osteoarthritis of lumbar spine|Osteoarthritis of lumbar spine
C1442878|T047|IS|388982007|SNOMEDCT_CORE|Panaritium of toe|Panaritium of toe
C1442903|T047|PT|416189003|SNOMEDCT_CORE|Exostosis|Exostosis
C1442903|T047|FN|416189003|SNOMEDCT_CORE|Exostosis|Exostosis
C1442903|T047|SY|416189003|SNOMEDCT_CORE|Exostosis - disorder|Exostosis
C1442903|T047|SY|416189003|SNOMEDCT_CORE|Exostosis disorder|Exostosis
C1442913|T047|IS|79962008|SNOMEDCT_CORE|Barsony-Polgar syndrome|Barsony-Teschendorf syndrome
C1442913|T047|SY|79962008|SNOMEDCT_CORE|Barsony-Teschendorf syndrome|Barsony-Teschendorf syndrome
C1442915|T047|SY|79962008|SNOMEDCT_CORE|Corkscrew esophagus|Corkscrew esophagus
C1442915|T047|SYGB|79962008|SNOMEDCT_CORE|Corkscrew oesophagus|Corkscrew esophagus
C1442915|T047|SY|79962008|SNOMEDCT_CORE|Curling esophagus|Corkscrew esophagus
C1442915|T047|SYGB|79962008|SNOMEDCT_CORE|Curling oesophagus|Corkscrew esophagus
C1442915|T047|SY|79962008|SNOMEDCT_CORE|Curling of esophagus|Corkscrew esophagus
C1442915|T047|SYGB|79962008|SNOMEDCT_CORE|Curling of oesophagus|Corkscrew esophagus
C1442915|T047|SY|79962008|SNOMEDCT_CORE|Rosary bead esophagus|Corkscrew esophagus
C1442915|T047|SYGB|79962008|SNOMEDCT_CORE|Rosary bead oesophagus|Corkscrew esophagus
C1442916|T046|SY|79962008|SNOMEDCT_CORE|Pseudo-obstruction of the esophagus|Pseudo-obstruction of the esophagus
C1442916|T046|SYGB|79962008|SNOMEDCT_CORE|Pseudo-obstruction of the oesophagus|Pseudo-obstruction of the esophagus
C1442950|T047|SY|11049006|SNOMEDCT_CORE|Radicular syndrome of upper limbs|Radicular syndrome of upper limbs
C1442958|T047|IS|46795000|SNOMEDCT_CORE|Actinic porokeratosis|Actinic porokeratosis
C1442965|T047|SY|111255008|SNOMEDCT_CORE|Aseptic necrosis of capital femoral epiphysis|Avascular necrosis of the capital femoral epiphysis
C1442965|T047|PT|111255008|SNOMEDCT_CORE|Avascular necrosis of the capital femoral epiphysis|Avascular necrosis of the capital femoral epiphysis
C1442965|T047|FN|111255008|SNOMEDCT_CORE|Avascular necrosis of the capital femoral epiphysis|Avascular necrosis of the capital femoral epiphysis
C1442965|T047|SY|111255008|SNOMEDCT_CORE|Perthes disease|Avascular necrosis of the capital femoral epiphysis
C1442965|T047|SY|111255008|SNOMEDCT_CORE|Perthes disease of hip|Avascular necrosis of the capital femoral epiphysis
C1442978|T047|SY|128545000|SNOMEDCT_CORE|External abdominal hernia|Hernia of abdominal wall
C1442978|T047|PT|128545000|SNOMEDCT_CORE|Hernia of abdominal wall|Hernia of abdominal wall
C1442978|T047|FN|128545000|SNOMEDCT_CORE|Hernia of abdominal wall|Hernia of abdominal wall
C1442981|T047|PT|41309000|SNOMEDCT_CORE|Alcoholic liver damage|Alcoholic liver damage
C1442981|T047|FN|41309000|SNOMEDCT_CORE|Alcoholic liver damage|Alcoholic liver damage
C1442981|T047|IS|41309000|SNOMEDCT_CORE|Alcoholic liver damage, NOS|Alcoholic liver damage
C1442994|T047|SY|237037006|SNOMEDCT_CORE|Acute pelvic inflammatory disease of the female pelvic organs AND/OR tissues|Acute pelvic inflammatory disease of the female pelvic organs AND/OR tissues
C1443005|T047|IS|48194001|SNOMEDCT_CORE|Hypertension in the obstetric context|Hypertension in the obstetric context
C1443027|T037|SY|11196001|SNOMEDCT_CORE|Opiate agonist poisoning|Opiate poisoning
C1443027|T037|SY|11196001|SNOMEDCT_CORE|Opiate poisoning|Opiate poisoning
C1443028|T037|IS|11196001|SNOMEDCT_CORE|Poisoning by opiate or related narcotic, NOS|Poisoning by opiate or related narcotic, NOS
C1443030|T037|SY|11196001|SNOMEDCT_CORE|Opiate and narcotic poisoning|Opiate and narcotic poisoning
C1443290|T047|PT|408749000|SNOMEDCT_CORE|Complex regional pain syndrome, type II, lower limb|Complex regional pain syndrome, type II, lower limb
C1443290|T047|FN|408749000|SNOMEDCT_CORE|Complex regional pain syndrome, type II, lower limb|Complex regional pain syndrome, type II, lower limb
C1443291|T047|PT|408750000|SNOMEDCT_CORE|Complex regional pain syndrome, type II, upper limb|Complex regional pain syndrome, type II, upper limb
C1443291|T047|FN|408750000|SNOMEDCT_CORE|Complex regional pain syndrome, type II, upper limb|Complex regional pain syndrome, type II, upper limb
C1443978|T046|PT|409666003|SNOMEDCT_CORE|Pathological fracture of neck of femur|Pathological fracture of neck of femur
C1443978|T046|FN|409666003|SNOMEDCT_CORE|Pathological fracture of neck of femur|Pathological fracture of neck of femur
C1443979|T046|PT|409667007|SNOMEDCT_CORE|Pathological fracture of femur|Pathological fracture of femur
C1443979|T046|FN|409667007|SNOMEDCT_CORE|Pathological fracture of femur|Pathological fracture of femur
C1443982|T033|PT|409673008|SNOMEDCT_CORE|ALT level raised|ALT level raised
C1443982|T033|OF|409673008|SNOMEDCT_CORE|ALT level raised|ALT level raised
C1444093|T047|SY|409796004|SNOMEDCT_CORE|Infection caused by antimicrobial resistant bacteria|Infection due to resistant bacteria
C1444093|T047|FN|409796004|SNOMEDCT_CORE|Infection caused by antimicrobial resistant bacteria|Infection due to resistant bacteria
C1444093|T047|SY|409796004|SNOMEDCT_CORE|Infection caused by resistant bacteria|Infection due to resistant bacteria
C1444093|T047|OF|409796004|SNOMEDCT_CORE|Infection due to antimicrobial resistant bacteria|Infection due to resistant bacteria
C1444093|T047|SY|409796004|SNOMEDCT_CORE|Infection due to antimicrobial resistant bacteria|Infection due to resistant bacteria
C1444093|T047|PT|409796004|SNOMEDCT_CORE|Infection due to resistant bacteria|Infection due to resistant bacteria
C1444094|T047|SY|409797008|SNOMEDCT_CORE|Infection caused by antimicrobial resistant fungi|Infection due to resistant fungi
C1444094|T047|FN|409797008|SNOMEDCT_CORE|Infection caused by antimicrobial resistant fungi|Infection due to resistant fungi
C1444094|T047|SY|409797008|SNOMEDCT_CORE|Infection caused by resistant fungi|Infection due to resistant fungi
C1444094|T047|OF|409797008|SNOMEDCT_CORE|Infection due to antimicrobial resistant fungi|Infection due to resistant fungi
C1444094|T047|SY|409797008|SNOMEDCT_CORE|Infection due to antimicrobial resistant fungi|Infection due to resistant fungi
C1444094|T047|PT|409797008|SNOMEDCT_CORE|Infection due to resistant fungi|Infection due to resistant fungi
C1444095|T047|SY|409798003|SNOMEDCT_CORE|Infection caused by antimicrobial resistant virus|Infection due to resistant virus
C1444095|T047|FN|409798003|SNOMEDCT_CORE|Infection caused by antimicrobial resistant virus|Infection due to resistant virus
C1444095|T047|SY|409798003|SNOMEDCT_CORE|Infection caused by resistant virus|Infection due to resistant virus
C1444095|T047|OF|409798003|SNOMEDCT_CORE|Infection due to antimicrobial resistant virus|Infection due to resistant virus
C1444095|T047|SY|409798003|SNOMEDCT_CORE|Infection due to antimicrobial resistant virus|Infection due to resistant virus
C1444095|T047|PT|409798003|SNOMEDCT_CORE|Infection due to resistant virus|Infection due to resistant virus
C1444680|T047|OAS|410567004|SNOMEDCT_CORE|Cloudy posterior capsule|Posterior capsule opacification
C1444680|T047|OAS|410567004|SNOMEDCT_CORE|PCF - Posterior capsular fibrosis|Posterior capsule opacification
C1444680|T047|OAS|410567004|SNOMEDCT_CORE|PCO - Posterior capsule opacification|Posterior capsule opacification
C1444680|T047|OAS|410567004|SNOMEDCT_CORE|Posterior capsular fibrosis|Posterior capsule opacification
C1444680|T047|OAS|410567004|SNOMEDCT_CORE|Posterior capsular opacification|Posterior capsule opacification
C1444680|T047|OAS|410567004|SNOMEDCT_CORE|Posterior capsule fibrosis|Posterior capsule opacification
C1444680|T047|OAP|410567004|SNOMEDCT_CORE|Posterior capsule opacification|Posterior capsule opacification
C1444680|T047|OAF|410567004|SNOMEDCT_CORE|Posterior capsule opacification|Posterior capsule opacification
C1446377|T033|PT|413307004|SNOMEDCT_CORE|Mental health problem|Mental health problem
C1446377|T033|FN|413307004|SNOMEDCT_CORE|Mental health problem|Mental health problem
C1449563|T047|PT|53043001|SNOMEDCT_CORE|Primary idiopathic dilated cardiomyopathy|Primary idiopathic dilated cardiomyopathy
C1449563|T047|FN|53043001|SNOMEDCT_CORE|Primary idiopathic dilated cardiomyopathy|Primary idiopathic dilated cardiomyopathy
C1455742|T047|PT|78868004|SNOMEDCT_CORE|Chronic mucoid otitis media|Chronic mucoid otitis media
C1455742|T047|FN|78868004|SNOMEDCT_CORE|Chronic mucoid otitis media|Chronic mucoid otitis media
C1455742|T047|IS|78868004|SNOMEDCT_CORE|Chronic mucoid otitis media, NOS|Chronic mucoid otitis media
C1455742|T047|SY|78868004|SNOMEDCT_CORE|Simple chronic mucoid otitis media|Chronic mucoid otitis media
C1455742|T047|IS|78868004|SNOMEDCT_CORE|Simple chronic mucoid otitis media, NOS|Chronic mucoid otitis media
C1455748|T047|IS|4927003|SNOMEDCT_CORE|Acute cyclitis|Acute cyclitis
C1455749|T047|SY|4927003|SNOMEDCT_CORE|Acute iridocyclitis|Acute iridocyclitis
C1455780|T047|PT|67754003|SNOMEDCT_CORE|Aortic valve sclerosis|Aortic valve sclerosis
C1455780|T047|FN|67754003|SNOMEDCT_CORE|Aortic valve sclerosis|Aortic valve sclerosis
C1455889|T033|PT|441087007|SNOMEDCT_CORE|Atypical squamous cells of undetermined significance on cervical Papanicolaou smear|Atypical squamous cells of undetermined significance on cervical Papanicolaou smear
C1455889|T033|FN|441087007|SNOMEDCT_CORE|Atypical squamous cells of undetermined significance on cervical Papanicolaou smear|Atypical squamous cells of undetermined significance on cervical Papanicolaou smear
C1456132|T047|PT|427794001|SNOMEDCT_CORE|Primary focal hyperhidrosis|Primary focal hyperhidrosis
C1456132|T047|FN|427794001|SNOMEDCT_CORE|Primary focal hyperhidrosis|Primary focal hyperhidrosis
C1456141|T047|OAP|430949005|SNOMEDCT_CORE|Decubitus ulcer of lower back|Pressure ulcer of lower back
C1456141|T047|OAF|430949005|SNOMEDCT_CORE|Decubitus ulcer of lower back|Pressure ulcer of lower back
C1456141|T047|PT|699215008|SNOMEDCT_CORE|Pressure ulcer of lower back|Pressure ulcer of lower back
C1456141|T047|FN|699215008|SNOMEDCT_CORE|Pressure ulcer of lower back|Pressure ulcer of lower back
C1456248|T047|PT|423633003|SNOMEDCT_CORE|Midline cystocele|Midline cystocele
C1456248|T047|FN|423633003|SNOMEDCT_CORE|Midline cystocele|Midline cystocele
C1456332|T048|PT|441527004|SNOMEDCT_CORE|Stimulant abuse|Stimulant abuse
C1456332|T048|FN|441527004|SNOMEDCT_CORE|Stimulant abuse|Stimulant abuse
C1456496|T037|SY|127294003|SNOMEDCT_CORE|Brain damage|Traumatic AND/OR non-traumatic brain injury
C1456496|T037|PT|127294003|SNOMEDCT_CORE|Traumatic AND/OR non-traumatic brain injury|Traumatic AND/OR non-traumatic brain injury
C1456496|T037|FN|127294003|SNOMEDCT_CORE|Traumatic AND/OR non-traumatic brain injury|Traumatic AND/OR non-traumatic brain injury
C1456771|T048|PT|64386003|SNOMEDCT_CORE|Sedative abuse|Sedative abuse
C1456771|T048|FN|64386003|SNOMEDCT_CORE|Sedative abuse|Sedative abuse
C1456771|T048|SY|64386003|SNOMEDCT_CORE|Tranquilizer abuse|Sedative abuse
C1456771|T048|SYGB|64386003|SNOMEDCT_CORE|Tranquilliser abuse|Sedative abuse
C1456771|T048|IS|64386003|SNOMEDCT_CORE|Tranquillizer abuse|Sedative abuse
C1456781|T191|SYGB|400010006|SNOMEDCT_CORE|Benign melanocytic naevus of skin|Benign melanocytic nevus of skin
C1456781|T191|SY|400010006|SNOMEDCT_CORE|Benign melanocytic nevus of skin|Benign melanocytic nevus of skin
C1456784|T048|IS|48500005|SNOMEDCT_CORE|Paranoia|Paranoid disorder
C1456784|T048|SY|191667009|SNOMEDCT_CORE|Paranoia|Paranoid disorder
C1456784|T048|IS|48500005|SNOMEDCT_CORE|Paranoia, NOS|Paranoid disorder
C1456784|T048|IS|48500005|SNOMEDCT_CORE|Paranoid disorder|Paranoid disorder
C1456784|T048|PT|191667009|SNOMEDCT_CORE|Paranoid disorder|Paranoid disorder
C1456784|T048|FN|191667009|SNOMEDCT_CORE|Paranoid disorder|Paranoid disorder
C1456784|T048|IS|48500005|SNOMEDCT_CORE|Paranoid disorder, NOS|Paranoid disorder
C1456784|T048|IS|48500005|SNOMEDCT_CORE|Paranoid psychosis|Paranoid disorder
C1456784|T048|SY|191667009|SNOMEDCT_CORE|Paranoid psychosis|Paranoid disorder
C1456822|T033|OAF|275520000|SNOMEDCT_CORE|Claudication|Claudication
C1456822|T033|OAP|275520000|SNOMEDCT_CORE|Claudication|Claudication
C1456868|T047|PT|371087003|SNOMEDCT_CORE|Diabetic foot ulcer|Diabetic foot ulcer
C1456868|T047|OF|371087003|SNOMEDCT_CORE|Diabetic foot ulcer|Diabetic foot ulcer
C1456868|T047|SY|371087003|SNOMEDCT_CORE|Ulcer of foot due to diabetes mellitus|Diabetic foot ulcer
C1456868|T047|FN|371087003|SNOMEDCT_CORE|Ulcer of foot due to diabetes mellitus|Diabetic foot ulcer
C1456876|T033|SY|39406005|SNOMEDCT_CORE|Legal abortion|Legal termination of pregnancy
C1456876|T033|PT|39406005|SNOMEDCT_CORE|Legal termination of pregnancy|Legal termination of pregnancy
C1456876|T033|SY|39406005|SNOMEDCT_CORE|Legally induced abortion|Legal termination of pregnancy
C1456876|T033|FN|39406005|SNOMEDCT_CORE|Legally induced abortion|Legal termination of pregnancy
C1456876|T033|SY|39406005|SNOMEDCT_CORE|Legally induced abortion - TOP|Legal termination of pregnancy
C1458140|T046|SY|64779008|SNOMEDCT_CORE|Bleeding diathesis|Bleeding tendency
C1458140|T046|SY|64779008|SNOMEDCT_CORE|Bleeding disorder|Bleeding tendency
C1458140|T046|SY|64779008|SNOMEDCT_CORE|Bleeding tendency|Bleeding tendency
C1458155|T191|SY|126926005|SNOMEDCT_CORE|Breast tumor|Neoplasm of breast
C1458155|T191|SYGB|126926005|SNOMEDCT_CORE|Breast tumour|Neoplasm of breast
C1458155|T191|PT|126926005|SNOMEDCT_CORE|Neoplasm of breast|Neoplasm of breast
C1458155|T191|FN|126926005|SNOMEDCT_CORE|Neoplasm of breast|Neoplasm of breast
C1458155|T191|SY|126926005|SNOMEDCT_CORE|Tumor of breast|Neoplasm of breast
C1458155|T191|SYGB|126926005|SNOMEDCT_CORE|Tumour of breast|Neoplasm of breast
C1510412|T046|SYGB|22036004|SNOMEDCT_CORE|Aneurysmal haematoma|Pseudoaneurysm
C1510412|T046|SY|22036004|SNOMEDCT_CORE|Aneurysmal hematoma|Pseudoaneurysm
C1510412|T046|SY|22036004|SNOMEDCT_CORE|False aneurysm|Pseudoaneurysm
C1510412|T046|PT|443089001|SNOMEDCT_CORE|Pseudoaneurysm|Pseudoaneurysm
C1510412|T046|PT|22036004|SNOMEDCT_CORE|Pseudoaneurysm|Pseudoaneurysm
C1510412|T046|FN|22036004|SNOMEDCT_CORE|Pseudoaneurysm|Pseudoaneurysm
C1510412|T046|FN|443089001|SNOMEDCT_CORE|Pseudoaneurysm|Pseudoaneurysm
C1510412|T046|SYGB|22036004|SNOMEDCT_CORE|Pulsatile haematoma|Pseudoaneurysm
C1510412|T046|SY|22036004|SNOMEDCT_CORE|Pulsatile hematoma|Pseudoaneurysm
C1510428|T047|PT|60404007|SNOMEDCT_CORE|Cerebral abscess|Cerebral abscess
C1510428|T047|FN|60404007|SNOMEDCT_CORE|Cerebral abscess|Cerebral abscess
C1510428|T047|SY|60404007|SNOMEDCT_CORE|Parenchymal intracranial abscess|Cerebral abscess
C1510429|T047|SY|45781009|SNOMEDCT_CORE|Compression neuropathy|Peripheral nerve entrapment syndrome
C1510429|T047|SY|45781009|SNOMEDCT_CORE|Entrapment neuropathy|Peripheral nerve entrapment syndrome
C1510429|T047|IS|45781009|SNOMEDCT_CORE|Entrapment neuropathy, NOS|Peripheral nerve entrapment syndrome
C1510429|T047|IS|45781009|SNOMEDCT_CORE|Entrapment syndrome, NOS|Peripheral nerve entrapment syndrome
C1510429|T047|SY|45781009|SNOMEDCT_CORE|Nerve entrapment syndrome|Peripheral nerve entrapment syndrome
C1510429|T047|FN|45781009|SNOMEDCT_CORE|Peripheral nerve entrapment syndrome|Peripheral nerve entrapment syndrome
C1510429|T047|PT|45781009|SNOMEDCT_CORE|Peripheral nerve entrapment syndrome|Peripheral nerve entrapment syndrome
C1510429|T047|SY|45781009|SNOMEDCT_CORE|Trapped nerve|Peripheral nerve entrapment syndrome
C1510431|T047|PT|2477008|SNOMEDCT_CORE|Superficial thrombophlebitis|Superficial thrombophlebitis
C1510431|T047|FN|2477008|SNOMEDCT_CORE|Superficial thrombophlebitis|Superficial thrombophlebitis
C1510431|T047|IS|2477008|SNOMEDCT_CORE|Superficial thrombophlebitis, NOS|Superficial thrombophlebitis
C1510446|T047|PTGB|413439005|SNOMEDCT_CORE|Acute ischaemic heart disease|Acute ischemic heart disease
C1510446|T047|PT|413439005|SNOMEDCT_CORE|Acute ischemic heart disease|Acute ischemic heart disease
C1510446|T047|FN|413439005|SNOMEDCT_CORE|Acute ischemic heart disease|Acute ischemic heart disease
C1510449|T047|IS|398155003|SNOMEDCT_CORE|Chronic iridocyclitis|Chronic iridocyclitis
C1510472|T048|SY|2403008|SNOMEDCT_CORE|Dependence syndrome|Psychoactive substance dependence
C1510472|T048|IS|191816009|SNOMEDCT_CORE|Drug addiction|Psychoactive substance dependence
C1510472|T048|IS|2403008|SNOMEDCT_CORE|Drug dependence|Psychoactive substance dependence
C1510472|T048|PT|191816009|SNOMEDCT_CORE|Drug dependence|Psychoactive substance dependence
C1510472|T048|FN|191816009|SNOMEDCT_CORE|Drug dependence|Psychoactive substance dependence
C1510472|T048|IS|2403008|SNOMEDCT_CORE|Drug dependence, NOS|Psychoactive substance dependence
C1510472|T048|PT|2403008|SNOMEDCT_CORE|Psychoactive substance dependence|Psychoactive substance dependence
C1510472|T048|FN|2403008|SNOMEDCT_CORE|Psychoactive substance dependence|Psychoactive substance dependence
C1510472|T048|IS|2403008|SNOMEDCT_CORE|Psychoactive substance dependence, NOS|Psychoactive substance dependence
C1510479|T047|IS|3548001|SNOMEDCT_CORE|Neuralgic amyotrophy|Neuralgic amyotrophy
C1510497|T033|SY|193570009|SNOMEDCT_CORE|Lens opacity|Lenticular opacity
C1510497|T033|SY|193570009|SNOMEDCT_CORE|Lenticular opacity|Lenticular opacity
C1510654|T047|SYGB|271737000|SNOMEDCT_CORE|Absolute anaemia|Absolute anemia
C1510654|T047|SY|271737000|SNOMEDCT_CORE|Absolute anemia|Absolute anemia
C1519353|T033|PT|271757001|SNOMEDCT_CORE|Papular eruption|Papular eruption
C1519353|T033|FN|271757001|SNOMEDCT_CORE|Papular eruption|Papular eruption
C1519353|T033|IS|271757001|SNOMEDCT_CORE|Papular rash|Papular eruption
C1521728|T047|IS|266257000|SNOMEDCT_CORE|Intermittent cerebral ischaemia|Intermittent cerebral ischemia
C1521728|T047|IS|266257000|SNOMEDCT_CORE|Intermittent cerebral ischemia|Intermittent cerebral ischemia
C1522512|T048|IS|17226007|SNOMEDCT_CORE|Transient situational disturbance|Transient situational disturbance
C1522512|T048|SY|192041001|SNOMEDCT_CORE|Transient situational disturbance|Transient situational disturbance
C1522512|T048|IS|17226007|SNOMEDCT_CORE|Transient situational disturbance, NOS|Transient situational disturbance
C1522520|T048|SY|17226007|SNOMEDCT_CORE|Adaptation reaction|Adaptation reaction
C1522520|T048|IS|17226007|SNOMEDCT_CORE|Adaptation reaction, NOS|Adaptation reaction
C1522522|T047|SY|111496009|SNOMEDCT_CORE|Hydrosyringomyelia|Hydrosyringomyelia
C1527168|T047|SY|38804009|SNOMEDCT_CORE|Bonnevie-Ullrich syndrome|Bonnevie-Ullrich syndrome
C1527226|T047|SY|62382002|SNOMEDCT_CORE|Calcinosis cutis, Raynaud's, sclerodactyly AND telangiectasia|CRST syndrome
C1527226|T047|IS|62382002|SNOMEDCT_CORE|Calcinosis cutis, Raynaud's, sclerodactyly and telangiectasia|CRST syndrome
C1527226|T047|SY|62382002|SNOMEDCT_CORE|Calcinosis, Raynaud phenomenon, sclerodactyly, and telangiectasia syndrome|CRST syndrome
C1527226|T047|SY|62382002|SNOMEDCT_CORE|Calcinosis, Raynaud's phenomenon, sclerodactyly, and telangiectasia syndrome|CRST syndrome
C1527226|T047|FN|62382002|SNOMEDCT_CORE|Calcinosis, Raynaud's phenomenon, sclerodactyly, and telangiectasia syndrome|CRST syndrome
C1527226|T047|OF|62382002|SNOMEDCT_CORE|Calcinosis, Raynaud's phenomenon, sclerodactyly, and telangiectasia syndrome|CRST syndrome
C1527226|T047|SY|62382002|SNOMEDCT_CORE|Calcinosis, Raynaud's phenomenon, sclerodactyly, telangiectasia syndrome|CRST syndrome
C1527226|T047|IS|62382002|SNOMEDCT_CORE|Calcinosis, Raynaud's phenomenon, sclerodactyly, telangiectasia syndrome|CRST syndrome
C1527226|T047|SY|62382002|SNOMEDCT_CORE|CRST - Calcinosis, Raynaud's phenomenon, sclerodactyly, telangiectasia syndrome|CRST syndrome
C1527226|T047|PT|62382002|SNOMEDCT_CORE|CRST syndrome|CRST syndrome
C1527226|T047|OF|62382002|SNOMEDCT_CORE|CRST syndrome|CRST syndrome
C1527303|T047|SY|13645005|SNOMEDCT_CORE|CAO - Chronic airflow obstruction|CAO - Chronic airflow obstruction
C1527303|T047|SY|13645005|SNOMEDCT_CORE|Chronic airflow obstruction|CAO - Chronic airflow obstruction
C1527310|T047|SY|39021009|SNOMEDCT_CORE|Ametropia|Ametropia
C1527311|T046|SY|2032001|SNOMEDCT_CORE|Intracranial swelling|Intracranial swelling
C1527320|T047|SY|13445001|SNOMEDCT_CORE|Aural vertigo|Aural vertigo
C1527336|T047|SY|83901003|SNOMEDCT_CORE|Sjögren syndrome|Sjögren's syndrome
C1527336|T047|SY|83901003|SNOMEDCT_CORE|Sjögren's disease|Sjögren's syndrome
C1527336|T047|IS|83901003|SNOMEDCT_CORE|Sjogren's disease|Sjögren's syndrome
C1527336|T047|SY|83901003|SNOMEDCT_CORE|Sjogren's syndrome|Sjögren's syndrome
C1527336|T047|PT|83901003|SNOMEDCT_CORE|Sjögren's syndrome|Sjögren's syndrome
C1527336|T047|FN|83901003|SNOMEDCT_CORE|Sjögren's syndrome|Sjögren's syndrome
C1527336|T047|SY|83901003|SNOMEDCT_CORE|Sjogrens syndrome|Sjögren's syndrome
C1527340|T033|PT|38160000|SNOMEDCT_CORE|Abnormal voice|Abnormal voice
C1527340|T033|FN|38160000|SNOMEDCT_CORE|Abnormal voice|Abnormal voice
C1527340|T033|IS|47004009|SNOMEDCT_CORE|Voice disturbance|Abnormal voice
C1527340|T033|IS|47004009|SNOMEDCT_CORE|Voice disturbance, NOS|Abnormal voice
C1527344|T048|IS|47004009|SNOMEDCT_CORE|Dysphonia|Dysphonia
C1527344|T048|IS|47004009|SNOMEDCT_CORE|Dysphonia, NOS|Dysphonia
C1527344|T048|IS|47004009|SNOMEDCT_CORE|Phonation disorder|Dysphonia
C1527347|T033|OAP|47004009|SNOMEDCT_CORE|Difficulty speaking|Difficulty speaking
C1527347|T033|OAF|47004009|SNOMEDCT_CORE|Difficulty speaking|Difficulty speaking
C1527347|T033|IS|47004009|SNOMEDCT_CORE|Disorder of speech|Difficulty speaking
C1527347|T033|IS|47004009|SNOMEDCT_CORE|Speech disorder|Difficulty speaking
C1527351|T047|PT|72274001|SNOMEDCT_CORE|Nerve root disorder|Nerve root disorder
C1527351|T047|FN|72274001|SNOMEDCT_CORE|Nerve root disorder|Nerve root disorder
C1527351|T047|IS|72274001|SNOMEDCT_CORE|Nerve root disorder, NOS|Nerve root disorder
C1527375|T047|SY|27431007|SNOMEDCT_CORE|Cystic disease of breast|Cystic disease of breast
C1527384|T184|SY|26079004|SNOMEDCT_CORE|Involuntary quiver|Quivering
C1527384|T184|SY|26079004|SNOMEDCT_CORE|Quivering|Quivering
C1527395|T047|SY|35065006|SNOMEDCT_CORE|Acute pseudo-obstruction of colon|Acute pseudo-obstruction of colon
C1527395|T047|SY|35065006|SNOMEDCT_CORE|Ogilvie's syndrome|Acute pseudo-obstruction of colon
C1527405|T033|PT|127062003|SNOMEDCT_CORE|Erythrocytosis|Erythrocytosis
C1527405|T033|IS|44865000|SNOMEDCT_CORE|Erythrocytosis|Erythrocytosis
C1527405|T033|FN|127062003|SNOMEDCT_CORE|Erythrocytosis|Erythrocytosis
C1527406|T047|SY|65323003|SNOMEDCT_CORE|Rhizomelic pseudopolyarthritis|Rhizomelic pseudopolyarthritis
C1527410|T047|SY|16726004|SNOMEDCT_CORE|Renal rickets|Renal rickets
C1532235|T047|PTGB|414027002|SNOMEDCT_CORE|Disorder of haematopoietic structure|Disorder of hematopoietic structure
C1532235|T047|PT|414027002|SNOMEDCT_CORE|Disorder of hematopoietic structure|Disorder of hematopoietic structure
C1532235|T047|FN|414027002|SNOMEDCT_CORE|Disorder of hematopoietic structure|Disorder of hematopoietic structure
C1532240|T047|PT|414033006|SNOMEDCT_CORE|Disorder of rotator cuff|Disorder of rotator cuff
C1532240|T047|FN|414033006|SNOMEDCT_CORE|Disorder of rotator cuff|Disorder of rotator cuff
C1532285|T020|OAF|414477008|SNOMEDCT_CORE|Incisional hernia of anterior abdominal wall without obstruction AND without gangrene|Ventral incisional hernia of anterior abdominal wall without obstruction AND without gangrene
C1532285|T020|OAS|414477008|SNOMEDCT_CORE|Incisional hernia of anterior abdominal wall without obstruction AND without gangrene|Ventral incisional hernia of anterior abdominal wall without obstruction AND without gangrene
C1532285|T020|OAP|414477008|SNOMEDCT_CORE|Ventral incisional hernia of anterior abdominal wall without obstruction AND without gangrene|Ventral incisional hernia of anterior abdominal wall without obstruction AND without gangrene
C1532320|T033|PT|414205003|SNOMEDCT_CORE|Family history of prostate cancer|Family history of prostate cancer
C1532320|T033|OF|414205003|SNOMEDCT_CORE|Family history of prostate cancer|Family history of prostate cancer
C1532320|T033|FN|414205003|SNOMEDCT_CORE|Family history of prostate cancer|Family history of prostate cancer
C1532381|T033|PT|414861001|SNOMEDCT_CORE|No evidence of recurrence of cancer|No evidence of recurrence of cancer
C1532381|T033|OF|414861001|SNOMEDCT_CORE|No evidence of recurrence of cancer|No evidence of recurrence of cancer
C1532381|T033|FN|414861001|SNOMEDCT_CORE|No evidence of recurrence of cancer|No evidence of recurrence of cancer
C1532396|T033|SY|415086001|SNOMEDCT_CORE|H/O: malignant neoplasm of bladder|History of malignant neoplasm of bladder
C1532396|T033|PT|415086001|SNOMEDCT_CORE|History of malignant neoplasm of bladder|History of malignant neoplasm of bladder
C1532396|T033|OF|415086001|SNOMEDCT_CORE|Personal history of primary malignant neoplasm of urinary bladder|History of malignant neoplasm of bladder
C1532396|T033|SY|415086001|SNOMEDCT_CORE|Personal history of primary malignant neoplasm of urinary bladder|History of malignant neoplasm of bladder
C1532396|T033|FN|415086001|SNOMEDCT_CORE|Personal history of primary malignant neoplasm of urinary bladder|History of malignant neoplasm of bladder
C1533012|T190|OAF|414399004|SNOMEDCT_CORE|Hernia of anterior abdominal wall without obstruction AND without gangrene|Hernia of anterior abdominal wall without obstruction AND without gangrene
C1533012|T190|OAP|414399004|SNOMEDCT_CORE|Hernia of anterior abdominal wall without obstruction AND without gangrene|Hernia of anterior abdominal wall without obstruction AND without gangrene
C1533012|T190|IS|414477008|SNOMEDCT_CORE|Ventral hernia without obstruction AND without gangrene|Hernia of anterior abdominal wall without obstruction AND without gangrene
C1533012|T190|OAS|414399004|SNOMEDCT_CORE|Ventral hernia without obstruction AND without gangrene|Hernia of anterior abdominal wall without obstruction AND without gangrene
C1533849|T047|SY|86276007|SNOMEDCT_CORE|Bleeding of subgingival space|Bleeding of subgingival space
C1533849|T047|SY|86276007|SNOMEDCT_CORE|Crevicular bleeding of gum|Bleeding of subgingival space
C1533849|T047|SY|86276007|SNOMEDCT_CORE|Gingival crevice bleeding|Bleeding of subgingival space
C1533849|T047|SY|86276007|SNOMEDCT_CORE|Gingival crevicular bleeding|Bleeding of subgingival space
C1535939|T047|SY|415125002|SNOMEDCT_CORE|PCP - Pneumocystis pneumonia|Pneumocystosis pneumonia
C1535939|T047|OF|415125002|SNOMEDCT_CORE|Pneumocystosis jiroveci pneumonia|Pneumocystosis pneumonia
C1535939|T047|IS|415125002|SNOMEDCT_CORE|Pneumocystosis jiroveci pneumonia|Pneumocystosis pneumonia
C1535939|T047|SY|415125002|SNOMEDCT_CORE|Pneumocystosis jirovecii pneumonia|Pneumocystosis pneumonia
C1535939|T047|FN|415125002|SNOMEDCT_CORE|Pneumocystosis jirovecii pneumonia|Pneumocystosis pneumonia
C1535939|T047|PT|415125002|SNOMEDCT_CORE|Pneumocystosis pneumonia|Pneumocystosis pneumonia
C1535939|T047|SY|415125002|SNOMEDCT_CORE|Pulmonary pneumocystosis|Pneumocystosis pneumonia
C1536114|T047|PT|426566004|SNOMEDCT_CORE|Central pain syndrome|Central pain syndrome
C1536114|T047|FN|426566004|SNOMEDCT_CORE|Central pain syndrome|Central pain syndrome
C1536148|T191|PT|237116001|SNOMEDCT_CORE|Chocolate cyst of ovary|Chocolate cyst of ovary
C1536148|T191|FN|237116001|SNOMEDCT_CORE|Chocolate cyst of ovary|Chocolate cyst of ovary
C1536148|T191|SY|237116001|SNOMEDCT_CORE|Endometrioma|Chocolate cyst of ovary
C1536148|T191|SY|237116001|SNOMEDCT_CORE|Endometriotic cyst of ovary|Chocolate cyst of ovary
C1536651|T047|OAS|238793001|SNOMEDCT_CORE|Arterial leg ulcer|Arterial leg ulcer
C1536885|T191|IS|93797001|SNOMEDCT_CORE|Malignant neoplasm of female genital organ|Primary malignant neoplasm of female genital organ
C1536885|T191|IS|93797001|SNOMEDCT_CORE|Malignant neoplasm of female genital organ, NOS|Primary malignant neoplasm of female genital organ
C1536885|T191|PT|93797001|SNOMEDCT_CORE|Primary malignant neoplasm of female genital organ|Primary malignant neoplasm of female genital organ
C1536885|T191|FN|93797001|SNOMEDCT_CORE|Primary malignant neoplasm of female genital organ|Primary malignant neoplasm of female genital organ
C1536978|T047|SY|12867002|SNOMEDCT_CORE|Abnormal fetal heart rate AND/OR rhythm affecting management of mother|Abnormal fetal heart rate AND/OR rhythm affecting management of mother
C1536978|T047|IS|12867002|SNOMEDCT_CORE|Abnormal fetal heart rate or rhythm affecting management of mother|Abnormal fetal heart rate AND/OR rhythm affecting management of mother
C1537189|T047|IS|13645005|SNOMEDCT_CORE|Chronic obstructive lung disease, NEC|Chronic obstructive lung disease, NEC
C1540802|T033|IS|44247006|SNOMEDCT_CORE|Fetus with birthweight of 1000-2499 grams and gestation of 28-37 weeks|Fetus with birthweight of 1000-2499 grams AND/OR gestation of 28-37 weeks
C1540802|T033|IS|44247006|SNOMEDCT_CORE|Fetus with birthweight of 1000-2499 grams AND/OR gestation of 28-37 weeks|Fetus with birthweight of 1000-2499 grams AND/OR gestation of 28-37 weeks
C1540912|T047|PT|128835008|SNOMEDCT_CORE|Hypereosinophilic syndrome|Hypereosinophilic syndrome
C1540912|T047|OF|128835008|SNOMEDCT_CORE|Hypereosinophilic syndrome|Hypereosinophilic syndrome
C1540912|T047|SY|128835008|SNOMEDCT_CORE|Hypereosinophilic syndrome/chronic eosinophilic leukemia|Hypereosinophilic syndrome
C1540912|T047|FN|128835008|SNOMEDCT_CORE|Hypereosinophilic syndrome/chronic eosinophilic leukemia|Hypereosinophilic syndrome
C1542178|T037|PT|414292006|SNOMEDCT_CORE|Fracture of lower leg|Fracture of lower leg
C1542178|T037|FN|414292006|SNOMEDCT_CORE|Fracture of lower leg|Fracture of lower leg
C1561613|T047|FN|441935006|SNOMEDCT_CORE|Acquired absence of all teeth|Acquired absence of all teeth
C1561613|T047|PT|441935006|SNOMEDCT_CORE|Acquired absence of all teeth|Acquired absence of all teeth
C1561613|T047|SY|441935006|SNOMEDCT_CORE|Complete edentulism|Acquired absence of all teeth
C1561643|T047|OAS|236425005|SNOMEDCT_CORE|Chronic kidney disease|Chronic kidney disease
C1561643|T047|PT|709044004|SNOMEDCT_CORE|Chronic kidney disease|Chronic kidney disease
C1561643|T047|FN|709044004|SNOMEDCT_CORE|Chronic kidney disease|Chronic kidney disease
C1561643|T047|OAS|236425005|SNOMEDCT_CORE|Chronic renal disease|Chronic kidney disease
C1561643|T047|SY|709044004|SNOMEDCT_CORE|Chronic renal disease|Chronic kidney disease
C1561643|T047|OAS|236425005|SNOMEDCT_CORE|CKD - chronic kidney disease|Chronic kidney disease
C1561643|T047|SY|709044004|SNOMEDCT_CORE|CKD - chronic kidney disease|Chronic kidney disease
C1561668|T033|PT|428942009|SNOMEDCT_CORE|History of fall|History of fall
C1561668|T033|FN|428942009|SNOMEDCT_CORE|History of fall|History of fall
C1561842|T048|SY|3972004|SNOMEDCT_CORE|Idiopathic insomnia|Idiopathic insomnia
C1561850|T048|PT|24121004|SNOMEDCT_CORE|Insomnia disorder related to another mental disorder|Insomnia disorder related to another mental disorder
C1561850|T048|FN|24121004|SNOMEDCT_CORE|Insomnia disorder related to another mental disorder|Insomnia disorder related to another mental disorder
C1561850|T048|SY|24121004|SNOMEDCT_CORE|Insomnia due to mental disorder|Insomnia disorder related to another mental disorder
C1561855|T047|PT|442292004|SNOMEDCT_CORE|Idiopathic hypersomnia without long sleep time|Idiopathic hypersomnia without long sleep time
C1561855|T047|FN|442292004|SNOMEDCT_CORE|Idiopathic hypersomnia without long sleep time|Idiopathic hypersomnia without long sleep time
C1562299|T047|PT|415992005|SNOMEDCT_CORE|Disorder of right cardiac ventricle|Disorder of right cardiac ventricle
C1562299|T047|FN|415992005|SNOMEDCT_CORE|Disorder of right cardiac ventricle|Disorder of right cardiac ventricle
C1562303|T033|SY|416030007|SNOMEDCT_CORE|Cervicovaginal cytology: LGSIL|Cervicovaginal cytology: Low grade squamous intraepithelial lesion
C1562303|T033|PT|416030007|SNOMEDCT_CORE|Cervicovaginal cytology: Low grade squamous intraepithelial lesion|Cervicovaginal cytology: Low grade squamous intraepithelial lesion
C1562303|T033|FN|416030007|SNOMEDCT_CORE|Cervicovaginal cytology: Low grade squamous intraepithelial lesion|Cervicovaginal cytology: Low grade squamous intraepithelial lesion
C1562303|T033|SY|416030007|SNOMEDCT_CORE|Cervicovaginal cytology: LSIL|Cervicovaginal cytology: Low grade squamous intraepithelial lesion
C1562305|T033|PT|416032004|SNOMEDCT_CORE|Cervicovaginal cytology normal or benign|Cervicovaginal cytology normal or benign
C1562305|T033|FN|416032004|SNOMEDCT_CORE|Cervicovaginal cytology normal or benign|Cervicovaginal cytology normal or benign
C1562306|T033|SY|416033009|SNOMEDCT_CORE|Cervicovaginal cytology: HGSIL or carcinoma|Cervicovaginal cytology: High grade squamous intraepithelial lesion or carcinoma
C1562306|T033|PT|416033009|SNOMEDCT_CORE|Cervicovaginal cytology: High grade squamous intraepithelial lesion or carcinoma|Cervicovaginal cytology: High grade squamous intraepithelial lesion or carcinoma
C1562306|T033|FN|416033009|SNOMEDCT_CORE|Cervicovaginal cytology: High grade squamous intraepithelial lesion or carcinoma|Cervicovaginal cytology: High grade squamous intraepithelial lesion or carcinoma
C1562306|T033|SY|416033009|SNOMEDCT_CORE|Cervicovaginal cytology: HSIL or carcinoma|Cervicovaginal cytology: High grade squamous intraepithelial lesion or carcinoma
C1562543|T047|PT|416770009|SNOMEDCT_CORE|Ocular histoplasmosis syndrome|Ocular histoplasmosis syndrome
C1562543|T047|FN|416770009|SNOMEDCT_CORE|Ocular histoplasmosis syndrome|Ocular histoplasmosis syndrome
C1562543|T047|SY|416770009|SNOMEDCT_CORE|OHS-ocular histoplasmosis syndrome|Ocular histoplasmosis syndrome
C1562890|T033|PT|416413003|SNOMEDCT_CORE|Advanced maternal age gravida|Advanced maternal age gravida
C1562890|T033|FN|416413003|SNOMEDCT_CORE|Advanced maternal age gravida|Advanced maternal age gravida
C1562890|T033|SY|416413003|SNOMEDCT_CORE|Advanced maternal age patient|Advanced maternal age gravida
C1562890|T033|SY|416413003|SNOMEDCT_CORE|AMA - advanced maternal age|Advanced maternal age gravida
C1563033|T033|SY|416519002|SNOMEDCT_CORE|Family history of kidney stone|Family history of renal stone
C1563033|T033|SY|416519002|SNOMEDCT_CORE|Family history of nephrolithiasis|Family history of renal stone
C1563033|T033|PT|416519002|SNOMEDCT_CORE|Family history of renal stone|Family history of renal stone
C1563033|T033|OF|416519002|SNOMEDCT_CORE|Family history of renal stone|Family history of renal stone
C1563033|T033|FN|416519002|SNOMEDCT_CORE|Family history of renal stone|Family history of renal stone
C1563292|T033|PT|160313009|SNOMEDCT_CORE|Family history of osteoporosis|Family history of osteoporosis
C1563292|T033|FN|160313009|SNOMEDCT_CORE|Family history of osteoporosis|Family history of osteoporosis
C1563292|T033|SY|160313009|SNOMEDCT_CORE|Family history: Osteoporosis|Family history of osteoporosis
C1563292|T033|OF|160313009|SNOMEDCT_CORE|Family history: Osteoporosis|Family history of osteoporosis
C1563292|T033|SY|160313009|SNOMEDCT_CORE|FH: Osteoporosis|Family history of osteoporosis
C1565489|T047|SY|236423003|SNOMEDCT_CORE|Impaired renal function|Renal impairment
C1565489|T047|SY|236423003|SNOMEDCT_CORE|Renal dysfunction|Renal impairment
C1565489|T047|PT|236423003|SNOMEDCT_CORE|Renal impairment|Renal impairment
C1565489|T047|FN|236423003|SNOMEDCT_CORE|Renal impairment|Renal impairment
C1565887|T184|PT|276549000|SNOMEDCT_CORE|Newborn physiological jaundice|Newborn physiological jaundice
C1565887|T184|OF|276549000|SNOMEDCT_CORE|Newborn physiological jaundice|Newborn physiological jaundice
C1565887|T184|FN|276549000|SNOMEDCT_CORE|Newborn physiological jaundice|Newborn physiological jaundice
C1565887|T184|SY|276549000|SNOMEDCT_CORE|Physiologic jaundice in newborn|Newborn physiological jaundice
C1578545|T033|SY|2314005|SNOMEDCT_CORE|Unprotected coitus|Unprotected sexual intercourse
C1578545|T033|SY|2314005|SNOMEDCT_CORE|Unprotected intercourse|Unprotected sexual intercourse
C1578545|T033|PT|2314005|SNOMEDCT_CORE|Unprotected sexual intercourse|Unprotected sexual intercourse
C1578545|T033|FN|2314005|SNOMEDCT_CORE|Unprotected sexual intercourse|Unprotected sexual intercourse
C1578594|T047|SYGB|1776003|SNOMEDCT_CORE|Renotubular acidaemia|Renotubular acidemia
C1578594|T047|SY|1776003|SNOMEDCT_CORE|Renotubular acidemia|Renotubular acidemia
C1579029|T047|SYGB|90688005|SNOMEDCT_CORE|Chronic uraemia|Chronic uremia
C1579029|T047|SY|90688005|SNOMEDCT_CORE|Chronic uremia|Chronic uremia
C1579688|T033|SY|270472006|SNOMEDCT_CORE|Anxious mother|Anxious mother
C1579830|T033|PT|417237009|SNOMEDCT_CORE|Blister|Blister
C1579830|T033|SY|417237009|SNOMEDCT_CORE|Blister of skin AND/OR mucosa|Blister
C1579830|T033|FN|417237009|SNOMEDCT_CORE|Blister of skin AND/OR mucosa|Blister
C1579830|T033|OF|417237009|SNOMEDCT_CORE|Blister of skin AND/OR mucosa|Blister
C1609538|T047|PT|11999007|SNOMEDCT_CORE|Inactive tuberculosis|Inactive tuberculosis
C1609538|T047|FN|11999007|SNOMEDCT_CORE|Inactive tuberculosis|Inactive tuberculosis
C1609538|T047|SY|11999007|SNOMEDCT_CORE|LTBI - Latent tuberculosis infection|Inactive tuberculosis
C1609538|T047|SY|11999007|SNOMEDCT_CORE|Tuberculosis infection latent|Inactive tuberculosis
C1610605|T047|PT|444547006|SNOMEDCT_CORE|Cutaneous graft-versus-host disease|Cutaneous graft-versus-host disease
C1610605|T047|SY|444547006|SNOMEDCT_CORE|Graft versus host disease of skin|Cutaneous graft-versus-host disease
C1610605|T047|FN|444547006|SNOMEDCT_CORE|Graft versus host disease of skin|Cutaneous graft-versus-host disease
C1611184|T046|PT|445512009|SNOMEDCT_CORE|Calcification of coronary artery|Calcification of coronary artery
C1611184|T046|FN|445512009|SNOMEDCT_CORE|Calcification of coronary artery|Calcification of coronary artery
C1621353|T047|IS|312956001|SNOMEDCT_CORE|Serous macular detachment|Serous macular detachment
C1621825|T047|SY|25924004|SNOMEDCT_CORE|Biliary calculus with cholecystitis|Biliary calculus with cholecystitis
C1621825|T047|IS|25924004|SNOMEDCT_CORE|Biliary calculus with cholecystitis, NOS|Biliary calculus with cholecystitis
C1621860|T033|IS|1855002|SNOMEDCT_CORE|Mental dullness|Mental dullness
C1621958|T191|SY|63634009|SNOMEDCT_CORE|GBM - Glioblastoma multiforme|Glioblastoma multiforme
C1621958|T191|SY|63634009|SNOMEDCT_CORE|Glioblastoma multiforme|Glioblastoma multiforme
C1621958|T191|OF|393563007|SNOMEDCT_CORE|Glioblastoma multiforme|Glioblastoma multiforme
C1621958|T191|PT|393563007|SNOMEDCT_CORE|Glioblastoma multiforme|Glioblastoma multiforme
C1621958|T191|FN|393563007|SNOMEDCT_CORE|Glioblastoma multiforme|Glioblastoma multiforme
C1621958|T191|SY|63634009|SNOMEDCT_CORE|GLM - Glioblastoma multiforme|Glioblastoma multiforme
C1621958|T191|SY|63634009|SNOMEDCT_CORE|Spongioblastoma multiforme|Glioblastoma multiforme
C1622502|T047|SY|419728003|SNOMEDCT_CORE|Laennec's cirrhosis|Portal cirrhosis
C1622502|T047|SY|419728003|SNOMEDCT_CORE|PC - Portal cirrhosis|Portal cirrhosis
C1622502|T047|PT|419728003|SNOMEDCT_CORE|Portal cirrhosis|Portal cirrhosis
C1622502|T047|FN|419728003|SNOMEDCT_CORE|Portal cirrhosis|Portal cirrhosis
C1641808|T047|PT|195474004|SNOMEDCT_CORE|Esophageal varices associated with another disorder|Esophageal varices associated with another disorder
C1641808|T047|FN|195474004|SNOMEDCT_CORE|Esophageal varices associated with another disorder|Esophageal varices associated with another disorder
C1641808|T047|PTGB|195474004|SNOMEDCT_CORE|Oesophageal varices associated with another disorder|Esophageal varices associated with another disorder
C1689817|T047|PT|195029002|SNOMEDCT_CORE|Cardiomyopathy associated with another disorder|Cardiomyopathy associated with another disorder
C1689817|T047|FN|195029002|SNOMEDCT_CORE|Cardiomyopathy associated with another disorder|Cardiomyopathy associated with another disorder
C1689817|T047|SY|195029002|SNOMEDCT_CORE|Cardiomyopathy, secondary|Cardiomyopathy associated with another disorder
C1689817|T047|SY|195029002|SNOMEDCT_CORE|Secondary cardiomyopathy|Cardiomyopathy associated with another disorder
C1691210|T033|OF|95922009|SNOMEDCT_CORE|Child sex abuse|Child sex abuse
C1691210|T033|PT|95922009|SNOMEDCT_CORE|Child sex abuse|Child sex abuse
C1691210|T033|FN|95922009|SNOMEDCT_CORE|Child sex abuse|Child sex abuse
C1691210|T033|SY|95922009|SNOMEDCT_CORE|Child sexual abuse|Child sex abuse
C1691210|T033|SY|95922009|SNOMEDCT_CORE|Sexual abuse of child|Child sex abuse
C1691215|T019|PT|204888000|SNOMEDCT_CORE|Hypospadias, penile|Hypospadias, penile
C1691215|T019|FN|204888000|SNOMEDCT_CORE|Hypospadias, penile|Hypospadias, penile
C1691215|T019|SY|204888000|SNOMEDCT_CORE|Urethral meatus underneath penis|Hypospadias, penile
C1691228|T047|OAP|236439005|SNOMEDCT_CORE|Cystic disease of kidney|Cystic disease of kidney
C1691228|T047|OAF|236439005|SNOMEDCT_CORE|Cystic disease of kidney|Cystic disease of kidney
C1691228|T047|OAS|236439005|SNOMEDCT_CORE|Cystic kidney disease|Cystic kidney disease
C1691779|T047|SY|85571008|SNOMEDCT_CORE|Cochlear hearing loss|Sensory hearing loss
C1691779|T047|SY|85571008|SNOMEDCT_CORE|Inner ear hearing loss|Sensory hearing loss
C1691779|T047|PT|85571008|SNOMEDCT_CORE|Sensory hearing loss|Sensory hearing loss
C1691779|T047|OF|85571008|SNOMEDCT_CORE|Sensory hearing loss|Sensory hearing loss
C1691779|T047|FN|85571008|SNOMEDCT_CORE|Sensory hearing loss|Sensory hearing loss
C1692340|T047|IS|58170007|SNOMEDCT_CORE|Viral meningitis, NEC|Viral meningitis, NEC
C1692871|T047|SY|417373000|SNOMEDCT_CORE|Inflammatory polyarthritis|Inflammatory polyarthritis
C1692872|T047|PT|416956002|SNOMEDCT_CORE|Undifferentiated inflammatory polyarthritis|Undifferentiated inflammatory polyarthritis
C1692872|T047|FN|416956002|SNOMEDCT_CORE|Undifferentiated inflammatory polyarthritis|Undifferentiated inflammatory polyarthritis
C1692886|T047|SY|48245008|SNOMEDCT_CORE|Arthritis due to bacterial infection|Bacterial arthritis
C1692886|T047|PT|48245008|SNOMEDCT_CORE|Bacterial arthritis|Bacterial arthritis
C1692886|T047|FN|48245008|SNOMEDCT_CORE|Bacterial arthritis|Bacterial arthritis
C1692886|T047|IS|48245008|SNOMEDCT_CORE|Bacterial arthritis, NOS|Bacterial arthritis
C1692886|T047|IS|48245008|SNOMEDCT_CORE|Pyogenic arthritis|Bacterial arthritis
C1692886|T047|IS|48245008|SNOMEDCT_CORE|Pyogenic bacterial arthritis|Bacterial arthritis
C1692886|T047|SY|48245008|SNOMEDCT_CORE|Septic arthritis|Bacterial arthritis
C1692886|T047|IS|48245008|SNOMEDCT_CORE|Septic arthritis, NOS|Bacterial arthritis
C1704231|T191|SY|230156002|SNOMEDCT_CORE|Neoplastic meningitis|Neoplastic meningitis
C1704272|T047|PT|266569009|SNOMEDCT_CORE|Benign prostatic hyperplasia|Benign prostatic hyperplasia
C1704272|T047|FN|266569009|SNOMEDCT_CORE|Benign prostatic hyperplasia|Benign prostatic hyperplasia
C1704272|T047|SY|266569009|SNOMEDCT_CORE|BPH - benign prostatic hyperplasia|Benign prostatic hyperplasia
C1704272|T047|SY|266569009|SNOMEDCT_CORE|Nodular hyperplasia of prostate gland|Benign prostatic hyperplasia
C1704273|T191|SY|11314008|SNOMEDCT_CORE|Endometrial polyp|Endometrial polyp
C1704330|T047|SY|234947003|SNOMEDCT_CORE|Dental disease|Disorder of teeth AND/OR supporting structures
C1704330|T047|SY|234947003|SNOMEDCT_CORE|Dental disorder|Disorder of teeth AND/OR supporting structures
C1704330|T047|OF|105995000|SNOMEDCT_CORE|Disease of teeth AND/OR supporting structures|Disorder of teeth AND/OR supporting structures
C1704330|T047|IS|105995000|SNOMEDCT_CORE|Disease of teeth AND/OR supporting structures|Disorder of teeth AND/OR supporting structures
C1704330|T047|FN|105995000|SNOMEDCT_CORE|Disorder of teeth AND/OR supporting structures|Disorder of teeth AND/OR supporting structures
C1704330|T047|PT|105995000|SNOMEDCT_CORE|Disorder of teeth AND/OR supporting structures|Disorder of teeth AND/OR supporting structures
C1704356|T191|PT|423699002|SNOMEDCT_CORE|Enchondroma|Enchondroma
C1704356|T191|FN|423699002|SNOMEDCT_CORE|Enchondroma|Enchondroma
C1704356|T191|SY|423699002|SNOMEDCT_CORE|True chondroma|Enchondroma
C1704417|T047|SYGB|238040008|SNOMEDCT_CORE|Familial hyperlipoproteinaemia type IIb|Familial hyperlipoproteinemia type IIb
C1704417|T047|SY|238040008|SNOMEDCT_CORE|Familial hyperlipoproteinemia type IIb|Familial hyperlipoproteinemia type IIb
C1704417|T047|SYGB|238040008|SNOMEDCT_CORE|FCHL - Familial combined hyperlipidaemia|Familial hyperlipoproteinemia type IIb
C1704417|T047|SY|238040008|SNOMEDCT_CORE|FCHL - Familial combined hyperlipidemia|Familial hyperlipoproteinemia type IIb
C1704417|T047|SYGB|238040008|SNOMEDCT_CORE|Fredrickson type IIb hyperlipoproteinaemia|Familial hyperlipoproteinemia type IIb
C1704417|T047|SY|238040008|SNOMEDCT_CORE|Fredrickson type IIb hyperlipoproteinemia|Familial hyperlipoproteinemia type IIb
C1704417|T047|SYGB|238040008|SNOMEDCT_CORE|Hyperapobetalipoproteinaemia|Familial hyperlipoproteinemia type IIb
C1704417|T047|SY|238040008|SNOMEDCT_CORE|Hyperapobetalipoproteinemia|Familial hyperlipoproteinemia type IIb
C1704429|T047|SY|15346004|SNOMEDCT_CORE|Familial high density lipoprotein deficiency|Familial hypoalphalipoproteinemia
C1704429|T047|PTGB|15346004|SNOMEDCT_CORE|Familial hypoalphalipoproteinaemia|Familial hypoalphalipoproteinemia
C1704429|T047|PT|15346004|SNOMEDCT_CORE|Familial hypoalphalipoproteinemia|Familial hypoalphalipoproteinemia
C1704429|T047|FN|15346004|SNOMEDCT_CORE|Familial hypoalphalipoproteinemia|Familial hypoalphalipoproteinemia
C1704436|T047|SY|399957001|SNOMEDCT_CORE|Peripheral arterial disease|Peripheral arterial disease
C1719455|T047|SY|428887009|SNOMEDCT_CORE|Asymmetric sensorineural hearing loss|Asymmetrical sensorineural hearing loss
C1719455|T047|PT|428887009|SNOMEDCT_CORE|Asymmetrical sensorineural hearing loss|Asymmetrical sensorineural hearing loss
C1719455|T047|FN|428887009|SNOMEDCT_CORE|Asymmetrical sensorineural hearing loss|Asymmetrical sensorineural hearing loss
C1719601|T033|SY|430933008|SNOMEDCT_CORE|Gravid uterus size for dates discrepancy|Uterine size for dates discrepancy
C1719601|T033|FN|430933008|SNOMEDCT_CORE|Gravid uterus size for dates discrepancy|Uterine size for dates discrepancy
C1719601|T033|SY|430933008|SNOMEDCT_CORE|Uterine size date discrepancy|Uterine size for dates discrepancy
C1719601|T033|PT|430933008|SNOMEDCT_CORE|Uterine size for dates discrepancy|Uterine size for dates discrepancy
C1719759|T047|IS|421893009|SNOMEDCT_CORE|Kidney disorder associated with juvenile-onset type diabetes mellitus|Renal disorder due to type 1 diabetes mellitus
C1719759|T047|SY|421893009|SNOMEDCT_CORE|Kidney disorder associated with type 1 diabetes mellitus|Renal disorder due to type 1 diabetes mellitus
C1719759|T047|IS|421893009|SNOMEDCT_CORE|Renal disorder associated with insulin dependent diabetes mellitus|Renal disorder due to type 1 diabetes mellitus
C1719759|T047|SY|421893009|SNOMEDCT_CORE|Renal disorder associated with type 1 diabetes mellitus|Renal disorder due to type 1 diabetes mellitus
C1719759|T047|OF|421893009|SNOMEDCT_CORE|Renal disorder associated with type I diabetes mellitus|Renal disorder due to type 1 diabetes mellitus
C1719759|T047|SY|421893009|SNOMEDCT_CORE|Renal disorder associated with type I diabetes mellitus|Renal disorder due to type 1 diabetes mellitus
C1719759|T047|PT|421893009|SNOMEDCT_CORE|Renal disorder due to type 1 diabetes mellitus|Renal disorder due to type 1 diabetes mellitus
C1719759|T047|FN|421893009|SNOMEDCT_CORE|Renal disorder due to type 1 diabetes mellitus|Renal disorder due to type 1 diabetes mellitus
C1719760|T047|SY|421895002|SNOMEDCT_CORE|Diabetic peripheral circulatory disorder|Peripheral vascular disorder due to diabetes mellitus
C1719760|T047|OF|421895002|SNOMEDCT_CORE|Peripheral circulatory disorder associated with diabetes mellitus|Peripheral vascular disorder due to diabetes mellitus
C1719760|T047|SY|421895002|SNOMEDCT_CORE|Peripheral circulatory disorder associated with diabetes mellitus|Peripheral vascular disorder due to diabetes mellitus
C1719760|T047|OF|421895002|SNOMEDCT_CORE|Peripheral vascular disorder co-occurrent and due to diabetes mellitus|Peripheral vascular disorder due to diabetes mellitus
C1719760|T047|IS|421895002|SNOMEDCT_CORE|Peripheral vascular disorder co-occurrent and due to diabetes mellitus|Peripheral vascular disorder due to diabetes mellitus
C1719760|T047|PT|421895002|SNOMEDCT_CORE|Peripheral vascular disorder due to diabetes mellitus|Peripheral vascular disorder due to diabetes mellitus
C1719760|T047|FN|421895002|SNOMEDCT_CORE|Peripheral vascular disorder due to diabetes mellitus|Peripheral vascular disorder due to diabetes mellitus
C1719783|T047|OP|420514000|SNOMEDCT_CORE|Persistent proteinuria associated with type 1 diabetes mellitus|Persistent proteinuria due to type 1 diabetes mellitus
C1719783|T047|OF|420514000|SNOMEDCT_CORE|Persistent proteinuria associated with type I diabetes mellitus|Persistent proteinuria due to type 1 diabetes mellitus
C1719783|T047|IS|420514000|SNOMEDCT_CORE|Persistent proteinuria associated with type I diabetes mellitus|Persistent proteinuria due to type 1 diabetes mellitus
C1719783|T047|PT|420514000|SNOMEDCT_CORE|Persistent proteinuria due to type 1 diabetes mellitus|Persistent proteinuria due to type 1 diabetes mellitus
C1719783|T047|FN|420514000|SNOMEDCT_CORE|Persistent proteinuria due to type 1 diabetes mellitus|Persistent proteinuria due to type 1 diabetes mellitus
C1719786|T191|PT|420519005|SNOMEDCT_CORE|Malignant lymphoma of the eye region|Malignant lymphoma of the eye region
C1719786|T191|FN|420519005|SNOMEDCT_CORE|Malignant lymphoma of the eye region|Malignant lymphoma of the eye region
C1719807|T047|OF|421920002|SNOMEDCT_CORE|Cataract co-occurrent and due to diabetes mellitus type 1|Cataract due to diabetes mellitus type 1
C1719807|T047|IS|421920002|SNOMEDCT_CORE|Cataract co-occurrent and due to diabetes mellitus type 1|Cataract due to diabetes mellitus type 1
C1719807|T047|PT|421920002|SNOMEDCT_CORE|Cataract due to diabetes mellitus type 1|Cataract due to diabetes mellitus type 1
C1719807|T047|FN|421920002|SNOMEDCT_CORE|Cataract of eye due to diabetes mellitus type 1|Cataract due to diabetes mellitus type 1
C1719807|T047|SY|421920002|SNOMEDCT_CORE|Cataract of eye due to diabetes mellitus type 1|Cataract due to diabetes mellitus type 1
C1719807|T047|SY|421920002|SNOMEDCT_CORE|Diabetes type 1 with cataract|Cataract due to diabetes mellitus type 1
C1719807|T047|SY|421920002|SNOMEDCT_CORE|Diabetic cataract associated with type 1 diabetes mellitus|Cataract due to diabetes mellitus type 1
C1719807|T047|OF|421920002|SNOMEDCT_CORE|Diabetic cataract associated with type I diabetes mellitus|Cataract due to diabetes mellitus type 1
C1719807|T047|SY|421920002|SNOMEDCT_CORE|Diabetic cataract associated with type I diabetes mellitus|Cataract due to diabetes mellitus type 1
C1719887|T047|OP|421986006|SNOMEDCT_CORE|Persistent proteinuria associated with type 2 diabetes mellitus|Persistent proteinuria due to type 2 diabetes mellitus
C1719887|T047|OF|421986006|SNOMEDCT_CORE|Persistent proteinuria associated with type II diabetes mellitus|Persistent proteinuria due to type 2 diabetes mellitus
C1719887|T047|IS|421986006|SNOMEDCT_CORE|Persistent proteinuria associated with type II diabetes mellitus|Persistent proteinuria due to type 2 diabetes mellitus
C1719887|T047|PT|421986006|SNOMEDCT_CORE|Persistent proteinuria due to type 2 diabetes mellitus|Persistent proteinuria due to type 2 diabetes mellitus
C1719887|T047|FN|421986006|SNOMEDCT_CORE|Persistent proteinuria due to type 2 diabetes mellitus|Persistent proteinuria due to type 2 diabetes mellitus
C1719929|T047|OP|421305000|SNOMEDCT_CORE|Persistent microalbuminuria associated with type 1 diabetes mellitus|Persistent microalbuminuria due to type 1 diabetes mellitus
C1719929|T047|OF|421305000|SNOMEDCT_CORE|Persistent microalbuminuria associated with type I diabetes mellitus|Persistent microalbuminuria due to type 1 diabetes mellitus
C1719929|T047|SY|421305000|SNOMEDCT_CORE|Persistent microalbuminuria associated with type I diabetes mellitus|Persistent microalbuminuria due to type 1 diabetes mellitus
C1719929|T047|PT|421305000|SNOMEDCT_CORE|Persistent microalbuminuria due to type 1 diabetes mellitus|Persistent microalbuminuria due to type 1 diabetes mellitus
C1719929|T047|FN|421305000|SNOMEDCT_CORE|Persistent microalbuminuria due to type 1 diabetes mellitus|Persistent microalbuminuria due to type 1 diabetes mellitus
C1719939|T047|IS|422014003|SNOMEDCT_CORE|Complication of adult-onset type diabetes mellitus|Disorder due to type 2 diabetes mellitus
C1719939|T047|IS|422014003|SNOMEDCT_CORE|Complication of type II diabetes mellitus|Disorder due to type 2 diabetes mellitus
C1719939|T047|OF|422014003|SNOMEDCT_CORE|Disorder associated with type 2 diabetes mellitus|Disorder due to type 2 diabetes mellitus
C1719939|T047|OP|422014003|SNOMEDCT_CORE|Disorder associated with type 2 diabetes mellitus|Disorder due to type 2 diabetes mellitus
C1719939|T047|OF|422014003|SNOMEDCT_CORE|Disorder associated with type II diabetes melliltus|Disorder due to type 2 diabetes mellitus
C1719939|T047|IS|422014003|SNOMEDCT_CORE|Disorder associated with type II diabetes melliltus|Disorder due to type 2 diabetes mellitus
C1719939|T047|IS|422014003|SNOMEDCT_CORE|Disorder associated with type II diabetes mellitus|Disorder due to type 2 diabetes mellitus
C1719939|T047|PT|422014003|SNOMEDCT_CORE|Disorder due to type 2 diabetes mellitus|Disorder due to type 2 diabetes mellitus
C1719939|T047|FN|422014003|SNOMEDCT_CORE|Disorder due to type 2 diabetes mellitus|Disorder due to type 2 diabetes mellitus
C1719939|T047|SY|422014003|SNOMEDCT_CORE|Disorder due to type II diabetes mellitus|Disorder due to type 2 diabetes mellitus
C1719988|T047|IS|421326000|SNOMEDCT_CORE|Diabetes type 2 with neurological disorder|Disorder of nervous system due to type 2 diabetes mellitus
C1719988|T047|PT|421326000|SNOMEDCT_CORE|Disorder of nervous system due to type 2 diabetes mellitus|Disorder of nervous system due to type 2 diabetes mellitus
C1719988|T047|FN|421326000|SNOMEDCT_CORE|Disorder of nervous system due to type 2 diabetes mellitus|Disorder of nervous system due to type 2 diabetes mellitus
C1719988|T047|IS|421326000|SNOMEDCT_CORE|Neurologic complication of adult-onset type diabetes mellitus|Disorder of nervous system due to type 2 diabetes mellitus
C1719988|T047|SY|421326000|SNOMEDCT_CORE|Neurologic disorder associated with type 2 diabetes mellitus|Disorder of nervous system due to type 2 diabetes mellitus
C1719988|T047|OF|421326000|SNOMEDCT_CORE|Neurologic disorder associated with type II diabetes mellitus|Disorder of nervous system due to type 2 diabetes mellitus
C1719988|T047|SY|421326000|SNOMEDCT_CORE|Neurologic disorder associated with type II diabetes mellitus|Disorder of nervous system due to type 2 diabetes mellitus
C1719988|T047|OF|421326000|SNOMEDCT_CORE|Neurological disorder co-occurrent and due to type 2 diabetes mellitus|Disorder of nervous system due to type 2 diabetes mellitus
C1719988|T047|IS|421326000|SNOMEDCT_CORE|Neurological disorder co-occurrent and due to type 2 diabetes mellitus|Disorder of nervous system due to type 2 diabetes mellitus
C1719988|T047|OP|421326000|SNOMEDCT_CORE|Neurological disorder with diabetes type 2|Disorder of nervous system due to type 2 diabetes mellitus
C1719988|T047|SY|421326000|SNOMEDCT_CORE|Neurological disorder with type 2 diabetes mellitus|Disorder of nervous system due to type 2 diabetes mellitus
C1720056|T047|IS|421365002|SNOMEDCT_CORE|Peripheral circulatory disorder associated with insulin-dependent diabetes mellitus|Peripheral circulatory disorder due to type 1 diabetes mellitus
C1720056|T047|IS|421365002|SNOMEDCT_CORE|Peripheral circulatory disorder associated with juvenile-onset type diabetes mellitus|Peripheral circulatory disorder due to type 1 diabetes mellitus
C1720056|T047|SY|421365002|SNOMEDCT_CORE|Peripheral circulatory disorder associated with type 1 diabetes mellitus|Peripheral circulatory disorder due to type 1 diabetes mellitus
C1720056|T047|OF|421365002|SNOMEDCT_CORE|Peripheral circulatory disorder associated with type I diabetes mellitus|Peripheral circulatory disorder due to type 1 diabetes mellitus
C1720056|T047|IS|421365002|SNOMEDCT_CORE|Peripheral circulatory disorder associated with type I diabetes mellitus|Peripheral circulatory disorder due to type 1 diabetes mellitus
C1720056|T047|PT|421365002|SNOMEDCT_CORE|Peripheral circulatory disorder due to type 1 diabetes mellitus|Peripheral circulatory disorder due to type 1 diabetes mellitus
C1720056|T047|FN|421365002|SNOMEDCT_CORE|Peripheral circulatory disorder due to type 1 diabetes mellitus|Peripheral circulatory disorder due to type 1 diabetes mellitus
C1720078|T047|SY|422088007|SNOMEDCT_CORE|Diabetic neurologic disease|Disorder of nervous system due to diabetes mellitus
C1720078|T047|IS|422088007|SNOMEDCT_CORE|Disorder of nervous system co-occurrent and due to diabetes mellitus|Disorder of nervous system due to diabetes mellitus
C1720078|T047|OF|422088007|SNOMEDCT_CORE|Disorder of nervous system co-occurrent and due to diabetes mellitus|Disorder of nervous system due to diabetes mellitus
C1720078|T047|PT|422088007|SNOMEDCT_CORE|Disorder of nervous system due to diabetes mellitus|Disorder of nervous system due to diabetes mellitus
C1720078|T047|FN|422088007|SNOMEDCT_CORE|Disorder of nervous system due to diabetes mellitus|Disorder of nervous system due to diabetes mellitus
C1720078|T047|SY|422088007|SNOMEDCT_CORE|Nervous system disorder due to diabetes mellitus|Disorder of nervous system due to diabetes mellitus
C1720078|T047|SY|422088007|SNOMEDCT_CORE|Neurologic complication of diabetes mellitus|Disorder of nervous system due to diabetes mellitus
C1720078|T047|OF|422088007|SNOMEDCT_CORE|Neurologic disorder associated with diabetes mellitus|Disorder of nervous system due to diabetes mellitus
C1720078|T047|SY|422088007|SNOMEDCT_CORE|Neurologic disorder associated with diabetes mellitus|Disorder of nervous system due to diabetes mellitus
C1720102|T047|IS|420715001|SNOMEDCT_CORE|Persistent microalbuminuria associated with adult-onset type diabetes mellitus|Persistent microalbuminuria due to type 2 diabetes mellitus
C1720102|T047|IS|420715001|SNOMEDCT_CORE|Persistent microalbuminuria associated with non-insulin dependent diabetes mellitus|Persistent microalbuminuria due to type 2 diabetes mellitus
C1720102|T047|OP|420715001|SNOMEDCT_CORE|Persistent microalbuminuria associated with type 2 diabetes mellitus|Persistent microalbuminuria due to type 2 diabetes mellitus
C1720102|T047|OF|420715001|SNOMEDCT_CORE|Persistent microalbuminuria associated with type II diabetes mellitus|Persistent microalbuminuria due to type 2 diabetes mellitus
C1720102|T047|SY|420715001|SNOMEDCT_CORE|Persistent microalbuminuria associated with type II diabetes mellitus|Persistent microalbuminuria due to type 2 diabetes mellitus
C1720102|T047|PT|420715001|SNOMEDCT_CORE|Persistent microalbuminuria due to type 2 diabetes mellitus|Persistent microalbuminuria due to type 2 diabetes mellitus
C1720102|T047|FN|420715001|SNOMEDCT_CORE|Persistent microalbuminuria due to type 2 diabetes mellitus|Persistent microalbuminuria due to type 2 diabetes mellitus
C1720165|T047|IS|422166005|SNOMEDCT_CORE|Peripheral circulatory disorder associated with adult-onset type diabetes mellitus|Peripheral circulatory disorder due to type 2 diabetes mellitus
C1720165|T047|IS|422166005|SNOMEDCT_CORE|Peripheral circulatory disorder associated with non-insulin dependent diabetes mellitus|Peripheral circulatory disorder due to type 2 diabetes mellitus
C1720165|T047|SY|422166005|SNOMEDCT_CORE|Peripheral circulatory disorder associated with type 2 diabetes mellitus|Peripheral circulatory disorder due to type 2 diabetes mellitus
C1720165|T047|OF|422166005|SNOMEDCT_CORE|Peripheral circulatory disorder associated with type II diabetes mellitus|Peripheral circulatory disorder due to type 2 diabetes mellitus
C1720165|T047|IS|422166005|SNOMEDCT_CORE|Peripheral circulatory disorder associated with type II diabetes mellitus|Peripheral circulatory disorder due to type 2 diabetes mellitus
C1720165|T047|PT|422166005|SNOMEDCT_CORE|Peripheral circulatory disorder due to type 2 diabetes mellitus|Peripheral circulatory disorder due to type 2 diabetes mellitus
C1720165|T047|FN|422166005|SNOMEDCT_CORE|Peripheral circulatory disorder due to type 2 diabetes mellitus|Peripheral circulatory disorder due to type 2 diabetes mellitus
C1720194|T047|SY|421468001|SNOMEDCT_CORE|Diabetes type 1 with neurological disorder|Disorder of nervous system due to type 1 diabetes mellitus
C1720194|T047|PT|421468001|SNOMEDCT_CORE|Disorder of nervous system due to type 1 diabetes mellitus|Disorder of nervous system due to type 1 diabetes mellitus
C1720194|T047|FN|421468001|SNOMEDCT_CORE|Disorder of nervous system due to type 1 diabetes mellitus|Disorder of nervous system due to type 1 diabetes mellitus
C1720194|T047|IS|421468001|SNOMEDCT_CORE|Neurologic complication of juvenile-onset diabetes mellitus|Disorder of nervous system due to type 1 diabetes mellitus
C1720194|T047|SY|421468001|SNOMEDCT_CORE|Neurological disorder associated with type 1 diabetes mellitus|Disorder of nervous system due to type 1 diabetes mellitus
C1720194|T047|OF|421468001|SNOMEDCT_CORE|Neurological disorder associated with type I diabetes mellitus|Disorder of nervous system due to type 1 diabetes mellitus
C1720194|T047|SY|421468001|SNOMEDCT_CORE|Neurological disorder associated with type I diabetes mellitus|Disorder of nervous system due to type 1 diabetes mellitus
C1720194|T047|IS|421468001|SNOMEDCT_CORE|Neurological disorder co-occurrent and due to type 1 diabetes mellitus|Disorder of nervous system due to type 1 diabetes mellitus
C1720194|T047|OF|421468001|SNOMEDCT_CORE|Neurological disorder co-occurrent and due to type 1 diabetes mellitus|Disorder of nervous system due to type 1 diabetes mellitus
C1720194|T047|SY|421468001|SNOMEDCT_CORE|Neurological disorder with type 1 diabetes mellitus|Disorder of nervous system due to type 1 diabetes mellitus
C1720297|T047|IS|420868002|SNOMEDCT_CORE|Complication of insulin-dependent diabetes mellitus|Disorder due to type 1 diabetes mellitus
C1720297|T047|IS|420868002|SNOMEDCT_CORE|Complication of juvenile-onset type diabetes mellitus|Disorder due to type 1 diabetes mellitus
C1720297|T047|IS|420868002|SNOMEDCT_CORE|Complication of type I diabetes mellitus|Disorder due to type 1 diabetes mellitus
C1720297|T047|OP|420868002|SNOMEDCT_CORE|Disorder associated with type 1 diabetes mellitus|Disorder due to type 1 diabetes mellitus
C1720297|T047|OF|420868002|SNOMEDCT_CORE|Disorder associated with type I diabetes mellitus|Disorder due to type 1 diabetes mellitus
C1720297|T047|SY|420868002|SNOMEDCT_CORE|Disorder associated with type I diabetes mellitus|Disorder due to type 1 diabetes mellitus
C1720297|T047|PT|420868002|SNOMEDCT_CORE|Disorder due to type 1 diabetes mellitus|Disorder due to type 1 diabetes mellitus
C1720297|T047|FN|420868002|SNOMEDCT_CORE|Disorder due to type 1 diabetes mellitus|Disorder due to type 1 diabetes mellitus
C1720457|T047|SY|420279001|SNOMEDCT_CORE|Diabetes type 2 with nephropathy|Renal disorder due to type 2 diabetes mellitus
C1720457|T047|IS|420279001|SNOMEDCT_CORE|Kidney disorder associated with adult-onset type diabetes mellitus|Renal disorder due to type 2 diabetes mellitus
C1720457|T047|SY|420279001|SNOMEDCT_CORE|Kidney disorder associated with type 2 diabetes mellitus|Renal disorder due to type 2 diabetes mellitus
C1720457|T047|IS|420279001|SNOMEDCT_CORE|Renal disorder associated with non-insulin dependent diabetes mellitus|Renal disorder due to type 2 diabetes mellitus
C1720457|T047|OP|420279001|SNOMEDCT_CORE|Renal disorder associated with type 2 diabetes mellitus|Renal disorder due to type 2 diabetes mellitus
C1720457|T047|OF|420279001|SNOMEDCT_CORE|Renal disorder associated with type II diabetes mellitus|Renal disorder due to type 2 diabetes mellitus
C1720457|T047|SY|420279001|SNOMEDCT_CORE|Renal disorder associated with type II diabetes mellitus|Renal disorder due to type 2 diabetes mellitus
C1720457|T047|PT|420279001|SNOMEDCT_CORE|Renal disorder due to type 2 diabetes mellitus|Renal disorder due to type 2 diabetes mellitus
C1720457|T047|FN|420279001|SNOMEDCT_CORE|Renal disorder due to type 2 diabetes mellitus|Renal disorder due to type 2 diabetes mellitus
C1720557|T047|OAS|421707005|SNOMEDCT_CORE|Diabetes type 2 with diabetic polyneuropathy|Polyneuropathy associated with type 2 diabetes mellitus
C1720557|T047|IS|421707005|SNOMEDCT_CORE|Polyneuropathy associated with adult-onset type diabetes mellitus|Polyneuropathy associated with type 2 diabetes mellitus
C1720557|T047|IS|421707005|SNOMEDCT_CORE|Polyneuropathy associated with non-insulin dependent diabetes mellitus|Polyneuropathy associated with type 2 diabetes mellitus
C1720557|T047|OAP|421707005|SNOMEDCT_CORE|Polyneuropathy associated with type 2 diabetes mellitus|Polyneuropathy associated with type 2 diabetes mellitus
C1720557|T047|OAF|421707005|SNOMEDCT_CORE|Polyneuropathy associated with type II diabetes mellitus|Polyneuropathy associated with type 2 diabetes mellitus
C1720557|T047|OAS|421707005|SNOMEDCT_CORE|Polyneuropathy associated with type II diabetes mellitus|Polyneuropathy associated with type 2 diabetes mellitus
C1720648|T047|IS|420436000|SNOMEDCT_CORE|Mononeuropathy associated with non-insulin dependent diabetes mellitus|Mononeuropathy due to type 2 diabetes mellitus
C1720648|T047|IS|420436000|SNOMEDCT_CORE|Mononeuropathy associated with type 2 diabetes mellitus|Mononeuropathy due to type 2 diabetes mellitus
C1720648|T047|OF|420436000|SNOMEDCT_CORE|Mononeuropathy associated with type II diabetes mellitus|Mononeuropathy due to type 2 diabetes mellitus
C1720648|T047|IS|420436000|SNOMEDCT_CORE|Mononeuropathy associated with type II diabetes mellitus|Mononeuropathy due to type 2 diabetes mellitus
C1720648|T047|IS|420436000|SNOMEDCT_CORE|Mononeuropathy co-occurrent and due to type 2 diabetes mellitus|Mononeuropathy due to type 2 diabetes mellitus
C1720648|T047|OF|420436000|SNOMEDCT_CORE|Mononeuropathy co-occurrent and due to type 2 diabetes mellitus|Mononeuropathy due to type 2 diabetes mellitus
C1720648|T047|PT|420436000|SNOMEDCT_CORE|Mononeuropathy due to type 2 diabetes mellitus|Mononeuropathy due to type 2 diabetes mellitus
C1720648|T047|FN|420436000|SNOMEDCT_CORE|Mononeuropathy due to type 2 diabetes mellitus|Mononeuropathy due to type 2 diabetes mellitus
C1720648|T047|SY|420436000|SNOMEDCT_CORE|Mononeuropathy with type 2 diabetes mellitus|Mononeuropathy due to type 2 diabetes mellitus
C1720717|T047|OAP|421165007|SNOMEDCT_CORE|Diabetic oculopathy associated with type 1 diabetes mellitus|Diabetic oculopathy associated with type 1 diabetes mellitus
C1720717|T047|OAF|421165007|SNOMEDCT_CORE|Diabetic oculopathy associated with type I diabetes mellitus|Diabetic oculopathy associated with type 1 diabetes mellitus
C1720717|T047|OAS|421165007|SNOMEDCT_CORE|Diabetic oculopathy associated with type I diabetes mellitus|Diabetic oculopathy associated with type 1 diabetes mellitus
C1720771|T019|PT|26614003|SNOMEDCT_CORE|Hydrocele of testis|Hydrocele of testis
C1720771|T019|FN|26614003|SNOMEDCT_CORE|Hydrocele of testis|Hydrocele of testis
C1735856|T047|SY|4473006|SNOMEDCT_CORE|Classical migraine|Migraine with typical aura
C1735856|T047|PT|230462002|SNOMEDCT_CORE|Migraine with typical aura|Migraine with typical aura
C1735856|T047|FN|230462002|SNOMEDCT_CORE|Migraine with typical aura|Migraine with typical aura
C1735914|T047|PT|438773007|SNOMEDCT_CORE|Recurrent pulmonary embolism|Recurrent pulmonary embolism
C1735914|T047|FN|438773007|SNOMEDCT_CORE|Recurrent pulmonary embolism|Recurrent pulmonary embolism
C1737329|T019|SY|276720006|SNOMEDCT_CORE|Birth defect|Dysmorphism
C1737329|T019|SY|276720006|SNOMEDCT_CORE|Dysmorphia|Dysmorphism
C1737329|T019|PT|276720006|SNOMEDCT_CORE|Dysmorphism|Dysmorphism
C1737329|T019|FN|276720006|SNOMEDCT_CORE|Dysmorphism|Dysmorphism
C1739363|T047|SY|266569009|SNOMEDCT_CORE|Prostatic area hypertrophy|Prostatic area hypertrophy
C1739363|T047|SY|266569009|SNOMEDCT_CORE|Prostatic hypertrophy|Prostatic area hypertrophy
C1740754|T047|PT|427603009|SNOMEDCT_CORE|Intermittent asthma|Intermittent asthma
C1740754|T047|FN|427603009|SNOMEDCT_CORE|Intermittent asthma|Intermittent asthma
C1800706|T047|SY|700250006|SNOMEDCT_CORE|Cryptogenic fibrosing alveolitis|Idiopathic pulmonary fibrosis
C1800706|T047|SY|700250006|SNOMEDCT_CORE|Idiopathic fibrosing alveolitis|Idiopathic pulmonary fibrosis
C1800706|T047|PT|700250006|SNOMEDCT_CORE|Idiopathic pulmonary fibrosis|Idiopathic pulmonary fibrosis
C1800706|T047|FN|700250006|SNOMEDCT_CORE|Idiopathic pulmonary fibrosis|Idiopathic pulmonary fibrosis
C1800706|T047|SY|700250006|SNOMEDCT_CORE|Usual interstitial pneumonia|Idiopathic pulmonary fibrosis
C1827052|T047|SY|423683008|SNOMEDCT_CORE|Classical migraine, intractable|Refractory migraine with aura
C1827052|T047|SY|423683008|SNOMEDCT_CORE|Intractable classical migraine|Refractory migraine with aura
C1827052|T047|SY|423683008|SNOMEDCT_CORE|Intractable migraine with aura|Refractory migraine with aura
C1827052|T047|PT|423683008|SNOMEDCT_CORE|Refractory migraine with aura|Refractory migraine with aura
C1827052|T047|FN|423683008|SNOMEDCT_CORE|Refractory migraine with aura|Refractory migraine with aura
C1827090|T033|PT|424959007|SNOMEDCT_CORE|Foreign body of neck|Foreign body of neck
C1827090|T033|FN|424959007|SNOMEDCT_CORE|Foreign body of neck|Foreign body of neck
C1827143|T191|SY|423700001|SNOMEDCT_CORE|Squamous cell carcinoma of auricle|Squamous cell carcinoma of auricle of ear
C1827143|T191|PT|423700001|SNOMEDCT_CORE|Squamous cell carcinoma of auricle of ear|Squamous cell carcinoma of auricle of ear
C1827143|T191|FN|423700001|SNOMEDCT_CORE|Squamous cell carcinoma of auricle of ear|Squamous cell carcinoma of auricle of ear
C1827143|T191|SY|423700001|SNOMEDCT_CORE|Squamous cell carcinoma of pinna|Squamous cell carcinoma of auricle of ear
C1827179|T047|OAS|424989000|SNOMEDCT_CORE|Diabetes type 2 with gastroparesis|Diabetic gastroparesis associated with type 2 diabetes mellitus
C1827179|T047|OAP|424989000|SNOMEDCT_CORE|Diabetic gastroparesis associated with type 2 diabetes mellitus|Diabetic gastroparesis associated with type 2 diabetes mellitus
C1827179|T047|OAF|424989000|SNOMEDCT_CORE|Diabetic gastroparesis associated with type 2 diabetes mellitus|Diabetic gastroparesis associated with type 2 diabetes mellitus
C1827190|T047|SY|425007008|SNOMEDCT_CORE|Common migraine, not intractable|Migraine without aura, not refractory
C1827190|T047|SY|425007008|SNOMEDCT_CORE|Migraine without aura, non-intractable|Migraine without aura, not refractory
C1827190|T047|PT|425007008|SNOMEDCT_CORE|Migraine without aura, not refractory|Migraine without aura, not refractory
C1827190|T047|FN|425007008|SNOMEDCT_CORE|Migraine without aura, not refractory|Migraine without aura, not refractory
C1827192|T047|PT|425011002|SNOMEDCT_CORE|Allergic fungal sinusitis|Allergic fungal sinusitis
C1827192|T047|FN|425011002|SNOMEDCT_CORE|Allergic fungal sinusitis|Allergic fungal sinusitis
C1827431|T191|PT|423812005|SNOMEDCT_CORE|Sarcoma of head and neck|Sarcoma of head and neck
C1827431|T191|FN|423812005|SNOMEDCT_CORE|Sarcoma of head and neck|Sarcoma of head and neck
C1827502|T191|PT|422572002|SNOMEDCT_CORE|Squamous cell carcinoma of chin|Squamous cell carcinoma of chin
C1827502|T191|FN|422572002|SNOMEDCT_CORE|Squamous cell carcinoma of chin|Squamous cell carcinoma of chin
C1827522|T047|PT|423226005|SNOMEDCT_CORE|Tendinitis of finger|Tendinitis of finger
C1827522|T047|FN|423226005|SNOMEDCT_CORE|Tendinitis of finger|Tendinitis of finger
C1827522|T047|SY|423226005|SNOMEDCT_CORE|Tendonitis of finger|Tendinitis of finger
C1827624|T047|SY|423279000|SNOMEDCT_CORE|Common migraine without aura, intractable|Refractory migraine without aura
C1827624|T047|SY|423279000|SNOMEDCT_CORE|Intractable common migraine|Refractory migraine without aura
C1827624|T047|SY|423279000|SNOMEDCT_CORE|Intractable migraine without aura|Refractory migraine without aura
C1827624|T047|PT|423279000|SNOMEDCT_CORE|Refractory migraine without aura|Refractory migraine without aura
C1827624|T047|FN|423279000|SNOMEDCT_CORE|Refractory migraine without aura|Refractory migraine without aura
C1827687|T046|OAP|425229001|SNOMEDCT_CORE|Chemotherapy-induced neutropenia|Chemotherapy-induced neutropenia
C1827687|T046|OAF|425229001|SNOMEDCT_CORE|Chemotherapy-induced neutropenia|Chemotherapy-induced neutropenia
C1827711|T191|SY|423284006|SNOMEDCT_CORE|Cancer of skin of neck, squamous cell|Squamous cell carcinoma of skin of neck
C1827711|T191|PT|423284006|SNOMEDCT_CORE|Squamous cell carcinoma of skin of neck|Squamous cell carcinoma of skin of neck
C1827711|T191|FN|423284006|SNOMEDCT_CORE|Squamous cell carcinoma of skin of neck|Squamous cell carcinoma of skin of neck
C1827851|T037|PT|424648000|SNOMEDCT_CORE|Closed fracture of base of fifth metatarsal bone|Closed fracture of base of fifth metatarsal bone
C1827851|T037|FN|424648000|SNOMEDCT_CORE|Closed fracture of base of fifth metatarsal bone|Closed fracture of base of fifth metatarsal bone
C1827966|T047|PT|424699007|SNOMEDCT_CORE|Migraine variants, not intractable|Migraine variants, not intractable
C1827966|T047|FN|424699007|SNOMEDCT_CORE|Migraine variants, not intractable|Migraine variants, not intractable
C1828009|T047|PT|423417009|SNOMEDCT_CORE|Tendinitis of hand|Tendinitis of hand
C1828009|T047|FN|423417009|SNOMEDCT_CORE|Tendinitis of hand|Tendinitis of hand
C1828009|T047|SY|423417009|SNOMEDCT_CORE|Tendonitis of hand|Tendinitis of hand
C1828079|T048|SY|425390006|SNOMEDCT_CORE|Dementia associated with Parkinson Disease|Dementia associated with Parkinson's Disease
C1828079|T048|PT|425390006|SNOMEDCT_CORE|Dementia associated with Parkinson's Disease|Dementia associated with Parkinson's Disease
C1828079|T048|FN|425390006|SNOMEDCT_CORE|Dementia associated with Parkinson's Disease|Dementia associated with Parkinson's Disease
C1828079|T048|SY|425390006|SNOMEDCT_CORE|Dementia in Parkinsons disease|Dementia associated with Parkinson's Disease
C1828173|T033|PT|422868009|SNOMEDCT_CORE|Unexplained weight loss|Unexplained weight loss
C1828173|T033|FN|422868009|SNOMEDCT_CORE|Unexplained weight loss|Unexplained weight loss
C1828213|T047|PT|424175006|SNOMEDCT_CORE|Nontraumatic rotator cuff tear|Nontraumatic rotator cuff tear
C1828213|T047|FN|424175006|SNOMEDCT_CORE|Nontraumatic rotator cuff tear|Nontraumatic rotator cuff tear
C1833142|T020|PT|239734000|SNOMEDCT_CORE|Contracture of elbow joint|Contracture of elbow joint
C1833142|T020|FN|239734000|SNOMEDCT_CORE|Contracture of elbow joint|Contracture of elbow joint
C1833142|T020|SY|239734000|SNOMEDCT_CORE|Elbow joint contracture|Contracture of elbow joint
C1840475|T047|SY|770626007|SNOMEDCT_CORE|Congenital Claude Bernard Horner syndrome|Congenital Horner syndrome
C1840475|T047|PT|770626007|SNOMEDCT_CORE|Congenital Horner syndrome|Congenital Horner syndrome
C1840475|T047|FN|770626007|SNOMEDCT_CORE|Congenital Horner syndrome|Congenital Horner syndrome
C1844383|T033|PT|428875002|SNOMEDCT_CORE|Recurrent bacterial infection|Recurrent bacterial infection
C1844383|T033|FN|428875002|SNOMEDCT_CORE|Recurrent bacterial infection|Recurrent bacterial infection
C1844820|T033|IS|298181000|SNOMEDCT_CORE|Hypermobility of joint|Range of joint movement increased
C1844820|T033|IS|298181000|SNOMEDCT_CORE|Joint hypermobility|Range of joint movement increased
C1844820|T033|PT|298181000|SNOMEDCT_CORE|Range of joint movement increased|Range of joint movement increased
C1844820|T033|FN|298181000|SNOMEDCT_CORE|Range of joint movement increased|Range of joint movement increased
C1848954|T033|PTGB|425492002|SNOMEDCT_CORE|Generalised dystonia|Generalized dystonia
C1848954|T033|PT|425492002|SNOMEDCT_CORE|Generalized dystonia|Generalized dystonia
C1848954|T033|FN|425492002|SNOMEDCT_CORE|Generalized dystonia|Generalized dystonia
C1850534|T046|PT|271808008|SNOMEDCT_CORE|Edema, generalized|Edema, generalized
C1850534|T046|FN|271808008|SNOMEDCT_CORE|Edema, generalized|Edema, generalized
C1850534|T046|PTGB|271808008|SNOMEDCT_CORE|Oedema, generalised|Edema, generalized
C1853729|T033|PT|445424004|SNOMEDCT_CORE|Weakness of vocal cord|Weakness of vocal cord
C1853729|T033|FN|445424004|SNOMEDCT_CORE|Weakness of vocal cord|Weakness of vocal cord
C1868851|T047|SY|445237003|SNOMEDCT_CORE|Portopulmonary hypertension|Pulmonary arterial hypertension associated with portal hypertension
C1868851|T047|FN|445237003|SNOMEDCT_CORE|Portopulmonary hypertension|Pulmonary arterial hypertension associated with portal hypertension
C1868851|T047|PT|445237003|SNOMEDCT_CORE|Pulmonary arterial hypertension associated with portal hypertension|Pulmonary arterial hypertension associated with portal hypertension
C1879321|T191|PTGB|359648001|SNOMEDCT_CORE|Acute myeloid leukaemia with maturation, FAB M2|Acute myeloid leukemia with maturation, FAB M2
C1879321|T191|FN|359648001|SNOMEDCT_CORE|Acute myeloid leukemia with maturation, FAB M2|Acute myeloid leukemia with maturation, FAB M2
C1879321|T191|PT|359648001|SNOMEDCT_CORE|Acute myeloid leukemia with maturation, FAB M2|Acute myeloid leukemia with maturation, FAB M2
C1879321|T191|SYGB|359648001|SNOMEDCT_CORE|M2 - Acute myeloblastic leukaemia with maturation|Acute myeloid leukemia with maturation, FAB M2
C1879321|T191|SY|359648001|SNOMEDCT_CORE|M2 - Acute myeloblastic leukemia with maturation|Acute myeloid leukemia with maturation, FAB M2
C1879328|T047|FN|193699007|SNOMEDCT_CORE|Blindness - both eyes|Blindness - both eyes
C1879328|T047|PT|193699007|SNOMEDCT_CORE|Blindness - both eyes|Blindness - both eyes
C1879328|T047|SY|193699007|SNOMEDCT_CORE|Both eyes total visual impairment|Blindness - both eyes
C1879338|T033|PT|74506000|SNOMEDCT_CORE|Bereavement|Bereavement
C1879338|T033|FN|74506000|SNOMEDCT_CORE|Bereavement due to life event|Bereavement
C1879338|T033|SY|74506000|SNOMEDCT_CORE|Bereavement due to life event|Bereavement
C1879338|T033|SY|74506000|SNOMEDCT_CORE|Bereavement reaction|Bereavement
C1879338|T033|OF|74506000|SNOMEDCT_CORE|Bereavement, life event|Bereavement
C1879338|T033|SY|74506000|SNOMEDCT_CORE|Mourning|Bereavement
C1882062|T191|SY|55342001|SNOMEDCT_CORE|Neoplasia|Neoplastic disease
C1882062|T191|SY|55342001|SNOMEDCT_CORE|Neoplasm|Neoplastic disease
C1882062|T191|PT|55342001|SNOMEDCT_CORE|Neoplastic disease|Neoplastic disease
C1882062|T191|FN|55342001|SNOMEDCT_CORE|Neoplastic disease|Neoplastic disease
C1882062|T191|IS|55342001|SNOMEDCT_CORE|Neoplastic disease, NOS|Neoplastic disease
C1882062|T191|SY|55342001|SNOMEDCT_CORE|Neoplastic growth|Neoplastic disease
C1882062|T191|IS|55342001|SNOMEDCT_CORE|Neoplastic syndrome|Neoplastic disease
C1882062|T191|IS|55342001|SNOMEDCT_CORE|Neoplastic syndrome, NOS|Neoplastic disease
C1882062|T191|SY|55342001|SNOMEDCT_CORE|New growth|Neoplastic disease
C1882062|T191|SY|55342001|SNOMEDCT_CORE|NG - Neoplastic growth|Neoplastic disease
C1882062|T191|SY|55342001|SNOMEDCT_CORE|NG - New growth|Neoplastic disease
C1956346|T047|SY|53741008|SNOMEDCT_CORE|CAD - Coronary artery disease|CAD - Coronary artery disease
C1956346|T047|SY|53741008|SNOMEDCT_CORE|Coronary artery disease|CAD - Coronary artery disease
C1956390|T047|SY|400130008|SNOMEDCT_CORE|Cranial arteritis|Cranial arteritis
C1956391|T047|SY|400130008|SNOMEDCT_CORE|Giant cell arteritis|Temporal arteritis
C1956391|T047|SY|400130008|SNOMEDCT_CORE|TA - Temporal arteritis|Temporal arteritis
C1956391|T047|PT|400130008|SNOMEDCT_CORE|Temporal arteritis|Temporal arteritis
C1956391|T047|FN|400130008|SNOMEDCT_CORE|Temporal arteritis|Temporal arteritis
C1956391|T047|SY|400130008|SNOMEDCT_CORE|Temporal giant cell arteritis|Temporal arteritis
C1956412|T019|IS|7484005|SNOMEDCT_CORE|Double outlet right ventricle with subpulmonary ventricular septal defect|Double outlet right ventricle with subpulmonary ventricular septal defect
C1956413|T019|SY|7484005|SNOMEDCT_CORE|Taussig-Bing defect|Taussig-Bing defect
C1956413|T019|SY|7484005|SNOMEDCT_CORE|Taussig-Bing syndrome|Taussig-Bing defect
C1959583|T047|SY|84114007|SNOMEDCT_CORE|Myocardial failure|Myocardial failure
C1959583|T047|IS|84114007|SNOMEDCT_CORE|Myocardial failure, NOS|Myocardial failure
C1959799|T047|PT|427649000|SNOMEDCT_CORE|Calcium renal calculus|Calcium renal calculus
C1959799|T047|FN|427649000|SNOMEDCT_CORE|Calcium renal calculus|Calcium renal calculus
C1959850|T047|PT|425772008|SNOMEDCT_CORE|Tendinitis of foot|Tendinitis of foot
C1959850|T047|FN|425772008|SNOMEDCT_CORE|Tendinitis of foot|Tendinitis of foot
C1959850|T047|SY|425772008|SNOMEDCT_CORE|Tendonitis of foot|Tendinitis of foot
C1960030|T047|PT|426014000|SNOMEDCT_CORE|Fistula of hard palate|Fistula of hard palate
C1960030|T047|FN|426014000|SNOMEDCT_CORE|Fistula of hard palate|Fistula of hard palate
C1960036|T048|PT|425832009|SNOMEDCT_CORE|Psychophysiologic insomnia|Psychophysiologic insomnia
C1960036|T048|FN|425832009|SNOMEDCT_CORE|Psychophysiologic insomnia|Psychophysiologic insomnia
C1960040|T047|PT|426033005|SNOMEDCT_CORE|Dysphagia as a late effect of cerebrovascular accident|Dysphagia as a late effect of cerebrovascular accident
C1960040|T047|FN|426033005|SNOMEDCT_CORE|Dysphagia as a late effect of cerebrovascular accident|Dysphagia as a late effect of cerebrovascular accident
C1960040|T047|SY|426033005|SNOMEDCT_CORE|Dysphagia, late effect of stroke|Dysphagia as a late effect of cerebrovascular accident
C1960045|T047|PT|427679007|SNOMEDCT_CORE|Mild intermittent asthma|Mild intermittent asthma
C1960045|T047|FN|427679007|SNOMEDCT_CORE|Mild intermittent asthma|Mild intermittent asthma
C1960046|T047|PT|426979002|SNOMEDCT_CORE|Mild persistent asthma|Mild persistent asthma
C1960046|T047|FN|426979002|SNOMEDCT_CORE|Mild persistent asthma|Mild persistent asthma
C1960047|T047|PT|427295004|SNOMEDCT_CORE|Moderate persistent asthma|Moderate persistent asthma
C1960047|T047|FN|427295004|SNOMEDCT_CORE|Moderate persistent asthma|Moderate persistent asthma
C1960048|T047|PT|426656000|SNOMEDCT_CORE|Severe persistent asthma|Severe persistent asthma
C1960048|T047|FN|426656000|SNOMEDCT_CORE|Severe persistent asthma|Severe persistent asthma
C1960052|T047|PT|426896000|SNOMEDCT_CORE|Chronic hypercapnic respiratory failure|Chronic hypercapnic respiratory failure
C1960052|T047|FN|426896000|SNOMEDCT_CORE|Chronic hypercapnic respiratory failure|Chronic hypercapnic respiratory failure
C1960052|T047|SY|426896000|SNOMEDCT_CORE|Chronic type 2 respiratory failure|Chronic hypercapnic respiratory failure
C1960052|T047|SY|426896000|SNOMEDCT_CORE|Chronic type II respiratory failure|Chronic hypercapnic respiratory failure
C1960174|T047|PT|426508001|SNOMEDCT_CORE|Ileal pouchitis|Ileal pouchitis
C1960174|T047|FN|426508001|SNOMEDCT_CORE|Ileal pouchitis|Ileal pouchitis
C1960195|T037|SY|426912003|SNOMEDCT_CORE|Splinter|Splinter foreign body
C1960195|T037|PT|426912003|SNOMEDCT_CORE|Splinter foreign body|Splinter foreign body
C1960195|T037|PT|443678007|SNOMEDCT_CORE|Splinter foreign body|Splinter foreign body
C1960195|T037|FN|426912003|SNOMEDCT_CORE|Splinter foreign body|Splinter foreign body
C1960195|T037|FN|443678007|SNOMEDCT_CORE|Splinter foreign body|Splinter foreign body
C1960453|T047|PT|427547007|SNOMEDCT_CORE|Female infertility due to diminished ovarian reserve|Female infertility due to diminished ovarian reserve
C1960453|T047|FN|427547007|SNOMEDCT_CORE|Female infertility due to diminished ovarian reserve|Female infertility due to diminished ovarian reserve
C1960678|T047|IS|712882000|SNOMEDCT_CORE|Autonomic neuropathy co-occurrent and due to type 1 diabetes mellitus|Autonomic neuropathy due to type 1 diabetes mellitus
C1960678|T047|OF|712882000|SNOMEDCT_CORE|Autonomic neuropathy co-occurrent and due to type 1 diabetes mellitus|Autonomic neuropathy due to type 1 diabetes mellitus
C1960678|T047|PT|712882000|SNOMEDCT_CORE|Autonomic neuropathy due to type 1 diabetes mellitus|Autonomic neuropathy due to type 1 diabetes mellitus
C1960678|T047|FN|712882000|SNOMEDCT_CORE|Autonomic neuropathy due to type 1 diabetes mellitus|Autonomic neuropathy due to type 1 diabetes mellitus
C1960678|T047|SY|712882000|SNOMEDCT_CORE|Autonomic neuropathy with type 1 diabetes mellitus|Autonomic neuropathy due to type 1 diabetes mellitus
C1960678|T047|SY|712882000|SNOMEDCT_CORE|Autonomic neuropathy with type I diabetes mellitus|Autonomic neuropathy due to type 1 diabetes mellitus
C1960678|T047|OAP|425442003|SNOMEDCT_CORE|Diabetic autonomic neuropathy associated with type 1 diabetes mellitus|Autonomic neuropathy due to type 1 diabetes mellitus
C1960678|T047|OAF|425442003|SNOMEDCT_CORE|Diabetic autonomic neuropathy associated with type 1 diabetes mellitus|Autonomic neuropathy due to type 1 diabetes mellitus
C1960678|T047|SY|712882000|SNOMEDCT_CORE|Diabetic autonomic neuropathy due to type 1 diabetes mellitus|Autonomic neuropathy due to type 1 diabetes mellitus
C1960678|T047|OF|712882000|SNOMEDCT_CORE|Diabetic autonomic neuropathy due to type 1 diabetes mellitus|Autonomic neuropathy due to type 1 diabetes mellitus
C1960678|T047|OAS|425442003|SNOMEDCT_CORE|Type 1 diabetic autonomic neuropathy|Autonomic neuropathy due to type 1 diabetes mellitus
C1960756|T033|PT|427589004|SNOMEDCT_CORE|Complicated grieving|Complicated grieving
C1960756|T033|FN|427589004|SNOMEDCT_CORE|Complicated grieving|Complicated grieving
C1960866|T047|PT|425771001|SNOMEDCT_CORE|Enlarging abdominal aortic aneurysm|Enlarging abdominal aortic aneurysm
C1960866|T047|FN|425771001|SNOMEDCT_CORE|Enlarging abdominal aortic aneurysm|Enlarging abdominal aortic aneurysm
C1960868|T046|PTGB|425957003|SNOMEDCT_CORE|Non-traumatic intracerebral ventricular haemorrhage|Non-traumatic intracerebral ventricular hemorrhage
C1960868|T046|PT|425957003|SNOMEDCT_CORE|Non-traumatic intracerebral ventricular hemorrhage|Non-traumatic intracerebral ventricular hemorrhage
C1960868|T046|FN|425957003|SNOMEDCT_CORE|Non-traumatic intracerebral ventricular hemorrhage|Non-traumatic intracerebral ventricular hemorrhage
C1960870|T047|IS|427419006|SNOMEDCT_CORE|Chronic migraine|Transformed migraine
C1960870|T047|SY|427419006|SNOMEDCT_CORE|Chronic migraine|Transformed migraine
C1960870|T047|PT|427419006|SNOMEDCT_CORE|Transformed migraine|Transformed migraine
C1960870|T047|FN|427419006|SNOMEDCT_CORE|Transformed migraine|Transformed migraine
C1960888|T184|PT|426702003|SNOMEDCT_CORE|Pain in female pelvis|Pain in female pelvis
C1960888|T184|FN|426702003|SNOMEDCT_CORE|Pain in female pelvis|Pain in female pelvis
C1961050|T047|PT|426263006|SNOMEDCT_CORE|Congestive heart failure due to left ventricular systolic dysfunction|Congestive heart failure due to left ventricular systolic dysfunction
C1961050|T047|FN|426263006|SNOMEDCT_CORE|Congestive heart failure due to left ventricular systolic dysfunction|Congestive heart failure due to left ventricular systolic dysfunction
C1961121|T019|SY|400159008|SNOMEDCT_CORE|Congenital vascular anomaly|Congenital vascular malformation
C1961121|T019|PT|400159008|SNOMEDCT_CORE|Congenital vascular malformation|Congenital vascular malformation
C1961121|T019|FN|400159008|SNOMEDCT_CORE|Congenital vascular malformation|Congenital vascular malformation
C1961121|T019|SY|400159008|SNOMEDCT_CORE|Vascular malformation|Congenital vascular malformation
C1961121|T019|SY|400159008|SNOMEDCT_CORE|VM - Vascular malformation|Congenital vascular malformation
C1962935|T033|SY|7293009|SNOMEDCT_CORE|Heavy for dates|Heavy-for-dates at birth regardless of gestation period
C1962935|T033|SY|7293009|SNOMEDCT_CORE|Heavy for gestation age infant|Heavy-for-dates at birth regardless of gestation period
C1962935|T033|PT|7293009|SNOMEDCT_CORE|Heavy-for-dates at birth regardless of gestation period|Heavy-for-dates at birth regardless of gestation period
C1962935|T033|FN|7293009|SNOMEDCT_CORE|Heavy-for-dates at birth regardless of gestation period|Heavy-for-dates at birth regardless of gestation period
C1962935|T033|OP|7293009|SNOMEDCT_CORE|Heavy-for-dates infant regardless of gestation period|Heavy-for-dates at birth regardless of gestation period
C1962935|T033|OF|7293009|SNOMEDCT_CORE|Heavy-for-dates infant regardless of gestation period|Heavy-for-dates at birth regardless of gestation period
C1962935|T033|SY|7293009|SNOMEDCT_CORE|Large-for-dates infant regardless of gestation period|Heavy-for-dates at birth regardless of gestation period
C1971019|T047|IS|89627008|SNOMEDCT_CORE|Na deficiency|Na deficiency
C1971019|T047|IS|89627008|SNOMEDCT_CORE|Na deficiency, NOS|Na deficiency
C1971021|T047|SY|43339004|SNOMEDCT_CORE|Potassium depletion|Potassium depletion
C1971624|T033|SY|79890006|SNOMEDCT_CORE|Anorexia|Loss of appetite
C1971624|T033|SY|79890006|SNOMEDCT_CORE|Anorexic|Loss of appetite
C1971624|T033|IS|79890006|SNOMEDCT_CORE|Lack of appetite|Loss of appetite
C1971624|T033|FN|79890006|SNOMEDCT_CORE|Loss of appetite|Loss of appetite
C1971624|T033|PT|79890006|SNOMEDCT_CORE|Loss of appetite|Loss of appetite
C1971624|T033|SY|79890006|SNOMEDCT_CORE|No appetite|Loss of appetite
C1971624|T033|SY|79890006|SNOMEDCT_CORE|Off food|Loss of appetite
C1971734|T047|PT|443820000|SNOMEDCT_CORE|Disorder of kidney and/or ureter|Disorder of kidney and/or ureter
C1971734|T047|FN|443820000|SNOMEDCT_CORE|Disorder of kidney and/or ureter|Disorder of kidney and/or ureter
C1971816|T019|IS|82525005|SNOMEDCT_CORE|Congenital fibrocystic kidney|Congenital fibrocystic kidney
C1971816|T047|IS|82525005|SNOMEDCT_CORE|Congenital fibrocystic kidney|Congenital fibrocystic kidney
C1971816|T019|IS|82525005|SNOMEDCT_CORE|Fibrocystic kidney|Congenital fibrocystic kidney
C1971816|T047|IS|82525005|SNOMEDCT_CORE|Fibrocystic kidney|Congenital fibrocystic kidney
C1996944|T047|SY|429447000|SNOMEDCT_CORE|Biceps tendon disorder|Disorder of tendon of biceps
C1996944|T047|SY|429447000|SNOMEDCT_CORE|Disorder of biceps tendon|Disorder of tendon of biceps
C1996944|T047|PT|429447000|SNOMEDCT_CORE|Disorder of tendon of biceps|Disorder of tendon of biceps
C1996944|T047|FN|429447000|SNOMEDCT_CORE|Disorder of tendon of biceps|Disorder of tendon of biceps
C1996954|T033|PT|427894009|SNOMEDCT_CORE|History of augmentation of breast|History of augmentation of breast
C1996954|T033|FN|427894009|SNOMEDCT_CORE|History of augmentation of breast|History of augmentation of breast
C1996954|T033|SY|427894009|SNOMEDCT_CORE|History of breast augmentation|History of augmentation of breast
C1996959|T047|SY|427788009|SNOMEDCT_CORE|Genital labial ulcer|Ulcer of genital labium
C1996959|T047|SY|427788009|SNOMEDCT_CORE|Labial ulceration|Ulcer of genital labium
C1996959|T047|PT|427788009|SNOMEDCT_CORE|Ulcer of genital labium|Ulcer of genital labium
C1996959|T047|FN|427788009|SNOMEDCT_CORE|Ulcer of genital labium|Ulcer of genital labium
C1996961|T184|PT|428171009|SNOMEDCT_CORE|Pain at rest due to peripheral vascular disease|Pain at rest due to peripheral vascular disease
C1996961|T184|FN|428171009|SNOMEDCT_CORE|Pain at rest due to peripheral vascular disease|Pain at rest due to peripheral vascular disease
C1996966|T033|PT|429479009|SNOMEDCT_CORE|History of radiation therapy|History of radiation therapy
C1996966|T033|FN|429479009|SNOMEDCT_CORE|History of radiation therapy|History of radiation therapy
C1996990|T033|PT|427858005|SNOMEDCT_CORE|Family history of malignant melanoma|Family history of malignant melanoma
C1996990|T033|FN|427858005|SNOMEDCT_CORE|Family history of malignant melanoma|Family history of malignant melanoma
C1997022|T033|SY|428283002|SNOMEDCT_CORE|History of colonic polyp|History of polyp of colon
C1997022|T033|FN|428283002|SNOMEDCT_CORE|History of polyp of colon|History of polyp of colon
C1997022|T033|PT|428283002|SNOMEDCT_CORE|History of polyp of colon|History of polyp of colon
C1997029|T033|SY|428071007|SNOMEDCT_CORE|History of coarctation of aorta repair|History of repair of coarctation of aorta
C1997029|T033|PT|428071007|SNOMEDCT_CORE|History of repair of coarctation of aorta|History of repair of coarctation of aorta
C1997029|T033|FN|428071007|SNOMEDCT_CORE|History of repair of coarctation of aorta|History of repair of coarctation of aorta
C1997034|T047|PT|427909005|SNOMEDCT_CORE|Chronic recurrent sinusitis|Chronic recurrent sinusitis
C1997034|T047|FN|427909005|SNOMEDCT_CORE|Chronic recurrent sinusitis|Chronic recurrent sinusitis
C1997037|T033|PTGB|428982002|SNOMEDCT_CORE|Dependence on haemodialysis due to end stage renal disease|Dependence on hemodialysis due to end stage renal disease
C1997037|T033|PT|428982002|SNOMEDCT_CORE|Dependence on hemodialysis due to end stage renal disease|Dependence on hemodialysis due to end stage renal disease
C1997037|T033|FN|428982002|SNOMEDCT_CORE|Dependence on hemodialysis due to end stage renal disease|Dependence on hemodialysis due to end stage renal disease
C1997091|T033|SY|429372004|SNOMEDCT_CORE|History of amputation of leg below knee|History of amputation of leg through tibia and fibula
C1997091|T033|PT|429372004|SNOMEDCT_CORE|History of amputation of leg through tibia and fibula|History of amputation of leg through tibia and fibula
C1997091|T033|FN|429372004|SNOMEDCT_CORE|History of amputation of leg through tibia and fibula|History of amputation of leg through tibia and fibula
C1997092|T047|PT|428163005|SNOMEDCT_CORE|Hypertensive left ventricular hypertrophy|Hypertensive left ventricular hypertrophy
C1997092|T047|FN|428163005|SNOMEDCT_CORE|Hypertensive left ventricular hypertrophy|Hypertensive left ventricular hypertrophy
C1997094|T033|PT|429487005|SNOMEDCT_CORE|Dependence on continuous positive airway pressure ventilation|Dependence on continuous positive airway pressure ventilation
C1997094|T033|FN|429487005|SNOMEDCT_CORE|Dependence on continuous positive airway pressure ventilation|Dependence on continuous positive airway pressure ventilation
C1997094|T033|SY|429487005|SNOMEDCT_CORE|Dependence on continuous positive airway pressure ventilation|Dependence on continuous positive airway pressure ventilation
C1997098|T033|PT|428882003|SNOMEDCT_CORE|History of cholecystectomy|History of cholecystectomy
C1997098|T033|FN|428882003|SNOMEDCT_CORE|History of cholecystectomy|History of cholecystectomy
C1997109|T046|IS|429673002|SNOMEDCT_CORE|Arteriosclerosis in coronary artery bypass graft|Arteriosclerosis of coronary artery bypass graft
C1997109|T046|OF|429673002|SNOMEDCT_CORE|Arteriosclerosis in coronary artery bypass graft|Arteriosclerosis of coronary artery bypass graft
C1997109|T046|PT|429673002|SNOMEDCT_CORE|Arteriosclerosis of coronary artery bypass graft|Arteriosclerosis of coronary artery bypass graft
C1997109|T046|FN|429673002|SNOMEDCT_CORE|Arteriosclerosis of coronary artery bypass graft|Arteriosclerosis of coronary artery bypass graft
C1997109|T046|SY|429673002|SNOMEDCT_CORE|Coronary arteriosclerosis of coronary artery bypass graft|Arteriosclerosis of coronary artery bypass graft
C1997146|T033|SY|428077006|SNOMEDCT_CORE|History of inguinal hernia surgery|History of repair of inguinal hernia
C1997146|T033|PT|428077006|SNOMEDCT_CORE|History of repair of inguinal hernia|History of repair of inguinal hernia
C1997146|T033|FN|428077006|SNOMEDCT_CORE|History of repair of inguinal hernia|History of repair of inguinal hernia
C1997157|T033|PT|428072000|SNOMEDCT_CORE|History of repair of musculotendinous cuff of shoulder|History of repair of musculotendinous cuff of shoulder
C1997157|T033|FN|428072000|SNOMEDCT_CORE|History of repair of musculotendinous cuff of shoulder|History of repair of musculotendinous cuff of shoulder
C1997157|T033|SY|428072000|SNOMEDCT_CORE|History of repair of rotator cuff|History of repair of musculotendinous cuff of shoulder
C1997165|T033|PT|428656009|SNOMEDCT_CORE|History of laser assisted in situ keratomileusis|History of laser assisted in situ keratomileusis
C1997165|T033|FN|428656009|SNOMEDCT_CORE|History of laser assisted in situ keratomileusis|History of laser assisted in situ keratomileusis
C1997165|T033|SY|428656009|SNOMEDCT_CORE|History of LASIK - laser assisted in situ keratomileusis|History of laser assisted in situ keratomileusis
C1997178|T033|SY|428835005|SNOMEDCT_CORE|History of amputation of great toe|History of amputation of hallux
C1997178|T033|PT|428835005|SNOMEDCT_CORE|History of amputation of hallux|History of amputation of hallux
C1997178|T033|FN|428835005|SNOMEDCT_CORE|History of amputation of hallux|History of amputation of hallux
C1997189|T033|SY|428848009|SNOMEDCT_CORE|History of carpal tunnel decompression|History of decompression of median nerve
C1997189|T033|PT|428848009|SNOMEDCT_CORE|History of decompression of median nerve|History of decompression of median nerve
C1997189|T033|FN|428848009|SNOMEDCT_CORE|History of decompression of median nerve|History of decompression of median nerve
C1997194|T046|PT|427793007|SNOMEDCT_CORE|Complication of urinary catheter|Complication of urinary catheter
C1997194|T046|FN|427793007|SNOMEDCT_CORE|Complication of urinary catheter|Complication of urinary catheter
C1997211|T047|SY|429350001|SNOMEDCT_CORE|Arthropathy of facet joint|Arthropathy of spinal facet joint
C1997211|T047|PT|429350001|SNOMEDCT_CORE|Arthropathy of spinal facet joint|Arthropathy of spinal facet joint
C1997211|T047|FN|429350001|SNOMEDCT_CORE|Arthropathy of spinal facet joint|Arthropathy of spinal facet joint
C1997258|T033|IS|428053000|SNOMEDCT_CORE|History of malignant basal cell neoplasm of of skin|History of malignant basal cell neoplasm of skin
C1997258|T033|OF|428053000|SNOMEDCT_CORE|History of malignant basal cell neoplasm of of skin|History of malignant basal cell neoplasm of skin
C1997258|T033|PT|428053000|SNOMEDCT_CORE|History of malignant basal cell neoplasm of skin|History of malignant basal cell neoplasm of skin
C1997258|T033|FN|428053000|SNOMEDCT_CORE|History of malignant basal cell neoplasm of skin|History of malignant basal cell neoplasm of skin
C1997258|T033|SY|428053000|SNOMEDCT_CORE|History of malignant basal cell tumor of skin|History of malignant basal cell neoplasm of skin
C1997258|T033|SYGB|428053000|SNOMEDCT_CORE|History of malignant basal cell tumour of skin|History of malignant basal cell neoplasm of skin
C1997282|T047|PT|427778008|SNOMEDCT_CORE|Incompetence of nasal valve|Incompetence of nasal valve
C1997282|T047|FN|427778008|SNOMEDCT_CORE|Incompetence of nasal valve|Incompetence of nasal valve
C1997282|T047|SY|427778008|SNOMEDCT_CORE|Nasal valve incompetence|Incompetence of nasal valve
C1997297|T033|PT|429254008|SNOMEDCT_CORE|History of malignant neoplasm of thyroid|History of malignant neoplasm of thyroid
C1997297|T033|FN|429254008|SNOMEDCT_CORE|History of malignant neoplasm of thyroid|History of malignant neoplasm of thyroid
C1997308|T033|PT|428079009|SNOMEDCT_CORE|History of transurethral prostatectomy|History of transurethral prostatectomy
C1997308|T033|FN|428079009|SNOMEDCT_CORE|History of transurethral prostatectomy|History of transurethral prostatectomy
C1997308|T033|SY|428079009|SNOMEDCT_CORE|History of transurethral resection of prostate|History of transurethral prostatectomy
C1997318|T047|PT|428173007|SNOMEDCT_CORE|Chronic hypoxemic respiratory failure|Chronic hypoxemic respiratory failure
C1997318|T047|FN|428173007|SNOMEDCT_CORE|Chronic hypoxemic respiratory failure|Chronic hypoxemic respiratory failure
C1997318|T047|SY|428173007|SNOMEDCT_CORE|Chronic type 1 respiratory failure|Chronic hypoxemic respiratory failure
C1997318|T047|SY|428173007|SNOMEDCT_CORE|Chronic type I respiratory failure|Chronic hypoxemic respiratory failure
C1997319|T033|PT|428912006|SNOMEDCT_CORE|History of placement of stent in anterior descending branch of left coronary artery|History of placement of stent in anterior descending branch of left coronary artery
C1997319|T033|FN|428912006|SNOMEDCT_CORE|History of placement of stent in anterior descending branch of left coronary artery|History of placement of stent in anterior descending branch of left coronary artery
C1997319|T033|SY|428912006|SNOMEDCT_CORE|History of stent placement in anterior descending branch of left coronary artery|History of placement of stent in anterior descending branch of left coronary artery
C1997347|T033|SY|429484003|SNOMEDCT_CORE|History of cancer of cervix|History of malignant neoplasm of cervix
C1997347|T033|PT|429484003|SNOMEDCT_CORE|History of malignant neoplasm of cervix|History of malignant neoplasm of cervix
C1997347|T033|FN|429484003|SNOMEDCT_CORE|History of malignant neoplasm of cervix|History of malignant neoplasm of cervix
C1997351|T047|PT|429589006|SNOMEDCT_CORE|Left ventricular cardiac dysfunction|Left ventricular cardiac dysfunction
C1997351|T047|FN|429589006|SNOMEDCT_CORE|Left ventricular cardiac dysfunction|Left ventricular cardiac dysfunction
C1997376|T047|SYGB|428383000|SNOMEDCT_CORE|Anaemia caused by medication|Anemia due to medication
C1997376|T047|PTGB|428383000|SNOMEDCT_CORE|Anaemia due to medication|Anemia due to medication
C1997376|T047|SY|428383000|SNOMEDCT_CORE|Anemia caused by medication|Anemia due to medication
C1997376|T047|FN|428383000|SNOMEDCT_CORE|Anemia caused by medication|Anemia due to medication
C1997376|T047|PT|428383000|SNOMEDCT_CORE|Anemia due to medication|Anemia due to medication
C1997376|T047|OF|428383000|SNOMEDCT_CORE|Anemia due to medication|Anemia due to medication
C1997376|T047|SYGB|428383000|SNOMEDCT_CORE|Drug induced anaemia|Anemia due to medication
C1997376|T047|SY|428383000|SNOMEDCT_CORE|Drug induced anemia|Anemia due to medication
C1997395|T033|SY|427749007|SNOMEDCT_CORE|History of knee surgery|History of operative procedure on knee
C1997395|T033|PT|427749007|SNOMEDCT_CORE|History of operative procedure on knee|History of operative procedure on knee
C1997395|T033|FN|427749007|SNOMEDCT_CORE|History of operative procedure on knee|History of operative procedure on knee
C1997419|T033|SY|428667005|SNOMEDCT_CORE|History of breast reduction|History of reduction of breast
C1997419|T033|PT|428667005|SNOMEDCT_CORE|History of reduction of breast|History of reduction of breast
C1997419|T033|FN|428667005|SNOMEDCT_CORE|History of reduction of breast|History of reduction of breast
C1997422|T033|PT|429016002|SNOMEDCT_CORE|History of medullary carcinoma of thyroid|History of medullary carcinoma of thyroid
C1997422|T033|FN|429016002|SNOMEDCT_CORE|History of medullary carcinoma of thyroid|History of medullary carcinoma of thyroid
C1997422|T033|SY|429016002|SNOMEDCT_CORE|History of medullary thyroid carcinoma|History of medullary carcinoma of thyroid
C1997428|T033|PT|428834009|SNOMEDCT_CORE|History of amputation of finger|History of amputation of finger
C1997428|T033|FN|428834009|SNOMEDCT_CORE|History of amputation of finger|History of amputation of finger
C1997520|T033|PT|428892006|SNOMEDCT_CORE|History of thyroidectomy|History of thyroidectomy
C1997520|T033|FN|428892006|SNOMEDCT_CORE|History of thyroidectomy|History of thyroidectomy
C1997535|T033|SY|428375006|SNOMEDCT_CORE|History of coronary artery disease with stent placement|History of placement of stent for coronary artery disease
C1997535|T033|PT|428375006|SNOMEDCT_CORE|History of placement of stent for coronary artery disease|History of placement of stent for coronary artery disease
C1997535|T033|FN|428375006|SNOMEDCT_CORE|History of placement of stent for coronary artery disease|History of placement of stent for coronary artery disease
C1997548|T033|PT|429255009|SNOMEDCT_CORE|History of papillary adenocarcinoma of thyroid|History of papillary adenocarcinoma of thyroid
C1997548|T033|FN|429255009|SNOMEDCT_CORE|History of papillary adenocarcinoma of thyroid|History of papillary adenocarcinoma of thyroid
C1997548|T033|SY|429255009|SNOMEDCT_CORE|History of papillary thyroid carcinoma|History of papillary adenocarcinoma of thyroid
C1997585|T047|PT|427921009|SNOMEDCT_CORE|Chronic ulcer of ankle|Chronic ulcer of ankle
C1997585|T047|FN|427921009|SNOMEDCT_CORE|Chronic ulcer of ankle|Chronic ulcer of ankle
C1997635|T033|FN|429696002|SNOMEDCT_CORE|Instability of femoropatellar joint|Patellar instability
C1997635|T033|SY|429696002|SNOMEDCT_CORE|Instability of femoropatellar joint|Patellar instability
C1997635|T033|SY|429696002|SNOMEDCT_CORE|Instability of patellofemoral joint|Patellar instability
C1997635|T033|PT|429696002|SNOMEDCT_CORE|Patellar instability|Patellar instability
C1997651|T047|IS|428007007|SNOMEDCT_CORE|Erectile dysfunction associated with type 2 diabetes mellitus|Erectile dysfunction due to type 2 diabetes mellitus
C1997651|T047|OF|428007007|SNOMEDCT_CORE|Erectile dysfunction associated with type 2 diabetes mellitus|Erectile dysfunction due to type 2 diabetes mellitus
C1997651|T047|OF|428007007|SNOMEDCT_CORE|Erectile dysfunction co-occurrent and due to type 2 diabetes mellitus|Erectile dysfunction due to type 2 diabetes mellitus
C1997651|T047|IS|428007007|SNOMEDCT_CORE|Erectile dysfunction co-occurrent and due to type 2 diabetes mellitus|Erectile dysfunction due to type 2 diabetes mellitus
C1997651|T047|PT|428007007|SNOMEDCT_CORE|Erectile dysfunction due to type 2 diabetes mellitus|Erectile dysfunction due to type 2 diabetes mellitus
C1997651|T047|FN|428007007|SNOMEDCT_CORE|Erectile dysfunction due to type 2 diabetes mellitus|Erectile dysfunction due to type 2 diabetes mellitus
C1997651|T047|SY|428007007|SNOMEDCT_CORE|Erectile dysfunction with type 2 diabetes mellitus|Erectile dysfunction due to type 2 diabetes mellitus
C1997686|T033|PT|429047008|SNOMEDCT_CORE|History of adenomatous polyp of colon|History of adenomatous polyp of colon
C1997686|T033|FN|429047008|SNOMEDCT_CORE|History of adenomatous polyp of colon|History of adenomatous polyp of colon
C1997701|T033|PT|428535004|SNOMEDCT_CORE|History of cataract extraction|History of cataract extraction
C1997701|T033|FN|428535004|SNOMEDCT_CORE|History of cataract extraction|History of cataract extraction
C1997711|T033|PT|428642007|SNOMEDCT_CORE|History of radical retropubic prostatectomy|History of radical retropubic prostatectomy
C1997711|T033|FN|428642007|SNOMEDCT_CORE|History of radical retropubic prostatectomy|History of radical retropubic prostatectomy
C1997752|T033|PT|428534000|SNOMEDCT_CORE|History of carotid endarterectomy|History of carotid endarterectomy
C1997752|T033|FN|428534000|SNOMEDCT_CORE|History of carotid endarterectomy|History of carotid endarterectomy
C1997795|T033|PT|427746000|SNOMEDCT_CORE|Mass of shoulder region|Mass of shoulder region
C1997795|T033|FN|427746000|SNOMEDCT_CORE|Mass of shoulder region|Mass of shoulder region
C1997820|T033|SY|429014004|SNOMEDCT_CORE|History of lymphoma|History of malignant lymphoma
C1997820|T033|PT|429014004|SNOMEDCT_CORE|History of malignant lymphoma|History of malignant lymphoma
C1997820|T033|FN|429014004|SNOMEDCT_CORE|History of malignant lymphoma|History of malignant lymphoma
C1997824|T033|SY|429410000|SNOMEDCT_CORE|History of cancer of esophagus|History of malignant neoplasm of esophagus
C1997824|T033|SYGB|429410000|SNOMEDCT_CORE|History of cancer of oesophagus|History of malignant neoplasm of esophagus
C1997824|T033|PT|429410000|SNOMEDCT_CORE|History of malignant neoplasm of esophagus|History of malignant neoplasm of esophagus
C1997824|T033|FN|429410000|SNOMEDCT_CORE|History of malignant neoplasm of esophagus|History of malignant neoplasm of esophagus
C1997824|T033|PTGB|429410000|SNOMEDCT_CORE|History of malignant neoplasm of oesophagus|History of malignant neoplasm of esophagus
C1997830|T033|PT|429290001|SNOMEDCT_CORE|History of radical hysterectomy|History of radical hysterectomy
C1997830|T033|FN|429290001|SNOMEDCT_CORE|History of radical hysterectomy|History of radical hysterectomy
C1997831|T033|SY|429164009|SNOMEDCT_CORE|History of decompressive lumbar laminectomy|History of excision of lamina of lumbar vertebra for decompression of spinal cord
C1997831|T033|PT|429164009|SNOMEDCT_CORE|History of excision of lamina of lumbar vertebra for decompression of spinal cord|History of excision of lamina of lumbar vertebra for decompression of spinal cord
C1997831|T033|FN|429164009|SNOMEDCT_CORE|History of excision of lamina of lumbar vertebra for decompression of spinal cord|History of excision of lamina of lumbar vertebra for decompression of spinal cord
C1997842|T033|PT|429046004|SNOMEDCT_CORE|History of sustained ventricular tachycardia|History of sustained ventricular tachycardia
C1997842|T033|FN|429046004|SNOMEDCT_CORE|History of sustained ventricular tachycardia|History of sustained ventricular tachycardia
C1997852|T033|PT|429280009|SNOMEDCT_CORE|History of amputation of foot|History of amputation of foot
C1997852|T033|FN|429280009|SNOMEDCT_CORE|History of amputation of foot|History of amputation of foot
C1997869|T033|PT|428540007|SNOMEDCT_CORE|History of mastectomy|History of mastectomy
C1997869|T033|FN|428540007|SNOMEDCT_CORE|History of mastectomy|History of mastectomy
C1997893|T047|PT|429192004|SNOMEDCT_CORE|Rheumatoid arthritis of foot|Rheumatoid arthritis of foot
C1997893|T047|FN|429192004|SNOMEDCT_CORE|Rheumatoid arthritis of foot|Rheumatoid arthritis of foot
C1997933|T033|SY|428941002|SNOMEDCT_CORE|History of cancer of uterine body|History of malignant neoplasm of uterine body
C1997933|T033|PT|428941002|SNOMEDCT_CORE|History of malignant neoplasm of uterine body|History of malignant neoplasm of uterine body
C1997933|T033|FN|428941002|SNOMEDCT_CORE|History of malignant neoplasm of uterine body|History of malignant neoplasm of uterine body
C1997946|T033|SY|428308007|SNOMEDCT_CORE|History of percutaneous transluminal angioplasty for coronary artery disease|History of percutaneous transluminal coronary angioplasty
C1997946|T033|PT|428308007|SNOMEDCT_CORE|History of percutaneous transluminal coronary angioplasty|History of percutaneous transluminal coronary angioplasty
C1997946|T033|FN|428308007|SNOMEDCT_CORE|History of percutaneous transluminal coronary angioplasty|History of percutaneous transluminal coronary angioplasty
C1997950|T033|SY|429090009|SNOMEDCT_CORE|History of cancer of ovary|History of malignant neoplasm of ovary
C1997950|T033|PT|429090009|SNOMEDCT_CORE|History of malignant neoplasm of ovary|History of malignant neoplasm of ovary
C1997950|T033|FN|429090009|SNOMEDCT_CORE|History of malignant neoplasm of ovary|History of malignant neoplasm of ovary
C1997954|T047|SY|428671008|SNOMEDCT_CORE|Arthropathy of lumbar facet|Arthropathy of lumbar facet joint
C1997954|T047|PT|428671008|SNOMEDCT_CORE|Arthropathy of lumbar facet joint|Arthropathy of lumbar facet joint
C1997954|T047|FN|428671008|SNOMEDCT_CORE|Arthropathy of lumbar facet joint|Arthropathy of lumbar facet joint
C1997972|T047|SY|427910000|SNOMEDCT_CORE|Diverticulitis of sigmoid|Diverticulitis of sigmoid colon
C1997972|T047|PT|427910000|SNOMEDCT_CORE|Diverticulitis of sigmoid colon|Diverticulitis of sigmoid colon
C1997972|T047|FN|427910000|SNOMEDCT_CORE|Diverticulitis of sigmoid colon|Diverticulitis of sigmoid colon
C1998033|T033|PT|429444007|SNOMEDCT_CORE|History of malignant neoplasm of ureter|History of malignant neoplasm of ureter
C1998033|T033|FN|429444007|SNOMEDCT_CORE|History of malignant neoplasm of ureter|History of malignant neoplasm of ureter
C1998045|T047|PT|427970008|SNOMEDCT_CORE|Subclinical hyperthyroidism|Subclinical hyperthyroidism
C1998045|T047|FN|427970008|SNOMEDCT_CORE|Subclinical hyperthyroidism|Subclinical hyperthyroidism
C1998051|T033|PT|429089000|SNOMEDCT_CORE|History of malignant neoplasm of endometrium|History of malignant neoplasm of endometrium
C1998051|T033|FN|429089000|SNOMEDCT_CORE|History of malignant neoplasm of endometrium|History of malignant neoplasm of endometrium
C1998103|T046|PT|429494008|SNOMEDCT_CORE|Postoperative seroma|Postoperative seroma
C1998103|T046|FN|429494008|SNOMEDCT_CORE|Postoperative seroma|Postoperative seroma
C1998121|T033|PT|427964002|SNOMEDCT_CORE|History of tympanostomy|History of tympanostomy
C1998121|T033|FN|427964002|SNOMEDCT_CORE|History of tympanostomy|History of tympanostomy
C1998127|T047|PT|429439000|SNOMEDCT_CORE|Complex cyst of uterine adnexa|Complex cyst of uterine adnexa
C1998127|T047|FN|429439000|SNOMEDCT_CORE|Complex cyst of uterine adnexa|Complex cyst of uterine adnexa
C1998127|T047|SY|429439000|SNOMEDCT_CORE|Complex uterine adnexal cyst|Complex cyst of uterine adnexa
C1998238|T033|SY|429409005|SNOMEDCT_CORE|History of cancer of the tongue|History of malignant neoplasm of tongue
C1998238|T033|PT|429409005|SNOMEDCT_CORE|History of malignant neoplasm of tongue|History of malignant neoplasm of tongue
C1998238|T033|FN|429409005|SNOMEDCT_CORE|History of malignant neoplasm of tongue|History of malignant neoplasm of tongue
C1998241|T033|PT|428251008|SNOMEDCT_CORE|History of appendectomy|History of appendectomy
C1998241|T033|FN|428251008|SNOMEDCT_CORE|History of appendectomy|History of appendectomy
C1998241|T033|PTGB|428251008|SNOMEDCT_CORE|History of appendicectomy|History of appendectomy
C1998255|T037|PT|428798001|SNOMEDCT_CORE|Closed fracture of tibial plateau|Closed fracture of tibial plateau
C1998255|T037|FN|428798001|SNOMEDCT_CORE|Closed fracture of tibial plateau|Closed fracture of tibial plateau
C1998257|T033|PT|428529004|SNOMEDCT_CORE|History of bilateral mastectomy|History of bilateral mastectomy
C1998257|T033|FN|428529004|SNOMEDCT_CORE|History of bilateral mastectomy|History of bilateral mastectomy
C1998265|T033|PT|429699009|SNOMEDCT_CORE|History of malignant neoplasm of colon|History of malignant neoplasm of colon
C1998265|T033|FN|429699009|SNOMEDCT_CORE|History of malignant neoplasm of colon|History of malignant neoplasm of colon
C1998267|T046|PT|428869006|SNOMEDCT_CORE|Mixed rhinitis|Mixed rhinitis
C1998267|T046|FN|428869006|SNOMEDCT_CORE|Mixed rhinitis|Mixed rhinitis
C1998270|T033|PT|427892008|SNOMEDCT_CORE|History of amputation of lesser toe|History of amputation of lesser toe
C1998270|T033|FN|427892008|SNOMEDCT_CORE|History of amputation of lesser toe|History of amputation of lesser toe
C1998270|T033|SY|427892008|SNOMEDCT_CORE|History of amputation of toe, other than great toe|History of amputation of lesser toe
C1998279|T033|SY|429285004|SNOMEDCT_CORE|History of anterior cruciate ligament tear reconstruction|History of reconstruction of anterior cruciate ligament tear
C1998279|T033|PT|429285004|SNOMEDCT_CORE|History of reconstruction of anterior cruciate ligament tear|History of reconstruction of anterior cruciate ligament tear
C1998279|T033|FN|429285004|SNOMEDCT_CORE|History of reconstruction of anterior cruciate ligament tear|History of reconstruction of anterior cruciate ligament tear
C1998298|T046|PT|427889009|SNOMEDCT_CORE|Hypertension associated with transplantation|Hypertension associated with transplantation
C1998298|T046|FN|427889009|SNOMEDCT_CORE|Hypertension associated with transplantation|Hypertension associated with transplantation
C1998329|T037|OAS|429564000|SNOMEDCT_CORE|Anaemia caused by chemotherapy|Anemia due to chemotherapy
C1998329|T037|OAP|429564000|SNOMEDCT_CORE|Anaemia due to chemotherapy|Anemia due to chemotherapy
C1998329|T037|OAS|429564000|SNOMEDCT_CORE|Anemia caused by chemotherapy|Anemia due to chemotherapy
C1998329|T037|OAF|429564000|SNOMEDCT_CORE|Anemia caused by chemotherapy|Anemia due to chemotherapy
C1998329|T037|OF|429564000|SNOMEDCT_CORE|Anemia due to chemotherapy|Anemia due to chemotherapy
C1998329|T037|OAP|429564000|SNOMEDCT_CORE|Anemia due to chemotherapy|Anemia due to chemotherapy
C1998334|T033|PT|428046009|SNOMEDCT_CORE|History of non-Hodgkins lymphoma|History of non-Hodgkins lymphoma
C1998334|T033|FN|428046009|SNOMEDCT_CORE|History of non-Hodgkins lymphoma|History of non-Hodgkins lymphoma
C1998380|T033|PTGB|428786006|SNOMEDCT_CORE|Localised superficial swelling of skin|Localized superficial swelling of skin
C1998380|T033|PT|428786006|SNOMEDCT_CORE|Localized superficial swelling of skin|Localized superficial swelling of skin
C1998380|T033|FN|428786006|SNOMEDCT_CORE|Localized superficial swelling of skin|Localized superficial swelling of skin
C1998384|T033|PT|429024007|SNOMEDCT_CORE|History of squamous cell carcinoma of skin|History of squamous cell carcinoma of skin
C1998384|T033|FN|429024007|SNOMEDCT_CORE|History of squamous cell carcinoma of skin|History of squamous cell carcinoma of skin
C1998388|T033|PT|429025008|SNOMEDCT_CORE|History of calculus of kidney|History of calculus of kidney
C1998388|T033|FN|429025008|SNOMEDCT_CORE|History of calculus of kidney|History of calculus of kidney
C1998388|T033|SY|429025008|SNOMEDCT_CORE|History of kidney stone|History of calculus of kidney
C1998388|T033|SY|429025008|SNOMEDCT_CORE|History of nephrolith|History of calculus of kidney
C1998388|T033|SY|429025008|SNOMEDCT_CORE|History of nephrolithiasis|History of calculus of kidney
C1998388|T033|SY|429025008|SNOMEDCT_CORE|History of renal calculus|History of calculus of kidney
C1998419|T033|PT|428078001|SNOMEDCT_CORE|History of total hysterectomy|History of total hysterectomy
C1998419|T033|FN|428078001|SNOMEDCT_CORE|History of total hysterectomy|History of total hysterectomy
C1998428|T048|SY|429672007|SNOMEDCT_CORE|Drug induced affective syndrome|Drug-induced mood disorder
C1998428|T048|SY|429672007|SNOMEDCT_CORE|Drug induced mood disorder|Drug-induced mood disorder
C1998428|T048|SY|429672007|SNOMEDCT_CORE|Drug-induced affective disorder|Drug-induced mood disorder
C1998428|T048|PT|429672007|SNOMEDCT_CORE|Drug-induced mood disorder|Drug-induced mood disorder
C1998428|T048|FN|429672007|SNOMEDCT_CORE|Drug-induced mood disorder|Drug-induced mood disorder
C1998449|T033|PT|428262008|SNOMEDCT_CORE|History of malignant neoplasm of prostate|History of malignant neoplasm of prostate
C1998449|T033|FN|428262008|SNOMEDCT_CORE|History of malignant neoplasm of prostate|History of malignant neoplasm of prostate
C1998978|T047|PT|129588001|SNOMEDCT_CORE|Adult failure to thrive syndrome|Adult failure to thrive syndrome
C1998978|T047|FN|129588001|SNOMEDCT_CORE|Adult failure to thrive syndrome|Adult failure to thrive syndrome
C1998986|T033|PT|54777007|SNOMEDCT_CORE|Deficient knowledge|Deficient knowledge
C1998986|T033|FN|54777007|SNOMEDCT_CORE|Deficient knowledge|Deficient knowledge
C1998986|T033|IS|54777007|SNOMEDCT_CORE|Deficient knowledge|Deficient knowledge
C1998986|T033|SY|54777007|SNOMEDCT_CORE|Knowledge deficit|Deficient knowledge
C1998986|T033|IS|54777007|SNOMEDCT_CORE|Knowledge deficit|Deficient knowledge
C1998986|T033|OF|54777007|SNOMEDCT_CORE|Knowledge deficit|Deficient knowledge
C2004435|T047|SYGB|82196007|SNOMEDCT_CORE|Intestinal ischaemia|Vascular insufficiency of intestine
C2004435|T047|SY|82196007|SNOMEDCT_CORE|Intestinal ischemia|Vascular insufficiency of intestine
C2004435|T047|SYGB|82196007|SNOMEDCT_CORE|Ischaemic bowel disease|Vascular insufficiency of intestine
C2004435|T047|IS|82196007|SNOMEDCT_CORE|Ischaemic bowel disease, NOS|Vascular insufficiency of intestine
C2004435|T047|SYGB|82196007|SNOMEDCT_CORE|Ischaemic disease of gut|Vascular insufficiency of intestine
C2004435|T047|SY|82196007|SNOMEDCT_CORE|Ischemic bowel disease|Vascular insufficiency of intestine
C2004435|T047|IS|82196007|SNOMEDCT_CORE|Ischemic bowel disease, NOS|Vascular insufficiency of intestine
C2004435|T047|SY|82196007|SNOMEDCT_CORE|Ischemic disease of gut|Vascular insufficiency of intestine
C2004435|T047|PT|82196007|SNOMEDCT_CORE|Vascular insufficiency of intestine|Vascular insufficiency of intestine
C2004435|T047|FN|82196007|SNOMEDCT_CORE|Vascular insufficiency of intestine|Vascular insufficiency of intestine
C2004435|T047|IS|82196007|SNOMEDCT_CORE|Vascular insufficiency of intestine, NOS|Vascular insufficiency of intestine
C2004435|T047|SY|82196007|SNOMEDCT_CORE|Vascular insufficiency of the intestine|Vascular insufficiency of intestine
C2004491|T046|PT|275322007|SNOMEDCT_CORE|Scar|Scar
C2004491|T046|FN|275322007|SNOMEDCT_CORE|Scar|Scar
C2004521|T047|MTH_SYGB|49472006|SNOMEDCT_CORE|Vitamin B<sub>12</sub> deficiency anaemia|Vitamin B>12< deficiency anemia
C2004521|T047|MTH_SY|49472006|SNOMEDCT_CORE|Vitamin B<sub>12</sub> deficiency anemia|Vitamin B>12< deficiency anemia
C2004521|T047|SYGB|49472006|SNOMEDCT_CORE|Vitamin B>12< deficiency anaemia|Vitamin B>12< deficiency anemia
C2004521|T047|SY|49472006|SNOMEDCT_CORE|Vitamin B>12< deficiency anemia|Vitamin B>12< deficiency anemia
C2004521|T047|MTH_SYGB|49472006|SNOMEDCT_CORE|Vitamin B12 deficiency anaemia|Vitamin B>12< deficiency anemia
C2004521|T047|MTH_SY|49472006|SNOMEDCT_CORE|Vitamin B12 deficiency anemia|Vitamin B>12< deficiency anemia
C2030468|T046|PT|442733008|SNOMEDCT_CORE|Hemiplegia as late effect of cerebrovascular accident|Hemiplegia as late effect of cerebrovascular accident
C2030468|T046|FN|442733008|SNOMEDCT_CORE|Hemiplegia as late effect of cerebrovascular accident|Hemiplegia as late effect of cerebrovascular accident
C2030469|T033|PT|442155009|SNOMEDCT_CORE|Hemiplegia of dominant side|Hemiplegia of dominant side
C2030469|T033|FN|442155009|SNOMEDCT_CORE|Hemiplegia of dominant side|Hemiplegia of dominant side
C2030470|T033|PT|441717007|SNOMEDCT_CORE|Hemiplegia of nondominant side|Hemiplegia of nondominant side
C2030470|T033|FN|441717007|SNOMEDCT_CORE|Hemiplegia of nondominant side|Hemiplegia of nondominant side
C2047520|T047|PTGB|267434003|SNOMEDCT_CORE|Mixed hyperlipidaemia|Mixed hyperlipidemia
C2047520|T047|FN|267434003|SNOMEDCT_CORE|Mixed hyperlipidemia|Mixed hyperlipidemia
C2047520|T047|PT|267434003|SNOMEDCT_CORE|Mixed hyperlipidemia|Mixed hyperlipidemia
C2047520|T047|SYGB|267434003|SNOMEDCT_CORE|Multiple-type hyperlipidaemia|Mixed hyperlipidemia
C2047520|T047|SY|267434003|SNOMEDCT_CORE|Multiple-type hyperlipidemia|Mixed hyperlipidemia
C2047937|T046|SY|74641007|SNOMEDCT_CORE|Ill defined condition|Ill-defined disease
C2047937|T046|SY|74641007|SNOMEDCT_CORE|Ill-defined condition|Ill-defined disease
C2047937|T046|PT|74641007|SNOMEDCT_CORE|Ill-defined disease|Ill-defined disease
C2047937|T046|FN|74641007|SNOMEDCT_CORE|Ill-defined disease|Ill-defined disease
C2063754|T047|PT|444548001|SNOMEDCT_CORE|Ulcerative pancolitis|Ulcerative pancolitis
C2063754|T047|FN|444548001|SNOMEDCT_CORE|Ulcerative pancolitis|Ulcerative pancolitis
C2063838|T020|PT|767679000|SNOMEDCT_CORE|Recurrent right inguinal hernia|Recurrent right inguinal hernia
C2063838|T020|FN|767679000|SNOMEDCT_CORE|Recurrent right inguinal hernia|Recurrent right inguinal hernia
C2076455|T037|PT|430984009|SNOMEDCT_CORE|Closed fracture of facial bone|Closed fracture of facial bone
C2076455|T037|FN|430984009|SNOMEDCT_CORE|Closed fracture of facial bone|Closed fracture of facial bone
C2081572|T033|PT|445122007|SNOMEDCT_CORE|Low lying placenta|Low lying placenta
C2081572|T033|FN|445122007|SNOMEDCT_CORE|Low lying placenta|Low lying placenta
C2088695|T037|PT|446314003|SNOMEDCT_CORE|Laceration of nail bed of finger|Laceration of nail bed of finger
C2088695|T037|FN|446314003|SNOMEDCT_CORE|Laceration of nail bed of finger|Laceration of nail bed of finger
C2089921|T037|PT|446896007|SNOMEDCT_CORE|Laceration of lower lip|Laceration of lower lip
C2089921|T037|FN|446896007|SNOMEDCT_CORE|Laceration of lower lip|Laceration of lower lip
C2108211|T037|OAP|262528003|SNOMEDCT_CORE|Bruise of head|Contusion of head
C2108211|T037|SY|735645009|SNOMEDCT_CORE|Bruise of head|Contusion of head
C2108211|T037|OAF|262528003|SNOMEDCT_CORE|Bruise of head|Contusion of head
C2108211|T037|PT|735645009|SNOMEDCT_CORE|Contusion of head|Contusion of head
C2108211|T037|FN|735645009|SNOMEDCT_CORE|Contusion of head|Contusion of head
C2108211|T037|OAS|262528003|SNOMEDCT_CORE|Superficial bruising of head|Contusion of head
C2141131|T047|PT|15971541000119105|SNOMEDCT_CORE|Left femoral hernia|Left femoral hernia
C2141131|T047|FN|15971541000119105|SNOMEDCT_CORE|Left femoral hernia|Left femoral hernia
C2145874|T037|PT|438505003|SNOMEDCT_CORE|Strain of trapezius muscle|Strain of trapezius muscle
C2145874|T037|FN|438505003|SNOMEDCT_CORE|Strain of trapezius muscle|Strain of trapezius muscle
C2171205|T047|OF|712883005|SNOMEDCT_CORE|Autonomic neuropathy co-occurrent and due to type 2 diabetes mellitus|Autonomic neuropathy due to type 2 diabetes mellitus
C2171205|T047|IS|712883005|SNOMEDCT_CORE|Autonomic neuropathy co-occurrent and due to type 2 diabetes mellitus|Autonomic neuropathy due to type 2 diabetes mellitus
C2171205|T047|PT|712883005|SNOMEDCT_CORE|Autonomic neuropathy due to type 2 diabetes mellitus|Autonomic neuropathy due to type 2 diabetes mellitus
C2171205|T047|FN|712883005|SNOMEDCT_CORE|Autonomic neuropathy due to type 2 diabetes mellitus|Autonomic neuropathy due to type 2 diabetes mellitus
C2171205|T047|SY|712883005|SNOMEDCT_CORE|Autonomic neuropathy with type 2 diabetes mellitus|Autonomic neuropathy due to type 2 diabetes mellitus
C2171205|T047|SY|712883005|SNOMEDCT_CORE|Autonomic neuropathy with type II diabetes mellitus|Autonomic neuropathy due to type 2 diabetes mellitus
C2171205|T047|OAF|423263001|SNOMEDCT_CORE|Diabetic autonomic neuropathy associated with type 2 diabetes mellitus|Autonomic neuropathy due to type 2 diabetes mellitus
C2171205|T047|OAP|423263001|SNOMEDCT_CORE|Diabetic autonomic neuropathy associated with type 2 diabetes mellitus|Autonomic neuropathy due to type 2 diabetes mellitus
C2171205|T047|OF|712883005|SNOMEDCT_CORE|Diabetic autonomic neuropathy due to type 2 diabetes mellitus|Autonomic neuropathy due to type 2 diabetes mellitus
C2171205|T047|SY|712883005|SNOMEDCT_CORE|Diabetic autonomic neuropathy due to type 2 diabetes mellitus|Autonomic neuropathy due to type 2 diabetes mellitus
C2174297|T033|PT|442098006|SNOMEDCT_CORE|Mass of foot|Mass of foot
C2174297|T033|FN|442098006|SNOMEDCT_CORE|Mass of foot|Mass of foot
C2201657|T020|PT|15971181000119105|SNOMEDCT_CORE|Right femoral hernia|Right femoral hernia
C2201657|T020|FN|15971181000119105|SNOMEDCT_CORE|Right femoral hernia|Right femoral hernia
C2229249|T033|SY|447071003|SNOMEDCT_CORE|Facial scar|Scar of face
C2229249|T033|PT|447071003|SNOMEDCT_CORE|Scar of face|Scar of face
C2229249|T033|FN|447071003|SNOMEDCT_CORE|Scar of face|Scar of face
C2239176|T191|SY|109841003|SNOMEDCT_CORE|HCC - Hepatocellular carcinoma|Liver cell carcinoma
C2239176|T191|SY|109841003|SNOMEDCT_CORE|Hepatocarcinoma|Liver cell carcinoma
C2239176|T191|SY|109841003|SNOMEDCT_CORE|Hepatocellular carcinoma|Liver cell carcinoma
C2239176|T191|IS|109841003|SNOMEDCT_CORE|Hepatocellular carcinoma|Liver cell carcinoma
C2239176|T191|SY|109841003|SNOMEDCT_CORE|LCC - Liver cell carcinoma|Liver cell carcinoma
C2239176|T191|SY|109841003|SNOMEDCT_CORE|Liver carcinoma|Liver cell carcinoma
C2239176|T191|PT|109841003|SNOMEDCT_CORE|Liver cell carcinoma|Liver cell carcinoma
C2239176|T191|IS|109841003|SNOMEDCT_CORE|Liver cell carcinoma|Liver cell carcinoma
C2239176|T191|FN|109841003|SNOMEDCT_CORE|Liver cell carcinoma|Liver cell carcinoma
C2239176|T191|SY|109841003|SNOMEDCT_CORE|Malignant hepatoma|Liver cell carcinoma
C2239176|T191|PT|187769009|SNOMEDCT_CORE|Primary carcinoma of liver|Liver cell carcinoma
C2239176|T191|FN|187769009|SNOMEDCT_CORE|Primary carcinoma of liver|Liver cell carcinoma
C2242769|T047|IS|24079001|SNOMEDCT_CORE|Besnier's prurigo|Besnier's prurigo
C2242769|T047|IS|24079001|SNOMEDCT_CORE|Prurigo of Besnier|Besnier's prurigo
C2242816|T047|SY|78868004|SNOMEDCT_CORE|Chronic MEE - Chronic middle ear effusion|Chronic secretory otitis media
C2242816|T047|SY|78868004|SNOMEDCT_CORE|Chronic middle ear effusion|Chronic secretory otitis media
C2242816|T047|SY|78868004|SNOMEDCT_CORE|Chronic non-suppurative otitis media with effusion|Chronic secretory otitis media
C2242816|T047|SY|78868004|SNOMEDCT_CORE|Chronic otitis media with effusion|Chronic secretory otitis media
C2242816|T047|SY|78868004|SNOMEDCT_CORE|Chronic secretory otitis media|Chronic secretory otitis media
C2242816|T047|SY|78868004|SNOMEDCT_CORE|Chronic secretory otitis media, mucoid|Chronic secretory otitis media
C2242816|T047|SY|78868004|SNOMEDCT_CORE|Chronic transudative otitis media|Chronic secretory otitis media
C2242996|T184|SY|62507009|SNOMEDCT_CORE|Tingling|Tingling sensation
C2242996|T184|IS|62507009|SNOMEDCT_CORE|Tingling sensation|Tingling sensation
C2243050|T033|OAP|161684005|SNOMEDCT_CORE|H/O: artificial opening|H/O: artificial opening
C2243050|T033|OF|161684005|SNOMEDCT_CORE|History of - artificial opening|H/O: artificial opening
C2243050|T033|IS|161684005|SNOMEDCT_CORE|History of - artificial opening|H/O: artificial opening
C2243050|T033|OAF|161684005|SNOMEDCT_CORE|History of artificial opening|H/O: artificial opening
C2243050|T033|OAS|161684005|SNOMEDCT_CORE|History of artificial opening|H/O: artificial opening
C2266788|T047|SY|254677004|SNOMEDCT_CORE|Follicular isthmus cyst|Trichilemmal cyst
C2266788|T047|SY|254677004|SNOMEDCT_CORE|Isthmus catagen cyst|Trichilemmal cyst
C2266788|T047|PT|254677004|SNOMEDCT_CORE|Trichilemmal cyst|Trichilemmal cyst
C2266788|T047|FN|254677004|SNOMEDCT_CORE|Trichilemmal cyst|Trichilemmal cyst
C2267227|T048|SY|78004001|SNOMEDCT_CORE|BN - Bulimia nervosa|Bulimia nervosa
C2267227|T048|PT|78004001|SNOMEDCT_CORE|Bulimia nervosa|Bulimia nervosa
C2267227|T048|FN|78004001|SNOMEDCT_CORE|Bulimia nervosa|Bulimia nervosa
C2314938|T033|SY|430954001|SNOMEDCT_CORE|Family history of cancer of genital system|Family history of malignant neoplasm of genital structure
C2314938|T033|PT|430954001|SNOMEDCT_CORE|Family history of malignant neoplasm of genital structure|Family history of malignant neoplasm of genital structure
C2314938|T033|FN|430954001|SNOMEDCT_CORE|Family history of malignant neoplasm of genital structure|Family history of malignant neoplasm of genital structure
C2315265|T047|PTGB|430348006|SNOMEDCT_CORE|Localised infection of skin AND/OR subcutaneous tissue|Localized infection of skin AND/OR subcutaneous tissue
C2315265|T047|PT|430348006|SNOMEDCT_CORE|Localized infection of skin AND/OR subcutaneous tissue|Localized infection of skin AND/OR subcutaneous tissue
C2315265|T047|FN|430348006|SNOMEDCT_CORE|Localized infection of skin AND/OR subcutaneous tissue|Localized infection of skin AND/OR subcutaneous tissue
C2315450|T047|PTGB|430347001|SNOMEDCT_CORE|Diverticulitis of caecum|Diverticulitis of cecum
C2315450|T047|PT|430347001|SNOMEDCT_CORE|Diverticulitis of cecum|Diverticulitis of cecum
C2315450|T047|FN|430347001|SNOMEDCT_CORE|Diverticulitis of cecum|Diverticulitis of cecum
C2315536|T047|PT|430725003|SNOMEDCT_CORE|Patellofemoral stress syndrome|Patellofemoral stress syndrome
C2315536|T047|FN|430725003|SNOMEDCT_CORE|Patellofemoral stress syndrome|Patellofemoral stress syndrome
C2315536|T047|SY|430725003|SNOMEDCT_CORE|Patellofemoral syndrome|Patellofemoral stress syndrome
C2315652|T047|PT|430959006|SNOMEDCT_CORE|Paralytic syndrome of dominant side as late effect of stroke|Paralytic syndrome of dominant side as late effect of stroke
C2315652|T047|FN|430959006|SNOMEDCT_CORE|Paralytic syndrome of dominant side as late effect of stroke|Paralytic syndrome of dominant side as late effect of stroke
C2315694|T047|PT|430985005|SNOMEDCT_CORE|Bilateral sensory hearing loss|Bilateral sensory hearing loss
C2315694|T047|FN|430985005|SNOMEDCT_CORE|Bilateral sensory hearing loss|Bilateral sensory hearing loss
C2315709|T047|PT|430031008|SNOMEDCT_CORE|Fetal hydronephrosis|Fetal hydronephrosis
C2315709|T047|FN|430031008|SNOMEDCT_CORE|Fetal hydronephrosis|Fetal hydronephrosis
C2315709|T047|SY|430031008|SNOMEDCT_CORE|Foetal hydronephrosis|Fetal hydronephrosis
C2315800|T047|PT|429975007|SNOMEDCT_CORE|Oral phase dysphagia|Oral phase dysphagia
C2315800|T047|FN|429975007|SNOMEDCT_CORE|Oral phase dysphagia|Oral phase dysphagia
C2315820|T019|PT|430166008|SNOMEDCT_CORE|Congenital anomaly of peripheral blood vessel|Congenital anomaly of peripheral blood vessel
C2315820|T019|FN|430166008|SNOMEDCT_CORE|Congenital anomaly of peripheral blood vessel|Congenital anomaly of peripheral blood vessel
C2315820|T019|SY|430166008|SNOMEDCT_CORE|Peripheral vascular congenital anomaly|Congenital anomaly of peripheral blood vessel
C2316134|T047|PT|431737008|SNOMEDCT_CORE|Acute lower urinary tract infection|Acute lower urinary tract infection
C2316134|T047|FN|431737008|SNOMEDCT_CORE|Acute lower urinary tract infection|Acute lower urinary tract infection
C2316134|T047|SY|431737008|SNOMEDCT_CORE|Lower urinary tract infection of sudden onset AND/OR short duration|Acute lower urinary tract infection
C2316203|T033|SY|429962007|SNOMEDCT_CORE|Family history of genetic disease|Family history of hereditary disease
C2316203|T033|PT|429962007|SNOMEDCT_CORE|Family history of hereditary disease|Family history of hereditary disease
C2316203|T033|FN|429962007|SNOMEDCT_CORE|Family history of hereditary disease|Family history of hereditary disease
C2316203|T033|SY|429962007|SNOMEDCT_CORE|Family history of heritable disorder|Family history of hereditary disease
C2316225|T047|PT|431237007|SNOMEDCT_CORE|Chronic headache disorder|Chronic headache disorder
C2316225|T047|FN|431237007|SNOMEDCT_CORE|Chronic headache disorder|Chronic headache disorder
C2316401|T047|PT|431855005|SNOMEDCT_CORE|Chronic kidney disease stage 1|Chronic kidney disease stage 1
C2316401|T047|FN|431855005|SNOMEDCT_CORE|Chronic kidney disease stage 1|Chronic kidney disease stage 1
C2316401|T047|SY|431855005|SNOMEDCT_CORE|CKD stage 1|Chronic kidney disease stage 1
C2316626|T047|SY|430474001|SNOMEDCT_CORE|Acquired adhesive capsulitis|Secondary adhesive capsulitis
C2316626|T047|PT|430474001|SNOMEDCT_CORE|Secondary adhesive capsulitis|Secondary adhesive capsulitis
C2316626|T047|FN|430474001|SNOMEDCT_CORE|Secondary adhesive capsulitis|Secondary adhesive capsulitis
C2316650|T033|SY|432615008|SNOMEDCT_CORE|Chronic facial pain|Chronic pain in face
C2316650|T033|PT|432615008|SNOMEDCT_CORE|Chronic pain in face|Chronic pain in face
C2316650|T033|FN|432615008|SNOMEDCT_CORE|Chronic pain in face|Chronic pain in face
C2316723|T047|PT|431481001|SNOMEDCT_CORE|Chronic pain due to injury|Chronic pain due to injury
C2316723|T047|FN|431481001|SNOMEDCT_CORE|Chronic pain due to injury|Chronic pain due to injury
C2316757|T033|SY|432352001|SNOMEDCT_CORE|Elevated creatine kinase level|Increased creatine kinase level
C2316757|T033|SY|432352001|SNOMEDCT_CORE|Increased CK level|Increased creatine kinase level
C2316757|T033|PT|432352001|SNOMEDCT_CORE|Increased creatine kinase level|Increased creatine kinase level
C2316757|T033|FN|432352001|SNOMEDCT_CORE|Increased creatine kinase level|Increased creatine kinase level
C2316757|T033|SY|432352001|SNOMEDCT_CORE|Increased phosphokinase|Increased creatine kinase level
C2316757|T033|SY|432352001|SNOMEDCT_CORE|Raised creatine kinase level|Increased creatine kinase level
C2316786|T047|PT|431856006|SNOMEDCT_CORE|Chronic kidney disease stage 2|Chronic kidney disease stage 2
C2316786|T047|FN|431856006|SNOMEDCT_CORE|Chronic kidney disease stage 2|Chronic kidney disease stage 2
C2316786|T047|SY|431856006|SNOMEDCT_CORE|CKD stage 2|Chronic kidney disease stage 2
C2316787|T047|PT|433144002|SNOMEDCT_CORE|Chronic kidney disease stage 3|Chronic kidney disease stage 3
C2316787|T047|FN|433144002|SNOMEDCT_CORE|Chronic kidney disease stage 3|Chronic kidney disease stage 3
C2316787|T047|SY|433144002|SNOMEDCT_CORE|CKD stage 3|Chronic kidney disease stage 3
C2316810|T047|PT|433146000|SNOMEDCT_CORE|Chronic kidney disease stage 5|Chronic kidney disease stage 5
C2316810|T047|FN|433146000|SNOMEDCT_CORE|Chronic kidney disease stage 5|Chronic kidney disease stage 5
C2316810|T047|SY|433146000|SNOMEDCT_CORE|CKD stage 5|Chronic kidney disease stage 5
C2316860|T046|SY|430947007|SNOMEDCT_CORE|Paralytic syndrome of non-dominant side as late effect of stroke|Paralytic syndrome of nondominant side as late effect of stroke
C2316860|T046|PT|430947007|SNOMEDCT_CORE|Paralytic syndrome of nondominant side as late effect of stroke|Paralytic syndrome of nondominant side as late effect of stroke
C2316860|T046|FN|430947007|SNOMEDCT_CORE|Paralytic syndrome of nondominant side as late effect of stroke|Paralytic syndrome of nondominant side as late effect of stroke
C2317045|T047|OAP|432083006|SNOMEDCT_CORE|Occlusive disease of artery of lower extremity|Occlusive disease of artery of lower extremity
C2317045|T047|OAF|432083006|SNOMEDCT_CORE|Occlusive disease of artery of lower extremity|Occlusive disease of artery of lower extremity
C2317404|T033|PT|429969003|SNOMEDCT_CORE|Family history of polyp of colon|Family history of polyp of colon
C2317404|T033|FN|429969003|SNOMEDCT_CORE|Family history of polyp of colon|Family history of polyp of colon
C2317445|T033|PT|429993008|SNOMEDCT_CORE|History of cerebrovascular accident without residual deficits|History of cerebrovascular accident without residual deficits
C2317445|T033|FN|429993008|SNOMEDCT_CORE|History of cerebrovascular accident without residual deficits|History of cerebrovascular accident without residual deficits
C2317473|T047|PT|431857002|SNOMEDCT_CORE|Chronic kidney disease stage 4|Chronic kidney disease stage 4
C2317473|T047|FN|431857002|SNOMEDCT_CORE|Chronic kidney disease stage 4|Chronic kidney disease stage 4
C2317473|T047|SY|431857002|SNOMEDCT_CORE|CKD stage 4|Chronic kidney disease stage 4
C2317516|T033|PT|431109006|SNOMEDCT_CORE|Carrier of vancomycin resistant enterococcus|Carrier of vancomycin resistant enterococcus
C2317516|T033|FN|431109006|SNOMEDCT_CORE|Carrier of vancomycin resistant enterococcus|Carrier of vancomycin resistant enterococcus
C2317516|T033|OF|431109006|SNOMEDCT_CORE|Carrier of vancomycin resistant enterococus|Carrier of vancomycin resistant enterococcus
C2317516|T033|IS|431109006|SNOMEDCT_CORE|Carrier of vancomycin resistant enterococus|Carrier of vancomycin resistant enterococcus
C2317549|T033|FN|432415000|SNOMEDCT_CORE|Methicillin resistant staphylococcus aureus carrier|Methicillin resistant staphylococcus aureus carrier
C2317549|T033|PT|432415000|SNOMEDCT_CORE|Methicillin resistant staphylococcus aureus carrier|Methicillin resistant staphylococcus aureus carrier
C2347126|T047|SY|239928004|SNOMEDCT_CORE|Microscopic polyangiitis|Microscopic polyarteritis nodosa
C2347126|T047|PT|239928004|SNOMEDCT_CORE|Microscopic polyarteritis nodosa|Microscopic polyarteritis nodosa
C2347126|T047|FN|239928004|SNOMEDCT_CORE|Microscopic polyarteritis nodosa|Microscopic polyarteritis nodosa
C2349195|T047|SY|54329005|SNOMEDCT_CORE|Acute anterior myocardial infarction|Acute myocardial infarction of anterior wall
C2349195|T047|PT|54329005|SNOMEDCT_CORE|Acute myocardial infarction of anterior wall|Acute myocardial infarction of anterior wall
C2349195|T047|FN|54329005|SNOMEDCT_CORE|Acute myocardial infarction of anterior wall|Acute myocardial infarction of anterior wall
C2349195|T047|IS|54329005|SNOMEDCT_CORE|Acute myocardial infarction of anterior wall, NOS|Acute myocardial infarction of anterior wall
C2349685|T033|PT|441099000|SNOMEDCT_CORE|Atypical squamous cells of undetermined significance on vaginal Papanicolaou smear|Atypical squamous cells of undetermined significance on vaginal Papanicolaou smear
C2349685|T033|FN|441099000|SNOMEDCT_CORE|Atypical squamous cells of undetermined significance on vaginal Papanicolaou smear|Atypical squamous cells of undetermined significance on vaginal Papanicolaou smear
C2350019|T191|FN|427359005|SNOMEDCT_CORE|Solitary nodule of lung|Solitary nodule of lung
C2350019|T191|PT|427359005|SNOMEDCT_CORE|Solitary nodule of lung|Solitary nodule of lung
C2350019|T191|SY|427359005|SNOMEDCT_CORE|Solitary pulmonary nodule|Solitary nodule of lung
C2350236|T047|OAP|45157009|SNOMEDCT_CORE|Idiopathic interstitial pneumonia|Idiopathic interstitial pneumonia
C2350242|T047|SY|8847002|SNOMEDCT_CORE|OA - Osteoarthritis of spine|OA - Osteoarthritis of the spine
C2350242|T047|SY|8847002|SNOMEDCT_CORE|OA - Osteoarthritis of the spine|OA - Osteoarthritis of the spine
C2350242|T047|SY|8847002|SNOMEDCT_CORE|Osteoarthritis of spine|OA - Osteoarthritis of the spine
C2355576|T191|SY|307651005|SNOMEDCT_CORE|Megakaryocytic myelosclerosis|Megakaryocytic myelosclerosis
C2363068|T037|PT|431307001|SNOMEDCT_CORE|Intentional poisoning by drug|Intentional poisoning by drug
C2363068|T037|OF|431307001|SNOMEDCT_CORE|Intentional poisoning by drug|Intentional poisoning by drug
C2363068|T037|FN|431307001|SNOMEDCT_CORE|Intentional poisoning caused by drug|Intentional poisoning by drug
C2363068|T037|SY|431307001|SNOMEDCT_CORE|Intentional poisoning caused by drug|Intentional poisoning by drug
C2364040|T033|PT|85623003|SNOMEDCT_CORE|Ineffective thermoregulation|Ineffective thermoregulation
C2364040|T033|FN|85623003|SNOMEDCT_CORE|Ineffective thermoregulation|Ineffective thermoregulation
C2364040|T033|SY|85623003|SNOMEDCT_CORE|Thermoregulation impairment|Ineffective thermoregulation
C2364164|T033|SY|1860003|SNOMEDCT_CORE|Disorder of fluid balance|Fluid volume disorder
C2364164|T033|PT|1860003|SNOMEDCT_CORE|Fluid volume disorder|Fluid volume disorder
C2364164|T033|FN|1860003|SNOMEDCT_CORE|Fluid volume disorder|Fluid volume disorder
C2364164|T033|IS|1860003|SNOMEDCT_CORE|Fluid volume disorder, NOS|Fluid volume disorder
C2364378|T033|PT|129831005|SNOMEDCT_CORE|Noncompliance with diagnostic testing|Noncompliance with diagnostic testing
C2364378|T033|FN|129831005|SNOMEDCT_CORE|Noncompliance with diagnostic testing|Noncompliance with diagnostic testing
C2364378|T033|SY|129831005|SNOMEDCT_CORE|Noncompliance: diagnostic testing|Noncompliance with diagnostic testing
C2364379|T033|PT|129832003|SNOMEDCT_CORE|Noncompliance with dietary regimen|Noncompliance with dietary regimen
C2364379|T033|FN|129832003|SNOMEDCT_CORE|Noncompliance with dietary regimen|Noncompliance with dietary regimen
C2364379|T033|SY|129832003|SNOMEDCT_CORE|Noncompliance with recommended nutrition plan|Noncompliance with dietary regimen
C2364379|T033|SY|129832003|SNOMEDCT_CORE|Noncompliance: dietary regimen|Noncompliance with dietary regimen
C2364379|T033|SY|129832003|SNOMEDCT_CORE|Noncompliance: recommended nutrition plan|Noncompliance with dietary regimen
C2367273|T047|PT|442073005|SNOMEDCT_CORE|Infection by methicillin sensitive Staphylococcus aureus|Infection by methicillin sensitive Staphylococcus aureus
C2367273|T047|SY|442073005|SNOMEDCT_CORE|Infection by methicillin susceptible Staphylococcus aureus|Infection by methicillin sensitive Staphylococcus aureus
C2367273|T047|OF|442073005|SNOMEDCT_CORE|Infection by methicillin susceptible Staphylococcus aureus|Infection by methicillin sensitive Staphylococcus aureus
C2367273|T047|SY|442073005|SNOMEDCT_CORE|Infection caused by methicillin sensitive Staphylococcus aureus|Infection by methicillin sensitive Staphylococcus aureus
C2367273|T047|SY|442073005|SNOMEDCT_CORE|Infection caused by methicillin susceptible Staphylococcus aureus|Infection by methicillin sensitive Staphylococcus aureus
C2367273|T047|FN|442073005|SNOMEDCT_CORE|Infection caused by methicillin susceptible Staphylococcus aureus|Infection by methicillin sensitive Staphylococcus aureus
C2584400|T033|PT|439590007|SNOMEDCT_CORE|Cardiovascular stress test abnormal|Cardiovascular stress test abnormal
C2584400|T033|FN|439590007|SNOMEDCT_CORE|Cardiovascular stress test abnormal|Cardiovascular stress test abnormal
C2584620|T047|SY|439698008|SNOMEDCT_CORE|Hereditary hypercoagulable disorder|Hereditary thrombophilia
C2584620|T047|PT|439698008|SNOMEDCT_CORE|Hereditary thrombophilia|Hereditary thrombophilia
C2584620|T047|FN|439698008|SNOMEDCT_CORE|Hereditary thrombophilia|Hereditary thrombophilia
C2584620|T047|SY|439698008|SNOMEDCT_CORE|Primary thrombophilia|Hereditary thrombophilia
C2584688|T033|IS|87860000|SNOMEDCT_CORE|Swollen testis|Testicular swelling
C2584688|T033|IS|87860000|SNOMEDCT_CORE|Testicular swelling|Testicular swelling
C2584688|T033|IS|87860000|SNOMEDCT_CORE|Testicular swelling, NOS|Testicular swelling
C2584784|T033|PT|441377000|SNOMEDCT_CORE|Thallium stress test abnormal|Thallium stress test abnormal
C2584784|T033|FN|441377000|SNOMEDCT_CORE|Thallium stress test abnormal|Thallium stress test abnormal
C2584975|T037|PT|438582003|SNOMEDCT_CORE|Acute injury of anterior cruciate ligament|Acute injury of anterior cruciate ligament
C2584975|T037|FN|438582003|SNOMEDCT_CORE|Acute injury of anterior cruciate ligament|Acute injury of anterior cruciate ligament
C2585886|T047|PT|439162001|SNOMEDCT_CORE|Embolism from thrombosis of vein of distal lower extremity|Embolism from thrombosis of vein of distal lower extremity
C2585886|T047|FN|439162001|SNOMEDCT_CORE|Embolism from thrombosis of vein of distal lower extremity|Embolism from thrombosis of vein of distal lower extremity
C2585886|T047|SY|439162001|SNOMEDCT_CORE|Embolism from venous thrombosis of lower leg|Embolism from thrombosis of vein of distal lower extremity
C2586056|T046|PT|440028005|SNOMEDCT_CORE|Permanent atrial fibrillation|Permanent atrial fibrillation
C2586056|T046|FN|440028005|SNOMEDCT_CORE|Permanent atrial fibrillation|Permanent atrial fibrillation
C2586286|T033|PT|438759003|SNOMEDCT_CORE|History of tonsillectomy|History of tonsillectomy
C2586286|T033|FN|438759003|SNOMEDCT_CORE|History of tonsillectomy|History of tonsillectomy
C2586308|T033|PT|439956007|SNOMEDCT_CORE|History of abnormal cervical Papanicolaou smear|History of abnormal cervical Papanicolaou smear
C2586308|T033|FN|439956007|SNOMEDCT_CORE|History of abnormal cervical Papanicolaou smear|History of abnormal cervical Papanicolaou smear
C2603353|T033|PT|440299000|SNOMEDCT_CORE|Mass of thoracic structure|Mass of thoracic structure
C2603353|T033|FN|440299000|SNOMEDCT_CORE|Mass of thoracic structure|Mass of thoracic structure
C2607914|T047|FN|61582004|SNOMEDCT_CORE|Allergic rhinitis|Allergic rhinitis
C2607914|T047|PT|61582004|SNOMEDCT_CORE|Allergic rhinitis|Allergic rhinitis
C2607914|T047|SY|61582004|SNOMEDCT_CORE|Allergic rhinitis due to allergen|Allergic rhinitis
C2607914|T047|IS|61582004|SNOMEDCT_CORE|Allergic rhinitis, NOS|Allergic rhinitis
C2607914|T047|SY|61582004|SNOMEDCT_CORE|AR - Allergic rhinitis|Allergic rhinitis
C2607914|T047|SY|61582004|SNOMEDCT_CORE|Atopic rhinitis|Allergic rhinitis
C2607928|T020|SY|399305009|SNOMEDCT_CORE|Non age related cataract|Nonsenile cataract
C2607928|T020|SY|399305009|SNOMEDCT_CORE|Non age-related cataract|Nonsenile cataract
C2607928|T020|PT|399305009|SNOMEDCT_CORE|Nonsenile cataract|Nonsenile cataract
C2607928|T020|FN|399305009|SNOMEDCT_CORE|Nonsenile cataract|Nonsenile cataract
C2711057|T047|SY|441794001|SNOMEDCT_CORE|Incomplete quadriplegia due to lesion at C5-C7 level|Incomplete tetraplegia due to lesion at C5-C7 level
C2711057|T047|FN|441794001|SNOMEDCT_CORE|Incomplete quadriplegia due to spinal cord lesion between fifth and seventh cervical vertebra|Incomplete tetraplegia due to lesion at C5-C7 level
C2711057|T047|SY|441794001|SNOMEDCT_CORE|Incomplete quadriplegia due to spinal cord lesion between fifth and seventh cervical vertebra|Incomplete tetraplegia due to lesion at C5-C7 level
C2711057|T047|PT|441794001|SNOMEDCT_CORE|Incomplete tetraplegia due to lesion at C5-C7 level|Incomplete tetraplegia due to lesion at C5-C7 level
C2711176|T047|SY|441705005|SNOMEDCT_CORE|Complete quadriplegia due to lesion at C1-C4 level|Complete tetraplegia due to lesion at C1-C4 level
C2711176|T047|FN|441705005|SNOMEDCT_CORE|Complete quadriplegia due to spinal cord lesion between first and fourth cervical vertebra|Complete tetraplegia due to lesion at C1-C4 level
C2711176|T047|SY|441705005|SNOMEDCT_CORE|Complete quadriplegia due to spinal cord lesion between first and fourth cervical vertebra|Complete tetraplegia due to lesion at C1-C4 level
C2711176|T047|PT|441705005|SNOMEDCT_CORE|Complete tetraplegia due to lesion at C1-C4 level|Complete tetraplegia due to lesion at C1-C4 level
C2711180|T047|SY|442438000|SNOMEDCT_CORE|Influenza caused by Influenza A virus|Influenza due to Influenza A virus
C2711180|T047|FN|442438000|SNOMEDCT_CORE|Influenza caused by Influenza A virus|Influenza due to Influenza A virus
C2711180|T047|PT|442438000|SNOMEDCT_CORE|Influenza due to Influenza A virus|Influenza due to Influenza A virus
C2711180|T047|OF|442438000|SNOMEDCT_CORE|Influenza due to Influenza A virus|Influenza due to Influenza A virus
C2711227|T047|PT|197321007|SNOMEDCT_CORE|Steatosis of liver|Steatosis of liver
C2711227|T047|FN|197321007|SNOMEDCT_CORE|Steatosis of liver|Steatosis of liver
C2711230|T047|SY|441688003|SNOMEDCT_CORE|Incomplete quadriplegia due to spinal cord lesion at C1-C4 level|Incomplete tetraplegia due to spinal cord lesion at C1-C4 level
C2711230|T047|FN|441688003|SNOMEDCT_CORE|Incomplete quadriplegia due to spinal cord lesion between first and fourth cervical vertebra|Incomplete tetraplegia due to spinal cord lesion at C1-C4 level
C2711230|T047|SY|441688003|SNOMEDCT_CORE|Incomplete quadriplegia due to spinal cord lesion between first and fourth cervical vertebra|Incomplete tetraplegia due to spinal cord lesion at C1-C4 level
C2711230|T047|PT|441688003|SNOMEDCT_CORE|Incomplete tetraplegia due to spinal cord lesion at C1-C4 level|Incomplete tetraplegia due to spinal cord lesion at C1-C4 level
C2711237|T047|SY|441574008|SNOMEDCT_CORE|Atherosclerosis artery|Atherosclerosis of artery
C2711237|T047|PT|441574008|SNOMEDCT_CORE|Atherosclerosis of artery|Atherosclerosis of artery
C2711237|T047|FN|441574008|SNOMEDCT_CORE|Atherosclerosis of artery|Atherosclerosis of artery
C2711273|T033|PT|441769002|SNOMEDCT_CORE|Cardiac defibrillator in situ|Cardiac defibrillator in situ
C2711273|T033|FN|441769002|SNOMEDCT_CORE|Cardiac defibrillator in situ|Cardiac defibrillator in situ
C2711374|T033|PT|441547007|SNOMEDCT_CORE|History of chronic urinary tract infection|History of chronic urinary tract infection
C2711374|T033|FN|441547007|SNOMEDCT_CORE|History of chronic urinary tract infection|History of chronic urinary tract infection
C2711399|T037|PT|442205007|SNOMEDCT_CORE|Stress fracture of tibia|Stress fracture of tibia
C2711399|T037|FN|442205007|SNOMEDCT_CORE|Stress fracture of tibia|Stress fracture of tibia
C2711434|T033|PTGB|442423001|SNOMEDCT_CORE|Single liveborn born in hospital by caesarean section|Single liveborn born in hospital by cesarean section
C2711434|T033|PT|442423001|SNOMEDCT_CORE|Single liveborn born in hospital by cesarean section|Single liveborn born in hospital by cesarean section
C2711434|T033|FN|442423001|SNOMEDCT_CORE|Single liveborn born in hospital by cesarean section|Single liveborn born in hospital by cesarean section
C2711438|T046|PT|442212003|SNOMEDCT_CORE|Residual cognitive deficit as late effect of cerebrovascular accident|Residual cognitive deficit as late effect of cerebrovascular accident
C2711438|T046|FN|442212003|SNOMEDCT_CORE|Residual cognitive deficit as late effect of cerebrovascular accident|Residual cognitive deficit as late effect of cerebrovascular accident
C2711438|T046|SY|442212003|SNOMEDCT_CORE|Residual cognitive deficit, late effect of stroke|Residual cognitive deficit as late effect of cerebrovascular accident
C2711480|T047|PT|441530006|SNOMEDCT_CORE|Chronic diastolic heart failure|Chronic diastolic heart failure
C2711480|T047|FN|441530006|SNOMEDCT_CORE|Chronic diastolic heart failure|Chronic diastolic heart failure
C2711482|T037|OAF|441702008|SNOMEDCT_CORE|Strain of muscle and/or tendon of wrist|Strain of muscle and/or tendon of wrist
C2711482|T037|OAP|441702008|SNOMEDCT_CORE|Strain of muscle and/or tendon of wrist|Strain of muscle and/or tendon of wrist
C2711482|T037|OAS|441702008|SNOMEDCT_CORE|Strain of wrist|Strain of muscle and/or tendon of wrist
C2711595|T033|PTGB|442365008|SNOMEDCT_CORE|Liveborn born in hospital by caesarean section|Liveborn born in hospital by cesarean section
C2711595|T033|PT|442365008|SNOMEDCT_CORE|Liveborn born in hospital by cesarean section|Liveborn born in hospital by cesarean section
C2711595|T033|FN|442365008|SNOMEDCT_CORE|Liveborn born in hospital by cesarean section|Liveborn born in hospital by cesarean section
C2711606|T047|SY|441980007|SNOMEDCT_CORE|Complete quadriplegia due to lesion at C5-C7 level|Complete tetraplegia due to lesion at C5-C7 level
C2711606|T047|FN|441980007|SNOMEDCT_CORE|Complete quadriplegia due to spinal cord lesion between fifth and seventh cervical vertebra|Complete tetraplegia due to lesion at C5-C7 level
C2711606|T047|SY|441980007|SNOMEDCT_CORE|Complete quadriplegia due to spinal cord lesion between fifth and seventh cervical vertebra|Complete tetraplegia due to lesion at C5-C7 level
C2711606|T047|PT|441980007|SNOMEDCT_CORE|Complete tetraplegia due to lesion at C5-C7 level|Complete tetraplegia due to lesion at C5-C7 level
C2711653|T047|PTGB|442481002|SNOMEDCT_CORE|Epilepsy characterised by intractable complex partial seizures|Epilepsy characterized by intractable complex partial seizures
C2711653|T047|PT|442481002|SNOMEDCT_CORE|Epilepsy characterized by intractable complex partial seizures|Epilepsy characterized by intractable complex partial seizures
C2711653|T047|FN|442481002|SNOMEDCT_CORE|Epilepsy characterized by intractable complex partial seizures|Epilepsy characterized by intractable complex partial seizures
C2711657|T033|PT|441667007|SNOMEDCT_CORE|Abnormal cervical Papanicolaou smear with positive human papillomavirus deoxyribonucleic acid test|Abnormal cervical Papanicolaou smear with positive human papillomavirus deoxyribonucleic acid test
C2711657|T033|SY|441667007|SNOMEDCT_CORE|Abnormal cervical Papanicolaou smear with positive human papillomavirus deoxyribonucleic acid test|Abnormal cervical Papanicolaou smear with positive human papillomavirus deoxyribonucleic acid test
C2711657|T033|FN|441667007|SNOMEDCT_CORE|Abnormal cervical Papanicolaou smear with positive human papillomavirus deoxyribonucleic acid test|Abnormal cervical Papanicolaou smear with positive human papillomavirus deoxyribonucleic acid test
C2711670|T048|SY|442351006|SNOMEDCT_CORE|Mental disorder caused by drug|Mental disorder due to drug
C2711670|T048|FN|442351006|SNOMEDCT_CORE|Mental disorder caused by drug|Mental disorder due to drug
C2711670|T048|PT|442351006|SNOMEDCT_CORE|Mental disorder due to drug|Mental disorder due to drug
C2711670|T048|OF|442351006|SNOMEDCT_CORE|Mental disorder due to drug|Mental disorder due to drug
C2711680|T033|PT|442234001|SNOMEDCT_CORE|Serum cholesterol borderline high|Serum cholesterol borderline high
C2711680|T033|FN|442234001|SNOMEDCT_CORE|Serum cholesterol borderline high|Serum cholesterol borderline high
C2711691|T033|PT|442646005|SNOMEDCT_CORE|Imaging of lung abnormal|Imaging of lung abnormal
C2711691|T033|FN|442646005|SNOMEDCT_CORE|Imaging of lung abnormal|Imaging of lung abnormal
C2711736|T047|PTGB|441678004|SNOMEDCT_CORE|Refractory generalised nonconvulsive epilepsy|Refractory generalized nonconvulsive epilepsy
C2711736|T047|PT|441678004|SNOMEDCT_CORE|Refractory generalized nonconvulsive epilepsy|Refractory generalized nonconvulsive epilepsy
C2711736|T047|FN|441678004|SNOMEDCT_CORE|Refractory generalized nonconvulsive epilepsy|Refractory generalized nonconvulsive epilepsy
C2711804|T033|SY|442342003|SNOMEDCT_CORE|Twin birth, in hospital, delivered by cesarean section|Twin liveborn born in hospital by cesarean section
C2711804|T033|PTGB|442342003|SNOMEDCT_CORE|Twin liveborn born in hospital by caesarean section|Twin liveborn born in hospital by cesarean section
C2711804|T033|PT|442342003|SNOMEDCT_CORE|Twin liveborn born in hospital by cesarean section|Twin liveborn born in hospital by cesarean section
C2711804|T033|FN|442342003|SNOMEDCT_CORE|Twin liveborn born in hospital by cesarean section|Twin liveborn born in hospital by cesarean section
C2711812|T033|PT|441924001|SNOMEDCT_CORE|Gestational age unknown|Gestational age unknown
C2711812|T033|FN|441924001|SNOMEDCT_CORE|Gestational age unknown|Gestational age unknown
C2711849|T046|PT|442024001|SNOMEDCT_CORE|Hemiplegia as late effect of cerebrovascular disease|Hemiplegia as late effect of cerebrovascular disease
C2711849|T046|FN|442024001|SNOMEDCT_CORE|Hemiplegia as late effect of cerebrovascular disease|Hemiplegia as late effect of cerebrovascular disease
C2711885|T047|PT|442439008|SNOMEDCT_CORE|Atherosclerosis of bypass graft of limb|Atherosclerosis of bypass graft of limb
C2711885|T047|FN|442439008|SNOMEDCT_CORE|Atherosclerosis of bypass graft of limb|Atherosclerosis of bypass graft of limb
C2711886|T047|PT|442693003|SNOMEDCT_CORE|Atherosclerosis of autologous vein bypass graft of limb|Atherosclerosis of autologous vein bypass graft of limb
C2711886|T047|FN|442693003|SNOMEDCT_CORE|Atherosclerosis of autologous vein bypass graft of limb|Atherosclerosis of autologous vein bypass graft of limb
C2711898|T033|SY|442327001|SNOMEDCT_CORE|Twin live born in hospital|Twin liveborn born in hospital
C2711898|T033|PT|442327001|SNOMEDCT_CORE|Twin liveborn born in hospital|Twin liveborn born in hospital
C2711898|T033|FN|442327001|SNOMEDCT_CORE|Twin liveborn born in hospital|Twin liveborn born in hospital
C2711966|T033|PT|442311008|SNOMEDCT_CORE|Liveborn born in hospital|Liveborn born in hospital
C2711966|T033|FN|442311008|SNOMEDCT_CORE|Liveborn born in hospital|Liveborn born in hospital
C2712998|T033|PT|441509002|SNOMEDCT_CORE|Cardiac pacemaker in situ|Cardiac pacemaker in situ
C2712998|T033|FN|441509002|SNOMEDCT_CORE|Cardiac pacemaker in situ|Cardiac pacemaker in situ
C2717899|T046|PT|128054009|SNOMEDCT_CORE|Deep venous thrombosis of upper extremity|Deep venous thrombosis of upper extremity
C2717899|T046|FN|128054009|SNOMEDCT_CORE|Deep venous thrombosis of upper extremity|Deep venous thrombosis of upper extremity
C2717961|T047|IS|78129009|SNOMEDCT_CORE|Thrombotic microangiopathy|Thrombotic microangiopathy
C2720436|T047|IS|73725006|SNOMEDCT_CORE|Fibrosis of pleura|Fibrosis of pleura
C2720436|T047|IS|73725006|SNOMEDCT_CORE|Pleural fibrosis|Fibrosis of pleura
C2724209|T047|IS|73725006|SNOMEDCT_CORE|Fibrothorax|Fibrothorax
C2732281|T047|IS|1679003|SNOMEDCT_CORE|Secondary osteoarthritis|Secondary osteoarthritis
C2732337|T046|PT|443760008|SNOMEDCT_CORE|Sleep hypoventilation|Sleep hypoventilation
C2732337|T046|FN|443760008|SNOMEDCT_CORE|Sleep hypoventilation|Sleep hypoventilation
C2732337|T046|SY|443760008|SNOMEDCT_CORE|Sleep related hypoventilation|Sleep hypoventilation
C2732402|T033|OAS|190371008|SNOMEDCT_CORE|Insulin-dependent diabetes mellitus - poor control|Type 1 diabetes mellitus uncontrolled
C2732402|T033|OAP|190371008|SNOMEDCT_CORE|Type 1 diabetes mellitus - poor control|Type 1 diabetes mellitus uncontrolled
C2732402|T033|PT|444073006|SNOMEDCT_CORE|Type 1 diabetes mellitus uncontrolled|Type 1 diabetes mellitus uncontrolled
C2732402|T033|OAF|190371008|SNOMEDCT_CORE|Type I diabetes mellitus - poor control|Type 1 diabetes mellitus uncontrolled
C2732402|T033|OAS|190371008|SNOMEDCT_CORE|Type I diabetes mellitus - poor control|Type 1 diabetes mellitus uncontrolled
C2732402|T033|SY|444073006|SNOMEDCT_CORE|Type I diabetes mellitus poorly controlled|Type 1 diabetes mellitus uncontrolled
C2732402|T033|SY|444073006|SNOMEDCT_CORE|Type I diabetes mellitus uncontrolled|Type 1 diabetes mellitus uncontrolled
C2732402|T033|FN|444073006|SNOMEDCT_CORE|Type I diabetes mellitus uncontrolled|Type 1 diabetes mellitus uncontrolled
C2732426|T037|PT|444491009|SNOMEDCT_CORE|Exposure to viral hepatitis|Exposure to viral hepatitis
C2732426|T037|FN|444491009|SNOMEDCT_CORE|Exposure to viral hepatitis|Exposure to viral hepatitis
C2732692|T033|PT|443460007|SNOMEDCT_CORE|Multigravida of advanced maternal age|Multigravida of advanced maternal age
C2732692|T033|FN|443460007|SNOMEDCT_CORE|Multigravida of advanced maternal age|Multigravida of advanced maternal age
C2732728|T033|IS|71781005|SNOMEDCT_CORE|Decreased body height|Short stature for age
C2732728|T033|IS|71781005|SNOMEDCT_CORE|Short for age|Short stature for age
C2732728|T033|IS|71781005|SNOMEDCT_CORE|Short stature for age|Short stature for age
C2732774|T191|IS|94022001|SNOMEDCT_CORE|Malignant neoplasm of skin of face|Malignant neoplasm of skin of face
C2732774|T191|IS|94022001|SNOMEDCT_CORE|Malignant neoplasm of skin of face, NOS|Malignant neoplasm of skin of face
C2732789|T037|PT|444507004|SNOMEDCT_CORE|Exposure to Mycobacterium tuberculosis|Exposure to Mycobacterium tuberculosis
C2732789|T037|FN|444507004|SNOMEDCT_CORE|Exposure to Mycobacterium tuberculosis|Exposure to Mycobacterium tuberculosis
C2732900|T033|PT|444412001|SNOMEDCT_CORE|Willing to be donor of liver|Willing to be donor of liver
C2732900|T033|FN|444412001|SNOMEDCT_CORE|Willing to be donor of liver|Willing to be donor of liver
C2732928|T037|PT|443786003|SNOMEDCT_CORE|Injury while engaged in sports activity|Injury while engaged in sports activity
C2732928|T037|FN|443786003|SNOMEDCT_CORE|Injury while engaged in sports activity|Injury while engaged in sports activity
C2732928|T037|PTGB|443786003|SNOMEDCT_CORE|Injury whilst engaged in sports activity|Injury while engaged in sports activity
C2732961|T037|FN|444107005|SNOMEDCT_CORE|Exposure to communicable disease|Exposure to communicable disease
C2732961|T037|PT|444107005|SNOMEDCT_CORE|Exposure to communicable disease|Exposure to communicable disease
C2733085|T046|PT|443165006|SNOMEDCT_CORE|Pathological fracture due to osteoporosis|Pathological fracture due to osteoporosis
C2733085|T046|FN|443165006|SNOMEDCT_CORE|Pathological fracture due to osteoporosis|Pathological fracture due to osteoporosis
C2733101|T037|PT|444486008|SNOMEDCT_CORE|Exposure to Hepatitis B virus|Exposure to Hepatitis B virus
C2733101|T037|FN|444486008|SNOMEDCT_CORE|Exposure to Hepatitis B virus|Exposure to Hepatitis B virus
C2733132|T037|PT|444387000|SNOMEDCT_CORE|Exposure to Bordetella pertussis|Exposure to Bordetella pertussis
C2733132|T037|FN|444387000|SNOMEDCT_CORE|Exposure to Bordetella pertussis|Exposure to Bordetella pertussis
C2733132|T037|SY|444387000|SNOMEDCT_CORE|Exposure to whooping cough|Exposure to Bordetella pertussis
C2733146|T033|SY|443694000|SNOMEDCT_CORE|Type 2 diabetes mellitus uncontrolled|Type II diabetes mellitus uncontrolled
C2733146|T033|SY|443694000|SNOMEDCT_CORE|Type II diabetes mellitus poorly controlled|Type II diabetes mellitus uncontrolled
C2733146|T033|PT|443694000|SNOMEDCT_CORE|Type II diabetes mellitus uncontrolled|Type II diabetes mellitus uncontrolled
C2733146|T033|FN|443694000|SNOMEDCT_CORE|Type II diabetes mellitus uncontrolled|Type II diabetes mellitus uncontrolled
C2733179|T046|PT|443762000|SNOMEDCT_CORE|Hypertrophic cardiomegaly|Hypertrophic cardiomegaly
C2733179|T046|FN|443762000|SNOMEDCT_CORE|Hypertrophic cardiomegaly|Hypertrophic cardiomegaly
C2733206|T047|PT|444003007|SNOMEDCT_CORE|Disorder of joint of shoulder region|Disorder of joint of shoulder region
C2733206|T047|FN|444003007|SNOMEDCT_CORE|Disorder of joint of shoulder region|Disorder of joint of shoulder region
C2733397|T047|IS|8186001|SNOMEDCT_CORE|Cor bovinum|Cor bovinum
C2733398|T191|PT|443496006|SNOMEDCT_CORE|Enchondroma of bone|Enchondroma of bone
C2733398|T191|FN|443496006|SNOMEDCT_CORE|Enchondroma of bone|Enchondroma of bone
C2733399|T191|PT|443495005|SNOMEDCT_CORE|Neoplasm of lymphoid system structure|Neoplasm of lymphoid system structure
C2733399|T191|FN|443495005|SNOMEDCT_CORE|Neoplasm of lymphoid system structure|Neoplasm of lymphoid system structure
C2733447|T047|SY|444197004|SNOMEDCT_CORE|Multiple system atrophy, Parkinson variant|Multiple system atrophy, Parkinson's variant
C2733447|T047|FN|444197004|SNOMEDCT_CORE|Multiple system atrophy, Parkinson variant|Multiple system atrophy, Parkinson's variant
C2733447|T047|PT|444197004|SNOMEDCT_CORE|Multiple system atrophy, Parkinson's variant|Multiple system atrophy, Parkinson's variant
C2748388|T046|PT|473023007|SNOMEDCT_CORE|Complication associated with device|Complication associated with device
C2748388|T046|FN|473023007|SNOMEDCT_CORE|Complication associated with device|Complication associated with device
C2830004|T048|SY|271782001|SNOMEDCT_CORE|Somnolence|Somnolence
C2854114|T191|SYGB|277571004|SNOMEDCT_CORE|Mature B-cell leukaemia Burkitt-type|Mature B-cell leukemia Burkitt-type
C2854114|T191|SY|277571004|SNOMEDCT_CORE|Mature B-cell leukemia Burkitt-type|Mature B-cell leukemia Burkitt-type
C2887088|T047|FN|448417001|SNOMEDCT_CORE|Sepsis caused by Staphylococcus aureus|Sepsis due to Staphylococcus aureus
C2887088|T047|SY|448417001|SNOMEDCT_CORE|Sepsis caused by Staphylococcus aureus|Sepsis due to Staphylococcus aureus
C2887088|T047|PT|448417001|SNOMEDCT_CORE|Sepsis due to Staphylococcus aureus|Sepsis due to Staphylococcus aureus
C2887088|T047|OF|448417001|SNOMEDCT_CORE|Sepsis due to Staphylococcus aureus|Sepsis due to Staphylococcus aureus
C2911574|T033|PT|444932008|SNOMEDCT_CORE|Dependence on ventilator|Dependence on ventilator
C2911574|T033|FN|444932008|SNOMEDCT_CORE|Dependence on ventilator|Dependence on ventilator
C2919021|T047|PT|199227004|SNOMEDCT_CORE|Diabetes mellitus during pregnancy - baby not yet delivered|Diabetes mellitus during pregnancy - baby not yet delivered
C2919021|T047|FN|199227004|SNOMEDCT_CORE|Diabetes mellitus during pregnancy - baby not yet delivered|Diabetes mellitus during pregnancy - baby not yet delivered
C2919140|T033|FN|75148009|SNOMEDCT_CORE|Employment problem|Employment problem
C2919140|T033|PT|75148009|SNOMEDCT_CORE|Employment problem|Employment problem
C2919160|T033|FN|445201008|SNOMEDCT_CORE|Carcinoembryonic antigen above reference range|High carcinoembryonic antigen level
C2919160|T033|SY|445201008|SNOMEDCT_CORE|Carcinoembryonic antigen above reference range|High carcinoembryonic antigen level
C2919160|T033|PT|445201008|SNOMEDCT_CORE|High carcinoembryonic antigen level|High carcinoembryonic antigen level
C2919177|T033|PT|444767004|SNOMEDCT_CORE|Fussy toddler|Fussy toddler
C2919177|T033|FN|444767004|SNOMEDCT_CORE|Fussy toddler|Fussy toddler
C2919178|T033|PT|445585003|SNOMEDCT_CORE|Livebirth born before admission to hospital|Livebirth born before admission to hospital
C2919178|T033|FN|445585003|SNOMEDCT_CORE|Livebirth born before admission to hospital|Livebirth born before admission to hospital
C2919187|T033|PT|445140006|SNOMEDCT_CORE|Periodic leg movements of sleep|Periodic leg movements of sleep
C2919187|T033|FN|445140006|SNOMEDCT_CORE|Periodic leg movements of sleep|Periodic leg movements of sleep
C2919204|T047|PT|445478004|SNOMEDCT_CORE|Degenerative joint disease of pelvis|Degenerative joint disease of pelvis
C2919204|T047|FN|445478004|SNOMEDCT_CORE|Degenerative joint disease of pelvis|Degenerative joint disease of pelvis
C2919204|T047|SY|445478004|SNOMEDCT_CORE|Osteoarthritis of pelvis|Degenerative joint disease of pelvis
C2919216|T033|PT|445179000|SNOMEDCT_CORE|Excessive self-criticism|Excessive self-criticism
C2919216|T033|FN|445179000|SNOMEDCT_CORE|Excessive self-criticism|Excessive self-criticism
C2919216|T033|OF|445179000|SNOMEDCT_CORE|Excessive selfcriticism|Excessive self-criticism
C2919216|T033|OP|445179000|SNOMEDCT_CORE|Excessive selfcriticism|Excessive self-criticism
C2919237|T047|PT|444769001|SNOMEDCT_CORE|Anovulatory amenorrhea|Anovulatory amenorrhea
C2919237|T047|FN|444769001|SNOMEDCT_CORE|Anovulatory amenorrhea|Anovulatory amenorrhea
C2919237|T047|PTGB|444769001|SNOMEDCT_CORE|Anovulatory amenorrhoea|Anovulatory amenorrhea
C2919296|T033|PT|445164007|SNOMEDCT_CORE|Clotting time above reference range|Clotting time above reference range
C2919296|T033|FN|445164007|SNOMEDCT_CORE|Clotting time above reference range|Clotting time above reference range
C2919331|T047|PT|444897001|SNOMEDCT_CORE|Hypoplasia of mandibular bone|Hypoplasia of mandibular bone
C2919331|T047|FN|444897001|SNOMEDCT_CORE|Hypoplasia of mandibular bone|Hypoplasia of mandibular bone
C2919376|T047|PT|445378003|SNOMEDCT_CORE|Acute exacerbation of bronchiectasis|Acute exacerbation of bronchiectasis
C2919376|T047|FN|445378003|SNOMEDCT_CORE|Acute exacerbation of bronchiectasis|Acute exacerbation of bronchiectasis
C2919377|T046|PT|444816006|SNOMEDCT_CORE|Embolism from thrombosis of vein of lower extremity|Embolism from thrombosis of vein of lower extremity
C2919377|T046|FN|444816006|SNOMEDCT_CORE|Embolism from thrombosis of vein of lower extremity|Embolism from thrombosis of vein of lower extremity
C2919395|T047|PT|444661007|SNOMEDCT_CORE|High risk pregnancy due to history of preterm labor|High risk pregnancy due to history of preterm labor
C2919395|T047|FN|444661007|SNOMEDCT_CORE|High risk pregnancy due to history of preterm labor|High risk pregnancy due to history of preterm labor
C2919395|T047|PTGB|444661007|SNOMEDCT_CORE|High risk pregnancy due to history of preterm labour|High risk pregnancy due to history of preterm labor
C2919404|T033|FN|445445006|SNOMEDCT_CORE|Low density lipoprotein cholesterol above reference range|Raised low density lipoprotein cholesterol
C2919404|T033|SY|445445006|SNOMEDCT_CORE|Low density lipoprotein cholesterol above reference range|Raised low density lipoprotein cholesterol
C2919404|T033|PT|445445006|SNOMEDCT_CORE|Raised low density lipoprotein cholesterol|Raised low density lipoprotein cholesterol
C2919431|T047|PT|444552001|SNOMEDCT_CORE|Hyperplasia of mandibular bone|Hyperplasia of mandibular bone
C2919431|T047|FN|444552001|SNOMEDCT_CORE|Hyperplasia of mandibular bone|Hyperplasia of mandibular bone
C2919460|T184|OAF|445422000|SNOMEDCT_CORE|Joint pain in ankle and foot|Joint pain in ankle and foot
C2919460|T184|OAP|445422000|SNOMEDCT_CORE|Joint pain in ankle and foot|Joint pain in ankle and foot
C2919545|T033|PT|444702007|SNOMEDCT_CORE|Irregular bowel habits|Irregular bowel habits
C2919545|T033|FN|444702007|SNOMEDCT_CORE|Irregular bowel habits|Irregular bowel habits
C2919575|T046|PT|444658006|SNOMEDCT_CORE|Nonsustained ventricular tachycardia|Nonsustained ventricular tachycardia
C2919575|T046|FN|444658006|SNOMEDCT_CORE|Nonsustained ventricular tachycardia|Nonsustained ventricular tachycardia
C2919576|T047|PT|445243001|SNOMEDCT_CORE|Left sided ulcerative colitis|Left sided ulcerative colitis
C2919576|T047|FN|445243001|SNOMEDCT_CORE|Left sided ulcerative colitis|Left sided ulcerative colitis
C2919577|T047|PT|444620007|SNOMEDCT_CORE|Male urinary stress incontinence|Male urinary stress incontinence
C2919577|T047|FN|444620007|SNOMEDCT_CORE|Male urinary stress incontinence|Male urinary stress incontinence
C2919578|T033|PT|445456006|SNOMEDCT_CORE|Mass of submandibular region|Mass of submandibular region
C2919578|T033|FN|445456006|SNOMEDCT_CORE|Mass of submandibular region|Mass of submandibular region
C2919586|T047|PT|444735002|SNOMEDCT_CORE|Instability of pelvic floor|Instability of pelvic floor
C2919586|T047|FN|444735002|SNOMEDCT_CORE|Instability of pelvic floor|Instability of pelvic floor
C2919587|T033|FN|444551008|SNOMEDCT_CORE|Antinuclear antibody above reference range|Raised antinuclear antibody
C2919587|T033|SY|444551008|SNOMEDCT_CORE|Antinuclear antibody above reference range|Raised antinuclear antibody
C2919587|T033|PT|444551008|SNOMEDCT_CORE|Raised antinuclear antibody|Raised antinuclear antibody
C2919588|T033|SY|445514005|SNOMEDCT_CORE|Helicobacter pylori antibody above reference range|Raised Helicobacter pylori antibody
C2919588|T033|FN|445514005|SNOMEDCT_CORE|Helicobacter pylori antibody above reference range|Raised Helicobacter pylori antibody
C2919588|T033|SY|445514005|SNOMEDCT_CORE|Helicobacter pylori antibody elevation|Raised Helicobacter pylori antibody
C2919588|T033|PT|445514005|SNOMEDCT_CORE|Raised Helicobacter pylori antibody|Raised Helicobacter pylori antibody
C2919618|T037|PT|444563003|SNOMEDCT_CORE|Exposure to Hepatitis C virus|Exposure to Hepatitis C virus
C2919618|T037|FN|444563003|SNOMEDCT_CORE|Exposure to Hepatitis C virus|Exposure to Hepatitis C virus
C2919631|T191|SY|444597005|SNOMEDCT_CORE|Extranodal marginal zone lymphoma of mucosa-associated lymphoid tissue of stomach|Mucosa-associated lymphoid tissue lymphoma of stomach
C2919631|T191|FN|444597005|SNOMEDCT_CORE|Extranodal marginal zone lymphoma of mucosa-associated lymphoid tissue of stomach|Mucosa-associated lymphoid tissue lymphoma of stomach
C2919631|T191|PT|444597005|SNOMEDCT_CORE|Mucosa-associated lymphoid tissue lymphoma of stomach|Mucosa-associated lymphoid tissue lymphoma of stomach
C2919754|T047|PT|445018004|SNOMEDCT_CORE|Spondylolysis of cervical spine|Spondylolysis of cervical spine
C2919754|T047|FN|445018004|SNOMEDCT_CORE|Spondylolysis of cervical spine|Spondylolysis of cervical spine
C2919828|T047|IS|64766004|SNOMEDCT_CORE|Chronic ulcerative colitis|Chronic ulcerative colitis
C2919828|T047|IS|64766004|SNOMEDCT_CORE|Chronic ulcerative colitis, NOS|Chronic ulcerative colitis
C2919898|T047|PT|445457002|SNOMEDCT_CORE|Hyperplasia of maxillary bone|Hyperplasia of maxillary bone
C2919898|T047|FN|445457002|SNOMEDCT_CORE|Hyperplasia of maxillary bone|Hyperplasia of maxillary bone
C2919899|T047|PT|444967008|SNOMEDCT_CORE|Hypoplasia of maxillary bone|Hypoplasia of maxillary bone
C2919899|T047|FN|444967008|SNOMEDCT_CORE|Hypoplasia of maxillary bone|Hypoplasia of maxillary bone
C2930812|T047|SYGB|58588007|SNOMEDCT_CORE|Generalised elastolysis|Generalized elastolysis
C2930812|T047|SY|58588007|SNOMEDCT_CORE|Generalized elastolysis|Generalized elastolysis
C2930898|T047|SY|59026006|SNOMEDCT_CORE|Benign essential blepharospasm|Benign essential blepharospasm
C2930898|T047|SY|59026006|SNOMEDCT_CORE|Essential blepharospasm|Benign essential blepharospasm
C2931404|T047|IS|58976002|SNOMEDCT_CORE|Albright hereditary osteodystrophy|Albright hereditary osteodystrophy
C2931404|T047|IS|58976002|SNOMEDCT_CORE|Albright hereditary osteodystrophy, NOS|Albright hereditary osteodystrophy, NOS
C2931822|T191|IS|187692001|SNOMEDCT_CORE|Nasopharyngeal carcinoma|Nasopharyngeal carcinoma
C2931838|T047|SY|15346004|SNOMEDCT_CORE|Familial HDL deficiency|Familial HDL deficiency
C2931914|T047|PT|34781003|SNOMEDCT_CORE|Vertebral artery syndrome|Vertebral artery syndrome
C2931914|T047|FN|34781003|SNOMEDCT_CORE|Vertebral artery syndrome|Vertebral artery syndrome
C2936664|T047|SYGB|23238000|SNOMEDCT_CORE|Acquired hypogammaglobulinaemia|Acquired hypogammaglobulinemia
C2936664|T047|SY|23238000|SNOMEDCT_CORE|Acquired hypogammaglobulinemia|Acquired hypogammaglobulinemia
C2936897|T047|SY|72275000|SNOMEDCT_CORE|Meyenburg-Altherr-Uehlinger syndrome|Meyenburg-Altherr-Uehlinger syndrome
C2937217|T047|PT|85225000|SNOMEDCT_CORE|Cyst of nasal sinus|Cyst of nasal sinus
C2937217|T047|FN|85225000|SNOMEDCT_CORE|Cyst of nasal sinus|Cyst of nasal sinus
C2937217|T047|IS|85225000|SNOMEDCT_CORE|Mucocele of nasal sinus|Cyst of nasal sinus
C2937217|T047|IS|85225000|SNOMEDCT_CORE|Mucous cyst of nasal sinus|Cyst of nasal sinus
C2937217|T047|SY|85225000|SNOMEDCT_CORE|Nasal sinus cyst|Cyst of nasal sinus
C2937260|T048|PT|191636007|SNOMEDCT_CORE|Mixed bipolar affective disorder|Mixed bipolar affective disorder
C2937260|T048|FN|191636007|SNOMEDCT_CORE|Mixed bipolar affective disorder|Mixed bipolar affective disorder
C2937358|T046|PTGB|274100004|SNOMEDCT_CORE|Cerebral haemorrhage|Cerebral hemorrhage
C2937358|T046|PT|274100004|SNOMEDCT_CORE|Cerebral hemorrhage|Cerebral hemorrhage
C2937358|T046|FN|274100004|SNOMEDCT_CORE|Cerebral hemorrhage|Cerebral hemorrhage
C2937358|T046|SYGB|274100004|SNOMEDCT_CORE|ICH - intracerebral haemorrhage|Cerebral hemorrhage
C2937358|T046|SY|274100004|SNOMEDCT_CORE|ICH - intracerebral hemorrhage|Cerebral hemorrhage
C2937358|T046|SYGB|274100004|SNOMEDCT_CORE|Intracerebral haemorrhage|Cerebral hemorrhage
C2937358|T046|IS|274100004|SNOMEDCT_CORE|Intracerebral haemorrhage|Cerebral hemorrhage
C2937358|T046|SY|274100004|SNOMEDCT_CORE|Intracerebral hemorrhage|Cerebral hemorrhage
C2937358|T046|IS|274100004|SNOMEDCT_CORE|Intracerebral hemorrhage|Cerebral hemorrhage
C2937421|T047|IS|266569009|SNOMEDCT_CORE|Hyperplasia of prostate|Hyperplasia of prostate
C2937421|T047|PT|433234005|SNOMEDCT_CORE|Hyperplasia of prostate|Hyperplasia of prostate
C2937421|T047|FN|433234005|SNOMEDCT_CORE|Hyperplasia of prostate|Hyperplasia of prostate
C2939419|T191|SY|128462008|SNOMEDCT_CORE|CA - Secondary cancer|Secondary malignant neoplastic disease
C2939419|T191|SY|128462008|SNOMEDCT_CORE|Metastases|Secondary malignant neoplastic disease
C2939419|T191|SY|128462008|SNOMEDCT_CORE|Metastatic cancer|Secondary malignant neoplastic disease
C2939419|T191|SY|128462008|SNOMEDCT_CORE|Metastatic malignant disease|Secondary malignant neoplastic disease
C2939419|T191|SY|128462008|SNOMEDCT_CORE|Metastatic neoplasm|Secondary malignant neoplastic disease
C2939419|T191|SY|128462008|SNOMEDCT_CORE|Secondaries|Secondary malignant neoplastic disease
C2939419|T191|SY|128462008|SNOMEDCT_CORE|Secondary cancer|Secondary malignant neoplastic disease
C2939419|T191|SY|128462008|SNOMEDCT_CORE|Secondary malignant deposit|Secondary malignant neoplastic disease
C2939419|T191|FN|128462008|SNOMEDCT_CORE|Secondary malignant neoplastic disease|Secondary malignant neoplastic disease
C2939419|T191|PT|128462008|SNOMEDCT_CORE|Secondary malignant neoplastic disease|Secondary malignant neoplastic disease
C2939419|T191|SY|128462008|SNOMEDCT_CORE|Secondary tumor|Secondary malignant neoplastic disease
C2939419|T191|SYGB|128462008|SNOMEDCT_CORE|Secondary tumour|Secondary malignant neoplastic disease
C2939419|T191|SY|128462008|SNOMEDCT_CORE|Tumor metastasis|Secondary malignant neoplastic disease
C2939419|T191|SYGB|128462008|SNOMEDCT_CORE|Tumour metastasis|Secondary malignant neoplastic disease
C2939447|T047|SY|367363000|SNOMEDCT_CORE|Right heart failure|Right ventricular failure
C2939447|T047|PT|367363000|SNOMEDCT_CORE|Right ventricular failure|Right ventricular failure
C2939447|T047|FN|367363000|SNOMEDCT_CORE|Right ventricular failure|Right ventricular failure
C2939465|T047|SY|124134002|SNOMEDCT_CORE|Deficiency of G-6PD|Deficiency of glucose-6-phosphate dehydrogenase
C2939465|T047|PT|124134002|SNOMEDCT_CORE|Deficiency of glucose-6-phosphate dehydrogenase|Deficiency of glucose-6-phosphate dehydrogenase
C2939465|T047|FN|124134002|SNOMEDCT_CORE|Deficiency of glucose-6-phosphate dehydrogenase|Deficiency of glucose-6-phosphate dehydrogenase
C2939465|T047|SY|124134002|SNOMEDCT_CORE|G6PD - Glucose-6-phosphate dehydrogenase deficiency|Deficiency of glucose-6-phosphate dehydrogenase
C2945552|T048|SY|31177006|SNOMEDCT_CORE|Attention deficit hyperactivity disorder combined|Attention deficit hyperactivity disorder, combined type
C2945552|T048|SY|31177006|SNOMEDCT_CORE|Attention deficit hyperactivity disorder combined type|Attention deficit hyperactivity disorder, combined type
C2945552|T048|PT|31177006|SNOMEDCT_CORE|Attention deficit hyperactivity disorder, combined type|Attention deficit hyperactivity disorder, combined type
C2945552|T048|FN|31177006|SNOMEDCT_CORE|Attention deficit hyperactivity disorder, combined type|Attention deficit hyperactivity disorder, combined type
C2945561|T047|IS|87688009|SNOMEDCT_CORE|Cholesterolosis of middle ear|Cholesterolosis of middle ear
C2945568|T047|PT|19399000|SNOMEDCT_CORE|Acute exudative otitis media|Acute exudative otitis media
C2945568|T047|FN|19399000|SNOMEDCT_CORE|Acute exudative otitis media|Acute exudative otitis media
C2945606|T047|FN|302690004|SNOMEDCT_CORE|Encopresis|Encopresis
C2945606|T047|PT|302690004|SNOMEDCT_CORE|Encopresis|Encopresis
C2945606|T047|OF|302690004|SNOMEDCT_CORE|Encopresis|Encopresis
C2959575|T033|PT|446653004|SNOMEDCT_CORE|Foreign body in lower limb|Foreign body in lower limb
C2959575|T033|FN|446653004|SNOMEDCT_CORE|Foreign body in lower limb|Foreign body in lower limb
C2959624|T047|SY|447043009|SNOMEDCT_CORE|Calculus of lower third of ureter|Ureteric stone of lower third of ureter
C2959624|T047|FN|447043009|SNOMEDCT_CORE|Calculus of lower third of ureter|Ureteric stone of lower third of ureter
C2959624|T047|PT|447043009|SNOMEDCT_CORE|Ureteric stone of lower third of ureter|Ureteric stone of lower third of ureter
C2959624|T047|SY|447043009|SNOMEDCT_CORE|Ureterolithiasis of lower third of ureter|Ureteric stone of lower third of ureter
C2959957|T037|PT|446859003|SNOMEDCT_CORE|Laceration of nail bed of toe|Laceration of nail bed of toe
C2959957|T037|FN|446859003|SNOMEDCT_CORE|Laceration of nail bed of toe|Laceration of nail bed of toe
C2979982|T046|OAP|399221001|SNOMEDCT_CORE|Bleeding from vagina|Vaginal bleeding
C2979982|T046|SY|289530006|SNOMEDCT_CORE|Bleeding from vagina|Vaginal bleeding
C2979982|T046|OAF|399221001|SNOMEDCT_CORE|Bleeding from vagina|Vaginal bleeding
C2979982|T046|FN|289530006|SNOMEDCT_CORE|Bleeding from vagina|Vaginal bleeding
C2979982|T046|OAS|399221001|SNOMEDCT_CORE|BVP - Vaginal bleeding|Vaginal bleeding
C2979982|T046|IS|289530006|SNOMEDCT_CORE|Finding of vaginal bleeding|Vaginal bleeding
C2979982|T046|OP|289530006|SNOMEDCT_CORE|Finding of vaginal bleeding|Vaginal bleeding
C2979982|T046|OAS|399221001|SNOMEDCT_CORE|Haemorrhage of vagina|Vaginal bleeding
C2979982|T046|OAS|399221001|SNOMEDCT_CORE|Hemorrhage of vagina|Vaginal bleeding
C2979982|T046|SY|289530006|SNOMEDCT_CORE|Observations of vaginal bleeding|Vaginal bleeding
C2979982|T046|OAS|399221001|SNOMEDCT_CORE|PV - Vaginal bleeding|Vaginal bleeding
C2979982|T046|OAS|399221001|SNOMEDCT_CORE|PV - Vaginal blood loss|Vaginal bleeding
C2979982|T046|OAS|399221001|SNOMEDCT_CORE|Vaginal bleeding|Vaginal bleeding
C2979982|T046|PT|289530006|SNOMEDCT_CORE|Vaginal bleeding|Vaginal bleeding
C2979982|T046|OAS|399221001|SNOMEDCT_CORE|Vaginal blood loss|Vaginal bleeding
C2980104|T047|IS|47382004|SNOMEDCT_CORE|Superficial mycosis|Superficial mycosis
C2980105|T047|IS|40603000|SNOMEDCT_CORE|Furunculosis of skin and subcutaneous tissue, NOS|Furunculosis of skin AND/OR subcutaneous tissue
C2980105|T047|OAP|40603000|SNOMEDCT_CORE|Furunculosis of skin AND/OR subcutaneous tissue|Furunculosis of skin AND/OR subcutaneous tissue
C2980105|T047|OAF|40603000|SNOMEDCT_CORE|Furunculosis of skin AND/OR subcutaneous tissue|Furunculosis of skin AND/OR subcutaneous tissue
C2980105|T047|OAS|40603000|SNOMEDCT_CORE|Recurring furuncles of skin|Furunculosis of skin AND/OR subcutaneous tissue
C2980105|T047|OAS|40603000|SNOMEDCT_CORE|Recurring skin boils|Furunculosis of skin AND/OR subcutaneous tissue
C2980106|T047|IS|55608001|SNOMEDCT_CORE|Prurigo mitis|Prurigo mitis
C2980107|T047|IS|55608001|SNOMEDCT_CORE|Hebra's prurigo|Hebra's prurigo
C2980107|T047|SY|55608001|SNOMEDCT_CORE|Urticaria papulosa of Hebra|Hebra's prurigo
C2981140|T047|SY|71111008|SNOMEDCT_CORE|Developmental glaucoma|Glaucoma of childhood
C2981140|T047|PT|71111008|SNOMEDCT_CORE|Glaucoma of childhood|Glaucoma of childhood
C2981140|T047|FN|71111008|SNOMEDCT_CORE|Glaucoma of childhood|Glaucoma of childhood
C2981140|T047|SY|71111008|SNOMEDCT_CORE|Infantile glaucoma|Glaucoma of childhood
C2981140|T047|SY|71111008|SNOMEDCT_CORE|Juvenile glaucoma|Glaucoma of childhood
C2981142|T047|SY|109996008|SNOMEDCT_CORE|Erythrodysplasia|Refractory anemia
C2981142|T047|SYGB|109996008|SNOMEDCT_CORE|Myelodysplastic syndrome: Refractory anaemia, without ringed sideroblasts, without excess blasts|Refractory anemia
C2981142|T047|FN|109996008|SNOMEDCT_CORE|Myelodysplastic syndrome: Refractory anemia, without ringed sideroblasts, without excess blasts|Refractory anemia
C2981142|T047|SY|109996008|SNOMEDCT_CORE|Myelodysplastic syndrome: Refractory anemia, without ringed sideroblasts, without excess blasts|Refractory anemia
C2981142|T047|SYGB|109996008|SNOMEDCT_CORE|RA - Refractory anaemia|Refractory anemia
C2981142|T047|SY|109996008|SNOMEDCT_CORE|RA - Refractory anemia|Refractory anemia
C2981142|T047|SYGB|109996008|SNOMEDCT_CORE|Refractory anaemia|Refractory anemia
C2981142|T047|PTGB|109996008|SNOMEDCT_CORE|Refractory anaemia|Refractory anemia
C2981142|T047|SY|109996008|SNOMEDCT_CORE|Refractory anemia|Refractory anemia
C2981142|T047|PT|109996008|SNOMEDCT_CORE|Refractory anemia|Refractory anemia
C3163829|T047|SY|449082003|SNOMEDCT_CORE|Sepsis caused by Gram negative bacteria|Sepsis due to Gram negative bacteria
C3163829|T047|FN|449082003|SNOMEDCT_CORE|Sepsis caused by Gram negative bacteria|Sepsis due to Gram negative bacteria
C3163829|T047|PT|449082003|SNOMEDCT_CORE|Sepsis due to Gram negative bacteria|Sepsis due to Gram negative bacteria
C3163829|T047|OF|449082003|SNOMEDCT_CORE|Sepsis due to Gram negative bacteria|Sepsis due to Gram negative bacteria
C3164125|T047|FN|448418006|SNOMEDCT_CORE|Sepsis caused by Streptococcus|Sepsis due to Streptococcus
C3164125|T047|SY|448418006|SNOMEDCT_CORE|Sepsis caused by Streptococcus|Sepsis due to Streptococcus
C3164125|T047|PT|448418006|SNOMEDCT_CORE|Sepsis due to Streptococcus|Sepsis due to Streptococcus
C3164125|T047|OF|448418006|SNOMEDCT_CORE|Sepsis due to Streptococcus|Sepsis due to Streptococcus
C3164130|T047|SY|449505005|SNOMEDCT_CORE|Sepsis caused by coagulase negative Staphylococcus|Sepsis due to coagulase negative Staphylococcus
C3164130|T047|FN|449505005|SNOMEDCT_CORE|Sepsis caused by coagulase negative Staphylococcus|Sepsis due to coagulase negative Staphylococcus
C3164130|T047|PT|449505005|SNOMEDCT_CORE|Sepsis due to coagulase negative Staphylococcus|Sepsis due to coagulase negative Staphylococcus
C3164130|T047|OF|449505005|SNOMEDCT_CORE|Sepsis due to coagulase negative Staphylococcus|Sepsis due to coagulase negative Staphylococcus
C3164254|T047|FN|447894003|SNOMEDCT_CORE|Sepsis caused by Staphylococcus|Sepsis due to Staphylococcus
C3164254|T047|SY|447894003|SNOMEDCT_CORE|Sepsis caused by Staphylococcus|Sepsis due to Staphylococcus
C3164254|T047|PT|447894003|SNOMEDCT_CORE|Sepsis due to Staphylococcus|Sepsis due to Staphylococcus
C3164254|T047|OF|447894003|SNOMEDCT_CORE|Sepsis due to Staphylococcus|Sepsis due to Staphylococcus
C3164258|T047|FN|447899008|SNOMEDCT_CORE|Sepsis caused by Escherichia coli|Sepsis due to Escherichia coli
C3164258|T047|SY|447899008|SNOMEDCT_CORE|Sepsis caused by Escherichia coli|Sepsis due to Escherichia coli
C3164258|T047|PT|447899008|SNOMEDCT_CORE|Sepsis due to Escherichia coli|Sepsis due to Escherichia coli
C3164258|T047|OF|447899008|SNOMEDCT_CORE|Sepsis due to Escherichia coli|Sepsis due to Escherichia coli
C3165209|T047|PT|448834003|SNOMEDCT_CORE|High density lipoprotein deficiency|High density lipoprotein deficiency
C3165209|T047|FN|448834003|SNOMEDCT_CORE|High density lipoprotein deficiency|High density lipoprotein deficiency
C3165526|T047|PT|217710005|SNOMEDCT_CORE|Congenital iodine deficiency syndrome|Congenital iodine deficiency syndrome
C3165526|T047|FN|217710005|SNOMEDCT_CORE|Congenital iodine deficiency syndrome|Congenital iodine deficiency syndrome
C3165526|T047|SY|217710005|SNOMEDCT_CORE|Fetal iodine deficiency syndrome|Congenital iodine deficiency syndrome
C3165526|T047|SYGB|217710005|SNOMEDCT_CORE|Foetal iodine deficiency syndrome|Congenital iodine deficiency syndrome
C3178801|T047|SY|230698000|SNOMEDCT_CORE|Lacunar stroke|Lacunar stroke
C3179349|T191|SY|420120006|SNOMEDCT_CORE|Gastrointestinal stromal sarcoma|Gastrointestinal stromal sarcoma
C3179349|T191|PT|128756002|SNOMEDCT_CORE|Gastrointestinal stromal sarcoma|Gastrointestinal stromal sarcoma
C3179349|T191|FN|128756002|SNOMEDCT_CORE|Gastrointestinal stromal sarcoma|Gastrointestinal stromal sarcoma
C3179349|T191|SY|128756002|SNOMEDCT_CORE|Gastrointestinal stromal tumor, malignant|Gastrointestinal stromal sarcoma
C3179349|T191|SYGB|128756002|SNOMEDCT_CORE|Gastrointestinal stromal tumour, malignant|Gastrointestinal stromal sarcoma
C3179349|T191|SY|128756002|SNOMEDCT_CORE|GIST, malignant|Gastrointestinal stromal sarcoma
C3203102|T047|PT|697898008|SNOMEDCT_CORE|Idiopathic pulmonary arterial hypertension|Idiopathic pulmonary arterial hypertension
C3203102|T047|FN|697898008|SNOMEDCT_CORE|Idiopathic pulmonary arterial hypertension|Idiopathic pulmonary arterial hypertension
C3203358|T046|PT|15993004|SNOMEDCT_CORE|Alveolar hypoventilation|Alveolar hypoventilation
C3203358|T046|FN|15993004|SNOMEDCT_CORE|Alveolar hypoventilation|Alveolar hypoventilation
C3241936|T046|IS|67782005|SNOMEDCT_CORE|Non-cardiogenic pulmonary edema|Non-cardiogenic pulmonary edema
C3241936|T046|IS|67782005|SNOMEDCT_CORE|Non-cardiogenic pulmonary oedema|Non-cardiogenic pulmonary edema
C3241944|T047|IS|6475002|SNOMEDCT_CORE|Alzheimer's disease with early onset|Primary degenerative dementia of the Alzheimer type, presenile onset, uncomplicated
C3241944|T047|IS|6475002|SNOMEDCT_CORE|Dementia in Alzheimer's disease - type 2|Primary degenerative dementia of the Alzheimer type, presenile onset, uncomplicated
C3241944|T047|IS|6475002|SNOMEDCT_CORE|Dementia in Alzheimer's disease with early onset|Primary degenerative dementia of the Alzheimer type, presenile onset, uncomplicated
C3241944|T047|SY|6475002|SNOMEDCT_CORE|Dementia of the Alzheimer's type, with early onset, uncomplicated|Primary degenerative dementia of the Alzheimer type, presenile onset, uncomplicated
C3241944|T047|IS|6475002|SNOMEDCT_CORE|Presenile dementia, Alzheimer's type|Primary degenerative dementia of the Alzheimer type, presenile onset, uncomplicated
C3241944|T047|PT|6475002|SNOMEDCT_CORE|Primary degenerative dementia of the Alzheimer type, presenile onset, uncomplicated|Primary degenerative dementia of the Alzheimer type, presenile onset, uncomplicated
C3241944|T047|FN|6475002|SNOMEDCT_CORE|Primary degenerative dementia of the Alzheimer type, presenile onset, uncomplicated|Primary degenerative dementia of the Alzheimer type, presenile onset, uncomplicated
C3241966|T033|SY|77176002|SNOMEDCT_CORE|Current smoker|Current smoker
C3249880|T033|SY|403194002|SNOMEDCT_CORE|Erythema solare|Solar erythema
C3249880|T033|SY|403194002|SNOMEDCT_CORE|Solar dermatitis|Solar erythema
C3249880|T033|PT|403194002|SNOMEDCT_CORE|Solar erythema|Solar erythema
C3249880|T033|FN|403194002|SNOMEDCT_CORE|Solar erythema|Solar erythema
C3249880|T033|SY|403194002|SNOMEDCT_CORE|Sunburn|Solar erythema
C3251816|T020|IS|74883004|SNOMEDCT_CORE|Aneurysm of thoracic aorta|Thoracic aortic aneurysm without rupture
C3251816|T020|IS|74883004|SNOMEDCT_CORE|Thoracic aortic aneurysm without mention of rupture|Thoracic aortic aneurysm without rupture
C3251816|T020|PT|74883004|SNOMEDCT_CORE|Thoracic aortic aneurysm without rupture|Thoracic aortic aneurysm without rupture
C3251816|T020|FN|74883004|SNOMEDCT_CORE|Thoracic aortic aneurysm without rupture|Thoracic aortic aneurysm without rupture
C3251825|T047|IS|238107002|SNOMEDCT_CORE|Dystrophy due to malnutrition|Dystrophy due to malnutrition
C3251829|T047|IS|58193001|SNOMEDCT_CORE|Congenital paraplegia|Congenital paraplegia
C3257803|T184|IS|193982009|SNOMEDCT_CORE|Watering eye|Watering eye
C3257803|T184|IS|193982009|SNOMEDCT_CORE|Watery eye|Watering eye
C3263722|T037|SY|417163006|SNOMEDCT_CORE|Injury|Traumatic AND/OR non-traumatic injury
C3263722|T037|PT|417163006|SNOMEDCT_CORE|Traumatic AND/OR non-traumatic injury|Traumatic AND/OR non-traumatic injury
C3263722|T037|FN|417163006|SNOMEDCT_CORE|Traumatic AND/OR non-traumatic injury|Traumatic AND/OR non-traumatic injury
C3263723|T037|IS|417746004|SNOMEDCT_CORE|Injury|Traumatic injury
C3263723|T037|SY|417746004|SNOMEDCT_CORE|Injury - disorder|Traumatic injury
C3263723|T037|SY|417746004|SNOMEDCT_CORE|Trauma|Traumatic injury
C3263723|T037|PT|417746004|SNOMEDCT_CORE|Traumatic injury|Traumatic injury
C3263723|T037|FN|417746004|SNOMEDCT_CORE|Traumatic injury|Traumatic injury
C3266014|T047|PT|449717009|SNOMEDCT_CORE|Cellulitis and abscess of upper limb|Cellulitis and abscess of upper limb
C3266014|T047|FN|449717009|SNOMEDCT_CORE|Cellulitis and abscess of upper limb|Cellulitis and abscess of upper limb
C3266180|T184|PT|449918009|SNOMEDCT_CORE|Cramp in lower leg|Cramp in lower leg
C3266180|T184|FN|449918009|SNOMEDCT_CORE|Cramp in lower leg|Cramp in lower leg
C3266685|T033|OP|591000119102|SNOMEDCT_CORE|Vaccine refused by patient|Vaccine refused by patient
C3266685|T033|PT|591000119102|SNOMEDCT_CORE|Vaccine refused by patient|Vaccine refused by patient
C3266685|T033|FN|591000119102|SNOMEDCT_CORE|Vaccine refused by patient|Vaccine refused by patient
C3463824|T191|SY|109995007|SNOMEDCT_CORE|MDS - Myelodysplastic syndrome|Myelodysplastic syndrome
C3463824|T191|SY|109995007|SNOMEDCT_CORE|Myelodysplastic syndrome|Myelodysplastic syndrome
C3463824|T191|PT|109995007|SNOMEDCT_CORE|Myelodysplastic syndrome|Myelodysplastic syndrome
C3463824|T191|FN|109995007|SNOMEDCT_CORE|Myelodysplastic syndrome|Myelodysplastic syndrome
C3472668|T037|PT|481000119104|SNOMEDCT_CORE|Strain of hamstring muscle|Strain of hamstring muscle
C3472668|T037|FN|481000119104|SNOMEDCT_CORE|Strain of hamstring muscle|Strain of hamstring muscle
C3472701|T047|PT|331000119106|SNOMEDCT_CORE|Tendinitis of elbow or forearm|Tendinitis of elbow or forearm
C3472701|T047|FN|331000119106|SNOMEDCT_CORE|Tendinitis of elbow or forearm|Tendinitis of elbow or forearm
C3489393|T047|IS|84089009|SNOMEDCT_CORE|Bergmann's syndrome|Hiatal hernia
C3489393|T047|SY|84089009|SNOMEDCT_CORE|Esophageal hiatal hernia|Hiatal hernia
C3489393|T047|SY|84089009|SNOMEDCT_CORE|Esophageal hiatus hernia|Hiatal hernia
C3489393|T047|SY|84089009|SNOMEDCT_CORE|HH - Hiatus hernia|Hiatal hernia
C3489393|T047|PT|84089009|SNOMEDCT_CORE|Hiatal hernia|Hiatal hernia
C3489393|T047|FN|84089009|SNOMEDCT_CORE|Hiatal hernia|Hiatal hernia
C3489393|T047|SY|84089009|SNOMEDCT_CORE|Hiatus hernia|Hiatal hernia
C3489393|T047|SYGB|84089009|SNOMEDCT_CORE|Oesophageal hiatal hernia|Hiatal hernia
C3489393|T047|SYGB|84089009|SNOMEDCT_CORE|Oesophageal hiatus hernia|Hiatal hernia
C3495439|T047|SY|266579006|SNOMEDCT_CORE|Inflammatory breast disease|Inflammatory disorder of breast
C3495439|T047|PT|266579006|SNOMEDCT_CORE|Inflammatory disorder of breast|Inflammatory disorder of breast
C3495439|T047|FN|266579006|SNOMEDCT_CORE|Inflammatory disorder of breast|Inflammatory disorder of breast
C3495439|T047|SY|266579006|SNOMEDCT_CORE|Mastitis|Inflammatory disorder of breast
C3495559|T047|SY|239796000|SNOMEDCT_CORE|JCA - Juvenile chronic arthritis|Juvenile chronic arthritis
C3495559|T047|SY|239796000|SNOMEDCT_CORE|Juvenile arthritis|Juvenile chronic arthritis
C3495559|T047|PT|239796000|SNOMEDCT_CORE|Juvenile chronic arthritis|Juvenile chronic arthritis
C3495559|T047|FN|239796000|SNOMEDCT_CORE|Juvenile chronic arthritis|Juvenile chronic arthritis
C3495801|T047|PT|195353004|SNOMEDCT_CORE|Granulomatosis with polyangiitis|Granulomatosis with polyangiitis
C3495801|T047|FN|195353004|SNOMEDCT_CORE|Granulomatosis with polyangiitis|Granulomatosis with polyangiitis
C3495801|T047|SYGB|195353004|SNOMEDCT_CORE|Necrotising respiratory granulomatosis|Granulomatosis with polyangiitis
C3495801|T047|SY|195353004|SNOMEDCT_CORE|Necrotizing respiratory granulomatosis|Granulomatosis with polyangiitis
C3495801|T047|IS|195353004|SNOMEDCT_CORE|Wegener granulomatosis|Granulomatosis with polyangiitis
C3495801|T047|IS|195353004|SNOMEDCT_CORE|Wegener's granulomatosis|Granulomatosis with polyangiitis
C3495801|T047|OF|195353004|SNOMEDCT_CORE|Wegener's granulomatosis|Granulomatosis with polyangiitis
C3532651|T033|PT|473158006|SNOMEDCT_CORE|History of live donor partial hepatectomy|History of live donor partial hepatectomy
C3532651|T033|FN|473158006|SNOMEDCT_CORE|History of live donor partial hepatectomy|History of live donor partial hepatectomy
C3532651|T033|SY|473158006|SNOMEDCT_CORE|History of liver donation|History of live donor partial hepatectomy
C3532651|T033|SY|473158006|SNOMEDCT_CORE|History of partial hepatectomy for liver donation|History of live donor partial hepatectomy
C3532655|T033|PT|473162000|SNOMEDCT_CORE|History of harvesting of stem cells for allotransplant|History of harvesting of stem cells for allotransplant
C3532655|T033|FN|473162000|SNOMEDCT_CORE|History of harvesting of stem cells for allotransplant|History of harvesting of stem cells for allotransplant
C3532655|T033|SY|473162000|SNOMEDCT_CORE|History of stem cell donation|History of harvesting of stem cells for allotransplant
C3536741|T019|SY|26146002|SNOMEDCT_CORE|Discordant ventriculoarterial connection with concordant atrioventricular connection|Discordant ventriculoarterial connection with concordant atrioventricular connection
C3537055|T046|IS|85224001|SNOMEDCT_CORE|Pilonidal abscess|Pilonidal cyst with abscess
C3537055|T046|PT|85224001|SNOMEDCT_CORE|Pilonidal cyst with abscess|Pilonidal cyst with abscess
C3537055|T046|FN|85224001|SNOMEDCT_CORE|Pilonidal cyst with abscess|Pilonidal cyst with abscess
C3537241|T033|IS|75148009|SNOMEDCT_CORE|Occupational problem|Occupational problem
C3539909|T033|PT|609328004|SNOMEDCT_CORE|Allergic disposition|Allergic disposition
C3539909|T033|OF|609328004|SNOMEDCT_CORE|Allergic disposition|Allergic disposition
C3539909|T033|FN|609328004|SNOMEDCT_CORE|Allergic disposition|Allergic disposition
C3539909|T033|SY|609328004|SNOMEDCT_CORE|Allergy|Allergic disposition
C3541213|T046|IS|12729009|SNOMEDCT_CORE|Delayed delivery after rupture of membranes|Prolonged rupture of membranes
C3541213|T046|IS|12729009|SNOMEDCT_CORE|Delayed delivery after spontaneous or unspecified rupture of membranes|Prolonged rupture of membranes
C3541213|T046|PT|12729009|SNOMEDCT_CORE|Prolonged rupture of membranes|Prolonged rupture of membranes
C3541213|T046|FN|12729009|SNOMEDCT_CORE|Prolonged rupture of membranes|Prolonged rupture of membranes
C3541213|T046|SY|12729009|SNOMEDCT_CORE|Rupture of amniotic sac 24 OR more hours before labor|Prolonged rupture of membranes
C3541213|T046|IS|12729009|SNOMEDCT_CORE|Rupture of amniotic sac 24 or more hours before labor|Prolonged rupture of membranes
C3541213|T046|SYGB|12729009|SNOMEDCT_CORE|Rupture of amniotic sac 24 OR more hours before labour|Prolonged rupture of membranes
C3541437|T033|OAP|268808004|SNOMEDCT_CORE|Fetal or neonatal effect of breech delivery and extraction|Fetal or neonatal effect of breech delivery and extraction
C3541437|T033|PT|4787007|SNOMEDCT_CORE|Fetal or neonatal effect of breech delivery and extraction|Fetal or neonatal effect of breech delivery and extraction
C3541437|T033|OAF|268808004|SNOMEDCT_CORE|Fetal or neonatal effect of breech delivery and extraction|Fetal or neonatal effect of breech delivery and extraction
C3541437|T033|FN|4787007|SNOMEDCT_CORE|Fetal or neonatal effect of breech delivery and extraction|Fetal or neonatal effect of breech delivery and extraction
C3541437|T033|OAP|268808004|SNOMEDCT_CORE|Foetal or neonatal effect of breech delivery and extraction|Fetal or neonatal effect of breech delivery and extraction
C3541437|T033|SY|4787007|SNOMEDCT_CORE|Foetal or neonatal effect of breech delivery and extraction|Fetal or neonatal effect of breech delivery and extraction
C3542501|T047|SY|40956001|SNOMEDCT_CORE|Acute idiopathic polyneuritis|Ascending paralysis
C3542501|T047|SY|40956001|SNOMEDCT_CORE|Acute idiopathic polyradiculoneuritis|Ascending paralysis
C3542501|T047|IS|40956001|SNOMEDCT_CORE|Acute infective polyneuritis|Ascending paralysis
C3542501|T047|IS|40956001|SNOMEDCT_CORE|Acute inflammatory demyelinating polyradiculoneuropathy|Ascending paralysis
C3542501|T047|SY|40956001|SNOMEDCT_CORE|Acute inflammatory neuropathy|Ascending paralysis
C3542501|T047|SY|40956001|SNOMEDCT_CORE|Acute post-infective radiculoneuropathy|Ascending paralysis
C3542501|T047|SY|40956001|SNOMEDCT_CORE|Ascending paralysis|Ascending paralysis
C3542501|T047|IS|40956001|SNOMEDCT_CORE|Infectious neuronitis|Ascending paralysis
C3542501|T047|IS|40956001|SNOMEDCT_CORE|PNS neuronitis|Ascending paralysis
C3543847|T047|IS|61628006|SNOMEDCT_CORE|Drug withdrawal syndrome in infant of dependent mother|Drug withdrawal syndrome in neonate of dependent mother
C3543847|T047|SY|609439002|SNOMEDCT_CORE|Drug withdrawal syndrome in infant of dependent mother|Drug withdrawal syndrome in neonate of dependent mother
C3543847|T047|FN|609439002|SNOMEDCT_CORE|Drug withdrawal syndrome in neonate of dependent mother|Drug withdrawal syndrome in neonate of dependent mother
C3543847|T047|PT|609439002|SNOMEDCT_CORE|Drug withdrawal syndrome in neonate of dependent mother|Drug withdrawal syndrome in neonate of dependent mother
C3650625|T046|PT|44991000119100|SNOMEDCT_CORE|Abnormal uterine bleeding|Abnormal uterine bleeding
C3650625|T046|FN|44991000119100|SNOMEDCT_CORE|Abnormal uterine bleeding|Abnormal uterine bleeding
C3650625|T046|SY|44991000119100|SNOMEDCT_CORE|Dysfunctional uterine bleeding|Abnormal uterine bleeding
C3662149|T046|PT|609496007|SNOMEDCT_CORE|Complication occurring during pregnancy|Complication occurring during pregnancy
C3662149|T046|FN|609496007|SNOMEDCT_CORE|Complication occurring during pregnancy|Complication occurring during pregnancy
C3662220|T047|OAP|18001006|SNOMEDCT_CORE|Fetal or neonatal effect of multiple pregnancy|Fetal or neonatal effect of multiple pregnancy
C3662220|T047|PT|206046007|SNOMEDCT_CORE|Fetal or neonatal effect of multiple pregnancy|Fetal or neonatal effect of multiple pregnancy
C3662220|T047|OAF|18001006|SNOMEDCT_CORE|Fetal or neonatal effect of multiple pregnancy|Fetal or neonatal effect of multiple pregnancy
C3662220|T047|FN|206046007|SNOMEDCT_CORE|Fetal or neonatal effect of multiple pregnancy|Fetal or neonatal effect of multiple pregnancy
C3662220|T047|SY|206046007|SNOMEDCT_CORE|Foetal or neonatal effect of multiple pregnancy|Fetal or neonatal effect of multiple pregnancy
C3662223|T046|SY|268798004|SNOMEDCT_CORE|Fetal effect of hydramnios|Fetal or neonatal effect of maternal polyhydramnios
C3662223|T046|PT|268798004|SNOMEDCT_CORE|Fetal or neonatal effect of maternal polyhydramnios|Fetal or neonatal effect of maternal polyhydramnios
C3662223|T046|FN|268798004|SNOMEDCT_CORE|Fetal or neonatal effect of maternal polyhydramnios|Fetal or neonatal effect of maternal polyhydramnios
C3662223|T046|SY|268798004|SNOMEDCT_CORE|Foetal effect of hydramnios|Fetal or neonatal effect of maternal polyhydramnios
C3662223|T046|SY|268798004|SNOMEDCT_CORE|Foetal or neonatal effect of maternal polyhydramnios|Fetal or neonatal effect of maternal polyhydramnios
C3662231|T033|PTGB|206065004|SNOMEDCT_CORE|Fetal or neonatal effect of placenta praevia|Fetal or neonatal effect of placenta previa
C3662231|T033|PT|206065004|SNOMEDCT_CORE|Fetal or neonatal effect of placenta previa|Fetal or neonatal effect of placenta previa
C3662231|T033|FN|206065004|SNOMEDCT_CORE|Fetal or neonatal effect of placenta previa|Fetal or neonatal effect of placenta previa
C3662231|T033|IS|206065004|SNOMEDCT_CORE|Fetus or neonate affected by placenta praevia|Fetal or neonatal effect of placenta previa
C3662231|T033|OP|206065004|SNOMEDCT_CORE|Fetus or neonate affected by placenta previa|Fetal or neonatal effect of placenta previa
C3662231|T033|OF|206065004|SNOMEDCT_CORE|Fetus or neonate affected by placenta previa|Fetal or neonatal effect of placenta previa
C3662231|T033|SYGB|206065004|SNOMEDCT_CORE|Foetal or neonatal effect of placenta praevia|Fetal or neonatal effect of placenta previa
C3662231|T033|OP|206065004|SNOMEDCT_CORE|Foetus or neonate affected by placenta praevia|Fetal or neonatal effect of placenta previa
C3662241|T033|OAF|73890002|SNOMEDCT_CORE|Fetal or neonatal effect of delivery by vacuum extractor|Fetal or neonatal effect of vacuum extraction delivery
C3662241|T033|OAP|73890002|SNOMEDCT_CORE|Fetal or neonatal effect of delivery by vacuum extractor|Fetal or neonatal effect of vacuum extraction delivery
C3662241|T033|SY|206122002|SNOMEDCT_CORE|Fetal or neonatal effect of delivery by vacuum extractor|Fetal or neonatal effect of vacuum extraction delivery
C3662241|T033|PT|206122002|SNOMEDCT_CORE|Fetal or neonatal effect of vacuum extraction delivery|Fetal or neonatal effect of vacuum extraction delivery
C3662241|T033|FN|206122002|SNOMEDCT_CORE|Fetal or neonatal effect of vacuum extraction delivery|Fetal or neonatal effect of vacuum extraction delivery
C3662241|T033|SY|206122002|SNOMEDCT_CORE|Foetal or neonatal effect of delivery by vacuum extractor|Fetal or neonatal effect of vacuum extraction delivery
C3662241|T033|SY|206122002|SNOMEDCT_CORE|Foetal or neonatal effect of vacuum extraction delivery|Fetal or neonatal effect of vacuum extraction delivery
C3662294|T190|PT|609380008|SNOMEDCT_CORE|Bowing deformity of lower limb|Bowing deformity of lower limb
C3662294|T190|FN|609380008|SNOMEDCT_CORE|Bowing deformity of lower limb|Bowing deformity of lower limb
C3665332|T047|IS|233873004|SNOMEDCT_CORE|Primary hypertrophic cardiomyopathy|Primary hypertrophic cardiomyopathy
C3665347|T033|IS|7973008|SNOMEDCT_CORE|Decreased vision|Visual impairment
C3665347|T033|SY|7973008|SNOMEDCT_CORE|Difficulty seeing|Visual impairment
C3665347|T033|IS|7973008|SNOMEDCT_CORE|Impaired vision|Visual impairment
C3665347|T033|SY|397540003|SNOMEDCT_CORE|Impaired vision|Visual impairment
C3665347|T033|SY|7973008|SNOMEDCT_CORE|Poor vision|Visual impairment
C3665347|T033|SY|7973008|SNOMEDCT_CORE|Reduced ability to see|Visual impairment
C3665347|T033|SY|7973008|SNOMEDCT_CORE|Sight impaired|Visual impairment
C3665347|T033|SY|397540003|SNOMEDCT_CORE|Visual difficulty|Visual impairment
C3665347|T033|IS|7973008|SNOMEDCT_CORE|Visual impairment|Visual impairment
C3665347|T033|PT|397540003|SNOMEDCT_CORE|Visual impairment|Visual impairment
C3665347|T033|FN|397540003|SNOMEDCT_CORE|Visual impairment|Visual impairment
C3665349|T047|SY|82598004|SNOMEDCT_CORE|Hypothyrotropic hypothyroidism|Secondary hypothyroidism
C3665349|T047|SY|82598004|SNOMEDCT_CORE|Pituitary hypothyroidism|Secondary hypothyroidism
C3665349|T047|PT|82598004|SNOMEDCT_CORE|Secondary hypothyroidism|Secondary hypothyroidism
C3665349|T047|FN|82598004|SNOMEDCT_CORE|Secondary hypothyroidism|Secondary hypothyroidism
C3665349|T047|SY|82598004|SNOMEDCT_CORE|TSH - Thyroid stimulating hormone deficiency|Secondary hypothyroidism
C3665349|T047|SY|82598004|SNOMEDCT_CORE|TSH deficiency|Secondary hypothyroidism
C3665357|T184|SY|9991008|SNOMEDCT_CORE|Intestinal colic|Intestinal colic
C3665386|T033|PT|7973008|SNOMEDCT_CORE|Abnormal vision|Abnormal vision
C3665386|T033|FN|7973008|SNOMEDCT_CORE|Abnormal vision|Abnormal vision
C3665386|T033|SY|7973008|SNOMEDCT_CORE|Partial sight|Abnormal vision
C3665386|T033|SY|7973008|SNOMEDCT_CORE|Problem seeing|Abnormal vision
C3665386|T033|SY|7973008|SNOMEDCT_CORE|Problem sight|Abnormal vision
C3665418|T047|OAP|276789009|SNOMEDCT_CORE|Labile hypertension|Labile hypertension
C3665418|T047|OAF|276789009|SNOMEDCT_CORE|Labile hypertension|Labile hypertension
C3665418|T047|OAS|276789009|SNOMEDCT_CORE|White coat hypertension|Labile hypertension
C3665419|T191|OAS|254937005|SNOMEDCT_CORE|Glioma of brain|Intracranial glioma
C3665419|T191|OAP|254937005|SNOMEDCT_CORE|Intracranial glioma|Intracranial glioma
C3665419|T191|OAF|254937005|SNOMEDCT_CORE|Intracranial glioma|Intracranial glioma
C3665447|T037|IS|10132008|SNOMEDCT_CORE|Burns of multiple specified sites|Burns of multiple specified sites
C3665497|T048|SY|66214007|SNOMEDCT_CORE|Nondependent abuse of drugs|Nondependent abuse of drugs
C3665593|T191|PTGB|400010006|SNOMEDCT_CORE|Melanocytic naevus of skin|Melanocytic nevus of skin
C3665593|T191|PT|400010006|SNOMEDCT_CORE|Melanocytic nevus of skin|Melanocytic nevus of skin
C3665593|T191|FN|400010006|SNOMEDCT_CORE|Melanocytic nevus of skin|Melanocytic nevus of skin
C3665593|T191|SY|400010006|SNOMEDCT_CORE|Mole of skin|Melanocytic nevus of skin
C3665593|T191|SYGB|400010006|SNOMEDCT_CORE|Pigmented naevus of skin|Melanocytic nevus of skin
C3665593|T191|SY|400010006|SNOMEDCT_CORE|Pigmented nevus of skin|Melanocytic nevus of skin
C3665595|T047|SY|57019003|SNOMEDCT_CORE|Mosaic wart|Mosaic wart
C3665596|T191|SY|57019003|SNOMEDCT_CORE|Wart|Wart
C3665608|T046|PTGB|396544001|SNOMEDCT_CORE|Caesarean wound disruption|Cesarean wound disruption
C3665608|T046|PT|396544001|SNOMEDCT_CORE|Cesarean wound disruption|Cesarean wound disruption
C3665608|T046|FN|396544001|SNOMEDCT_CORE|Cesarean wound disruption|Cesarean wound disruption
C3665667|T048|SY|46244001|SNOMEDCT_CORE|Recurrent major depression in complete remission|Recurrent major depression in full remission
C3665667|T048|OF|46244001|SNOMEDCT_CORE|Recurrent major depression in complete remission|Recurrent major depression in full remission
C3665667|T048|PT|46244001|SNOMEDCT_CORE|Recurrent major depression in full remission|Recurrent major depression in full remission
C3665667|T048|FN|46244001|SNOMEDCT_CORE|Recurrent major depression in full remission|Recurrent major depression in full remission
C3669043|T047|FN|697929007|SNOMEDCT_CORE|Intermittent hypertension|Intermittent hypertension
C3669043|T047|PT|697929007|SNOMEDCT_CORE|Intermittent hypertension|Intermittent hypertension
C3695127|T191|SY|254938000|SNOMEDCT_CORE|Astrocytic tumor of brain|Astrocytoma of brain
C3695127|T191|SYGB|254938000|SNOMEDCT_CORE|Astrocytic tumour of brain|Astrocytoma of brain
C3695127|T191|PT|254938000|SNOMEDCT_CORE|Astrocytoma of brain|Astrocytoma of brain
C3695127|T191|FN|254938000|SNOMEDCT_CORE|Astrocytoma of brain|Astrocytoma of brain
C3714509|T047|SY|2492009|SNOMEDCT_CORE|Disorder of nutrition|Nutritional disorder
C3714509|T047|SY|2492009|SNOMEDCT_CORE|Nutritional disease|Nutritional disorder
C3714509|T047|IS|2492009|SNOMEDCT_CORE|Nutritional disease, NOS|Nutritional disorder
C3714509|T047|PT|2492009|SNOMEDCT_CORE|Nutritional disorder|Nutritional disorder
C3714509|T047|FN|2492009|SNOMEDCT_CORE|Nutritional disorder|Nutritional disorder
C3714509|T047|IS|2492009|SNOMEDCT_CORE|Nutritional disorder, NOS|Nutritional disorder
C3714552|T184|SY|13791008|SNOMEDCT_CORE|Debility|Weakness
C3714552|T184|SY|13791008|SNOMEDCT_CORE|Feeling weak|Weakness
C3714552|T184|SY|13791008|SNOMEDCT_CORE|General weakness|Weakness
C3714552|T184|SY|13791008|SNOMEDCT_CORE|Lassitude|Weakness
C3714552|T184|SY|13791008|SNOMEDCT_CORE|Weakness|Weakness
C3714552|T184|SY|13791008|SNOMEDCT_CORE|Weakness - general|Weakness
C3714581|T047|SY|82525005|SNOMEDCT_CORE|Multicystic dysplastic kidney|Multicystic dysplastic kidney
C3714619|T047|IS|48606007|SNOMEDCT_CORE|Insulin resistance syndrome|Insulin resistance syndrome
C3714625|T033|PT|247398009|SNOMEDCT_CORE|Neuropathic pain|Neuropathic pain
C3714625|T033|FN|247398009|SNOMEDCT_CORE|Neuropathic pain|Neuropathic pain
C3714636|T047|PT|205237003|SNOMEDCT_CORE|Pneumonitis|Pneumonitis
C3714636|T047|FN|205237003|SNOMEDCT_CORE|Pneumonitis|Pneumonitis
C3714744|T048|PT|268637002|SNOMEDCT_CORE|Psychosexual dysfunction|Psychosexual dysfunction
C3714744|T048|FN|268637002|SNOMEDCT_CORE|Psychosexual dysfunction|Psychosexual dysfunction
C3714756|T048|SY|110359009|SNOMEDCT_CORE|Intellectual developmental disorder|Intellectual functioning disability
C3714756|T048|IS|228156007|SNOMEDCT_CORE|Intellectual disability|Intellectual functioning disability
C3714756|T048|IS|1855002|SNOMEDCT_CORE|Intellectual disability|Intellectual functioning disability
C3714756|T048|OF|110359009|SNOMEDCT_CORE|Intellectual disability|Intellectual functioning disability
C3714756|T048|PT|110359009|SNOMEDCT_CORE|Intellectual disability|Intellectual functioning disability
C3714756|T048|FN|110359009|SNOMEDCT_CORE|Intellectual disability|Intellectual functioning disability
C3714756|T048|PT|228156007|SNOMEDCT_CORE|Intellectual functioning disability|Intellectual functioning disability
C3714756|T048|FN|228156007|SNOMEDCT_CORE|Intellectual functioning disability|Intellectual functioning disability
C3714756|T048|IS|110359009|SNOMEDCT_CORE|Intellectual limitation|Intellectual functioning disability
C3714756|T048|IS|1855002|SNOMEDCT_CORE|Intellectual limitation|Intellectual functioning disability
C3714756|T048|SY|228156007|SNOMEDCT_CORE|Intellectual limitation|Intellectual functioning disability
C3714756|T048|SY|110359009|SNOMEDCT_CORE|Mental retardation|Intellectual functioning disability
C3714757|T047|SY|410795001|SNOMEDCT_CORE|JRA - Juvenile rheumatoid arthritis|Juvenile rheumatoid arthritis
C3714757|T047|PT|410795001|SNOMEDCT_CORE|Juvenile rheumatoid arthritis|Juvenile rheumatoid arthritis
C3714757|T047|FN|410795001|SNOMEDCT_CORE|Juvenile rheumatoid arthritis|Juvenile rheumatoid arthritis
C3714760|T047|SY|102449007|SNOMEDCT_CORE|Drug-induced tardive dyskinesia|Tardive dyskinesia
C3714760|T047|PT|102449007|SNOMEDCT_CORE|Tardive dyskinesia|Tardive dyskinesia
C3714760|T047|FN|102449007|SNOMEDCT_CORE|Tardive dyskinesia|Tardive dyskinesia
C3714760|T047|SY|102449007|SNOMEDCT_CORE|TD - Tardive dyskinesia|Tardive dyskinesia
C3853727|T033|SY|110483000|SNOMEDCT_CORE|Tobacco use|Tobacco user
C3853727|T033|PT|110483000|SNOMEDCT_CORE|Tobacco user|Tobacco user
C3853727|T033|FN|110483000|SNOMEDCT_CORE|Tobacco user|Tobacco user
C3853727|T033|OF|110483000|SNOMEDCT_CORE|Tobacco user|Tobacco user
C3854304|T019|IS|77945009|SNOMEDCT_CORE|Congenital renal cyst, single|Congenital renal cyst, single
C3875321|T047|PT|703938007|SNOMEDCT_CORE|Inflammatory dermatosis|Inflammatory dermatosis
C3875321|T047|FN|703938007|SNOMEDCT_CORE|Inflammatory dermatosis|Inflammatory dermatosis
C3887337|T019|PT|767002009|SNOMEDCT_CORE|Congenital dislocation of left hip|Congenital dislocation of left hip
C3887337|T019|FN|767002009|SNOMEDCT_CORE|Congenital dislocation of left hip|Congenital dislocation of left hip
C3887338|T019|PT|767003004|SNOMEDCT_CORE|Congenital dislocation of right hip|Congenital dislocation of right hip
C3887338|T019|FN|767003004|SNOMEDCT_CORE|Congenital dislocation of right hip|Congenital dislocation of right hip
C3887499|T047|PT|722223000|SNOMEDCT_CORE|Cyst of kidney|Cyst of kidney
C3887499|T047|FN|722223000|SNOMEDCT_CORE|Cyst of kidney|Cyst of kidney
C3887499|T047|SY|722223000|SNOMEDCT_CORE|Renal cyst|Cyst of kidney
C3887506|T047|SY|44548000|SNOMEDCT_CORE|Hyperkinesia|Hyperkinesia
C3887506|T047|IS|44548000|SNOMEDCT_CORE|Hyperkinesia, NOS|Hyperkinesia
C3887506|T047|IS|44548000|SNOMEDCT_CORE|Hyperkinesis, NOS|Hyperkinesia
C3887524|T047|SY|93448009|SNOMEDCT_CORE|Erosion of skin|Erosion of skin
C3887547|T047|SY|27405005|SNOMEDCT_CORE|Central sleep apnea|Central sleep apnea syndrome
C3887547|T047|PT|27405005|SNOMEDCT_CORE|Central sleep apnea syndrome|Central sleep apnea syndrome
C3887547|T047|FN|27405005|SNOMEDCT_CORE|Central sleep apnea syndrome|Central sleep apnea syndrome
C3887547|T047|SYGB|27405005|SNOMEDCT_CORE|Central sleep apnoea|Central sleep apnea syndrome
C3887547|T047|PTGB|27405005|SNOMEDCT_CORE|Central sleep apnoea syndrome|Central sleep apnea syndrome
C3887547|T047|SY|27405005|SNOMEDCT_CORE|CSA - Central sleep apnea|Central sleep apnea syndrome
C3887547|T047|SYGB|27405005|SNOMEDCT_CORE|CSA - Central sleep apnoea|Central sleep apnea syndrome
C3887551|T048|SY|386807006|SNOMEDCT_CORE|Memory dysfunction|Memory dysfunction
C3887597|T020|PT|1539003|SNOMEDCT_CORE|Acquired trigger finger|Acquired trigger finger
C3887597|T020|FN|1539003|SNOMEDCT_CORE|Acquired trigger finger|Acquired trigger finger
C3887597|T020|SY|1539003|SNOMEDCT_CORE|Nodular tendinous disease of finger|Acquired trigger finger
C3887597|T020|SY|1539003|SNOMEDCT_CORE|Trigger finger|Acquired trigger finger
C3887597|T020|SY|1539003|SNOMEDCT_CORE|Triggering of finger|Acquired trigger finger
C3887611|T184|IS|24199005|SNOMEDCT_CORE|Restless|Restlessness
C3887611|T184|IS|24199005|SNOMEDCT_CORE|Restlessness|Restlessness
C3887639|T047|SY|84568007|SNOMEDCT_CORE|Autoimmune gastritis|Autoimmune gastritis
C3887875|T033|SY|12184005|SNOMEDCT_CORE|VFD - Visual field defect|Visual field defect
C3887875|T033|PT|12184005|SNOMEDCT_CORE|Visual field defect|Visual field defect
C3887875|T033|FN|12184005|SNOMEDCT_CORE|Visual field defect|Visual field defect
C3887875|T033|IS|12184005|SNOMEDCT_CORE|Visual field defect, NOS|Visual field defect
C4039208|T046|PT|709493000|SNOMEDCT_CORE|Digestive system reflux|Digestive system reflux
C4039208|T046|FN|709493000|SNOMEDCT_CORE|Digestive system reflux|Digestive system reflux
C4040007|T047|PT|712537009|SNOMEDCT_CORE|Complex regional pain syndrome of upper limb|Complex regional pain syndrome of upper limb
C4040007|T047|FN|712537009|SNOMEDCT_CORE|Complex regional pain syndrome of upper limb|Complex regional pain syndrome of upper limb
C4040007|T047|OAS|2103002|SNOMEDCT_CORE|Reflex sympathetic dystrophy of upper extremity|Complex regional pain syndrome of upper limb
C4040007|T047|OAF|2103002|SNOMEDCT_CORE|Reflex sympathetic dystrophy of upper extremity|Complex regional pain syndrome of upper limb
C4040007|T047|SY|712537009|SNOMEDCT_CORE|Reflex sympathetic dystrophy of upper limb|Complex regional pain syndrome of upper limb
C4040007|T047|OAP|2103002|SNOMEDCT_CORE|Shoulder-hand syndrome|Complex regional pain syndrome of upper limb
C4040007|T047|OAS|2103002|SNOMEDCT_CORE|Steinbrocker's syndrome|Complex regional pain syndrome of upper limb
C4041032|T191|PT|708921005|SNOMEDCT_CORE|Carcinoma of central portion of breast|Carcinoma of central portion of breast
C4041032|T191|FN|708921005|SNOMEDCT_CORE|Carcinoma of central portion of breast|Carcinoma of central portion of breast
C4048328|T191|IS|363354003|SNOMEDCT_CORE|Ca cervix|Cancer of cervix
C4048328|T191|SY|363354003|SNOMEDCT_CORE|Cancer of cervix|Cancer of cervix
C4075133|T047|FN|714751007|SNOMEDCT_CORE|Inflammatory disorder of bone of jaw|Residual osteitis
C4075133|T047|SY|714751007|SNOMEDCT_CORE|Inflammatory disorder of bone of jaw|Residual osteitis
C4075133|T047|PT|714751007|SNOMEDCT_CORE|Residual osteitis|Residual osteitis
C4075825|T047|OF|713706002|SNOMEDCT_CORE|Polyneuropathy co-occurrent and due to type 2 diabetes mellitus|Polyneuropathy due to type 2 diabetes mellitus
C4075825|T047|IS|713706002|SNOMEDCT_CORE|Polyneuropathy co-occurrent and due to type 2 diabetes mellitus|Polyneuropathy due to type 2 diabetes mellitus
C4075825|T047|SY|713706002|SNOMEDCT_CORE|Polyneuropathy due to diabetes mellitus type II|Polyneuropathy due to type 2 diabetes mellitus
C4075825|T047|PT|713706002|SNOMEDCT_CORE|Polyneuropathy due to type 2 diabetes mellitus|Polyneuropathy due to type 2 diabetes mellitus
C4075825|T047|FN|713706002|SNOMEDCT_CORE|Polyneuropathy due to type 2 diabetes mellitus|Polyneuropathy due to type 2 diabetes mellitus
C4075839|T047|OF|713703005|SNOMEDCT_CORE|Gastroparesis co-occurrent and due to type 2 diabetes mellitus|Gastroparesis due to type 2 diabetes mellitus
C4075839|T047|IS|713703005|SNOMEDCT_CORE|Gastroparesis co-occurrent and due to type 2 diabetes mellitus|Gastroparesis due to type 2 diabetes mellitus
C4075839|T047|SY|713703005|SNOMEDCT_CORE|Gastroparesis due to diabetes mellitus type II|Gastroparesis due to type 2 diabetes mellitus
C4075839|T047|PT|713703005|SNOMEDCT_CORE|Gastroparesis due to type 2 diabetes mellitus|Gastroparesis due to type 2 diabetes mellitus
C4075839|T047|FN|713703005|SNOMEDCT_CORE|Gastroparesis due to type 2 diabetes mellitus|Gastroparesis due to type 2 diabetes mellitus
C4075839|T047|SY|713703005|SNOMEDCT_CORE|Gastroparesis with type 2 diabetes mellitus|Gastroparesis due to type 2 diabetes mellitus
C4082762|T047|SY|402134005|SNOMEDCT_CORE|Dermatophytosis of nail|Onychomycosis due to dermatophyte
C4082762|T047|SY|402134005|SNOMEDCT_CORE|Onychomycosis caused by dermatophyte|Onychomycosis due to dermatophyte
C4082762|T047|FN|402134005|SNOMEDCT_CORE|Onychomycosis caused by dermatophyte|Onychomycosis due to dermatophyte
C4082762|T047|OF|402134005|SNOMEDCT_CORE|Onychomycosis due to dermatophyte|Onychomycosis due to dermatophyte
C4082762|T047|PT|402134005|SNOMEDCT_CORE|Onychomycosis due to dermatophyte|Onychomycosis due to dermatophyte
C4082762|T047|SY|402134005|SNOMEDCT_CORE|Tinea of nail|Onychomycosis due to dermatophyte
C4082762|T047|SY|402134005|SNOMEDCT_CORE|Tinea unguium|Onychomycosis due to dermatophyte
C4082764|T047|PT|715852004|SNOMEDCT_CORE|Gastrointestinal infection|Gastrointestinal infection
C4082764|T047|SY|715852004|SNOMEDCT_CORE|Infection of gastrointestinal tract|Gastrointestinal infection
C4082764|T047|FN|715852004|SNOMEDCT_CORE|Infection of gastrointestinal tract|Gastrointestinal infection
C4082974|T047|SY|410812005|SNOMEDCT_CORE|Dupuytren disease|Dupuytren's disease
C4082974|T047|PT|410812005|SNOMEDCT_CORE|Dupuytren's disease|Dupuytren's disease
C4082974|T047|FN|410812005|SNOMEDCT_CORE|Dupuytren's disease|Dupuytren's disease
C4083212|T047|SY|87872006|SNOMEDCT_CORE|Androgenetic alopecia|Male pattern alopecia
C4083212|T047|SY|87872006|SNOMEDCT_CORE|Androgenic alopecia|Male pattern alopecia
C4083212|T047|SY|87872006|SNOMEDCT_CORE|Common baldness|Male pattern alopecia
C4083212|T047|SY|87872006|SNOMEDCT_CORE|Hereditary alopecia|Male pattern alopecia
C4083212|T047|PT|87872006|SNOMEDCT_CORE|Male pattern alopecia|Male pattern alopecia
C4083212|T047|FN|87872006|SNOMEDCT_CORE|Male pattern alopecia|Male pattern alopecia
C4083212|T047|SY|87872006|SNOMEDCT_CORE|Male pattern baldness|Male pattern alopecia
C4083212|T047|SY|87872006|SNOMEDCT_CORE|Pattern baldness|Male pattern alopecia
C4280951|T033|PT|762898005|SNOMEDCT_CORE|Swelling of bilateral lower limbs|Swelling of bilateral lower limbs
C4280951|T033|FN|762898005|SNOMEDCT_CORE|Swelling of bilateral lower limbs|Swelling of bilateral lower limbs
C4282032|T191|IS|398838000|SNOMEDCT_CORE|Basal cell papilloma|Senile hyperkeratosis
C4282032|T191|IS|398838000|SNOMEDCT_CORE|BCP - Basal cell papilloma|Senile hyperkeratosis
C4282032|T191|SY|398838000|SNOMEDCT_CORE|Keratosis senilis|Senile hyperkeratosis
C4282032|T191|IS|398838000|SNOMEDCT_CORE|Pigmented basal cell papilloma|Senile hyperkeratosis
C4282032|T191|IS|398838000|SNOMEDCT_CORE|Seborrheic wart|Senile hyperkeratosis
C4282032|T191|IS|398838000|SNOMEDCT_CORE|Seborrhoeic wart|Senile hyperkeratosis
C4282032|T191|PT|398838000|SNOMEDCT_CORE|Senile hyperkeratosis|Senile hyperkeratosis
C4282032|T191|FN|398838000|SNOMEDCT_CORE|Senile hyperkeratosis|Senile hyperkeratosis
C4282032|T191|SY|398838000|SNOMEDCT_CORE|Senile keratosis|Senile hyperkeratosis
C4282032|T191|SY|398838000|SNOMEDCT_CORE|Senile wart|Senile hyperkeratosis
C4302291|T037|PT|722813003|SNOMEDCT_CORE|Strain of tendon of wrist|Strain of tendon of wrist
C4302291|T037|FN|722813003|SNOMEDCT_CORE|Strain of tendon of wrist|Strain of tendon of wrist
C4302760|T037|PT|10850741000119108|SNOMEDCT_CORE|Accidental needle stick injury|Accidental needle stick injury
C4302760|T037|FN|10850741000119108|SNOMEDCT_CORE|Accidental needle stick injury|Accidental needle stick injury
C4304130|T033|PT|12275351000119103|SNOMEDCT_CORE|Breast cancer screening declined|Breast cancer screening declined
C4304130|T033|FN|12275351000119103|SNOMEDCT_CORE|Breast cancer screening declined|Breast cancer screening declined
C4304387|T047|PT|719860006|SNOMEDCT_CORE|Acute infectious conjunctivitis|Acute infectious conjunctivitis
C4304387|T047|FN|719860006|SNOMEDCT_CORE|Acute infectious conjunctivitis|Acute infectious conjunctivitis
C4317009|T047|SY|397881000|SNOMEDCT_CORE|DD - Diverticular disease|Diverticular disease
C4317009|T047|PT|397881000|SNOMEDCT_CORE|Diverticular disease|Diverticular disease
C4317009|T047|FN|397881000|SNOMEDCT_CORE|Diverticular disease|Diverticular disease
C4317009|T047|IS|397881000|SNOMEDCT_CORE|Diverticulosis|Diverticular disease
C4317109|T047|SY|313307000|SNOMEDCT_CORE|Epileptic attack|Epileptic seizure
C4317109|T047|SY|313307000|SNOMEDCT_CORE|Epileptic convulsion|Epileptic seizure
C4317109|T047|SY|313307000|SNOMEDCT_CORE|Epileptic fit|Epileptic seizure
C4317109|T047|PT|313307000|SNOMEDCT_CORE|Epileptic seizure|Epileptic seizure
C4317109|T047|FN|313307000|SNOMEDCT_CORE|Epileptic seizure|Epileptic seizure
C4509972|T033|PT|723620004|SNOMEDCT_CORE|Requires vaccination|Requires vaccination
C4509972|T033|FN|723620004|SNOMEDCT_CORE|Requires vaccination|Requires vaccination
C4520843|T047|PT|77489003|SNOMEDCT_CORE|Pterygium|Pterygium
C4520843|T047|FN|77489003|SNOMEDCT_CORE|Pterygium|Pterygium
C4520843|T047|IS|77489003|SNOMEDCT_CORE|Pterygium, NOS|Pterygium
C4520843|T047|SY|77489003|SNOMEDCT_CORE|Web eye|Pterygium
C4520847|T033|SY|123785006|SNOMEDCT_CORE|IgG subclass deficiency|Immunoglobulin G subclass deficiency
C4520847|T033|OF|123785006|SNOMEDCT_CORE|Immunoglobin G subclass deficiency|Immunoglobulin G subclass deficiency
C4520847|T033|SY|123785006|SNOMEDCT_CORE|Immunoglobin G subclass deficiency|Immunoglobulin G subclass deficiency
C4520847|T033|FN|123785006|SNOMEDCT_CORE|Immunoglobulin G subclass deficiency|Immunoglobulin G subclass deficiency
C4520847|T033|PT|123785006|SNOMEDCT_CORE|Immunoglobulin G subclass deficiency|Immunoglobulin G subclass deficiency
C4543483|T047|SY|734986006|SNOMEDCT_CORE|Complex regional pain syndrome of lower extremity|Complex regional pain syndrome of lower limb
C4543483|T047|PT|734986006|SNOMEDCT_CORE|Complex regional pain syndrome of lower limb|Complex regional pain syndrome of lower limb
C4543483|T047|FN|734986006|SNOMEDCT_CORE|Complex regional pain syndrome of lower limb|Complex regional pain syndrome of lower limb
C4544405|T047|PT|736499003|SNOMEDCT_CORE|Polyp of nasal cavity and/or nasal sinus|Polyp of nasal cavity and/or nasal sinus
C4544405|T047|FN|736499003|SNOMEDCT_CORE|Polyp of nasal cavity and/or nasal sinus|Polyp of nasal cavity and/or nasal sinus
C4545499|T047|SY|739681000|SNOMEDCT_CORE|Diabetic oculopathy due to type 1 diabetes mellitus|Disorder of eye due to type 1 diabetes mellitus
C4545499|T047|OF|739681000|SNOMEDCT_CORE|Diabetic oculopathy due to type I diabetes mellitus|Disorder of eye due to type 1 diabetes mellitus
C4545499|T047|SY|739681000|SNOMEDCT_CORE|Diabetic oculopathy due to type I diabetes mellitus|Disorder of eye due to type 1 diabetes mellitus
C4545499|T047|OF|739681000|SNOMEDCT_CORE|Disorder of eye co-occurrent and due to type 1 diabetes mellitus|Disorder of eye due to type 1 diabetes mellitus
C4545499|T047|IS|739681000|SNOMEDCT_CORE|Disorder of eye co-occurrent and due to type 1 diabetes mellitus|Disorder of eye due to type 1 diabetes mellitus
C4545499|T047|PT|739681000|SNOMEDCT_CORE|Disorder of eye due to type 1 diabetes mellitus|Disorder of eye due to type 1 diabetes mellitus
C4545499|T047|FN|739681000|SNOMEDCT_CORE|Disorder of eye due to type 1 diabetes mellitus|Disorder of eye due to type 1 diabetes mellitus
C4545499|T047|SY|739681000|SNOMEDCT_CORE|Disorder of eye with type 1 diabetes mellitus|Disorder of eye due to type 1 diabetes mellitus
C4545715|T047|OAP|746009000|SNOMEDCT_CORE|Left femoral hernia without obstruction and without gangrene|Left femoral hernia without obstruction and without gangrene
C4545715|T047|OAF|746009000|SNOMEDCT_CORE|Left femoral hernia without obstruction and without gangrene|Left femoral hernia without obstruction and without gangrene
C4545718|T047|OAP|746010005|SNOMEDCT_CORE|Right femoral hernia without obstruction and without gangrene|Right femoral hernia without obstruction and without gangrene
C4545718|T047|OAF|746010005|SNOMEDCT_CORE|Right femoral hernia without obstruction and without gangrene|Right femoral hernia without obstruction and without gangrene
C4546414|T019|SY|762907005|SNOMEDCT_CORE|Agenesis of left kidney|Left renal agenesis
C4546414|T019|FN|762907005|SNOMEDCT_CORE|Agenesis of left kidney|Left renal agenesis
C4546414|T019|PT|762907005|SNOMEDCT_CORE|Left renal agenesis|Left renal agenesis
C4546415|T019|FN|762908000|SNOMEDCT_CORE|Agenesis of right kidney|Right renal agenesis
C4546415|T019|SY|762908000|SNOMEDCT_CORE|Agenesis of right kidney|Right renal agenesis
C4546415|T019|PT|762908000|SNOMEDCT_CORE|Right renal agenesis|Right renal agenesis
C4551518|T046|PT|71897006|SNOMEDCT_CORE|Venous stasis|Venous stasis
C4551518|T046|FN|71897006|SNOMEDCT_CORE|Venous stasis|Venous stasis
C4551518|T046|IS|71897006|SNOMEDCT_CORE|Venous stasis, NOS|Venous stasis
C4551520|T184|SY|30721006|SNOMEDCT_CORE|Cerebellar tremor|Intention tremor
C4551520|T184|IS|30721006|SNOMEDCT_CORE|Hunt's tremor|Intention tremor
C4551520|T184|PT|30721006|SNOMEDCT_CORE|Intention tremor|Intention tremor
C4551520|T184|FN|30721006|SNOMEDCT_CORE|Intention tremor|Intention tremor
C4551520|T184|SY|30721006|SNOMEDCT_CORE|Volitional tremor|Intention tremor
C4551521|T184|SY|30721006|SNOMEDCT_CORE|Kinetic tremor|Kinetic tremor
C4551636|T047|IS|42513006|SNOMEDCT_CORE|Thygeson's superficial punctate keratitis|Thygeson's superficial punctate keratitis
C4551650|T047|SY|63305008|SNOMEDCT_CORE|Esophageal stricture|Stricture of esophagus
C4551650|T047|SYGB|63305008|SNOMEDCT_CORE|Oesophageal stricture|Stricture of esophagus
C4551650|T047|PT|63305008|SNOMEDCT_CORE|Stricture of esophagus|Stricture of esophagus
C4551650|T047|FN|63305008|SNOMEDCT_CORE|Stricture of esophagus|Stricture of esophagus
C4551650|T047|PTGB|63305008|SNOMEDCT_CORE|Stricture of oesophagus|Stricture of esophagus
C4551651|T047|IS|47639008|SNOMEDCT_CORE|Coccygeal fistula|Coccygeal fistula
C4551651|T047|IS|47639008|SNOMEDCT_CORE|Pilonidal fistula|Coccygeal fistula
C4551659|T047|SYGB|28998008|SNOMEDCT_CORE|Intraretinal haemorrhage|Intraretinal hemorrhage
C4551659|T047|SY|28998008|SNOMEDCT_CORE|Intraretinal hemorrhage|Intraretinal hemorrhage
C4551677|T019|IS|414667000|SNOMEDCT_CORE|Myelocystocele|Myelocystocele
C4551685|T033|SY|64228003|SNOMEDCT_CORE|Diaphragmatic paralysis|Paralysis of diaphragm
C4551685|T033|PT|64228003|SNOMEDCT_CORE|Paralysis of diaphragm|Paralysis of diaphragm
C4551685|T033|FN|64228003|SNOMEDCT_CORE|Paralysis of diaphragm|Paralysis of diaphragm
C4551691|T047|PT|76618002|SNOMEDCT_CORE|Urethral stricture|Urethral stricture
C4551691|T047|FN|76618002|SNOMEDCT_CORE|Urethral stricture|Urethral stricture
C4551691|T047|IS|76618002|SNOMEDCT_CORE|Urethral stricture, NOS|Urethral stricture
C4551754|T033|SY|165746003|SNOMEDCT_CORE|Rh negative|RhD negative
C4551754|T033|OF|165746003|SNOMEDCT_CORE|Rh negative|RhD negative
C4551754|T033|PT|165746003|SNOMEDCT_CORE|RhD negative|RhD negative
C4551754|T033|FN|165746003|SNOMEDCT_CORE|RhD negative|RhD negative
C4551754|T033|SY|165746003|SNOMEDCT_CORE|Rhesus negative|RhD negative
C4551827|T047|IS|73297009|SNOMEDCT_CORE|Hereditary progressive muscular dystrophy|Hereditary progressive muscular dystrophy
C4551862|T047|SY|28978003|SNOMEDCT_CORE|Nuchal dystonia-dementia syndrome|Progressive supranuclear ophthalmoplegia
C4551862|T047|PT|28978003|SNOMEDCT_CORE|Progressive supranuclear ophthalmoplegia|Progressive supranuclear ophthalmoplegia
C4551862|T047|FN|28978003|SNOMEDCT_CORE|Progressive supranuclear ophthalmoplegia|Progressive supranuclear ophthalmoplegia
C4551862|T047|IS|28978003|SNOMEDCT_CORE|Steele-Richardson-Olszewski syndrome|Progressive supranuclear ophthalmoplegia
C4552097|T047|SYGB|52298009|SNOMEDCT_CORE|Linear sebaceous naevus|Linear sebaceous nevus sequence
C4552097|T047|PTGB|52298009|SNOMEDCT_CORE|Linear sebaceous naevus sequence|Linear sebaceous nevus sequence
C4552097|T047|SY|52298009|SNOMEDCT_CORE|Linear sebaceous nevus|Linear sebaceous nevus sequence
C4552097|T047|PT|52298009|SNOMEDCT_CORE|Linear sebaceous nevus sequence|Linear sebaceous nevus sequence
C4552097|T047|FN|52298009|SNOMEDCT_CORE|Linear sebaceous nevus sequence|Linear sebaceous nevus sequence
C4552097|T047|IS|52298009|SNOMEDCT_CORE|Naevus sebaceous of Jadassohn|Linear sebaceous nevus sequence
C4552097|T047|IS|52298009|SNOMEDCT_CORE|Naevus sebaceus of Jadassohn|Linear sebaceous nevus sequence
C4552097|T047|IS|52298009|SNOMEDCT_CORE|Nevus sebaceous of Jadassohn|Linear sebaceous nevus sequence
C4552097|T047|IS|52298009|SNOMEDCT_CORE|Nevus sebaceus of Jadassohn|Linear sebaceous nevus sequence
C4552097|T047|IS|52298009|SNOMEDCT_CORE|Organoid naevus|Linear sebaceous nevus sequence
C4552097|T047|IS|52298009|SNOMEDCT_CORE|Organoid nevus|Linear sebaceous nevus sequence
C4552097|T047|IS|52298009|SNOMEDCT_CORE|Sebaceous nevus|Linear sebaceous nevus sequence
C4552100|T047|OP|315058005|SNOMEDCT_CORE|Lynch syndrome|Lynch syndrome
C4707419|T033|PT|765378003|SNOMEDCT_CORE|History of primary malignant neoplasm of skin|History of primary malignant neoplasm of skin
C4707419|T033|FN|765378003|SNOMEDCT_CORE|History of primary malignant neoplasm of skin|History of primary malignant neoplasm of skin
C4707862|T033|PT|766877008|SNOMEDCT_CORE|Constantly crying infant|Constantly crying infant
C4707862|T033|FN|766877008|SNOMEDCT_CORE|Constantly crying infant|Constantly crying infant
C4708167|T047|PTGB|767657005|SNOMEDCT_CORE|Anaemia due to and following chemotherapy|Anemia due to and following chemotherapy
C4708167|T047|PT|767657005|SNOMEDCT_CORE|Anemia due to and following chemotherapy|Anemia due to and following chemotherapy
C4708167|T047|FN|767657005|SNOMEDCT_CORE|Anemia due to and following chemotherapy|Anemia due to and following chemotherapy
C4708168|T047|PTGB|767658000|SNOMEDCT_CORE|Neutropaenia due to and following chemotherapy|Neutropenia due to and following chemotherapy
C4708168|T047|PT|767658000|SNOMEDCT_CORE|Neutropenia due to and following chemotherapy|Neutropenia due to and following chemotherapy
C4708168|T047|FN|767658000|SNOMEDCT_CORE|Neutropenia due to and following chemotherapy|Neutropenia due to and following chemotherapy
C4708188|T190|OAP|767690005|SNOMEDCT_CORE|Obstruction without gangrene co-occurrent and due to right inguinal hernia|Obstruction without gangrene co-occurrent and due to right inguinal hernia
C4708188|T190|OAF|767690005|SNOMEDCT_CORE|Obstruction without gangrene co-occurrent and due to right inguinal hernia|Obstruction without gangrene co-occurrent and due to right inguinal hernia
C4708189|T190|OAP|767691009|SNOMEDCT_CORE|Obstruction without gangrene co-occurrent and due to left inguinal hernia|Obstruction without gangrene co-occurrent and due to left inguinal hernia
C4708189|T190|OAF|767691009|SNOMEDCT_CORE|Obstruction without gangrene co-occurrent and due to left inguinal hernia|Obstruction without gangrene co-occurrent and due to left inguinal hernia
C4708260|T047|OAP|767746007|SNOMEDCT_CORE|Obstruction without gangrene co-occurrent and due to recurrent left inguinal hernia|Obstruction without gangrene co-occurrent and due to recurrent left inguinal hernia
C4708260|T047|OAF|767746007|SNOMEDCT_CORE|Obstruction without gangrene co-occurrent and due to recurrent left inguinal hernia|Obstruction without gangrene co-occurrent and due to recurrent left inguinal hernia
C4708261|T047|OAP|767747003|SNOMEDCT_CORE|Obstruction without gangrene co-occurrent and due to recurrent right inguinal hernia|Obstruction without gangrene co-occurrent and due to recurrent right inguinal hernia
C4708261|T047|OAF|767747003|SNOMEDCT_CORE|Obstruction without gangrene co-occurrent and due to recurrent right inguinal hernia|Obstruction without gangrene co-occurrent and due to recurrent right inguinal hernia
C4721411|T046|PT|203522001|SNOMEDCT_CORE|Osteolysis|Osteolysis
C4721411|T046|FN|203522001|SNOMEDCT_CORE|Osteolysis|Osteolysis
C4721414|T191|PT|443487006|SNOMEDCT_CORE|Mantle cell lymphoma|Mantle cell lymphoma
C4721414|T191|FN|443487006|SNOMEDCT_CORE|Mantle cell lymphoma|Mantle cell lymphoma
C4721444|T191|PTGB|277571004|SNOMEDCT_CORE|B-cell acute lymphoblastic leukaemia|B-cell acute lymphoblastic leukaemia
C4721444|T191|SYGB|277571004|SNOMEDCT_CORE|Burkitt's leukaemia|Burkitt's leukaemia
C4721444|T191|SY|277571004|SNOMEDCT_CORE|Burkitt's leukemia|Burkitt's leukemia
C4721453|T047|PT|42658009|SNOMEDCT_CORE|Disorder of the peripheral nervous system|Peripheral nerve disease
C4721453|T047|FN|42658009|SNOMEDCT_CORE|Disorder of the peripheral nervous system|Peripheral nerve disease
C4721453|T047|IS|42658009|SNOMEDCT_CORE|Disorder of the peripheral nervous system, NOS|Peripheral nerve disease
C4721453|T047|PT|302226006|SNOMEDCT_CORE|Peripheral nerve disease|Peripheral nerve disease
C4721453|T047|FN|302226006|SNOMEDCT_CORE|Peripheral nerve disease|Peripheral nerve disease
C4721453|T047|IS|42658009|SNOMEDCT_CORE|Peripheral nerve disorder|Peripheral nerve disease
C4721453|T047|IS|42658009|SNOMEDCT_CORE|Peripheral nerve disorder, NOS|Peripheral nerve disease
C4721453|T047|IS|42658009|SNOMEDCT_CORE|Peripheral neuropathy|Peripheral nerve disease
C4721453|T047|SY|302226006|SNOMEDCT_CORE|Peripheral neuropathy|Peripheral nerve disease
C4721453|T047|IS|42658009|SNOMEDCT_CORE|Peripheral neuropathy, NOS|Peripheral nerve disease
C4721453|T047|IS|42658009|SNOMEDCT_CORE|PN - Peripheral neuropathy|Peripheral nerve disease
C4721508|T047|IS|45157009|SNOMEDCT_CORE|Hamman-Rich disease|Hamman-Rich disease
C4721555|T047|PT|408335007|SNOMEDCT_CORE|Autoimmune hepatitis|Autoimmune hepatitis
C4721555|T047|FN|408335007|SNOMEDCT_CORE|Autoimmune hepatitis|Autoimmune hepatitis
C4721579|T191|IS|94365007|SNOMEDCT_CORE|Metastatic colorectal cancer|Metastatic colorectal cancer
C4721806|T191|PT|254701007|SNOMEDCT_CORE|Basal cell carcinoma of skin|Basal cell carcinoma of skin
C4721806|T191|FN|254701007|SNOMEDCT_CORE|Basal cell carcinoma of skin|Basal cell carcinoma of skin
C4721806|T191|SY|254701007|SNOMEDCT_CORE|Basalioma|Basal cell carcinoma of skin
C4721806|T191|SY|254701007|SNOMEDCT_CORE|BCC - Basal cell carcinoma of skin|Basal cell carcinoma of skin
C4721806|T191|SY|254701007|SNOMEDCT_CORE|Cancer of skin, basal cell|Basal cell carcinoma of skin
C4721806|T191|SY|254701007|SNOMEDCT_CORE|Rodent ulcer|Basal cell carcinoma of skin
C4721806|T191|SY|254701007|SNOMEDCT_CORE|RU - Rodent ulcer|Basal cell carcinoma of skin
C4722157|T046|PT|771113001|SNOMEDCT_CORE|Sodium retention|Sodium retention
C4722157|T046|FN|771113001|SNOMEDCT_CORE|Sodium retention|Sodium retention
C4750120|T033|SY|772005003|SNOMEDCT_CORE|Failed delivery by vacuum extraction|Failed ventouse delivery
C4750120|T033|PT|772005003|SNOMEDCT_CORE|Failed ventouse delivery|Failed ventouse delivery
C4750120|T033|FN|772005003|SNOMEDCT_CORE|Failed ventouse delivery|Failed ventouse delivery
C4750323|T047|PT|772139001|SNOMEDCT_CORE|Obstruction co-occurrent and due to left femoral hernia|Obstruction co-occurrent and due to left femoral hernia
C4750323|T047|FN|772139001|SNOMEDCT_CORE|Obstruction co-occurrent and due to left femoral hernia|Obstruction co-occurrent and due to left femoral hernia
C4750324|T047|PT|772140004|SNOMEDCT_CORE|Obstruction co-occurrent and due to right femoral hernia|Obstruction co-occurrent and due to right femoral hernia
C4750324|T047|FN|772140004|SNOMEDCT_CORE|Obstruction co-occurrent and due to right femoral hernia|Obstruction co-occurrent and due to right femoral hernia
C4750325|T047|PT|772141000|SNOMEDCT_CORE|Obstruction co-occurrent and due to recurrent right inguinal hernia|Obstruction co-occurrent and due to recurrent right inguinal hernia
C4750325|T047|FN|772141000|SNOMEDCT_CORE|Obstruction co-occurrent and due to recurrent right inguinal hernia|Obstruction co-occurrent and due to recurrent right inguinal hernia
C4750326|T047|PT|772142007|SNOMEDCT_CORE|Obstruction co-occurrent and due to recurrent left inguinal hernia|Obstruction co-occurrent and due to recurrent left inguinal hernia
C4750326|T047|FN|772142007|SNOMEDCT_CORE|Obstruction co-occurrent and due to recurrent left inguinal hernia|Obstruction co-occurrent and due to recurrent left inguinal hernia
C4750327|T047|PT|772143002|SNOMEDCT_CORE|Obstruction co-occurrent and due to left inguinal hernia|Obstruction co-occurrent and due to left inguinal hernia
C4750327|T047|FN|772143002|SNOMEDCT_CORE|Obstruction co-occurrent and due to left inguinal hernia|Obstruction co-occurrent and due to left inguinal hernia
C4750328|T047|PT|772144008|SNOMEDCT_CORE|Obstruction co-occurrent and due to right inguinal hernia|Obstruction co-occurrent and due to right inguinal hernia
C4750328|T047|FN|772144008|SNOMEDCT_CORE|Obstruction co-occurrent and due to right inguinal hernia|Obstruction co-occurrent and due to right inguinal hernia
C4758660|T047|PT|782594005|SNOMEDCT_CORE|Allergy to soy protein|Allergy to soy protein
C4758660|T047|FN|782594005|SNOMEDCT_CORE|Allergy to soy protein|Allergy to soy protein
C4759705|T047|SY|310387003|SNOMEDCT_CORE|Diabetic intracapillary glomerulosclerosis|Intracapillary glomerulosclerosis of kidney due to diabetes mellitus
C4759705|T047|OF|310387003|SNOMEDCT_CORE|Diabetic intracapillary glomerulosclerosis|Intracapillary glomerulosclerosis of kidney due to diabetes mellitus
C4759705|T047|OF|310387003|SNOMEDCT_CORE|Intracapillary glomerulosclerosis due to diabetes mellitus|Intracapillary glomerulosclerosis of kidney due to diabetes mellitus
C4759705|T047|SY|310387003|SNOMEDCT_CORE|Intracapillary glomerulosclerosis due to diabetes mellitus|Intracapillary glomerulosclerosis of kidney due to diabetes mellitus
C4759705|T047|PT|310387003|SNOMEDCT_CORE|Intracapillary glomerulosclerosis of kidney due to diabetes mellitus|Intracapillary glomerulosclerosis of kidney due to diabetes mellitus
C4759705|T047|FN|310387003|SNOMEDCT_CORE|Intracapillary glomerulosclerosis of kidney due to diabetes mellitus|Intracapillary glomerulosclerosis of kidney due to diabetes mellitus
C4759727|T047|SY|402863005|SNOMEDCT_CORE|Gravitational ulcer|Venous stasis ulcer of leg
C4759727|T047|SY|402863005|SNOMEDCT_CORE|Stasis ulcer of leg|Venous stasis ulcer of leg
C4759727|T047|PT|402863005|SNOMEDCT_CORE|Venous stasis ulcer of leg|Venous stasis ulcer of leg
C4759727|T047|FN|402863005|SNOMEDCT_CORE|Venous stasis ulcer of leg|Venous stasis ulcer of leg
C4759727|T047|SY|402863005|SNOMEDCT_CORE|Venous ulcer of leg|Venous stasis ulcer of leg
C4759727|T047|OF|402863005|SNOMEDCT_CORE|Venous ulcer of leg|Venous stasis ulcer of leg
C4761312|T047|SY|70241007|SNOMEDCT_CORE|Dietary deficiency|Nutritional deficiency disorder
C4761312|T047|SY|70241007|SNOMEDCT_CORE|Nutritional deficiencies|Nutritional deficiency disorder
C4761312|T047|SY|70241007|SNOMEDCT_CORE|Nutritional deficiency|Nutritional deficiency disorder
C4761312|T047|OF|70241007|SNOMEDCT_CORE|Nutritional deficiency|Nutritional deficiency disorder
C4761312|T047|PT|70241007|SNOMEDCT_CORE|Nutritional deficiency disorder|Nutritional deficiency disorder
C4761312|T047|FN|70241007|SNOMEDCT_CORE|Nutritional deficiency disorder|Nutritional deficiency disorder
C4761312|T047|IS|70241007|SNOMEDCT_CORE|Nutritional deficiency disorder, NOS|Nutritional deficiency disorder
C4761312|T047|IS|70241007|SNOMEDCT_CORE|Nutritional deficiency, NOS|Nutritional deficiency disorder
C5190995|T033|PT|783572008|SNOMEDCT_CORE|Has special educational needs|Has special educational needs
C5190995|T033|FN|783572008|SNOMEDCT_CORE|Has special educational needs|Has special educational needs
C5191627|T047|PT|785696007|SNOMEDCT_CORE|Malabsorption syndrome due to intolerance to lactose|Malabsorption syndrome due to intolerance to lactose
C5191627|T047|FN|785696007|SNOMEDCT_CORE|Malabsorption syndrome due to intolerance to lactose|Malabsorption syndrome due to intolerance to lactose
C5191648|T047|PT|785744001|SNOMEDCT_CORE|Bronchitis co-occurrent with acute wheeze|Bronchitis co-occurrent with acute wheeze
C5191648|T047|FN|785744001|SNOMEDCT_CORE|Bronchitis co-occurrent with acute wheeze|Bronchitis co-occurrent with acute wheeze
C5191649|T047|PT|785745000|SNOMEDCT_CORE|Acute bronchitis co-occurrent with wheeze|Acute bronchitis co-occurrent with wheeze
C5191649|T047|FN|785745000|SNOMEDCT_CORE|Acute bronchitis co-occurrent with wheeze|Acute bronchitis co-occurrent with wheeze
C5192274|T048|PT|786919007|SNOMEDCT_CORE|Sexually assaultive behavior|Sexually assaultive behavior
C5192274|T048|FN|786919007|SNOMEDCT_CORE|Sexually assaultive behavior|Sexually assaultive behavior
C5192274|T048|PTGB|786919007|SNOMEDCT_CORE|Sexually assaultive behaviour|Sexually assaultive behavior
C5200920|T048|PT|29212009|SNOMEDCT_CORE|Alcohol-induced organic mental disorder|Alcohol-induced organic mental disorder
C5200920|T048|FN|29212009|SNOMEDCT_CORE|Alcohol-induced organic mental disorder|Alcohol-induced organic mental disorder
C5200920|T048|IS|29212009|SNOMEDCT_CORE|Alcohol-induced organic mental disorder, NOS|Alcohol-induced organic mental disorder
C5200920|T048|SY|29212009|SNOMEDCT_CORE|Alcohol-related disorder|Alcohol-induced organic mental disorder
C5200920|T048|IS|29212009|SNOMEDCT_CORE|Alcohol-related disorder, NOS|Alcohol-induced organic mental disorder
C5200931|T033|IS|192007009|SNOMEDCT_CORE|"Short-sleeper"|Short-sleeper
C5200931|T033|PT|192007009|SNOMEDCT_CORE|Short-sleeper|Short-sleeper
C5200931|T033|FN|192007009|SNOMEDCT_CORE|Short-sleeper|Short-sleeper
C5200931|T033|OF|192007009|SNOMEDCT_CORE|Short-sleeper|Short-sleeper
