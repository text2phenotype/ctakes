C0019683|T034||LNC|HIV AB
C0019683|T034||LNC|HIV ANTIBODIES
C3714540|T034||LNC|HIV ANTIBODY TEST
C3714540|T034||LNC|HIV ANTIBODY MEASUREMENT
C0019683|T034||LNC|ANTIBODIES, AIDS
C0019683|T034||LNC|ANTIBODIES, HIV
C0019683|T034||LNC|ANTIBODIES, HIV ASSOCIATED
C0019683|T034||LNC|ANTIBODIES, HIV-ASSOCIATED
C0019683|T034||LNC| THIS IS THE OLD NAME FOR HIV, BUT NOW REFERS TO A NEW AND DIFFERENT VIRUS. THERE'S A CHANCE YOU MIGHT MISS SOME PEOPLE WHO WERE DIAGNOSED A LONG TIME AGO BY EXCLUDING IT, BUT IT SEEMS UNLIKELY TO ME
C0019683|T034||LNC|ANTIBODIES, HTLV-III
C0019683|T034||LNC|THIS IS AN OLD BUT SPECIFIC NAME FOR HIV, SAFE TO INCLUDE
C0019683|T034||LNC|ANTIBODIES, LAV
C0019683|T034||LNC|ANTIBODIES, LYMPHADENOPATHY ASSOCIATED
C0019683|T034||LNC|ANTIBODIES, LYMPHADENOPATHY-ASSOCIATED
C0019683|T034||LNC|HIV ANTIBODIES
C0019683|T034||LNC|HTLV WIII ANTIBODIES
C0019683|T034||LNC|HTLV WIII LAV ANTIBODIES
C0019683|T034||LNC|LYMPHOTROPIC VIRUS TYPE III ANTIBODIES HUMAN T
C0019683|T034||LNC|HTLV-III ANTIBODIES
C0019683|T034||LNC|HIV ANTIBODIES [CHEMICAL/INGREDIENT]
C0019683|T034||LNC|HTLV III ANTIBODIES
C0019683|T034||LNC|LAV ANTIBODIES
C0019683|T034||LNC|LYMPHADENOPATHY ASSOCIATED ANTIBODIES
C0019683|T034||LNC|T LYMPHOTROPIC VIRUS TYPE III ANTIBODIES, HUMAN
C0019683|T034||LNC|AIDS ANTIBODIES
C0019683|T034||LNC|HIV ASSOCIATED ANTIBODIES
C0019683|T034||LNC|T-LYMPHOTROPIC VIRUS TYPE III ANTIBODIES, HUMAN
C0019683|T034||LNC|HIV-ASSOCIATED ANTIBODIES
C0019683|T034||LNC|HTLV-III-LAV ANTIBODIES
C0019683|T034||LNC|HTLV III LAV ANTIBODIES
C0019683|T034||LNC|LYMPHADENOPATHY-ASSOCIATED ANTIBODIES
C0019683|T034||LNC|HIV ANTIBODY
C0019683|T034||LNC|HIV - HUMAN IMMUNODEFICIENCY VIRUS ANTIBODY
C0019683|T034||LNC|HUMAN IMMUNODEFICIENCY VIRUS ANTIBODY
C0019683|T034||LNC|HUMAN IMMUNODEFICIENCY VIRUS ANTIBODY 
C0019683|T034||LNC|HTLV-III ANTIBODY
C0474652|T034||LNC|HUMAN IMMUNODEFICIENCY VIRUS ANTIBODY TITER MEASUREMENT
C0474652|T034||LNC|HUMAN IMMUNODEFICIENCY VIRUS ANTIBODY LEVEL 
C0474652|T034||LNC|HUMAN IMMUNODEFICIENCY VIRUS ANTIBODY LEVEL
C0474652|T034||LNC|HUMAN IMMUNODEFICIENCY VIRUS ANTIBODY LEVEL 
C0474652|T034||LNC|HIV - HUMAN IMMUNODEFICIENCY VIRUS ANTIBODY TITER
C0474652|T034||LNC|HIV - HUMAN IMMUNODEFICIENCY VIRUS ANTIBODY TITRE
C0474652|T034||LNC|HUMAN IMMUNODEFICIENCY VIRUS ANTIBODY TITER
C0474652|T034||LNC|HUMAN IMMUNODEFICIENCY VIRUS ANTIBODY TITRE
C0474652|T034||LNC|HUMAN IMMUNODEFICIENCY VIRUS ANTIBODY TITER MEASUREMENT 
C0474652|T034||LNC|HUMAN IMMUNODEFICIENCY VIRUS ANTIBODY TITRE MEASUREMENT
C0474652|T034||LNC|HUMAN IMMUNODEFICIENCY VIRUS ANTIBODY ASSAY
C3181597|T034||LNC|4E10 MAB
C3181597|T034||LNC|MAB 4E10
C3181597|T034||LNC|4E10 MONOCLONAL ANTIBODY
C4043370|T034||LNC|I'M NOT SURE THIS IS A COMMON ANTIBODY USED IN THE ELISA, BUT I CAN'T IMAGINE YOU'D SEE IT IN A CHART IN ANY OTHER CONTEXT, SO I DONT HTINK IT WILL GENERATE NOISE
C0369497|T034|MTHU002639|LNC|HUMAN IMMUNODEFICIENCY VIRUS, TYPE I ANTIBODY|HIV 1 AB
C0369497|T034|MTHU002639|LNC|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 ANTIBODY|HIV 1 AB
C0369497|T034|MTHU002639|LNC|HIV 1 AB|HIV 1 AB
C0369497|T034|MTHU002639|LNC|HUMAN IMMUNODEFICIENCY VIRUS 1 ANTIBODY|HIV 1 AB
C0369497|T034|MTHU002639|LNC|HUMAN IMMUNODEFICIENCY VIRUS, TYPE I ANTIBODY |HIV 1 AB
C0369497|T034|MTHU002639|LNC|HIV-1 ANTIBODY|HIV 1 AB
C0369497|T034|MTHU002639|LNC|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 ANTIBODY |HIV 1 AB
C0369497|T034|MTHU002639|LNC|LAV-1 ANTIBODY|HIV 1 AB
C0369500|T034|MTHU010597|LNC|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 (HIV-2) ANTIBODY|HIV 2 AB
C0369500|T034|MTHU010597|LNC|HIV 2 AB|HIV 2 AB
C0369500|T034|MTHU010597|LNC|HUMAN IMMUNODEFICIENCY VIRUS 2 ANTIBODY|HIV 2 AB
C0369500|T034|MTHU010597|LNC|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 ANTIBODY|HIV 2 AB
C0369500|T034|MTHU010597|LNC|HUMAN IMMUNODEFICIENCY VIRUS, TYPE II ANTIBODY |HIV 2 AB
C0369500|T034|MTHU010597|LNC|HUMAN IMMUNODEFICIENCY VIRUS, TYPE II ANTIBODY|HIV 2 AB
C3714540|T034||LNC|HIV ANTIBODY
C3714540|T034||LNC|HIV ANTIBODY MEASUREMENT
C3714540|T034||LNC|HIVAB
