C2910651|T053||SNOMEDCT_US|UNKNOWN ROUTE OF HCV TRANSMISSION
C2910651|T053||SNOMEDCT_US|UNKNOWN ROUTE OF HCV INFECTION
C2910651|T053||SNOMEDCT_US|UNKNOWN ROUTE OF INFECTION
C2910651|T053||SNOMEDCT_US|CONTACT WITH AND (SUSPECTED) EXPOSURE TO VIRAL HEPATITIS
C2910651|T053||SNOMEDCT_US|CONTACT WITH VIRAL HEPATITIS
C2910651|T053||SNOMEDCT_US|CONTACT WITH HEPATITIS C VIRUS
C2910651|T053||SNOMEDCT_US|CONTACT WITH VIRAL HEPATITIS
C2910651|T053||SNOMEDCT_US|CONTACT WITH HCV
C2919618|T053|444563003|SNOMEDCT_US|EXPOSURE TO HCV|EXPOSURE TO HEPATITIS C VIRUS (EVENT)
C2919618|T053|444563003|SNOMEDCT_US|EXPOSURE TO HEPATITIS C|EXPOSURE TO HEPATITIS C VIRUS (EVENT)
C2919618|T053|444563003|SNOMEDCT_US|EXPOSURE TO HEPATITIS C VIRUS|EXPOSURE TO HEPATITIS C VIRUS (EVENT)
C2910651|T053||SNOMEDCT_US|CONTACT WITH AND (SUSPECTED) EXPOSURE TO VIRAL HEPATITIS
C1096517|T053||SNOMEDCT_US|EXPOSURE TO HEPATITIS C 
C1096517|T053||SNOMEDCT_US|EXPOSURE TO HEPATITIS C
C1096517|T053||SNOMEDCT_US|HEPATITIS C EXPOSURE
