C0035078|T047|156092003|SNOMEDCT_US|KIDNEY FAILURE|RENAL FAILURE (DISORDER)
C1565489|T047|236423003|SNOMEDCT_US|RENAL INSUFFICIENCY|RENAL DYSFUNCTION
C0022660|T047|14669001|SNOMEDCT_US|KIDNEY FAILURE, ACUTE|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|ACUTE RENAL FAILURE|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|ACUTE RENAL FAILURE, UNSPECIFIED|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|ARF|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|ACUTE RENAL FAILURE |ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|ARF (ACUTE RENAL FAILURE)|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|ACUTE KIDNEY FAILURE|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|ACUTE KIDNEY FAILURE NOS|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|ACUTE KIDNEY FAILURE, UNSPECIFIED|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|ACUTE AND UNSPECIFIED RENAL FAILURE|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|RENAL FAILURE, ACUTE|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|KIDNEY FAILURE, ACUTE [DISEASE/FINDING]|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|KIDNEY FAILURES, ACUTE|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|ACUTE KIDNEY FAILURES|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|ACUTE RENAL FAILURES|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|RENAL FAILURES, ACUTE|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|FAILURE;RENAL;ACUTE|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|ACUTE RENAL FAILURE NOS |ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|ACUTE RENAL FAILURE |ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|ACUTE RENAL FAILURE NOS|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|AKI|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|ACUTE KIDNEY INJURY|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|FAILURE KIDNEY ACUTE|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|KIDNEY FAILURE ACUTE|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|RENAL SHUTDOWN ACUTE|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|RENAL FAILURE ACUTE|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|ACUTE RENAL FAILURE SYNDROME|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|ARF - ACUTE RENAL FAILURE|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|ACUTE RENAL FAILURE SYNDROME |ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022660|T047|14669001|SNOMEDCT_US|ACUTE RENAL FAILURE SYNDROME, NOS|ACUTE RENAL FAILURE SYNDROME (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|KIDNEY FAILURE, CHRONIC|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|CHRONIC RENAL FAILURE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|DISEASE, END-STAGE KIDNEY|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|DISEASE, END-STAGE RENAL|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|END-STAGE RENAL FAILURE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|KIDNEY DISEASE, END-STAGE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|RENAL DISEASE, END STAGE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|RENAL FAILURE, END STAGE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|END STAGE KIDNEY DISEASE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|END STAGE RENAL DISEASE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|CRF|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|CHRONIC RENAL FAILURE, UNSPECIFIED|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|END-STAGE RENAL DISEASE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|END STAGE CHRONIC RENAL FAILURE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|END STAGE CHRONC RENAL FAILURE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|END STAGE KIDNEY DIS|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|RENAL DIS END STAGE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|END STAGE RENAL DIS|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|END STAGE RENAL FAILURE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|END STAGE RENAL DISEASE |END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|CHRONIC RENAL FAILURE |END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|ESRD (END STAGE RENAL DISEASE)|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|CRF - CHRONIC RENAL FAILURE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|CHRONIC RENAL DISEASE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|CHRONIC RENAL FAILURE NOS|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|END-STAGE KIDNEY DISEASE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|RENAL FAILURE, CHRONIC|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|ESRD|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|RENAL FAILURE, END-STAGE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|CHRONIC KIDNEY FAILURE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|KIDNEY FAILURE, CHRONIC [DISEASE/FINDING]|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|RENAL DISEASE, END-STAGE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|FAILURE;RENAL;CHRONIC|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|RENAL FAILURE - CHRONIC|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|RENAL FAILURE (CHRONIC)|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|END STAGE RENAL FAILURE |END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|FAILURE, RENAL -CHRONIC|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|CHRONIC RENAL FAILURE SYNDROME|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|KIDNEY FAILURE CHRONIC|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|END STAGE RENAL DISEASE (ESRD)|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|RENAL FAILURE CHRONIC|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|ESCRF - END STAGE CHRONIC RENAL FAILURE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|ESRD - END STAGE RENAL DISEASE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|ESRF - END STAGE RENAL FAILURE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|CHRONIC RENAL FAILURE SYNDROME |END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|END STAGE RENAL DISEASE |END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|DISEASE (OR DISORDER); KIDNEY, END-STAGE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|DISEASE (OR DISORDER); RENAL, END-STAGE|END STAGE RENAL FAILURE (DISORDER)
C0022661|T047|197755007|SNOMEDCT_US|CHRONIC RENAL FAILURE SYNDROME, NOS|END STAGE RENAL FAILURE (DISORDER)
C0041948|T047|44730006|SNOMEDCT_US|UREMIA OF RENAL ORIGIN|UREMIA (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|KIDNEY FAILURE|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|RENAL FAILURE|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|UNSPECIFIED RENAL FAILURE|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|RENAL FAILURE |RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|RENAL FAILURE NOS|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|UNSPECIFIED KIDNEY FAILURE|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|KIDNEY FAILURE [DISEASE/FINDING]|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|KIDNEY FAILURES|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|FAILURE, RENAL|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|FAILURE, KIDNEY|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|FAILURES, KIDNEY|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|FAILURES, RENAL|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|RENAL FAILURES|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|RENAL INSUFFICIENCY|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|ESRD|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|RENAL FAILURE UNSPECIFIED|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|RENAL FAILURE UNSPECIFIED |RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|RENAL FAILURE |RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|RENAL FAILURE SYNDROME|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|FAILURE KIDNEY|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|RENAL FAILURE, UNSPECIFIED|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|RENAL INSUFFICIENCY SYNDROME|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|RF - RENAL FAILURE|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|RENAL FAILURE SYNDROME |RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|FAILURE; RENAL|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|KIDNEY; FAILURE|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|RENAL; FAILURE|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|RENAL FAILURE SYNDROME, NOS|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|RENAL INSUFFICIENCY SYNDROME, NOS|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|RENAL FAILURE NOT OTHERWISE SPECIFIED|RENAL FAILURE (DISORDER)
C0035078|T047|156092003|SNOMEDCT_US|FAILURE;RENAL;NOS|RENAL FAILURE (DISORDER)
C0403462|T047|236433006|SNOMEDCT_US|ACUTE ON CHRONIC RENAL FAILURE|ACUTE-ON-CHRONIC RENAL FAILURE (DISORDER)
C0403462|T047|236433006|SNOMEDCT_US|RENAL FAILURE ACUTE ON CHRONIC|ACUTE-ON-CHRONIC RENAL FAILURE (DISORDER)
C0403462|T047|236433006|SNOMEDCT_US|ACUTE-ON-CHRONIC RENAL FAILURE |ACUTE-ON-CHRONIC RENAL FAILURE (DISORDER)
C0403462|T047|236433006|SNOMEDCT_US|ACUTE-ON-CHRONIC RENAL FAILURE|ACUTE-ON-CHRONIC RENAL FAILURE (DISORDER)
C2919930|T047|445120004|SNOMEDCT_US|URAEMIA DUE TO INADEQUATE RENAL PERFUSION|UREMIA DUE TO INADEQUATE RENAL PERFUSION (DISORDER)
C2919930|T047|445120004|SNOMEDCT_US|UREMIA DUE TO INADEQUATE RENAL PERFUSION |UREMIA DUE TO INADEQUATE RENAL PERFUSION (DISORDER)
C2919930|T047|445120004|SNOMEDCT_US|UREMIA DUE TO INADEQUATE RENAL PERFUSION|UREMIA DUE TO INADEQUATE RENAL PERFUSION (DISORDER)
C0574786|T047|298015003|SNOMEDCT_US|ACUTE RENAL FAILURE WITH MEDULLARY NECROSIS|ACUTE RENAL PAPILLARY NECROSIS WITH RENAL FAILURE (DISORDER)
C0574786|T047|298015003|SNOMEDCT_US|ACUTE KIDNEY FAILURE WITH MEDULLARY NECROSIS|ACUTE RENAL PAPILLARY NECROSIS WITH RENAL FAILURE (DISORDER)
C0574786|T047|298015003|SNOMEDCT_US|ACUTE RENAL FAILURE WITH LESION OF RENAL MEDULLARY (PAPILLARY) NECROSIS|ACUTE RENAL PAPILLARY NECROSIS WITH RENAL FAILURE (DISORDER)
C0574786|T047|298015003|SNOMEDCT_US|ACUTE RENAL PAPILLARY NECROSIS WITH RENAL FAILURE|ACUTE RENAL PAPILLARY NECROSIS WITH RENAL FAILURE (DISORDER)
C0574786|T047|298015003|SNOMEDCT_US|ACUTE RENAL PAPILLARY NECROSIS WITH RENAL FAILURE |ACUTE RENAL PAPILLARY NECROSIS WITH RENAL FAILURE (DISORDER)
C0574786|T047|298015003|SNOMEDCT_US|INSUFFICIENCY; RENAL, ACUTE, WITH NECROSIS, MEDULLARY, MEDULLARY|ACUTE RENAL PAPILLARY NECROSIS WITH RENAL FAILURE (DISORDER)
C0574786|T047|298015003|SNOMEDCT_US|KIDNEY; INSUFFICIENCY, ACUTE, WITH NECROSIS, MEDULLARY, MEDULLARY|ACUTE RENAL PAPILLARY NECROSIS WITH RENAL FAILURE (DISORDER)
C0574786|T047|298015003|SNOMEDCT_US|ACUTE RENAL FAILURE WITH RENAL PAPILLARY NECROSIS|ACUTE RENAL PAPILLARY NECROSIS WITH RENAL FAILURE (DISORDER)
C0574786|T047|298015003|SNOMEDCT_US|ACUTE RENAL FAILURE WITH LESION OF RENAL MEDULLARY NECROSIS|ACUTE RENAL PAPILLARY NECROSIS WITH RENAL FAILURE (DISORDER)
C0495124|T047||SNOMEDCT_US|POSTPROCEDURAL RENAL FAILURE
C0495124|T047||SNOMEDCT_US|POSTPROCEDURAL RENAL INSUFFICIENCY 
C0495124|T047||SNOMEDCT_US|POSTPROCEDURAL RENAL INSUFFICIENCY
C0495124|T047||SNOMEDCT_US|POSTPROCEDURAL RENAL FAILURE 
C0495124|T047||SNOMEDCT_US|INSUFFICIENCY; RENAL, POSTPROCEDURAL
C0495124|T047||SNOMEDCT_US|KIDNEY; INSUFFICIENCY, POSTPROCEDURAL
C0495124|T047||SNOMEDCT_US|NECROSIS; TUBULAR, POSTPROCEDURAL
C0495124|T047||SNOMEDCT_US|TUBULAR; NECROSIS, POSTPROCEDURAL
C0410932|T047|268854008|SNOMEDCT_US|CONGENITAL RENAL FAILURE|CONGENITAL RENAL FAILURE (DISORDER)
C0410932|T047|268854008|SNOMEDCT_US|RENAL FAILURE CONGENITAL|CONGENITAL RENAL FAILURE (DISORDER)
C0410932|T047|268854008|SNOMEDCT_US|CONGENITAL RENAL FAILURE |CONGENITAL RENAL FAILURE (DISORDER)
C0410932|T047|268854008|SNOMEDCT_US|CONGENITAL RENAL FAILURE |CONGENITAL RENAL FAILURE (DISORDER)
C0410932|T047|268854008|SNOMEDCT_US|INSUFFICIENCY; RENAL, CONGENITAL|CONGENITAL RENAL FAILURE (DISORDER)
C0410932|T047|268854008|SNOMEDCT_US|KIDNEY; INSUFFICIENCY, CONGENITAL|CONGENITAL RENAL FAILURE (DISORDER)
C2316810|T047|433146000|SNOMEDCT_US|ESRD|CKD STAGE 5
C2316810|T047|433146000|SNOMEDCT_US|END STAGE KIDNEY DISEASE|CKD STAGE 5
C2316810|T047|433146000|SNOMEDCT_US|END STAGE KIDNEY FAILURE|CKD STAGE 5
C2316810|T047|433146000|SNOMEDCT_US|END STAGE RENAL FAILURE|CKD STAGE 5
C2316810|T047|433146000|SNOMEDCT_US|CHRONIC KIDNEY DISEASE STAGE 5 |CKD STAGE 5
C2316810|T047|433146000|SNOMEDCT_US|CHRONIC KIDNEY DISEASE STAGE 5|CKD STAGE 5
C2316810|T047|433146000|SNOMEDCT_US|CHRONIC KIDNEY DISEASE STAGE 5 |CKD STAGE 5
C2316810|T047|433146000|SNOMEDCT_US|CHRONIC KIDNEY DISEASE, STAGE 5|CKD STAGE 5
C2316810|T047|433146000|SNOMEDCT_US|END STAGE RENAL DISEASE|CKD STAGE 5
C2316810|T047|433146000|SNOMEDCT_US|CKD STAGE 5|CKD STAGE 5
C2316810|T047|433146000|SNOMEDCT_US|END-STAGE RENAL DISEASE|CKD STAGE 5
C2316810|T047|433146000|SNOMEDCT_US|RENAL FAILURE, ENDSTAGE|CKD STAGE 5
C2316810|T047|433146000|SNOMEDCT_US|ESRD, END STAGE RENAL DISEASE|CKD STAGE 5
C2316810|T047|433146000|SNOMEDCT_US|RENAL DISEASE (ESRD), END STAGE|CKD STAGE 5
C2316810|T047|433146000|SNOMEDCT_US|RENAL DISEASE, END STAGE|CKD STAGE 5
C2316810|T047|433146000|SNOMEDCT_US|END STAGE RENAL DISEASE (ESRD)|CKD STAGE 5
C2316810|T047|433146000|SNOMEDCT_US|DISEASE (ESRD), END STAGE RENAL|CKD STAGE 5
C2316810|T047|433146000|SNOMEDCT_US|CHRONIC RENAL FAILURE|CKD STAGE 5
C2316810|T047|433146000|SNOMEDCT_US|STAGE 5 CHRONIC KIDNEY DISEASE|CKD STAGE 5
C2316810|T047|433146000|SNOMEDCT_US|END-STAGE RENAL FAILURE|CKD STAGE 5
C0404974|T047|198844003|SNOMEDCT_US|RENAL SHUTDOWN FOLLOWING ABORTIVE PREGNANCY |RENAL SHUTDOWN FOLLOWING ABORTIVE PREGNANCY (DISORDER)
C0404974|T047|198844003|SNOMEDCT_US|RENAL SHUTDOWN FOLLOWING ABORTIVE PREGNANCY|RENAL SHUTDOWN FOLLOWING ABORTIVE PREGNANCY (DISORDER)
C1534552|T047|266616000|SNOMEDCT_US|(RENAL FAILURE NOS) OR (URAEMIA NOS)|(RENAL FAILURE NOS) OR (URAEMIA NOS) (DISORDER)
C1534552|T047|266616000|SNOMEDCT_US|(RENAL FAILURE NOS) OR (UREMIA NOS)|(RENAL FAILURE NOS) OR (URAEMIA NOS) (DISORDER)
C1534552|T047|266616000|SNOMEDCT_US|(RENAL FAILURE NOS) OR (URAEMIA NOS) |(RENAL FAILURE NOS) OR (URAEMIA NOS) (DISORDER)
C1534552|T047|266616000|SNOMEDCT_US|(RENAL FAILURE UNSPECIFIED) OR (URAEMIA NOS) |(RENAL FAILURE NOS) OR (URAEMIA NOS) (DISORDER)
C1534552|T047|266616000|SNOMEDCT_US|(RENAL FAILURE UNSPECIFIED) OR (URAEMIA NOS)|(RENAL FAILURE NOS) OR (URAEMIA NOS) (DISORDER)
C1534552|T047|266616000|SNOMEDCT_US|(RENAL FAILURE UNSPECIFIED) OR (UREMIA NOS)|(RENAL FAILURE NOS) OR (URAEMIA NOS) (DISORDER)
C3662191|T047|609452007|SNOMEDCT_US|INDUCED TERMINATION OF PREGNANCY COMPLICATED BY RENAL FAILURE|INDUCED TERMINATION OF PREGNANCY COMPLICATED BY RENAL FAILURE (DISORDER)
C3662191|T047|609452007|SNOMEDCT_US|INDUCED TERMINATION OF PREGNANCY COMPLICATED BY RENAL FAILURE |INDUCED TERMINATION OF PREGNANCY COMPLICATED BY RENAL FAILURE (DISORDER)
C3662191|T047|609452007|SNOMEDCT_US|TERMINATION OF PREGNANCY COMPLICATED BY RENAL FAILURE|INDUCED TERMINATION OF PREGNANCY COMPLICATED BY RENAL FAILURE (DISORDER)
C1565662|T047|236424009|SNOMEDCT_US|ACUTE RENAL INSUFFICIENCY |ACUTE RENAL IMPAIRMENT (DISORDER)
C1565662|T047|236424009|SNOMEDCT_US|ACUTE RENAL INSUFFICIENCY|ACUTE RENAL IMPAIRMENT (DISORDER)
C1565662|T047|236424009|SNOMEDCT_US|RENAL INSUFFICIENCY (ACUTE)|ACUTE RENAL IMPAIRMENT (DISORDER)
C1565662|T047|236424009|SNOMEDCT_US|ACUTE RENAL INSUFFICIENCIES|ACUTE RENAL IMPAIRMENT (DISORDER)
C1565662|T047|236424009|SNOMEDCT_US|RENAL INSUFFICIENCIES, ACUTE|ACUTE RENAL IMPAIRMENT (DISORDER)
C1565662|T047|236424009|SNOMEDCT_US|KIDNEY INSUFFICIENCIES, ACUTE|ACUTE RENAL IMPAIRMENT (DISORDER)
C1565662|T047|236424009|SNOMEDCT_US|ACUTE KIDNEY INSUFFICIENCIES|ACUTE RENAL IMPAIRMENT (DISORDER)
C1565662|T047|236424009|SNOMEDCT_US|ACUTE KIDNEY INSUFFICIENCY|ACUTE RENAL IMPAIRMENT (DISORDER)
C1565662|T047|236424009|SNOMEDCT_US|RENAL INSUFFICIENCY, ACUTE|ACUTE RENAL IMPAIRMENT (DISORDER)
C1565662|T047|236424009|SNOMEDCT_US|KIDNEY INSUFFICIENCY, ACUTE|ACUTE RENAL IMPAIRMENT (DISORDER)
C1565662|T047|236424009|SNOMEDCT_US|ACUTE RENAL IMPAIRMENT|ACUTE RENAL IMPAIRMENT (DISORDER)
C1565662|T047|236424009|SNOMEDCT_US|ACUTE RENAL IMPAIRMENT |ACUTE RENAL IMPAIRMENT (DISORDER)
C1565662|T047|236424009|SNOMEDCT_US|INSUFFICIENCY; RENAL, ACUTE|ACUTE RENAL IMPAIRMENT (DISORDER)
C0588179|T047|310647000|SNOMEDCT_US|ANAEMIA SECONDARY TO RENAL FAILURE|ANEMIA SECONDARY TO RENAL FAILURE (DISORDER)
C0588179|T047|310647000|SNOMEDCT_US|ANEMIA SECONDARY TO RENAL FAILURE|ANEMIA SECONDARY TO RENAL FAILURE (DISORDER)
C0588179|T047|310647000|SNOMEDCT_US|ANAEMIA SECONDARY TO RENAL FAILURE |ANEMIA SECONDARY TO RENAL FAILURE (DISORDER)
C0588179|T047|310647000|SNOMEDCT_US|ANEMIA SECONDARY TO RENAL FAILURE |ANEMIA SECONDARY TO RENAL FAILURE (DISORDER)
C1565489|T047|236423003|SNOMEDCT_US|RENAL INSUFFICIENCY|RENAL DYSFUNCTION
C1565489|T047|236423003|SNOMEDCT_US|IMPAIRED RENAL FUNCTION|RENAL DYSFUNCTION
C1565489|T047|236423003|SNOMEDCT_US|RENAL INSUFFICIENCY |RENAL DYSFUNCTION
C1565489|T047|236423003|SNOMEDCT_US|RENAL INSUFFICIENCY [DISEASE/FINDING]|RENAL DYSFUNCTION
C1565489|T047|236423003|SNOMEDCT_US|KIDNEY INSUFFICIENCY|RENAL DYSFUNCTION
C1565489|T047|236423003|SNOMEDCT_US|INSUFFICIENCY;RENAL|RENAL DYSFUNCTION
C1565489|T047|236423003|SNOMEDCT_US|RENAL IMPAIRMENT |RENAL DYSFUNCTION
C1565489|T047|236423003|SNOMEDCT_US|RENAL IMPAIRMENT|RENAL DYSFUNCTION
C1565489|T047|236423003|SNOMEDCT_US|RENAL DYSFUNCTION|RENAL DYSFUNCTION
C1565489|T047|236423003|SNOMEDCT_US|KIDNEY IMPAIRMENT|RENAL DYSFUNCTION
C1565489|T047|236423003|SNOMEDCT_US|INSUFFICIENCY RENAL|RENAL DYSFUNCTION
C1565489|T047|236423003|SNOMEDCT_US|RENAL IMPAIRMENT NOS|RENAL DYSFUNCTION
C1565489|T047|236423003|SNOMEDCT_US|INSUFFICIENCY; RENAL|RENAL DYSFUNCTION
C1565489|T047|236423003|SNOMEDCT_US|KIDNEY; INSUFFICIENCY|RENAL DYSFUNCTION
C1565489|T047|236423003|SNOMEDCT_US|KIDNEY INSUFFICIENCIES|RENAL DYSFUNCTION
C1565489|T047|236423003|SNOMEDCT_US|RENAL INSUFFICIENCIES|RENAL DYSFUNCTION
C1565489|T047|236423003|SNOMEDCT_US|INSUFFICIENCY, KIDNEY|RENAL DYSFUNCTION
C4075836|T047|713696000|SNOMEDCT_US|RENAL FAILURE SYNDROME CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|RENAL FAILURE SYNDROME CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075836|T047|713696000|SNOMEDCT_US|RENAL FAILURE SYNDROME CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |RENAL FAILURE SYNDROME CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C0348879|T047|194780003|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE, UNSPECIFIED, WITH RENAL FAILURE|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348879|T047|194780003|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348879|T047|194780003|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE |HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348879|T047|194780003|SNOMEDCT_US|HYPERTENSIVE HEART AND CHRONIC KIDNEY DISEASE WITH RENAL FAILURE|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348879|T047|194780003|SNOMEDCT_US|HY HT/KD NOS ST V W/O HF|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348879|T047|194780003|SNOMEDCT_US|HYPERTENSIVE HEART AND CHRONIC KIDNEY DISEASE, UNSPECIFIED, WITHOUT HEART FAILURE AND WITH CHRONIC KIDNEY DISEASE STAGE V OR END STAGE RENAL DISEASE|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348879|T047|194780003|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE |HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348879|T047|194780003|SNOMEDCT_US|FAILURE; CARDIORENAL, HYPERTENSIVE, WITH RENAL FAILURE|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348879|T047|194780003|SNOMEDCT_US|INSUFFICIENCY; RENAL, WITH HYPERTENSIVE HEART DISEASE|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348879|T047|194780003|SNOMEDCT_US|KIDNEY; INSUFFICIENCY, WITH HYPERTENSIVE HEART DISEASE|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|HYPERTENSIVE RENAL DISEASE, UNSPECIFIED, WITH RENAL FAILURE|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|HYP KID NOS W CR KID V|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|HYPERTENSIVE CHRONIC KIDNEY DISEASE, UNSPECIFIED, WITH CHRONIC KIDNEY DISEASE STAGE V OR END STAGE RENAL DISEASE|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|HYPERTENSIVE KIDNEY DISEASE WITH RENAL FAILURE |HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|HYPERTENSIVE KIDNEY DISEASE WITH RENAL FAILURE|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE |HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|HYPERTENSION; RENAL DISEASE, HYPERTENSIVE, WITH RENAL FAILURE|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|INSUFFICIENCY; RENAL, CHRONIC, HYPERTENSIVE|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|INSUFFICIENCY; RENAL, WITH HYPERTENSION|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|KIDNEY; HYPERTENSION, WITH RENAL FAILURE|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0494576|T047|194781004|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE, UNSPECIFIED, WITH CONGESTIVE HEART FAILURE AND RENAL FAILURE|HYPERTENSIVE HEART AND RENAL DISEASE WITH BOTH (CONGESTIVE) HEART FAILURE AND RENAL FAILURE (DISORDER)
C0494576|T047|194781004|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE WITH BOTH (CONGESTIVE) HEART FAILURE AND RENAL FAILURE|HYPERTENSIVE HEART AND RENAL DISEASE WITH BOTH (CONGESTIVE) HEART FAILURE AND RENAL FAILURE (DISORDER)
C0494576|T047|194781004|SNOMEDCT_US|HYP HT/KD NOS ST V W HF|HYPERTENSIVE HEART AND RENAL DISEASE WITH BOTH (CONGESTIVE) HEART FAILURE AND RENAL FAILURE (DISORDER)
C0494576|T047|194781004|SNOMEDCT_US|HYPERTENSIVE HEART AND CHRONIC KIDNEY DISEASE, UNSPECIFIED, WITH HEART FAILURE AND CHRONIC KIDNEY DISEASE STAGE V OR END STAGE RENAL DISEASE|HYPERTENSIVE HEART AND RENAL DISEASE WITH BOTH (CONGESTIVE) HEART FAILURE AND RENAL FAILURE (DISORDER)
C0494576|T047|194781004|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE, UNSPECIFIED, WITH HEART FAILURE AND RENAL FAILURE|HYPERTENSIVE HEART AND RENAL DISEASE WITH BOTH (CONGESTIVE) HEART FAILURE AND RENAL FAILURE (DISORDER)
C0494576|T047|194781004|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE WITH BOTH (CONGESTIVE) HEART FAILURE AND RENAL FAILURE |HYPERTENSIVE HEART AND RENAL DISEASE WITH BOTH (CONGESTIVE) HEART FAILURE AND RENAL FAILURE (DISORDER)
C0494576|T047|194781004|SNOMEDCT_US|INSUFFICIENCY; RENAL, WITH HYPERTENSIVE HEART DISEASE AND HEART FAILURE|HYPERTENSIVE HEART AND RENAL DISEASE WITH BOTH (CONGESTIVE) HEART FAILURE AND RENAL FAILURE (DISORDER)
C0494576|T047|194781004|SNOMEDCT_US|KIDNEY; INSUFFICIENCY, WITH HYPERTENSIVE HEART DISEASE AND HEART FAILURE|HYPERTENSIVE HEART AND RENAL DISEASE WITH BOTH (CONGESTIVE) HEART FAILURE AND RENAL FAILURE (DISORDER)
C0403448|T047|269301005|SNOMEDCT_US|KIDNEY FAILURE AS A COMPLICATION OF CARE|RENAL FAILURE AS A COMPLICATION OF CARE (DISORDER)
C0403448|T047|269301005|SNOMEDCT_US|RENAL FAILURE AS A COMPLICATION OF CARE|RENAL FAILURE AS A COMPLICATION OF CARE (DISORDER)
C0403448|T047|269301005|SNOMEDCT_US|RENAL FAILURE AS A COMPLICATION OF CARE |RENAL FAILURE AS A COMPLICATION OF CARE (DISORDER)
C0404973|T047|198847005|SNOMEDCT_US|RENAL FAILURE FOLLOWING ABORTION|RENAL FAILURE NOS FOLLOWING ABORTIVE PREGNANCY (FINDING)
C0404973|T047|198847005|SNOMEDCT_US|RENAL FAILURE FOLLOWING ABORTION |RENAL FAILURE NOS FOLLOWING ABORTIVE PREGNANCY (FINDING)
C0404973|T047|198847005|SNOMEDCT_US|RENAL FAILURE NOS FOLLOWING ABORTIVE PREGNANCY|RENAL FAILURE NOS FOLLOWING ABORTIVE PREGNANCY (FINDING)
C0404973|T047|198847005|SNOMEDCT_US|RENAL FAILURE FOLLOWING ABORTIVE PREGNANCY|RENAL FAILURE NOS FOLLOWING ABORTIVE PREGNANCY (FINDING)
C0404973|T047|198847005|SNOMEDCT_US|RENAL FAILURE NOS FOLLOWING ABORTIVE PREGNANCY |RENAL FAILURE NOS FOLLOWING ABORTIVE PREGNANCY (FINDING)
C0404973|T047|198847005|SNOMEDCT_US|RENAL FAILURE NOS FOLLOWING ABORTIVE PREGNANCY |RENAL FAILURE NOS FOLLOWING ABORTIVE PREGNANCY (FINDING)
C0404973|T047|198847005|SNOMEDCT_US|RENAL FAILURE FOLLOWING ABORTIVE PREGNANCY |RENAL FAILURE NOS FOLLOWING ABORTIVE PREGNANCY (FINDING)
C0477745|T047|198525004|SNOMEDCT_US|OTHER ACUTE RENAL FAILURE|[X]OTHER ACUTE RENAL FAILURE (DISORDER)
C0477745|T047|198525004|SNOMEDCT_US|OTHER ACUTE KIDNEY FAILURE|[X]OTHER ACUTE RENAL FAILURE (DISORDER)
C0477745|T047|198525004|SNOMEDCT_US|[X]OTHER ACUTE RENAL FAILURE|[X]OTHER ACUTE RENAL FAILURE (DISORDER)
C0477745|T047|198525004|SNOMEDCT_US|OTHER ACUTE RENAL FAILURE |[X]OTHER ACUTE RENAL FAILURE (DISORDER)
C0477745|T047|198525004|SNOMEDCT_US|[X]OTHER ACUTE RENAL FAILURE |[X]OTHER ACUTE RENAL FAILURE (DISORDER)
C0477746|T047|198526003|SNOMEDCT_US|OTHER CHRONIC RENAL FAILURE|[X]OTHER CHRONIC RENAL FAILURE (DISORDER)
C0477746|T047|198526003|SNOMEDCT_US|[X]OTHER CHRONIC RENAL FAILURE|[X]OTHER CHRONIC RENAL FAILURE (DISORDER)
C0477746|T047|198526003|SNOMEDCT_US|[X]OTHER CHRONIC RENAL FAILURE |[X]OTHER CHRONIC RENAL FAILURE (DISORDER)
C0542211|T047|275408006|SNOMEDCT_US|POSTOPERATIVE RENAL FAILURE|POSTOPERATIVE RENAL FAILURE (DISORDER)
C0542211|T047|275408006|SNOMEDCT_US|POSTOPERATIVE RENAL FAILURE |POSTOPERATIVE RENAL FAILURE (DISORDER)
C0156556|T047|10123006|SNOMEDCT_US|UNSPECIFIED ABORTION COMPLICATED BY RENAL FAILURE|ABORTION COMPLICATED BY RENAL FAILURE (DISORDER)
C0156556|T047|10123006|SNOMEDCT_US|UNSPECIFIED TYPE OF ABORTION, UNSPECIFIED, COMPLICATED BY RENAL FAILURE|ABORTION COMPLICATED BY RENAL FAILURE (DISORDER)
C0156556|T047|10123006|SNOMEDCT_US|ABORTION COMPLICATED BY RENAL FAILURE |ABORTION COMPLICATED BY RENAL FAILURE (DISORDER)
C0156556|T047|10123006|SNOMEDCT_US|ABORTION COMPLICATED BY RENAL FAILURE|ABORTION COMPLICATED BY RENAL FAILURE (DISORDER)
C0156556|T047|10123006|SNOMEDCT_US|ABORTION WITH RENAL FAILURE|ABORTION COMPLICATED BY RENAL FAILURE (DISORDER)
C0156556|T047|10123006|SNOMEDCT_US|AB NOS W RENAL FAIL-UNSP|ABORTION COMPLICATED BY RENAL FAILURE (DISORDER)
C0156556|T047|10123006|SNOMEDCT_US|UNSPECIFIED ABORTION, COMPLICATED BY RENAL FAILURE, UNSPECIFIED|ABORTION COMPLICATED BY RENAL FAILURE (DISORDER)
C0156556|T047|10123006|SNOMEDCT_US|ABORTION COMPLICATED BY RENAL FAILURE |ABORTION COMPLICATED BY RENAL FAILURE (DISORDER)
C2931783|T047|109477002|SNOMEDCT_US|AI1G|LUBINSKY SYNDROME
C2931783|T047|109477002|SNOMEDCT_US|AMELOGENESIS IMPERFECTA, TYPE IG|LUBINSKY SYNDROME
C2931783|T047|109477002|SNOMEDCT_US|AMELOGENESIS IMPERFECTA NEPHROCALCINOSIS|LUBINSKY SYNDROME
C2931783|T047|109477002|SNOMEDCT_US|ENAMEL RENAL SYNDROME|LUBINSKY SYNDROME
C2931783|T047|109477002|SNOMEDCT_US|GENERALIZED ENAMEL HYPOPLASIA AND RENAL DYSFUNCTION|LUBINSKY SYNDROME
C2931783|T047|109477002|SNOMEDCT_US|ABSENT ENAMEL, NEPHROCALCINOSIS AND APPARENTLY NORMAL CALCIUM METABOLISM|LUBINSKY SYNDROME
C2931783|T047|109477002|SNOMEDCT_US|AMELOGENESIS IMPERFECTA, HYPOPLASTIC, AND NEPHROCALCINOSIS|LUBINSKY SYNDROME
C2931783|T047|109477002|SNOMEDCT_US|ENAMEL-RENAL SYNDROME|LUBINSKY SYNDROME
C2931783|T047|109477002|SNOMEDCT_US|AMELOGENESIS IMPERFECTA AND GINGIVAL FIBROMATOSIS SYNDROME|LUBINSKY SYNDROME
C2931783|T047|109477002|SNOMEDCT_US|AIGFS|LUBINSKY SYNDROME
C2931783|T047|109477002|SNOMEDCT_US|AMELOGENESIS IMPERFECTA, HYPOPLASTIC, WITH NEPHROCALCINOSIS|LUBINSKY SYNDROME
C2931783|T047|109477002|SNOMEDCT_US|ENAMEL-RENAL-GINGIVAL SYNDROME|LUBINSKY SYNDROME
C2931783|T047|109477002|SNOMEDCT_US|AMELOGENESIS IMPERFECTA AND NEPHROCALCINOSIS|LUBINSKY SYNDROME
C2931783|T047|109477002|SNOMEDCT_US|MCGIBBON LUBINSKY SYNDROME|LUBINSKY SYNDROME
C2931783|T047|109477002|SNOMEDCT_US|ENAMEL-RENAL SYNDROME |LUBINSKY SYNDROME
C2931783|T047|109477002|SNOMEDCT_US|LUBINSKY SYNDROME|LUBINSKY SYNDROME
C2931783|T047|109477002|SNOMEDCT_US|AMELOGENESIS IMPERFECTA, NEPHROCALCINOSIS AND IMPAIRED RENAL CONCENTRATION|LUBINSKY SYNDROME
C0269314|T047|43629001|SNOMEDCT_US|RENAL FAILURE FOLLOWING MOLAR AND/OR ECTOPIC PREGNANCY |RENAL FAILURE FOLLOWING MOLAR AND/OR ECTOPIC PREGNANCY (DISORDER)
C0269314|T047|43629001|SNOMEDCT_US|RENAL FAILURE FOLLOWING MOLAR AND/OR ECTOPIC PREGNANCY|RENAL FAILURE FOLLOWING MOLAR AND/OR ECTOPIC PREGNANCY (DISORDER)
C0269314|T047|43629001|SNOMEDCT_US|RENAL FAILURE FOLLOWING MOLAR OR ECTOPIC PREGNANCY|RENAL FAILURE FOLLOWING MOLAR AND/OR ECTOPIC PREGNANCY (DISORDER)
C1386521|T047||SNOMEDCT_US|WHILE "UREMIA" CAN BE CAUSED BY PRE/POST RENAL CAUSES, THESE SEVERE COMPLICATIONS LIKELY INDICATE RENAL FAILURE
C1386521|T047||SNOMEDCT_US|APHASIA; UREMIC
C1390022|T047||SNOMEDCT_US|BLINDNESS; UREMIC
C1390022|T047||SNOMEDCT_US|UREMIC; BLINDNESS
C0151567|T047|95569006|SNOMEDCT_US|COMA URAEMIC|UREMIC COMA (DISORDER)
C0151567|T047|95569006|SNOMEDCT_US|URAEMIC COMA|UREMIC COMA (DISORDER)
C0151567|T047|95569006|SNOMEDCT_US|COMA UREMIC|UREMIC COMA (DISORDER)
C0151567|T047|95569006|SNOMEDCT_US|UREMIC COMA|UREMIC COMA (DISORDER)
C0151567|T047|95569006|SNOMEDCT_US|UREMIC COMA |UREMIC COMA (DISORDER)
C0151567|T047|95569006|SNOMEDCT_US|COMA; UREMIC|UREMIC COMA (DISORDER)
C0151567|T047|95569006|SNOMEDCT_US|UREMIC; COMA|UREMIC COMA (DISORDER)
C0234540|T047|49255002|SNOMEDCT_US|UREMIC CONVULSION|UREMIC CONVULSION (FINDING)
C0234540|T047|49255002|SNOMEDCT_US|URAEMIC CONVULSION|UREMIC CONVULSION (FINDING)
C0234540|T047|49255002|SNOMEDCT_US|UREMIC CONVULSION |UREMIC CONVULSION (FINDING)
C0234540|T047|49255002|SNOMEDCT_US|CONVULSIONS; UREMIC|UREMIC CONVULSION (FINDING)
C0234540|T047|49255002|SNOMEDCT_US|UREMIC; CONVULSIONS|UREMIC CONVULSION (FINDING)
C0748288|T047||SNOMEDCT_US|DECOMPENSATION; RENAL
C0748288|T047||SNOMEDCT_US|KIDNEY; DECOMPENSATION
C1395122|T047||SNOMEDCT_US|DELIRIUM; UREMIC
C1395122|T047||SNOMEDCT_US|UREMIC; DELIRIUM
C1395967|T047||SNOMEDCT_US|DYSPNEA; UREMIC
C1395967|T047||SNOMEDCT_US|UREMIC; DYSPNEA
C0232807|T047|76114004|SNOMEDCT_US|DECREASED RENAL FUNCTION|DECREASED RENAL FUNCTION (FINDING)
C0232807|T047|76114004|SNOMEDCT_US|DECREASED KIDNEY FUNCTION|DECREASED RENAL FUNCTION (FINDING)
C0232807|T047|76114004|SNOMEDCT_US|FUNCTION KIDNEY DECREASED|DECREASED RENAL FUNCTION (FINDING)
C0232807|T047|76114004|SNOMEDCT_US|DECREASED RENAL FUNCTION |DECREASED RENAL FUNCTION (FINDING)
C0232807|T047|76114004|SNOMEDCT_US|FUNCTION; LOW, KIDNEY|DECREASED RENAL FUNCTION (FINDING)
C0232807|T047|76114004|SNOMEDCT_US|LOW; FUNCTION, KIDNEY|DECREASED RENAL FUNCTION (FINDING)
C0151746|T047|39539005|SNOMEDCT_US|ABNORMAL RENAL FUNCTION|ABNORMAL RENAL FUNCTION (FINDING)
C0151746|T047|39539005|SNOMEDCT_US|RENAL FUNCTIONAL ABNORMALITY|ABNORMAL RENAL FUNCTION (FINDING)
C0151746|T047|39539005|SNOMEDCT_US|ABNORMAL RENAL PHYSIOLOGY|ABNORMAL RENAL FUNCTION (FINDING)
C0151746|T047|39539005|SNOMEDCT_US|ABNORMALITY OF RENAL PHYSIOLOGY|ABNORMAL RENAL FUNCTION (FINDING)
C0151746|T047|39539005|SNOMEDCT_US|DYSFUNCTION KIDNEY|ABNORMAL RENAL FUNCTION (FINDING)
C0151746|T047|39539005|SNOMEDCT_US|RENAL FUNCTION ABNORMAL|ABNORMAL RENAL FUNCTION (FINDING)
C0151746|T047|39539005|SNOMEDCT_US|FUNCTION KIDNEY ABNORMAL|ABNORMAL RENAL FUNCTION (FINDING)
C0151746|T047|39539005|SNOMEDCT_US|KIDNEY DYSFUNCTION|ABNORMAL RENAL FUNCTION (FINDING)
C0151746|T047|39539005|SNOMEDCT_US|KIDNEY FUNCTION ABNORMAL|ABNORMAL RENAL FUNCTION (FINDING)
C0151746|T047|39539005|SNOMEDCT_US|ABNORMAL RENAL FUNCTION |ABNORMAL RENAL FUNCTION (FINDING)
C0151746|T047|39539005|SNOMEDCT_US|DYSFUNCTION; KIDNEY|ABNORMAL RENAL FUNCTION (FINDING)
C1401758|T047||SNOMEDCT_US|FEVER; UREMIC
C1401758|T047||SNOMEDCT_US|UREMIC; FEVER
C1408265|T047||SNOMEDCT_US|KIDNEY; FUNCTIONAL DISTURBANCE
C0232808|T047|155876003|SNOMEDCT_US|NONFUNCTIONING KIDNEY |NON-FUNCTIONING KIDNEY (DISORDER)
C0232808|T047|155876003|SNOMEDCT_US|NONFUNCTIONING KIDNEY|NON-FUNCTIONING KIDNEY (DISORDER)
C0232808|T047|155876003|SNOMEDCT_US|NON-FUNCTIONING KIDNEY|NON-FUNCTIONING KIDNEY (DISORDER)
C0232808|T047|155876003|SNOMEDCT_US|NON-FUNCTIONING KIDNEY |NON-FUNCTIONING KIDNEY (DISORDER)
C0232808|T047|155876003|SNOMEDCT_US|NFK - NON-FUNCTIONING KIDNEY|NON-FUNCTIONING KIDNEY (DISORDER)
C0232808|T047|155876003|SNOMEDCT_US|SHUTDOWN RENAL|NON-FUNCTIONING KIDNEY (DISORDER)
C0232808|T047|155876003|SNOMEDCT_US|ABSENT RENAL FUNCTION|NON-FUNCTIONING KIDNEY (DISORDER)
C0232808|T047|155876003|SNOMEDCT_US|KIDNEY; NONFUNCTIONING|NON-FUNCTIONING KIDNEY (DISORDER)
C0232808|T047|155876003|SNOMEDCT_US|NONFUNCTIONING; KIDNEY|NON-FUNCTIONING KIDNEY (DISORDER)
C0232808|T047|155876003|SNOMEDCT_US|ABSENT RENAL FUNCTION |NON-FUNCTIONING KIDNEY (DISORDER)
C0232808|T047|155876003|SNOMEDCT_US|ABSENT RENAL FUNCTION |NON-FUNCTIONING KIDNEY (DISORDER)
C1407023|T047||SNOMEDCT_US|KIDNEY; TOXEMIA
C1407023|T047||SNOMEDCT_US|TOXEMIA; KIDNEY
C1406177|T047||SNOMEDCT_US|RENAL; SUPPRESSION
C1406177|T047||SNOMEDCT_US|SUPPRESSION; RENAL
C1407025|T047||SNOMEDCT_US|TOXEMIA; UREMIC
C1407025|T047||SNOMEDCT_US|UREMIC; TOXEMIA
C1407026|T047||SNOMEDCT_US|TOXEMIA; URINARY
C1407026|T047||SNOMEDCT_US|URINARY; TOXEMIA
C0235446|T047|371019009|SNOMEDCT_US|AZOTEMIA DUE TO INTRARENAL DISEASE|INTRARENAL AZOTEMIA
C0235446|T047|371019009|SNOMEDCT_US|RENAL AZOTEMIA|INTRARENAL AZOTEMIA
C0235446|T047|371019009|SNOMEDCT_US|RENAL AZOTEMIA |INTRARENAL AZOTEMIA
C0235446|T047|371019009|SNOMEDCT_US|INTRARENAL AZOTEMIA|INTRARENAL AZOTEMIA
C0235446|T047|371019009|SNOMEDCT_US|AZOTAEMIA DUE TO INTRARENAL DISEASE|INTRARENAL AZOTEMIA
C0235446|T047|371019009|SNOMEDCT_US|AZOTEMIA DUE TO INTRARENAL DISEASE |INTRARENAL AZOTEMIA
C0235446|T047|371019009|SNOMEDCT_US|INTRARENAL AZOTAEMIA|INTRARENAL AZOTEMIA
C0235446|T047|371019009|SNOMEDCT_US|RENAL AZOTAEMIA|INTRARENAL AZOTEMIA
C0235446|T047|371019009|SNOMEDCT_US|AZOTEMIA RENAL|INTRARENAL AZOTEMIA
C0235446|T047|371019009|SNOMEDCT_US|AZOTAEMIA RENAL|INTRARENAL AZOTEMIA
C0235446|T047|371019009|SNOMEDCT_US|AZOTEMIA OF RENAL ORIGIN|INTRARENAL AZOTEMIA
C0235446|T047|371019009|SNOMEDCT_US|AZOTAEMIA OF RENAL ORIGIN|INTRARENAL AZOTEMIA
C1278220|T047|144426008|SNOMEDCT_US|DETERIORATING RENAL FUNCTION|DETERIORATING RENAL FUNCTION (SITUATION)
C1278220|T047|144426008|SNOMEDCT_US|DETERIORATING RENAL FUNCTION |DETERIORATING RENAL FUNCTION (SITUATION)
C1278220|T047|144426008|SNOMEDCT_US|DETERIORATING RENAL FUNCTION |DETERIORATING RENAL FUNCTION (SITUATION)
C0456040|T047|276583007|SNOMEDCT_US|NEWBORN RENAL DYSFUNCTION|NEWBORN RENAL DYSFUNCTION (DISORDER)
C0456040|T047|276583007|SNOMEDCT_US|NEWBORN RENAL DYSFUNCTION |NEWBORN RENAL DYSFUNCTION (DISORDER)
C0403447|T047|236425005|SNOMEDCT_US|CHRONIC RENAL INSUFFICIENCY|CHRONIC RENAL IMPAIRMENT (DISORDER)
C0403447|T047|236425005|SNOMEDCT_US|CHRONIC RENAL INSUFFICIENCY |CHRONIC RENAL IMPAIRMENT (DISORDER)
C0403447|T047|236425005|SNOMEDCT_US|CHRONIC KIDNEY INSUFFICIENCY|CHRONIC RENAL IMPAIRMENT (DISORDER)
C0403447|T047|236425005|SNOMEDCT_US|RENAL INSUFFICIENCY, CHRONIC|CHRONIC RENAL IMPAIRMENT (DISORDER)
C0403447|T047|236425005|SNOMEDCT_US|RENAL INSUFFICIENCY, CHRONIC [DISEASE/FINDING]|CHRONIC RENAL IMPAIRMENT (DISORDER)
C0403447|T047|236425005|SNOMEDCT_US|KIDNEY INSUFFICIENCY, CHRONIC|CHRONIC RENAL IMPAIRMENT (DISORDER)
C0403447|T047|236425005|SNOMEDCT_US|CHRONIC RENAL IMPAIRMENT|CHRONIC RENAL IMPAIRMENT (DISORDER)
C0403447|T047|236425005|SNOMEDCT_US|CHRONIC RENAL IMPAIRMENT |CHRONIC RENAL IMPAIRMENT (DISORDER)
C0403447|T047|236425005|SNOMEDCT_US|INSUFFICIENCY; RENAL, CHRONIC, END STAGE RENAL DISEASE|CHRONIC RENAL IMPAIRMENT (DISORDER)
C0403447|T047|236425005|SNOMEDCT_US|INSUFFICIENCY; RENAL, CHRONIC|CHRONIC RENAL IMPAIRMENT (DISORDER)
C0403447|T047|236425005|SNOMEDCT_US|INSUFFICIENCY; RENAL, END STAGE|CHRONIC RENAL IMPAIRMENT (DISORDER)
C0403447|T047|236425005|SNOMEDCT_US|KIDNEY; INSUFFICIENCY, CHRONIC|CHRONIC RENAL IMPAIRMENT (DISORDER)
C0403447|T047|236425005|SNOMEDCT_US|CHRONIC KIDNEY INSUFFICIENCIES|CHRONIC RENAL IMPAIRMENT (DISORDER)
C0403447|T047|236425005|SNOMEDCT_US|CHRONIC RENAL INSUFFICIENCIES|CHRONIC RENAL IMPAIRMENT (DISORDER)
C0403447|T047|236425005|SNOMEDCT_US|KIDNEY INSUFFICIENCIES, CHRONIC|CHRONIC RENAL IMPAIRMENT (DISORDER)
C0403447|T047|236425005|SNOMEDCT_US|RENAL INSUFFICIENCIES, CHRONIC|CHRONIC RENAL IMPAIRMENT (DISORDER)
C0585398|T047|307532008|SNOMEDCT_US|ACUTE-ON-CHRONIC RENAL IMPAIRMENT |ACUTE-ON-CHRONIC RENAL IMPAIRMENT (DISORDER)
C0585398|T047|307532008|SNOMEDCT_US|ACUTE-ON-CHRONIC RENAL IMPAIRMENT|ACUTE-ON-CHRONIC RENAL IMPAIRMENT (DISORDER)
C2242703|T047|445236007|SNOMEDCT_US|CARDIORENAL SYNDROME|CARDIORENAL SYNDROME (DISORDER)
C2242703|T047|445236007|SNOMEDCT_US|CARDIORENAL SYNDROME |CARDIORENAL SYNDROME (DISORDER)
C2242703|T047|445236007|SNOMEDCT_US|CARDIO-RENAL SYNDROMES|CARDIORENAL SYNDROME (DISORDER)
C2242703|T047|445236007|SNOMEDCT_US|SYNDROME, RENOCARDIAC|CARDIORENAL SYNDROME (DISORDER)
C2242703|T047|445236007|SNOMEDCT_US|SYNDROME, CARDIORENAL|CARDIORENAL SYNDROME (DISORDER)
C2242703|T047|445236007|SNOMEDCT_US|CARDIO-RENAL SYNDROME|CARDIORENAL SYNDROME (DISORDER)
C2242703|T047|445236007|SNOMEDCT_US|SYNDROME, CARDIO-RENAL|CARDIORENAL SYNDROME (DISORDER)
C2242703|T047|445236007|SNOMEDCT_US|SYNDROMES, CARDIO-RENAL|CARDIORENAL SYNDROME (DISORDER)
C2242703|T047|445236007|SNOMEDCT_US|CARDIORENAL SYNDROMES|CARDIORENAL SYNDROME (DISORDER)
C2242703|T047|445236007|SNOMEDCT_US|SYNDROMES, CARDIORENAL|CARDIORENAL SYNDROME (DISORDER)
C2242703|T047|445236007|SNOMEDCT_US|RENO-CARDIAC SYNDROMES|CARDIORENAL SYNDROME (DISORDER)
C2242703|T047|445236007|SNOMEDCT_US|SYNDROMES, RENOCARDIAC|CARDIORENAL SYNDROME (DISORDER)
C2242703|T047|445236007|SNOMEDCT_US|CARDIO RENAL SYNDROME|CARDIORENAL SYNDROME (DISORDER)
C2242703|T047|445236007|SNOMEDCT_US|RENOCARDIAC SYNDROMES|CARDIORENAL SYNDROME (DISORDER)
C2242703|T047|445236007|SNOMEDCT_US|RENO CARDIAC SYNDROME|CARDIORENAL SYNDROME (DISORDER)
C2242703|T047|445236007|SNOMEDCT_US|SYNDROME, RENO-CARDIAC|CARDIORENAL SYNDROME (DISORDER)
C2242703|T047|445236007|SNOMEDCT_US|SYNDROMES, RENO-CARDIAC|CARDIORENAL SYNDROME (DISORDER)
C2242703|T047|445236007|SNOMEDCT_US|RENO-CARDIAC SYNDROME|CARDIORENAL SYNDROME (DISORDER)
C2242703|T047|445236007|SNOMEDCT_US|CARDIO-RENAL SYNDROME [DISEASE/FINDING]|CARDIORENAL SYNDROME (DISORDER)
C2242703|T047|445236007|SNOMEDCT_US|RENOCARDIAC SYNDROME|CARDIORENAL SYNDROME (DISORDER)
C1859722|T047|720513002|SNOMEDCT_US|ARC SYNDROME|ARTHROGRYPOSIS WITH RENAL DYSFUNCTION AND CHOLESTASIS SYNDROME (DISORDER)
C1859722|T047|720513002|SNOMEDCT_US|ARTHROGRYPOSIS RENAL DYSFUNCTION CHOLESTASIS SYNDROME|ARTHROGRYPOSIS WITH RENAL DYSFUNCTION AND CHOLESTASIS SYNDROME (DISORDER)
C1859722|T047|720513002|SNOMEDCT_US|ARTHROGRYPOSIS MULTIPLEX CONGENITA, RENAL DYSFUNCTION, AND CHOLESTASIS|ARTHROGRYPOSIS WITH RENAL DYSFUNCTION AND CHOLESTASIS SYNDROME (DISORDER)
C1859722|T047|720513002|SNOMEDCT_US|ARCS1|ARTHROGRYPOSIS WITH RENAL DYSFUNCTION AND CHOLESTASIS SYNDROME (DISORDER)
C1859722|T047|720513002|SNOMEDCT_US|ARTHROGRYPOSIS, RENAL DYSFUNCTION, AND CHOLESTASIS 1|ARTHROGRYPOSIS WITH RENAL DYSFUNCTION AND CHOLESTASIS SYNDROME (DISORDER)
C1859722|T047|720513002|SNOMEDCT_US|ARTHROGRYPOSIS, RENAL DYSFUNCTION, AND CHOLESTASIS|ARTHROGRYPOSIS WITH RENAL DYSFUNCTION AND CHOLESTASIS SYNDROME (DISORDER)
C1852759|T047|446449009|SNOMEDCT_US|PAPILLORENAL SYNDROME|RENAL COLOBOMA SYNDROME (DISORDER)
C1852759|T047|446449009|SNOMEDCT_US|OPTIC NERVE COLOBOMA WITH RENAL DISEASE|RENAL COLOBOMA SYNDROME (DISORDER)
C1852759|T047|446449009|SNOMEDCT_US|COLOBOMA OF OPTIC NERVE WITH RENAL DISEASE|RENAL COLOBOMA SYNDROME (DISORDER)
C1852759|T047|446449009|SNOMEDCT_US|RENAL-COLOBOMA SYNDROME|RENAL COLOBOMA SYNDROME (DISORDER)
C1852759|T047|446449009|SNOMEDCT_US|OPTIC COLOBOMA, VESICOURETERAL REFLUX, AND RENAL ANOMALIES|RENAL COLOBOMA SYNDROME (DISORDER)
C1852759|T047|446449009|SNOMEDCT_US|RENAL COLOBOMA SYNDROME |RENAL COLOBOMA SYNDROME (DISORDER)
C1852759|T047|446449009|SNOMEDCT_US|RENAL COLOBOMA SYNDROME|RENAL COLOBOMA SYNDROME (DISORDER)
C1852759|T047|446449009|SNOMEDCT_US|RENAL-COLOBOMA SYNDROME WITH MACULAR ABNORMALITIES|RENAL COLOBOMA SYNDROME (DISORDER)
C1852759|T047|446449009|SNOMEDCT_US|OPTIC NERVE COLOBOMA RENAL SYNDROME|RENAL COLOBOMA SYNDROME (DISORDER)
C1852759|T047|446449009|SNOMEDCT_US|COLOBOMA-URETERAL-RENAL SYNDROME|RENAL COLOBOMA SYNDROME (DISORDER)
C1852759|T047|446449009|SNOMEDCT_US|PAPRS|RENAL COLOBOMA SYNDROME (DISORDER)
C1852759|T047|446449009|SNOMEDCT_US|CONGENITAL ANOMALIES OF THE KIDNEY AND URINARY TRACT WITH OR WITHOUT OCULAR ABNORMALITIES|RENAL COLOBOMA SYNDROME (DISORDER)
C1852759|T047|446449009|SNOMEDCT_US|CAKUT WITH OR WITHOUT OCULAR ABNORMALITIES|RENAL COLOBOMA SYNDROME (DISORDER)
C0400972|T047|235914003|SNOMEDCT_US|BILIARY MALFORMATION WITH RENAL TUBULAR INSUFFICIENCY|BILIARY MALFORMATION ASSOCIATED WITH RENAL TUBULAR INSUFFICIENCY (DISORDER)
C0400972|T047|235914003|SNOMEDCT_US|CHOLESTATIC JAUNDICE AND RENAL TUBULAR INSUFFICIENCY|BILIARY MALFORMATION ASSOCIATED WITH RENAL TUBULAR INSUFFICIENCY (DISORDER)
C0400972|T047|235914003|SNOMEDCT_US|LUTZ RICHNER LANDOLT SYNDROME|BILIARY MALFORMATION ASSOCIATED WITH RENAL TUBULAR INSUFFICIENCY (DISORDER)
C0400972|T047|235914003|SNOMEDCT_US|RENAL TUBULAR INSUFFICIENCY, CHOLESTATIC JAUNDICE, AND MULTIPLE CONGENITAL ANOMALIES|BILIARY MALFORMATION ASSOCIATED WITH RENAL TUBULAR INSUFFICIENCY (DISORDER)
C0400972|T047|235914003|SNOMEDCT_US|BILIARY MALFORMATION ASSOCIATED WITH RENAL TUBULAR INSUFFICIENCY|BILIARY MALFORMATION ASSOCIATED WITH RENAL TUBULAR INSUFFICIENCY (DISORDER)
C0400972|T047|235914003|SNOMEDCT_US|BILIARY MALFORMATION ASSOCIATED WITH RENAL TUBULAR INSUFFICIENCY |BILIARY MALFORMATION ASSOCIATED WITH RENAL TUBULAR INSUFFICIENCY (DISORDER)
C2609414|T047|14350001000004108|SNOMEDCT_US|ACUTE KIDNEY INJURY|ACUTE INJURY OF KIDNEY (DISORDER)
C2609414|T047|14350001000004108|SNOMEDCT_US|ACUTE RENAL INJURIES|ACUTE INJURY OF KIDNEY (DISORDER)
C2609414|T047|14350001000004108|SNOMEDCT_US|RENAL INJURY, ACUTE|ACUTE INJURY OF KIDNEY (DISORDER)
C2609414|T047|14350001000004108|SNOMEDCT_US|ACUTE KIDNEY INJURIES|ACUTE INJURY OF KIDNEY (DISORDER)
C2609414|T047|14350001000004108|SNOMEDCT_US|RENAL INJURIES, ACUTE|ACUTE INJURY OF KIDNEY (DISORDER)
C2609414|T047|14350001000004108|SNOMEDCT_US|KIDNEY INJURY, ACUTE|ACUTE INJURY OF KIDNEY (DISORDER)
C2609414|T047|14350001000004108|SNOMEDCT_US|KIDNEY INJURIES, ACUTE|ACUTE INJURY OF KIDNEY (DISORDER)
C2609414|T047|14350001000004108|SNOMEDCT_US|ACUTE KIDNEY INJURY [DISEASE/FINDING]|ACUTE INJURY OF KIDNEY (DISORDER)
C2609414|T047|14350001000004108|SNOMEDCT_US|ACUTE RENAL INJURY|ACUTE INJURY OF KIDNEY (DISORDER)
C2609414|T047|14350001000004108|SNOMEDCT_US|ACUTE INJURY OF KIDNEY|ACUTE INJURY OF KIDNEY (DISORDER)
C2609414|T047|14350001000004108|SNOMEDCT_US|ACUTE INJURY OF KIDNEY |ACUTE INJURY OF KIDNEY (DISORDER)
C0403361|T047|197671004|SNOMEDCT_US|RENAL INSUFFICIENCY WITH GROWTH FAILURE|RENAL FUNCTION IMPAIRMENT WITH GROWTH FAILURE (DISORDER)
C0403361|T047|197671004|SNOMEDCT_US|RENAL INSUFFICIENCY WITH GROWTH FAILURE |RENAL FUNCTION IMPAIRMENT WITH GROWTH FAILURE (DISORDER)
C0403361|T047|197671004|SNOMEDCT_US|RENAL FUNCTION IMPAIRMENT WITH GROWTH FAILURE|RENAL FUNCTION IMPAIRMENT WITH GROWTH FAILURE (DISORDER)
C0403361|T047|197671004|SNOMEDCT_US|RENAL FUNCTION IMPAIRMENT WITH GROWTH FAILURE |RENAL FUNCTION IMPAIRMENT WITH GROWTH FAILURE (DISORDER)
C0403720|T047|236713006|SNOMEDCT_US|NEPHROLITHIASIS, X-LINKED RECESSIVE, WITH RENAL FAILURE|X-LINKED RECESSIVE NEPHROLITHIASIS WITH RENAL FAILURE (DISORDER)
C0403720|T047|236713006|SNOMEDCT_US|NPHL1|X-LINKED RECESSIVE NEPHROLITHIASIS WITH RENAL FAILURE (DISORDER)
C0403720|T047|236713006|SNOMEDCT_US|X-LINKED RECESSIVE NEPHROLITHIASIS WITH RENAL FAILURE|X-LINKED RECESSIVE NEPHROLITHIASIS WITH RENAL FAILURE (DISORDER)
C0403720|T047|236713006|SNOMEDCT_US|NEPHROLITHIASIS 1|X-LINKED RECESSIVE NEPHROLITHIASIS WITH RENAL FAILURE (DISORDER)
C0403720|T047|236713006|SNOMEDCT_US|NEPHROLITHIASIS, X-LINKED RECESSIVE, TYPE 1|X-LINKED RECESSIVE NEPHROLITHIASIS WITH RENAL FAILURE (DISORDER)
C0403720|T047|236713006|SNOMEDCT_US|UROLITHIASIS, X-LINKED RECESSIVE, TYPE 1|X-LINKED RECESSIVE NEPHROLITHIASIS WITH RENAL FAILURE (DISORDER)
C0403720|T047|236713006|SNOMEDCT_US|X-LINKED RECESSIVE NEPHROLITHIASIS WITH RENAL FAILURE |X-LINKED RECESSIVE NEPHROLITHIASIS WITH RENAL FAILURE (DISORDER)
C2751310|T047||SNOMEDCT_US|HNFJ2
C2751310|T047||SNOMEDCT_US|HYPERURICEMIC NEPHROPATHY, FAMILIAL JUVENILE, 2
C2751310|T047||SNOMEDCT_US|EARLY-ONSET HYPERURICEMIA, ANEMIA, AND PROGRESSIVE KIDNEY FAILURE
C2751310|T047||SNOMEDCT_US|HYPERURICEMIC NEPHROPATHY, FAMILIAL JUVENILE 2
C2751310|T047||SNOMEDCT_US|FAMILIAL JUVENILE HYPERURICEMIC NEPHROPATHY 2
C2751310|T047||SNOMEDCT_US|REN-RELATED KIDNEY DISEASE
C3854173|T047|129561000119108|SNOMEDCT_US|PRE-RENAL ACUTE KIDNEY INJURY |PRE-RENAL ACUTE KIDNEY INJURY (DISORDER)
C3854173|T047|129561000119108|SNOMEDCT_US|PRERENAL RENAL FAILURE|PRE-RENAL ACUTE KIDNEY INJURY (DISORDER)
C3854173|T047|129561000119108|SNOMEDCT_US|ACUTE RENAL FAILURE|PRE-RENAL ACUTE KIDNEY INJURY (DISORDER)
C3854173|T047|129561000119108|SNOMEDCT_US|PRE-RENAL ACUTE KIDNEY INJURY|PRE-RENAL ACUTE KIDNEY INJURY (DISORDER)
C1839604|T047||SNOMEDCT_US|RENAL FAILURE IN ADULTHOOD
C1561643|T047|709044004|SNOMEDCT_US|CHRONIC RENAL DISEASE|CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|CHRONIC KIDNEY DISEASE|CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|CHRONIC KIDNEY DIS NOS|CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|CKD - CHRONIC KIDNEY DISEASE|CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|CHRONIC KIDNEY DISEASE (CKD)|CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|CHRONIC KIDNEY DISEASE, UNSPECIFIED|CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|DISEASE, CHRONIC KIDNEY|CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|DISEASES, CHRONIC RENAL|CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|KIDNEY DISEASES, CHRONIC|CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|DISEASE, CHRONIC RENAL|CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|DISEASES, CHRONIC KIDNEY|CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|RENAL DISEASE, CHRONIC|CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|KIDNEY DISEASE, CHRONIC|CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|RENAL DISEASES, CHRONIC|CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|CKD|CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|CHRONIC KIDNEY DISEASES|CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|CHRONIC RENAL INSUFFICIENCY|CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|LOSS OF RENAL FUNCTION|CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|CHRONIC KIDNEY DISEASE |CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|CHRONIC RENAL FAILURE|CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|CHRONIC RENAL DISEASES|CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|DISEASE (OR DISORDER); KIDNEY, CHRONIC|CKD - CHRONIC KIDNEY DISEASE
C1561643|T047|709044004|SNOMEDCT_US|KIDNEY; DISEASE, CHRONIC|CKD - CHRONIC KIDNEY DISEASE
C1843276|T047||SNOMEDCT_US|RENAL FAILURE, REVERSIBLE
C1843276|T047||SNOMEDCT_US|REVERSIBLE RENAL FAILURE
C0184571|T047|130948000|SNOMEDCT_US|IMPAIRED KIDNEY FUNCTION|RENAL ALTERATION (FINDING)
C4076161|T047|713453003|SNOMEDCT_US|RENAL IMPAIRMENT CAUSED BY POLYOMAVIRUS |RENAL IMPAIRMENT CAUSED BY POLYOMAVIRUS (DISORDER)
C4076161|T047|713453003|SNOMEDCT_US|RENAL IMPAIRMENT CAUSED BY POLYOMAVIRUS|RENAL IMPAIRMENT CAUSED BY POLYOMAVIRUS (DISORDER)
C1285418|T047|363287001|SNOMEDCT_US|RENAL FAILURE ASSOCIATED WITH RENAL VASCULAR DISEASE |RENAL FAILURE ASSOCIATED WITH RENAL VASCULAR DISEASE (DISORDER)
C1285418|T047|363287001|SNOMEDCT_US|RENAL FAILURE ASSOCIATED WITH RENAL VASCULAR DISEASE|RENAL FAILURE ASSOCIATED WITH RENAL VASCULAR DISEASE (DISORDER)
