C0338831|T048|231494001|SNOMEDCT_US|MANIC|MANIA (DISORDER)
C0241934|T048|281257007|SNOMEDCT_US|HYPOMANIA|HYPOMANIC MOOD (FINDING)
C0154436|T048|191658009|SNOMEDCT_US|ATYPICAL MANIC DISORDER|ATYPICAL MANIC DISORDER (DISORDER)
C0154436|T048|191658009|SNOMEDCT_US|ATYPICAL MANIC DISORDER |ATYPICAL MANIC DISORDER (DISORDER)
C0154436|T048|191658009|SNOMEDCT_US|ATYPICAL MANIC DISORDER |ATYPICAL MANIC DISORDER (DISORDER)
C0338831|T048|231494001|SNOMEDCT_US|MANIA|MANIA (DISORDER)
C0338831|T048|231494001|SNOMEDCT_US|MANIC STATES|MANIA (DISORDER)
C0338831|T048|231494001|SNOMEDCT_US|STATE, MANIC|MANIA (DISORDER)
C0338831|T048|231494001|SNOMEDCT_US|STATES, MANIC|MANIA (DISORDER)
C0338831|T048|231494001|SNOMEDCT_US|MANIC|MANIA (DISORDER)
C0338831|T048|231494001|SNOMEDCT_US|MANIC STATE|MANIA (DISORDER)
C0338831|T048|231494001|SNOMEDCT_US|MANIA NOS|MANIA (DISORDER)
C0338831|T048|231494001|SNOMEDCT_US|MANIA |MANIA (DISORDER)
C0349208|T048|192354000|SNOMEDCT_US|MANIC EPISODE, UNSPECIFIED|[X] MANIA: [EPISODE, UNSPECIFIED] OR [NOS] (DISORDER)
C0349208|T048|192354000|SNOMEDCT_US|MANIC EPISODE|[X] MANIA: [EPISODE, UNSPECIFIED] OR [NOS] (DISORDER)
C0349208|T048|192354000|SNOMEDCT_US|MANIC EPISODE |[X] MANIA: [EPISODE, UNSPECIFIED] OR [NOS] (DISORDER)
C0349208|T048|192354000|SNOMEDCT_US|[X]MANIA NOS|[X] MANIA: [EPISODE, UNSPECIFIED] OR [NOS] (DISORDER)
C0349208|T048|192354000|SNOMEDCT_US|[X]MANIC EPISODE, UNSPECIFIED|[X] MANIA: [EPISODE, UNSPECIFIED] OR [NOS] (DISORDER)
C0349208|T048|192354000|SNOMEDCT_US|[X]MANIC EPISODE|[X] MANIA: [EPISODE, UNSPECIFIED] OR [NOS] (DISORDER)
C0349208|T048|192354000|SNOMEDCT_US|[X] MANIA: [EPISODE, UNSPECIFIED] OR [NOS]|[X] MANIA: [EPISODE, UNSPECIFIED] OR [NOS] (DISORDER)
C0349208|T048|192354000|SNOMEDCT_US|[X]MANIC EPISODE, UNSPECIFIED |[X] MANIA: [EPISODE, UNSPECIFIED] OR [NOS] (DISORDER)
C0349208|T048|192354000|SNOMEDCT_US|[X] MANIA: [EPISODE, UNSPECIFIED] OR [NOS] |[X] MANIA: [EPISODE, UNSPECIFIED] OR [NOS] (DISORDER)
C0349208|T048|192354000|SNOMEDCT_US|EPISODE; MANIC|[X] MANIA: [EPISODE, UNSPECIFIED] OR [NOS] (DISORDER)
C0349208|T048|192354000|SNOMEDCT_US|MANIC; EPISODE|[X] MANIA: [EPISODE, UNSPECIFIED] OR [NOS] (DISORDER)
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR DISORDERS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC DEPRESSIVE ILLNESS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR AFFECTIVE PSYCHOSIS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR DISORDER|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC DEPRESSIVE PSYCHOSIS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESSIVE PSYCHOSES|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|PSYCHOSES, BIPOLAR AFFECTIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|PSYCHOSES, MANIC DEPRESSIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|PSYCHOSIS, BIPOLAR AFFECTIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|PSYCHOSIS, MANIC DEPRESSIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR AFFECTIVE DISORDER|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|DISORDER, BIPOLAR|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESSIVE PSYCHOSIS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR AFFECTIVE DISORDER, UNSPECIFIED|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR DIS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESSION|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC DEPRESSIVE DISORDER|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BPAD|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|UNSPECIFIED BIPOLAR DISORDER|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|UNSPECIFIED BIPOLAR DISORDER |DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR DISORDER NOT OTHERWISE SPECIFIED|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC DEPRESSIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR DISORDER NOS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESSIVE REACTION|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESSIVE ILLNESS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR DISORDER, UNSPECIFIED|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|AFFECTIVE PSYCHOSIS, BIPOLAR|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR DISORDER [DISEASE/FINDING]|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|PSYCHOSES, MANIC-DEPRESSIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|PSYCHOSIS, MANIC-DEPRESSIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|DISORDER;BIPOLAR|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|DEPRESSION;MANIC|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|PSYCHOSIS;MANIC DEPRESSIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BI-POLAR DISORDER|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR DISORDER |DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|UNSPECIFIED BIPOLAR AFFECTIVE DISORDER|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|DEPRESSIVE-MANIC PSYCH.|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|UNSPECIFIED BIPOLAR AFFECTIVE DISORDER |DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|UNSPECIFIED BIPOLAR AFFECTIVE DISORDER, UNSPECIFIED|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|[X]BIPOLAR AFFECTIVE DISORDER, UNSPECIFIED|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|[X]BIPOLAR AFFECTIVE DISORDER, UNSPECIFIED |DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|UNSPECIFIED BIPOLAR AFFECTIVE DISORDER, UNSPECIFIED |DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|UNSPECIFIED BIPOLAR AFFECTIVE DISORDER, NOS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESS.PSYCHOSES|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|UNSPECIFIED BIPOLAR AFFECTIVE DISORDER, NOS |DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC DEPRESSION|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC DEPRESSIVE REACTION|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|REACTION MANIC-DEPRESSIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|PSYCHOSIS MANIC-DEPRESSIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MDI - MANIC-DEPRESSIVE ILLNESS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR; DISORDER, AFFECTIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR; DISORDER|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|DISORDER; BIPOLAR, AFFECTIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|DISORDER; BIPOLAR|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESSIVE; DISORDER|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESSIVE; PSYCHOSIS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESSIVE; SYNDROME|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|PSYCHOSIS; MANIC-DEPRESSIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|SYNDROME; MANIC-DEPRESSIVE|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR DISORDER, NOS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|BIPOLAR MOOD DISORDER|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESSIVE REACTION NOS|DEPRESSIVE-MANIC PSYCH.
C0005586|T048|268749008|SNOMEDCT_US|MANIC-DEPRESSIVE SYNDROME NOS|DEPRESSIVE-MANIC PSYCH.
C0236756|T048|191582005|SNOMEDCT_US|MANIC DISORDER, SINGLE EPISODE, UNSPECIFIED DEGREE|SINGLE MANIC EPISODE, UNSPECIFIED (DISORDER)
C0236756|T048|191582005|SNOMEDCT_US|BIPOLAR I DISORDER WITH SINGLE MANIC EPISODE |SINGLE MANIC EPISODE, UNSPECIFIED (DISORDER)
C0236756|T048|191582005|SNOMEDCT_US|BIPOLAR I DISORDER WITH SINGLE MANIC EPISODE|SINGLE MANIC EPISODE, UNSPECIFIED (DISORDER)
C0236756|T048|191582005|SNOMEDCT_US|BIPOL I SINGLE MANIC NOS|SINGLE MANIC EPISODE, UNSPECIFIED (DISORDER)
C0236756|T048|191582005|SNOMEDCT_US|BIPOLAR I DISORDER, SINGLE MANIC EPISODE, UNSPECIFIED|SINGLE MANIC EPISODE, UNSPECIFIED (DISORDER)
C0236756|T048|191582005|SNOMEDCT_US|BIPOLAR 1 DISORDER, SINGLE MANIC EPISODE|SINGLE MANIC EPISODE, UNSPECIFIED (DISORDER)
C0236756|T048|191582005|SNOMEDCT_US|MANIC DISORDER, SINGLE EPISODE NOS |SINGLE MANIC EPISODE, UNSPECIFIED (DISORDER)
C0236756|T048|191582005|SNOMEDCT_US|MANIC DISORDER, SINGLE EPISODE|SINGLE MANIC EPISODE, UNSPECIFIED (DISORDER)
C0236756|T048|191582005|SNOMEDCT_US|MANIC DISORDER, SINGLE EPISODE NOS|SINGLE MANIC EPISODE, UNSPECIFIED (DISORDER)
C0236756|T048|191582005|SNOMEDCT_US|SINGLE MANIC EPISODE, UNSPECIFIED|SINGLE MANIC EPISODE, UNSPECIFIED (DISORDER)
C0236756|T048|191582005|SNOMEDCT_US|SINGLE MANIC EPISODE, UNSPECIFIED |SINGLE MANIC EPISODE, UNSPECIFIED (DISORDER)
C0236756|T048|191582005|SNOMEDCT_US|MANIC DISORDER, SINGLE EPISODE |SINGLE MANIC EPISODE, UNSPECIFIED (DISORDER)
C0236756|T048|191582005|SNOMEDCT_US|MANIC EPISODE SINGLE|SINGLE MANIC EPISODE, UNSPECIFIED (DISORDER)
C0236756|T048|191582005|SNOMEDCT_US|BIPOLAR I DISORDER, SINGLE MANIC EPISODE|SINGLE MANIC EPISODE, UNSPECIFIED (DISORDER)
C0236756|T048|191582005|SNOMEDCT_US|MANIC DISORDER, SINGLE EPISODE |SINGLE MANIC EPISODE, UNSPECIFIED (DISORDER)
C0236756|T048|191582005|SNOMEDCT_US|BIPOLAR I DISORDER, SINGLE MANIC EPISODE |SINGLE MANIC EPISODE, UNSPECIFIED (DISORDER)
C0338846|T048|231495000|SNOMEDCT_US|MANIC STUPOR|MANIC STUPOR (DISORDER)
C0338846|T048|231495000|SNOMEDCT_US|MANIC STUPOR |MANIC STUPOR (DISORDER)
C0338846|T048|231495000|SNOMEDCT_US|MANIC EPISODE STUPOR|MANIC STUPOR (DISORDER)
C0338846|T048|231495000|SNOMEDCT_US|MANIC STUPOR |MANIC STUPOR (DISORDER)
C0338846|T048|231495000|SNOMEDCT_US|MANIC; STUPOR|MANIC STUPOR (DISORDER)
C0338846|T048|231495000|SNOMEDCT_US|STUPOR; MANIC|MANIC STUPOR (DISORDER)
C0338832|T048|192364009|SNOMEDCT_US|MANIC DISORDER WITH RECURRENT EPISODE|[X]RECURRENT MANIC EPISODES
C0338832|T048|192364009|SNOMEDCT_US|MANIC DISORDER, RECURRENT EPISODE|[X]RECURRENT MANIC EPISODES
C0338832|T048|192364009|SNOMEDCT_US|MANIC DISORDER WITH RECURRENT EPISODE |[X]RECURRENT MANIC EPISODES
C0338832|T048|192364009|SNOMEDCT_US|RECURRENT MANIC EPISODES NOS|[X]RECURRENT MANIC EPISODES
C0338832|T048|192364009|SNOMEDCT_US|RECURRENT MANIC EPISODE NOS |[X]RECURRENT MANIC EPISODES
C0338832|T048|192364009|SNOMEDCT_US|RECURRENT MANIC EPISODES, UNSPECIFIED |[X]RECURRENT MANIC EPISODES
C0338832|T048|192364009|SNOMEDCT_US|[X]RECURRENT MANIC EPISODES|[X]RECURRENT MANIC EPISODES
C0338832|T048|192364009|SNOMEDCT_US|RECURRENT MANIC EPISODE NOS|[X]RECURRENT MANIC EPISODES
C0338832|T048|192364009|SNOMEDCT_US|RECURRENT MANIC EPISODES, UNSPECIFIED|[X]RECURRENT MANIC EPISODES
C0338832|T048|192364009|SNOMEDCT_US|RECURRENT MANIC EPISODES|[X]RECURRENT MANIC EPISODES
C0338832|T048|192364009|SNOMEDCT_US|RECURRENT MANIC EPISODES |[X]RECURRENT MANIC EPISODES
C0270601|T048|41932008|SNOMEDCT_US|MALAYSIAN CULTURE|AMOK (DISORDER)
C0270601|T048|41932008|SNOMEDCT_US|MANIC EPISODE AMOK|AMOK (DISORDER)
C0270601|T048|41932008|SNOMEDCT_US|AMOK |AMOK (DISORDER)
C0270601|T048|41932008|SNOMEDCT_US|CATHARD|AMOK (DISORDER)
C0270601|T048|41932008|SNOMEDCT_US|IICH'AA|AMOK (DISORDER)
C0270601|T048|41932008|SNOMEDCT_US|MAL DE PELEA|AMOK (DISORDER)
C0270601|T048|41932008|SNOMEDCT_US|AMOK |AMOK (DISORDER)
C0270601|T048|41932008|SNOMEDCT_US|AMUCK|AMOK (DISORDER)
C0241934|T048|281257007|SNOMEDCT_US|HYPOMANIA|HYPOMANIC MOOD (FINDING)
C0241934|T048|281257007|SNOMEDCT_US|HYPOMANIA |HYPOMANIC MOOD (FINDING)
C0241934|T048|281257007|SNOMEDCT_US|HYPOMANIA |HYPOMANIC MOOD (FINDING)
C0241934|T048|281257007|SNOMEDCT_US|MANIC EPISODE HYPOMANIA|HYPOMANIC MOOD (FINDING)
C0241934|T048|281257007|SNOMEDCT_US|HYPOMANIC MOOD|HYPOMANIC MOOD (FINDING)
C0241934|T048|281257007|SNOMEDCT_US|HYPOMANIC MOOD |HYPOMANIC MOOD (FINDING)
C0865308|T048||SNOMEDCT_US|MANIA NOS SINGLE EPISODE OR UNSPECIFIED
C0865309|T048||SNOMEDCT_US|MONOPOLAR MANIA NOS SINGLE EPISODE OR UNSPECIFIED
C2874863|T048||SNOMEDCT_US|MANIC EPISODE WITHOUT PSYCHOTIC SYMPTOMS
C2874863|T048||SNOMEDCT_US|MANIC EPISODE WITHOUT PSYCHOTIC SYMPTOMS, UNSPECIFIED
C2874863|T048||SNOMEDCT_US|MANIC EPISODE WITHOUT PSYCHOTIC SYMPTOMS 
C0564408|T048|405273008|SNOMEDCT_US|MANIC MOOD|MANIC MOOD (FINDING)
C0564408|T048|405273008|SNOMEDCT_US|MANIC|MANIC MOOD (FINDING)
C0564408|T048|405273008|SNOMEDCT_US|MANIC MOOD |MANIC MOOD (FINDING)
C0865305|T048||SNOMEDCT_US|HYPOMANIA NOS SINGLE EPISODE OR UNSPECIFIED
C0865306|T048||SNOMEDCT_US|MILD HYPOMANIA NOS SINGLE EPISODE OR UNSPECIFIED
C0865307|T048||SNOMEDCT_US|HYPOMANIC PSYCHOSIS SINGLE EPISODE OR UNSPECIFIED
C1389907|T048||SNOMEDCT_US|BIPOLAR; DISORDER, SINGLE MANIC EPISODE, MILD
C1389907|T048||SNOMEDCT_US|DISORDER; BIPOLAR, SINGLE MANIC EPISODE, MILD
C1396834|T048||SNOMEDCT_US|EPISODE; HYPOMANIC
C1396834|T048||SNOMEDCT_US|HYPOMANIC; EPISODE
C1400223|T048||SNOMEDCT_US|EXCITEMENT; HYPOMANIC
C1400223|T048||SNOMEDCT_US|HYPOMANIC; EXCITEMENT
C0683410|T048||SNOMEDCT_US|HYPOMANIC PSYCHOSES
C0683410|T048||SNOMEDCT_US|HYPOMANIC PSYCHOSIS
C0683410|T048||SNOMEDCT_US|HYPOMANIC; PSYCHOSIS
C0683410|T048||SNOMEDCT_US|PSYCHOSIS; HYPOMANIC
C1400224|T048||SNOMEDCT_US|HYPOMANIC; REACTION
C1400224|T048||SNOMEDCT_US|REACTION; HYPOMANIC
