C0023890|T047|19943007|SNOMEDCT_US|LIVER CIRRHOSIS|CIRRHOSIS OF LIVER (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|LIVER CIRRHOSIS, ALCOHOLIC|ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|ALCOHOLIC LIVER CIRRHOSIS|ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|LIVER CIRRHOSIS, ALCOHOLIC|ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|ALCOHOLIC CIRRHOSIS OF LIVER|ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|ALCOHOLIC CIRRHOSIS|ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|ALCOHOLIC CIRRHOSIS |ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|CIRRHOSIS ALCOHOLIC|ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|ALCOHOL CIRRHOSIS LIVER|ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|ALCOHOLIC CIRRHOSIS NOS|ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|HEPATIC CIRRHOSIS, ALCOHOLIC|ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|LIVER CIRRHOSIS, ALCOHOLIC [DISEASE/FINDING]|ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|ALCOHOLIC CIRRHOSIS OF LIVER |ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|LAENNEC; ALCOHOLIC|ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|LAENNEC; CIRRHOSIS, ALCOHOLIC|ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|CIRRHOSIS; LAENNEC, ALCOHOLIC|ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|CIRRHOSIS; ALCOHOLIC|ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|CIRRHOSIS; LIVER, ALCOHOLIC|ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|LIVER; CIRRHOSIS, ALCOHOLIC|ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|ALCOHOL; LAENNEC|ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|ALCOHOL; CIRRHOSIS|ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|ALCOHOLIC CIRRHOSIS OF LIVER  [AMBIGUOUS]|ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|ALCOHOLIC HEPATIC CIRRHOSIS|ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|LAENNEC'S CIRRHOSIS, ALCOHOLIC|ALCOHOLIC CIRRHOSIS (DISORDER)
C0023891|T047|420054005|SNOMEDCT_US|ALCOHOLIC CIRRHOSIS |ALCOHOLIC CIRRHOSIS (DISORDER)
C0023892|T047|1761006|SNOMEDCT_US|LIVER CIRRHOSES, BILIARY|BILIARY CIRRHOSIS (DISORDER)
C0023892|T047|1761006|SNOMEDCT_US|LIVER CIRRHOSIS, BILIARY|BILIARY CIRRHOSIS (DISORDER)
C0023892|T047|1761006|SNOMEDCT_US|CIRRHOSIS, BILIARY|BILIARY CIRRHOSIS (DISORDER)
C0023892|T047|1761006|SNOMEDCT_US|BILIARY CIRRHOSIS, UNSPECIFIED|BILIARY CIRRHOSIS (DISORDER)
C0023892|T047|1761006|SNOMEDCT_US|BILIARY CIRRHOSIS|BILIARY CIRRHOSIS (DISORDER)
C0023892|T047|1761006|SNOMEDCT_US|CIRRHOSIS BILARY|BILIARY CIRRHOSIS (DISORDER)
C0023892|T047|1761006|SNOMEDCT_US|BILIARY LIVER CIRRHOSIS|BILIARY CIRRHOSIS (DISORDER)
C0023892|T047|1761006|SNOMEDCT_US|LIVER CIRRHOSIS, BILIARY [DISEASE/FINDING]|BILIARY CIRRHOSIS (DISORDER)
C0023892|T047|1761006|SNOMEDCT_US|CIRRHOSIS BILIARY|BILIARY CIRRHOSIS (DISORDER)
C0023892|T047|1761006|SNOMEDCT_US|BILIARY CIRRHOSIS |BILIARY CIRRHOSIS (DISORDER)
C0023892|T047|1761006|SNOMEDCT_US|BILIARY CIRRHOSIS NOS |BILIARY CIRRHOSIS (DISORDER)
C0023892|T047|1761006|SNOMEDCT_US|BILIARY CIRRHOSIS NOS|BILIARY CIRRHOSIS (DISORDER)
C0023892|T047|1761006|SNOMEDCT_US|CHOLANGITIC CIRRHOSIS|BILIARY CIRRHOSIS (DISORDER)
C0023892|T047|1761006|SNOMEDCT_US|CHOLESTATIC CIRRHOSIS|BILIARY CIRRHOSIS (DISORDER)
C0023892|T047|1761006|SNOMEDCT_US|BILIARY CIRRHOSIS |BILIARY CIRRHOSIS (DISORDER)
C0023892|T047|1761006|SNOMEDCT_US|BILIARY; CIRRHOSIS|BILIARY CIRRHOSIS (DISORDER)
C0023892|T047|1761006|SNOMEDCT_US|CIRRHOSIS; BILIARY|BILIARY CIRRHOSIS (DISORDER)
C0023892|T047|1761006|SNOMEDCT_US|CIRRHOSIS, CHOLANGITIC|BILIARY CIRRHOSIS (DISORDER)
C0023892|T047|1761006|SNOMEDCT_US|CIRRHOSIS, CHOLESTATIC|BILIARY CIRRHOSIS (DISORDER)
C0023893|T047||SNOMEDCT_US|LIVER CIRRHOSIS, EXPERIMENTAL
C0023890|T047|19943007|SNOMEDCT_US|CIRRHOSES, HEPATIC|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|CIRRHOSES, LIVER|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|CIRRHOSIS, HEPATIC|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|HEPATIC CIRRHOSES|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|LIVER CIRRHOSES|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|LIVER CIRRHOSIS|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|CIRRHOSIS|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|HEPATIC CIRRHOSIS|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|CIRRHOSIS OF LIVER|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|HEPATIC CIRRHOSIS |CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|CIRRHOSIS (OF LIVER) NOS|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|LIVER CIRRHOSIS [DISEASE/FINDING]|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|CIRRHOSIS, LIVER|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|CIRRHOSIS (OF);LIVER|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|CIRRHOSIS OF LIVER NOS|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|CIRRHOSIS OF LIVER NOS |CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|LIVER--CIRRHOSIS|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|HEPATIC CIRRHOSIS NOS|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|CIRRHOSIS LIVER|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|CL - CIRRHOSIS OF LIVER|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|CIRRHOSIS OF LIVER |CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|CIRRHOSIS; LIVER|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|LIVER; CIRRHOSIS|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|CIRRHOSIS OF LIVER, NOS|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|HEPATIC CIRRHOSIS, NOS|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|CIRRHOSIS (LIVER)|CIRRHOSIS OF LIVER (DISORDER)
C0023890|T047|19943007|SNOMEDCT_US|CIRRHOSIS OF THE LIVER|CIRRHOSIS OF LIVER (DISORDER)
C0267809|T047|89580002|SNOMEDCT_US|CIRRHOSIS, CRYPTOGENIC|CRYPTOGENIC CIRRHOSIS (DISORDER)
C0267809|T047|89580002|SNOMEDCT_US|CRYPTOGENIC CIRRHOSIS|CRYPTOGENIC CIRRHOSIS (DISORDER)
C0267809|T047|89580002|SNOMEDCT_US|CRYPTOGENIC CIRRHOSIS |CRYPTOGENIC CIRRHOSIS (DISORDER)
C0267809|T047|89580002|SNOMEDCT_US|CRYPTOGENIC CIRRHOSIS (OF LIVER)|CRYPTOGENIC CIRRHOSIS (DISORDER)
C0267809|T047|89580002|SNOMEDCT_US|CRYPTOGENIC CIRRHOSIS OF LIVER|CRYPTOGENIC CIRRHOSIS (DISORDER)
C0267809|T047|89580002|SNOMEDCT_US|CRYPTOGENIC CIRRHOSIS |CRYPTOGENIC CIRRHOSIS (DISORDER)
C1442995|T047|399126000|SNOMEDCT_US|PIGMENTARY CIRRHOSIS |BRONZE CIRRHOSIS (DISORDER)
C1442995|T047|399126000|SNOMEDCT_US|PIGMENTARY CIRRHOSIS|BRONZE CIRRHOSIS (DISORDER)
C1442995|T047|399126000|SNOMEDCT_US|PIGMENTARY CIRRHOSIS (OF LIVER)|BRONZE CIRRHOSIS (DISORDER)
C1442995|T047|399126000|SNOMEDCT_US|BRONZE CIRRHOSIS|BRONZE CIRRHOSIS (DISORDER)
C1442995|T047|399126000|SNOMEDCT_US|PIGMENTARY CIRRHOSIS OF LIVER|BRONZE CIRRHOSIS (DISORDER)
C1442995|T047|399126000|SNOMEDCT_US|BRONZED CIRRHOSIS|BRONZE CIRRHOSIS (DISORDER)
C1442995|T047|399126000|SNOMEDCT_US|BRONZE CIRRHOSIS |BRONZE CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|POSTNECROTIC CIRRHOSIS |POSTNECROTIC CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|POSTNECROTIC CIRRHOSIS|POSTNECROTIC CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|MACRONODULAR CIRRHOSIS|POSTNECROTIC CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|MACRONODULAR CIRRHOSIS |POSTNECROTIC CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|MACRONODULAR CIRRHOSIS (OF LIVER)|POSTNECROTIC CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|POSTNECROTIC CIRRHOSIS (OF LIVER)|POSTNECROTIC CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|POSTNECROTIC CIRRHOSIS OF LIVER|POSTNECROTIC CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|HYPERTROPHIC PORTAL CIRRHOSIS|POSTNECROTIC CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|MACRONODULAR CIRRHOSIS OF LIVER|POSTNECROTIC CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|PNC - POSTNECROTIC CIRRHOSIS|POSTNECROTIC CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|MACRONODULAR CIRRHOSIS |POSTNECROTIC CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|CIRRHOSIS LIVER POSTNECROTIC|POSTNECROTIC CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|HEPATIC CIRRHOSIS POST NECROTIC|POSTNECROTIC CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|CIRRHOSIS LIVER POST NECROTIC|POSTNECROTIC CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|HEALED YELLOW ATROPHY OF LIVER|POSTNECROTIC CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|POSTNECROTIC CIRRHOSIS |POSTNECROTIC CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|CIRRHOSIS; MACRONODULAR|POSTNECROTIC CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|CIRRHOSIS; PERIPORTAL|POSTNECROTIC CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|CIRRHOSIS; POSTNECROTIC|POSTNECROTIC CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|MACRONODULAR; CIRRHOSIS|POSTNECROTIC CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|PERIPORTAL; CIRRHOSIS|POSTNECROTIC CIRRHOSIS (DISORDER)
C2004456|T047|86454000|SNOMEDCT_US|POSTNECROTIC; CIRRHOSIS|POSTNECROTIC CIRRHOSIS (DISORDER)
C0267812|T047|21861000|SNOMEDCT_US|MICRONODULAR CIRRHOSIS|MICRONODULAR CIRRHOSIS (DISORDER)
C0267812|T047|21861000|SNOMEDCT_US|MICRONODULAR CIRRHOSIS |MICRONODULAR CIRRHOSIS (DISORDER)
C0267812|T047|21861000|SNOMEDCT_US|MICRONODULAR CIRRHOSIS |MICRONODULAR CIRRHOSIS (DISORDER)
C0267812|T047|21861000|SNOMEDCT_US|CIRRHOSIS; MICRONODULAR|MICRONODULAR CIRRHOSIS (DISORDER)
C0267812|T047|21861000|SNOMEDCT_US|MICRONODULAR; CIRRHOSIS|MICRONODULAR CIRRHOSIS (DISORDER)
C0085699|T047|74669004|SNOMEDCT_US|CARDIAC CIRRHOSIS|CARDIAC CIRRHOSIS (DISORDER)
C0085699|T047|74669004|SNOMEDCT_US|CARDIAC CIRRHOSIS |CARDIAC CIRRHOSIS (DISORDER)
C0085699|T047|74669004|SNOMEDCT_US|CONGESTIVE CIRRHOSIS|CARDIAC CIRRHOSIS (DISORDER)
C0085699|T047|74669004|SNOMEDCT_US|CARDIAC CIRRHOSIS |CARDIAC CIRRHOSIS (DISORDER)
C0085699|T047|74669004|SNOMEDCT_US|CARDIAC; CIRRHOSIS|CARDIAC CIRRHOSIS (DISORDER)
C0085699|T047|74669004|SNOMEDCT_US|CIRRHOSE CARDIAQUE|CARDIAC CIRRHOSIS (DISORDER)
C0085699|T047|74669004|SNOMEDCT_US|CIRRHOSIS; CARDIAC|CARDIAC CIRRHOSIS (DISORDER)
C0085699|T047|74669004|SNOMEDCT_US|CIRRHOSIS; CONGESTIVE|CARDIAC CIRRHOSIS (DISORDER)
C0085699|T047|74669004|SNOMEDCT_US|CONGESTIVE; CIRRHOSIS|CARDIAC CIRRHOSIS (DISORDER)
C0085699|T047|74669004|SNOMEDCT_US|CARDIAC CIRRHOSIS, NOS|CARDIAC CIRRHOSIS (DISORDER)
C2062319|T047||SNOMEDCT_US|CIRRHOSIS, RARE TYPES
C2062319|T047||SNOMEDCT_US|RARE TYPES OF CIRRHOSIS
C2062319|T047||SNOMEDCT_US|RARE TYPES OF CIRRHOSIS 
C2075269|T047||SNOMEDCT_US|CIRRHOSIS DUE TO HEPATITIS A
C2075269|T047||SNOMEDCT_US|CIRRHOSIS DUE TO HEPATITIS A 
C2075270|T047||SNOMEDCT_US|CIRRHOSIS DUE TO HEPATITIS B
C2075270|T047||SNOMEDCT_US|CIRRHOSIS DUE TO HEPATITIS B 
C2075271|T047||SNOMEDCT_US|CIRRHOSIS DUE TO HEPATITIS C 
C2075271|T047||SNOMEDCT_US|CIRRHOSIS DUE TO HEPATITIS C
C1622502|T047|197308000|SNOMEDCT_US|PORTAL CIRRHOSIS (OF LIVER)|PORTAL CIRRHOSIS UNSPECIFIED (DISORDER)
C1622502|T047|197308000|SNOMEDCT_US|PORTAL CIRRHOSIS UNSPECIFIED|PORTAL CIRRHOSIS UNSPECIFIED (DISORDER)
C1622502|T047|197308000|SNOMEDCT_US|LAENNEC'S CIRRHOSIS|PORTAL CIRRHOSIS UNSPECIFIED (DISORDER)
C1622502|T047|197308000|SNOMEDCT_US|PORTAL CIRRHOSIS|PORTAL CIRRHOSIS UNSPECIFIED (DISORDER)
C1622502|T047|197308000|SNOMEDCT_US|PORTAL CIRRHOSIS |PORTAL CIRRHOSIS UNSPECIFIED (DISORDER)
C1622502|T047|197308000|SNOMEDCT_US|PORTAL CIRRHOSIS UNSPECIFIED |PORTAL CIRRHOSIS UNSPECIFIED (DISORDER)
C1622502|T047|197308000|SNOMEDCT_US|PC - PORTAL CIRRHOSIS|PORTAL CIRRHOSIS UNSPECIFIED (DISORDER)
C1622502|T047|197308000|SNOMEDCT_US|CIRRHOSIS PORTAL|PORTAL CIRRHOSIS UNSPECIFIED (DISORDER)
C1622502|T047|197308000|SNOMEDCT_US|PORTAL CIRRHOSIS |PORTAL CIRRHOSIS UNSPECIFIED (DISORDER)
C1622502|T047|197308000|SNOMEDCT_US|LAENNEC; CIRRHOSIS|PORTAL CIRRHOSIS UNSPECIFIED (DISORDER)
C1622502|T047|197308000|SNOMEDCT_US|CIRRHOSIS; LAENNEC|PORTAL CIRRHOSIS UNSPECIFIED (DISORDER)
C1622502|T047|197308000|SNOMEDCT_US|CIRRHOSIS; PORTAL|PORTAL CIRRHOSIS UNSPECIFIED (DISORDER)
C1622502|T047|197308000|SNOMEDCT_US|PORTAL; CIRRHOSIS|PORTAL CIRRHOSIS UNSPECIFIED (DISORDER)
C1622502|T047|197308000|SNOMEDCT_US|PORTAL CIRRHOSIS, NOS|PORTAL CIRRHOSIS UNSPECIFIED (DISORDER)
C0400947|T047|197293003|SNOMEDCT_US|CIRRHOSIS DIFFUSE NODULAR|DIFFUSE NODULAR CIRRHOSIS (DISORDER)
C0400947|T047|197293003|SNOMEDCT_US|CIRRHOSIS DIFFUSE NODULAR |DIFFUSE NODULAR CIRRHOSIS (DISORDER)
C0400947|T047|197293003|SNOMEDCT_US|DIFFUSE NODULAR CIRRHOSIS|DIFFUSE NODULAR CIRRHOSIS (DISORDER)
C0400947|T047|197293003|SNOMEDCT_US|DIFFUSE NODULAR CIRRHOSIS |DIFFUSE NODULAR CIRRHOSIS (DISORDER)
C0400951|T047|197304003|SNOMEDCT_US|CIRRHOSIS CARDITUBERCULOUS |CARDITUBERCULOUS CIRRHOSIS (DISORDER)
C0400951|T047|197304003|SNOMEDCT_US|CIRRHOSIS CARDITUBERCULOUS|CARDITUBERCULOUS CIRRHOSIS (DISORDER)
C0400951|T047|197304003|SNOMEDCT_US|CARDITUBERCULOUS CIRRHOSIS|CARDITUBERCULOUS CIRRHOSIS (DISORDER)
C0400951|T047|197304003|SNOMEDCT_US|CARDITUBERCULOUS CIRRHOSIS |CARDITUBERCULOUS CIRRHOSIS (DISORDER)
C0268074|T047|6183001|SNOMEDCT_US|INDIAN CHILDHOOD CIRRHOSIS|INDIAN CHILDHOOD CIRRHOSIS (DISORDER)
C0268074|T047|6183001|SNOMEDCT_US|CIRRHOSIS, FAMILIAL, WITH PULMONARY HYPERTENSION|INDIAN CHILDHOOD CIRRHOSIS (DISORDER)
C0268074|T047|6183001|SNOMEDCT_US|SEN SYNDROME|INDIAN CHILDHOOD CIRRHOSIS (DISORDER)
C0268074|T047|6183001|SNOMEDCT_US|CIRRHOSIS-FAMILIAL WITH PULMONARY HYPERTENSION|INDIAN CHILDHOOD CIRRHOSIS (DISORDER)
C0268074|T047|6183001|SNOMEDCT_US|ICC - INDIAN CHILDHOOD CIRRHOSIS|INDIAN CHILDHOOD CIRRHOSIS (DISORDER)
C0268074|T047|6183001|SNOMEDCT_US|INDIAN CHILDHOOD CIRRHOSIS |INDIAN CHILDHOOD CIRRHOSIS (DISORDER)
C0268074|T047|6183001|SNOMEDCT_US|INDIAN CHILDHOOD; CIRRHOSIS|INDIAN CHILDHOOD CIRRHOSIS (DISORDER)
C0268074|T047|6183001|SNOMEDCT_US|CIRRHOSIS; INDIAN CHILDHOOD|INDIAN CHILDHOOD CIRRHOSIS (DISORDER)
C1392670|T047||SNOMEDCT_US|CONGENITAL CIRRHOSIS (OF LIVER)
C1392670|T047||SNOMEDCT_US|CONGENITAL CIRRHOSIS LIVER
C1392670|T047||SNOMEDCT_US|CONGENITAL CIRRHOSIS OF LIVER
C1392670|T047||SNOMEDCT_US|CONGENITAL CIRRHOSIS OF LIVER 
C1392670|T047||SNOMEDCT_US|CIRRHOSIS; LIVER, CONGENITAL
C0239946|T047|197317000|SNOMEDCT_US|FIBROSES, LIVER|FIBROSIS OF LIVER (DISORDER)
C0239946|T047|197317000|SNOMEDCT_US|LIVER FIBROSES|FIBROSIS OF LIVER (DISORDER)
C0239946|T047|197317000|SNOMEDCT_US|HEPATIC FIBROSIS|FIBROSIS OF LIVER (DISORDER)
C0239946|T047|197317000|SNOMEDCT_US|HEPATIC FIBROSIS |FIBROSIS OF LIVER (DISORDER)
C0239946|T047|197317000|SNOMEDCT_US|LIVER FIBROSIS|FIBROSIS OF LIVER (DISORDER)
C0239946|T047|197317000|SNOMEDCT_US|FIBROSIS OF LIVER|FIBROSIS OF LIVER (DISORDER)
C0239946|T047|197317000|SNOMEDCT_US|FIBROSIS OF LIVER |FIBROSIS OF LIVER (DISORDER)
C0239946|T047|197317000|SNOMEDCT_US|FIBROSIS LIVER|FIBROSIS OF LIVER (DISORDER)
C0239946|T047|197317000|SNOMEDCT_US|HEPATIC FIBROSIS |FIBROSIS OF LIVER (DISORDER)
C0239946|T047|197317000|SNOMEDCT_US|FIBROSIS; LIVER|FIBROSIS OF LIVER (DISORDER)
C0239946|T047|197317000|SNOMEDCT_US|LIVER; FIBROSIS|FIBROSIS OF LIVER (DISORDER)
C0239946|T047|197317000|SNOMEDCT_US|HEPATIC FIBROSIS, NOS|FIBROSIS OF LIVER (DISORDER)
C0239946|T047|197317000|SNOMEDCT_US|FIBROSIS, LIVER|FIBROSIS OF LIVER (DISORDER)
C3662136|T047|831000119103|SNOMEDCT_US|CHRONIC HEPATITIS C WITH STAGE 4 FIBROSIS|CHRONIC HEPATITIS C WITH STAGE 4 FIBROSIS
C3662136|T047|831000119103|SNOMEDCT_US|CIRRHOSIS OF LIVER DUE TO CHRONIC HEPATITS C |CHRONIC HEPATITIS C WITH STAGE 4 FIBROSIS
C3662136|T047|831000119103|SNOMEDCT_US|CIRRHOSIS OF LIVER DUE TO CHRONIC HEPATITS C|CHRONIC HEPATITIS C WITH STAGE 4 FIBROSIS
C3662136|T047|831000119103|SNOMEDCT_US|CIRRHOSIS OF LIVER DUE TO CHRONIC HEPATITIS C|CHRONIC HEPATITIS C WITH STAGE 4 FIBROSIS
C3662136|T047|831000119103|SNOMEDCT_US|CIRRHOSIS OF LIVER DUE TO CHRONIC HEPATITIS C |CHRONIC HEPATITIS C WITH STAGE 4 FIBROSIS
C0275872|T047|16070004|SNOMEDCT_US|SYPHILITIC CIRRHOSIS|SYPHILITIC CIRRHOSIS (DISORDER)
C0275872|T047|16070004|SNOMEDCT_US|CIRRHOSIS SYPHILITIC|SYPHILITIC CIRRHOSIS (DISORDER)
C0275872|T047|16070004|SNOMEDCT_US|SYPHILITIC CIRRHOSIS |SYPHILITIC CIRRHOSIS (DISORDER)
C0275872|T047|16070004|SNOMEDCT_US|HEPAR LOBATUM|SYPHILITIC CIRRHOSIS (DISORDER)
C0275872|T047|16070004|SNOMEDCT_US|SYPHILITIC CIRRHOSIS |SYPHILITIC CIRRHOSIS (DISORDER)
C1861556|T047||SNOMEDCT_US|CIRRHOSIS, FAMILIAL
C0009714|T047|79607001|SNOMEDCT_US|CONGENITAL HEPATIC FIBROSIS|CONGENITAL HEPATIC FIBROSIS (DISORDER)
C0009714|T047|79607001|SNOMEDCT_US|HEPATIC FIBROSIS, CONGENITAL|CONGENITAL HEPATIC FIBROSIS (DISORDER)
C0009714|T047|79607001|SNOMEDCT_US|CONGENITAL HEPATIC FIBROSIS |CONGENITAL HEPATIC FIBROSIS (DISORDER)
C0009714|T047|79607001|SNOMEDCT_US|CONGENITAL FIBROSE LIVER|CONGENITAL HEPATIC FIBROSIS (DISORDER)
C0009714|T047|79607001|SNOMEDCT_US|CONGENITAL HEPATIC FIBROSIS |CONGENITAL HEPATIC FIBROSIS (DISORDER)
C1859088|T047||SNOMEDCT_US|COPPER TOXICOSIS, IDIOPATHIC
C1859088|T047||SNOMEDCT_US| CAN BE SEVERAL THINGS (INDUCTION CHEMOTHERAPY)
C3874483|T047|103611000119102|SNOMEDCT_US|CIRRHOSIS OF LIVER DUE TO HEPATITIS B |CIRRHOSIS OF LIVER DUE TO HEPATITIS B (DISORDER)
C3874483|T047|103611000119102|SNOMEDCT_US|CIRRHOSIS OF LIVER DUE TO HEPATITIS B|CIRRHOSIS OF LIVER DUE TO HEPATITIS B (DISORDER)
C1392669|T047||SNOMEDCT_US|MIXED CIRRHOSIS
C1392669|T047||SNOMEDCT_US|CIRRHOSIS; MIXED TYPE
C1392669|T047||SNOMEDCT_US|MIXED; CIRRHOSIS
C0010398|T047|45256007|SNOMEDCT_US|CRUVEILHIER BAUMGARTEN SYNDROME|CRUVEILHIER-BAUMGARTEN SYNDROME (DISORDER)
C0010398|T047|45256007|SNOMEDCT_US|SYNDROME, CRUVEILHIER-BAUMGARTEN|CRUVEILHIER-BAUMGARTEN SYNDROME (DISORDER)
C0010398|T047|45256007|SNOMEDCT_US|CRUVEILHIER-BAUMGARTEN SYNDROME|CRUVEILHIER-BAUMGARTEN SYNDROME (DISORDER)
C0010398|T047|45256007|SNOMEDCT_US|CRUVEILHIER-BAUMGARTEN SYNDROME |CRUVEILHIER-BAUMGARTEN SYNDROME (DISORDER)
C0010398|T047|45256007|SNOMEDCT_US|CIRRHOSIS; BAUMGARTEN-CRUVEILHIER|CRUVEILHIER-BAUMGARTEN SYNDROME (DISORDER)
C0010398|T047|45256007|SNOMEDCT_US|CIRRHOSIS; CRUVEILHIER-BAUMGARTEN|CRUVEILHIER-BAUMGARTEN SYNDROME (DISORDER)
C0010398|T047|45256007|SNOMEDCT_US|BAUMGARTEN-CRUVEILHIER; CIRRHOSIS|CRUVEILHIER-BAUMGARTEN SYNDROME (DISORDER)
C0010398|T047|45256007|SNOMEDCT_US|BAUMGARTEN-CRUVEILHIER|CRUVEILHIER-BAUMGARTEN SYNDROME (DISORDER)
C0010398|T047|45256007|SNOMEDCT_US|CRUVEILHIER-BAUMGARTEN; CIRRHOSIS|CRUVEILHIER-BAUMGARTEN SYNDROME (DISORDER)
C0010398|T047|45256007|SNOMEDCT_US|CRUVEILHIER-BAUMGARTEN|CRUVEILHIER-BAUMGARTEN SYNDROME (DISORDER)
C0267806|T047|76301009|SNOMEDCT_US|FLORID CIRRHOSIS|FLORID CIRRHOSIS (DISORDER)
C0267806|T047|76301009|SNOMEDCT_US|FLORID CIRRHOSIS |FLORID CIRRHOSIS (DISORDER)
C0267817|T047|536002|SNOMEDCT_US|GLISSONIAN CIRRHOSIS|GLISSONIAN CIRRHOSIS (DISORDER)
C0267817|T047|536002|SNOMEDCT_US|GLISSONIAN CIRRHOSIS |GLISSONIAN CIRRHOSIS (DISORDER)
C0267815|T047|78208005|SNOMEDCT_US|PIGMENT CIRRHOSIS|PIGMENT CIRRHOSIS (DISORDER)
C0267815|T047|78208005|SNOMEDCT_US|PIGMENT CIRRHOSIS |PIGMENT CIRRHOSIS (DISORDER)
C0267813|T047|27156006|SNOMEDCT_US|POSTHEPATITIC CIRRHOSIS|POSTHEPATITIC CIRRHOSIS (DISORDER)
C0267813|T047|27156006|SNOMEDCT_US|POSTHEPATITIC CIRRHOSIS |POSTHEPATITIC CIRRHOSIS (DISORDER)
C0267813|T047|27156006|SNOMEDCT_US|CIRRHOSIS; POSTHEPATITIC|POSTHEPATITIC CIRRHOSIS (DISORDER)
C0267813|T047|27156006|SNOMEDCT_US|POSTHEPATITIC; CIRRHOSIS|POSTHEPATITIC CIRRHOSIS (DISORDER)
C0156189|T047|197279005|SNOMEDCT_US|CHRONIC LIVER DISEASE AND CIRRHOSIS|CIRRHOSIS AND CHRONIC LIVER DISEASE (DISORDER)
C0156189|T047|197279005|SNOMEDCT_US|CIRRHOSIS/CHRONIC LIVER DIS.|CIRRHOSIS AND CHRONIC LIVER DISEASE (DISORDER)
C0156189|T047|197279005|SNOMEDCT_US|CIRRHOSIS AND CHRONIC LIVER DISEASE|CIRRHOSIS AND CHRONIC LIVER DISEASE (DISORDER)
C0156189|T047|197279005|SNOMEDCT_US|CIRRHOSIS AND CHRONIC LIVER DISEASE |CIRRHOSIS AND CHRONIC LIVER DISEASE (DISORDER)
C0341446|T047|235899008|SNOMEDCT_US|HEPATIC SCLEROSIS|HEPATIC SCLEROSIS (DISORDER)
C0341446|T047|235899008|SNOMEDCT_US|HEPATIC SCLEROSIS |HEPATIC SCLEROSIS (DISORDER)
C0341446|T047|235899008|SNOMEDCT_US|HEPATIC SCLEROSIS |HEPATIC SCLEROSIS (DISORDER)
C0341446|T047|235899008|SNOMEDCT_US|LIVER; SCLEROSIS|HEPATIC SCLEROSIS (DISORDER)
C0341446|T047|235899008|SNOMEDCT_US|SCLEROSIS; LIVER|HEPATIC SCLEROSIS (DISORDER)
C0348749|T047|197553002|SNOMEDCT_US|OTHER AND UNSPECIFIED CIRRHOSIS OF LIVER|[X]OTHER AND UNSPECIFIED CIRRHOSIS OF LIVER (DISORDER)
C0348749|T047|197553002|SNOMEDCT_US|[X]OTHER AND UNSPECIFIED CIRRHOSIS OF LIVER |[X]OTHER AND UNSPECIFIED CIRRHOSIS OF LIVER (DISORDER)
C0348749|T047|197553002|SNOMEDCT_US|[X]OTHER AND UNSPECIFIED CIRRHOSIS OF LIVER|[X]OTHER AND UNSPECIFIED CIRRHOSIS OF LIVER (DISORDER)
C0400941|T047|197296006|SNOMEDCT_US|PORTAL CIRRHOSIS CAPSULAR |CAPSULAR PORTAL CIRRHOSIS (DISORDER)
C0400941|T047|197296006|SNOMEDCT_US|PORTAL CIRRHOSIS CAPSULAR|CAPSULAR PORTAL CIRRHOSIS (DISORDER)
C0400941|T047|197296006|SNOMEDCT_US|CAPSULAR PORTAL CIRRHOSIS|CAPSULAR PORTAL CIRRHOSIS (DISORDER)
C0400941|T047|197296006|SNOMEDCT_US|CAPSULAR PORTAL CIRRHOSIS |CAPSULAR PORTAL CIRRHOSIS (DISORDER)
C0400957|T047|271440004|SNOMEDCT_US|CIRRHOSIS SECONDARY TO CHOLESTASIS |CIRRHOSIS SECONDARY TO CHOLESTASIS (DISORDER)
C0400957|T047|271440004|SNOMEDCT_US|CIRRHOSIS SECONDARY TO CHOLESTASIS|CIRRHOSIS SECONDARY TO CHOLESTASIS (DISORDER)
C0400942|T047|197294009|SNOMEDCT_US|PORTAL CIRRHOSIS FATTY|FATTY PORTAL CIRRHOSIS (DISORDER)
C0400942|T047|197294009|SNOMEDCT_US|PORTAL CIRRHOSIS FATTY |FATTY PORTAL CIRRHOSIS (DISORDER)
C0400942|T047|197294009|SNOMEDCT_US|FATTY PORTAL CIRRHOSIS|FATTY PORTAL CIRRHOSIS (DISORDER)
C0400942|T047|197294009|SNOMEDCT_US|FATTY PORTAL CIRRHOSIS |FATTY PORTAL CIRRHOSIS (DISORDER)
C0400961|T047|235901004|SNOMEDCT_US|HEPATIC FIBROSIS WITH HEPATIC SCLEROSIS|HEPATIC FIBROSIS WITH HEPATIC SCLEROSIS (DISORDER)
C0400961|T047|235901004|SNOMEDCT_US|HEPATIC FIBROSIS WITH HEPATIC SCLEROSIS |HEPATIC FIBROSIS WITH HEPATIC SCLEROSIS (DISORDER)
C0400961|T047|235901004|SNOMEDCT_US|HEPATIC FIBROSIS WITH HEPATIC SCLEROSIS |HEPATIC FIBROSIS WITH HEPATIC SCLEROSIS (DISORDER)
C0400961|T047|235901004|SNOMEDCT_US|FIBROSIS; LIVER, WITH SCLEROSIS|HEPATIC FIBROSIS WITH HEPATIC SCLEROSIS (DISORDER)
C0400961|T047|235901004|SNOMEDCT_US|SCLEROSIS; LIVER, WITH FIBROSIS|HEPATIC FIBROSIS WITH HEPATIC SCLEROSIS (DISORDER)
C0400949|T047|235896001|SNOMEDCT_US|INFECTIOUS CIRRHOSIS NOS |INFECTIOUS CIRRHOSIS (DISORDER)
C0400949|T047|235896001|SNOMEDCT_US|INFECTIOUS CIRRHOSIS NOS|INFECTIOUS CIRRHOSIS (DISORDER)
C0400949|T047|235896001|SNOMEDCT_US|INFECTIOUS CIRRHOSIS|INFECTIOUS CIRRHOSIS (DISORDER)
C0400949|T047|235896001|SNOMEDCT_US|INFECTIOUS CIRRHOSIS |INFECTIOUS CIRRHOSIS (DISORDER)
C0400940|T047|197299004|SNOMEDCT_US|PIGMENTARY PORTAL CIRRHOSIS|PIGMENTARY PORTAL CIRRHOSIS (DISORDER)
C0400940|T047|197299004|SNOMEDCT_US|PIGMENTARY PORTAL CIRRHOSIS |PIGMENTARY PORTAL CIRRHOSIS (DISORDER)
C0400956|T047|123604002|SNOMEDCT_US|TOXIC CIRRHOSIS|TOXIC CIRRHOSIS (DISORDER)
C0400956|T047|123604002|SNOMEDCT_US|TOXIC CIRRHOSIS |TOXIC CIRRHOSIS (DISORDER)
C0400939|T047|197301006|SNOMEDCT_US|PORTAL CIRRHOSIS TOXIC |TOXIC PORTAL CIRRHOSIS (DISORDER)
C0400939|T047|197301006|SNOMEDCT_US|PORTAL CIRRHOSIS TOXIC|TOXIC PORTAL CIRRHOSIS (DISORDER)
C0400939|T047|197301006|SNOMEDCT_US|TOXIC PORTAL CIRRHOSIS|TOXIC PORTAL CIRRHOSIS (DISORDER)
C0400939|T047|197301006|SNOMEDCT_US|TOXIC PORTAL CIRRHOSIS |TOXIC PORTAL CIRRHOSIS (DISORDER)
C0400938|T047|197291001|SNOMEDCT_US|PORTAL CIRRHOSIS UNILOBULAR |UNILOBULAR PORTAL CIRRHOSIS (DISORDER)
C0400938|T047|197291001|SNOMEDCT_US|PORTAL CIRRHOSIS UNILOBULAR|UNILOBULAR PORTAL CIRRHOSIS (DISORDER)
C0400938|T047|197291001|SNOMEDCT_US|UNILOBULAR PORTAL CIRRHOSIS|UNILOBULAR PORTAL CIRRHOSIS (DISORDER)
C0400938|T047|197291001|SNOMEDCT_US|UNILOBULAR PORTAL CIRRHOSIS |UNILOBULAR PORTAL CIRRHOSIS (DISORDER)
C0400943|T047|266468003|SNOMEDCT_US|CIRRHOSIS, NONALCOHOLIC|CIRRHOSIS - NON-ALCOHOLIC (DISORDER)
C0400943|T047|266468003|SNOMEDCT_US|NON-ALCOHOLIC CIRRHOSIS NOS|CIRRHOSIS - NON-ALCOHOLIC (DISORDER)
C0400943|T047|266468003|SNOMEDCT_US|CIRRHOSIS - NON ALCOHOLIC|CIRRHOSIS - NON-ALCOHOLIC (DISORDER)
C0400943|T047|266468003|SNOMEDCT_US|CIRRHOSIS - NON-ALCOHOLIC|CIRRHOSIS - NON-ALCOHOLIC (DISORDER)
C0400943|T047|266468003|SNOMEDCT_US|CIRRHOSIS - NON-ALCOHOLIC |CIRRHOSIS - NON-ALCOHOLIC (DISORDER)
C0400943|T047|266468003|SNOMEDCT_US|NON-ALCOHOLIC CIRRHOSIS NOS |CIRRHOSIS - NON-ALCOHOLIC (DISORDER)
C0400943|T047|266468003|SNOMEDCT_US|CIRRHOSIS OF LIVER NOT DUE TO ALCOHOL|CIRRHOSIS - NON-ALCOHOLIC (DISORDER)
C0400943|T047|266468003|SNOMEDCT_US|CIRRHOSIS OF LIVER NOT DUE TO ALCOHOL |CIRRHOSIS - NON-ALCOHOLIC (DISORDER)
C0400955|T047|235897005|SNOMEDCT_US|HYPOXIA-ASSOCIATED CIRRHOSIS|HYPOXIA-ASSOCIATED CIRRHOSIS (DISORDER)
C0400955|T047|235897005|SNOMEDCT_US|HYPOXIA-ASSOCIATED CIRRHOSIS |HYPOXIA-ASSOCIATED CIRRHOSIS (DISORDER)
C1263668|T047|123606000|SNOMEDCT_US|CHOLANGIOLITIC CIRRHOSIS |CHOLANGIOLITIC CIRRHOSIS (DISORDER)
C1263668|T047|123606000|SNOMEDCT_US|CHOLANGIOLITIC CIRRHOSIS|CHOLANGIOLITIC CIRRHOSIS (DISORDER)
C1263668|T047|123606000|SNOMEDCT_US|CHOLANGIOLITIC; CIRRHOSIS|CHOLANGIOLITIC CIRRHOSIS (DISORDER)
C1263668|T047|123606000|SNOMEDCT_US|CIRRHOSIS; CHOLANGIOLITIC|CHOLANGIOLITIC CIRRHOSIS (DISORDER)
C1299579|T047|371139006|SNOMEDCT_US|EARLY CIRRHOSIS |EARLY CIRRHOSIS (DISORDER)
C1299579|T047|371139006|SNOMEDCT_US|EARLY CIRRHOSIS|EARLY CIRRHOSIS (DISORDER)
C1263666|T047|123717006|SNOMEDCT_US|ADVANCED CIRRHOSIS |ADVANCED CIRRHOSIS (DISORDER)
C1263666|T047|123717006|SNOMEDCT_US|ADVANCED CIRRHOSIS|ADVANCED CIRRHOSIS (DISORDER)
C1263665|T047|123716002|SNOMEDCT_US|LATENT CIRRHOSIS |LATENT CIRRHOSIS (DISORDER)
C1263665|T047|123716002|SNOMEDCT_US|LATENT CIRRHOSIS|LATENT CIRRHOSIS (DISORDER)
C1263663|T047|123605001|SNOMEDCT_US|NUTRITIONAL CIRRHOSIS |NUTRITIONAL CIRRHOSIS (DISORDER)
C1263663|T047|123605001|SNOMEDCT_US|NUTRITIONAL CIRRHOSIS|NUTRITIONAL CIRRHOSIS (DISORDER)
C1263663|T047|123605001|SNOMEDCT_US|CIRRHOSIS; NUTRITIONAL|NUTRITIONAL CIRRHOSIS (DISORDER)
C1263663|T047|123605001|SNOMEDCT_US|NUTRITIONAL; CIRRHOSIS|NUTRITIONAL CIRRHOSIS (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|PRIMARY BILIARY CIRRHOSIS|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|PRIMARY BILIARY CIRRHOSIS |BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|BILIARY CIRRHOSIS PRIMARY|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|PBC|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|BILIARY CIRRHOSIS, PRIMARY, 1|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|PRIMARY BILARY CIRRHOSIS (PBC)|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|CHRONIC NONSUPPURATIVE DESTRUCTIVE CHOLANGITIS|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|BILIARY CIRRHOSIS (& [PRIMARY]) |BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|BILIARY CIRRHOSIS|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|BILIARY CIRRHOSIS (& [PRIMARY])|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|CHRONIC NON-SUPPURATIVE DESTRUCTIVE CHOLANGITIS|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|CHOLANGITIS, CHRONIC NONSUPPURATIVE DESTRUCTIVE|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|PBC- PRIMARY BILIARY CIRRHOSIS|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|PRIMARY BILIARY CIRRHOSIS |BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|BILIARY; CIRRHOSIS, PRIMARY|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|HANOT|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|CHOLANGITIS; CHRONIC NONSUPPURATIVE DESTRUCTIVE|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|CHRONIC; CHOLANGITIS, CHRONIC NONSUPPURATIVE DESTRUCTIVE, DESTRUCTIVE|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|CIRRHOSIS; BILIARY, PRIMARY|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|BILIARY CIRRHOSIS, PRIMARY|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0008312|T047|155815006|SNOMEDCT_US|CIRRHOSIS;BILIARY;PRIMARY|BILIARY CIRRHOSIS (& [PRIMARY]) (DISORDER)
C0238065|T047|12368000|SNOMEDCT_US|OBSTRUCTIVE LIVER CIRRHOSIS|SECONDARY BILIARY CIRRHOSIS (DISORDER)
C0238065|T047|12368000|SNOMEDCT_US|SECONDARY BILIARY CIRRHOSIS|SECONDARY BILIARY CIRRHOSIS (DISORDER)
C0238065|T047|12368000|SNOMEDCT_US|SECONDARY BILIARY CIRRHOSIS |SECONDARY BILIARY CIRRHOSIS (DISORDER)
C0238065|T047|12368000|SNOMEDCT_US|BILIARY CIRRHOSIS SECONDARY|SECONDARY BILIARY CIRRHOSIS (DISORDER)
C0238065|T047|12368000|SNOMEDCT_US|LIVER CIRRHOSIS, OBSTRUCTIVE|SECONDARY BILIARY CIRRHOSIS (DISORDER)
C0238065|T047|12368000|SNOMEDCT_US|CIRRHOSIS, SECONDARY BILIARY|SECONDARY BILIARY CIRRHOSIS (DISORDER)
C0238065|T047|12368000|SNOMEDCT_US|SECONDARY BILIARY CIRRHOSIS |SECONDARY BILIARY CIRRHOSIS (DISORDER)
C0238065|T047|12368000|SNOMEDCT_US|CIRRHOSIS; BILIARY, SECONDARY|SECONDARY BILIARY CIRRHOSIS (DISORDER)
C0238065|T047|12368000|SNOMEDCT_US|BILIARY CIRRHOSIS, SECONDARY|SECONDARY BILIARY CIRRHOSIS (DISORDER)
C0400935|T047|266471006|SNOMEDCT_US|JUVENILE PORTAL CIRRHOSIS|JUVENILE PORTAL CIRRHOSIS (DISORDER)
C0400935|T047|266471006|SNOMEDCT_US|CHILDHOOD FUNCTION CIRRHOSIS|JUVENILE PORTAL CIRRHOSIS (DISORDER)
C0400935|T047|266471006|SNOMEDCT_US|JUVENILE PORTAL CIRRHOSIS |JUVENILE PORTAL CIRRHOSIS (DISORDER)
C1960179|T047|425413006|SNOMEDCT_US|DRUG-INDUCED CIRRHOSIS OF LIVER |DRUG-INDUCED HEPATIC CIRRHOSIS
C1960179|T047|425413006|SNOMEDCT_US|DRUG-INDUCED HEPATIC CIRRHOSIS|DRUG-INDUCED HEPATIC CIRRHOSIS
C1960179|T047|425413006|SNOMEDCT_US|DRUG-INDUCED CIRRHOSIS OF LIVER|DRUG-INDUCED HEPATIC CIRRHOSIS
C0400925|T047|235880004|SNOMEDCT_US|ALCOHOLIC FIBROSIS AND SCLEROSIS OF LIVER|ALCOHOLIC FIBROSIS AND SCLEROSIS OF LIVER (DISORDER)
C0400925|T047|235880004|SNOMEDCT_US|ALCOHOLIC SCLEROSIS AND FIBROSIS OF LIVER |ALCOHOLIC FIBROSIS AND SCLEROSIS OF LIVER (DISORDER)
C0400925|T047|235880004|SNOMEDCT_US|ALCOHOLIC SCLEROSIS AND FIBROSIS OF LIVER|ALCOHOLIC FIBROSIS AND SCLEROSIS OF LIVER (DISORDER)
C0400925|T047|235880004|SNOMEDCT_US|ALCOHOLIC FIBROSIS AND SCLEROSIS OF LIVER |ALCOHOLIC FIBROSIS AND SCLEROSIS OF LIVER (DISORDER)
C2887912|T047||SNOMEDCT_US|ALCOHOLIC CIRRHOSIS OF LIVER WITHOUT ASCITES
C2887913|T047||SNOMEDCT_US|ALCOHOLIC CIRRHOSIS OF LIVER WITH ASCITES
C3509286|T047||SNOMEDCT_US|CIRRHOSIS ALCOHOLIC (LAENNEC'S) WITH ASCITES
C3509286|T047||SNOMEDCT_US|ALCOHOLIC CIRRHOSIS WITH ASCITES
C3509286|T047||SNOMEDCT_US|ALCOHOLIC CIRRHOSIS WITH ASCITES 
C3838604|T047||SNOMEDCT_US|ALCOHOLIC CIRRHOSIS WITHOUT ASCITES
C3838604|T047||SNOMEDCT_US|ALCOHOLIC CIRRHOSIS WITHOUT ASCITES 
C3838604|T047||SNOMEDCT_US|CIRRHOSIS ALCOHOLIC (LAENNEC'S) WITHOUT ASCITES
C3838604|T047||SNOMEDCT_US|ALCOHOLIC (LAENNEC'S) CIRRHOSIS WITHOUT ASCITES
C1392672|T047||SNOMEDCT_US|CIRRHOSIS; MACRONODULAR, ALCOHOLIC
C1392672|T047||SNOMEDCT_US|MACRONODULAR; CIRRHOSIS, ALCOHOLIC
C1392673|T047||SNOMEDCT_US|CIRRHOSIS; MICRONODULAR, ALCOHOLIC
C1392673|T047||SNOMEDCT_US|MICRONODULAR; CIRRHOSIS, ALCOHOLIC
C1392676|T047||SNOMEDCT_US|CIRRHOSIS; PORTAL, ALCOHOLIC
C1392676|T047||SNOMEDCT_US|PORTAL; CIRRHOSIS, ALCOHOLIC
C1392677|T047||SNOMEDCT_US|CIRRHOSIS; POSTNECROTIC, ALCOHOLIC
C1392677|T047||SNOMEDCT_US|POSTNECROTIC; CIRRHOSIS, ALCOHOLIC
C1392681|T047||SNOMEDCT_US|CIRRHOSIS; NUTRITIONAL, ALCOHOL
C1392681|T047||SNOMEDCT_US|NUTRITIONAL; CIRRHOSIS, ALCOHOL
