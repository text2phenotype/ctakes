C3160090|T121|N0000182638|NDFRT|HCV NS3/4A PROTEASE INHIBITORS [MOA]|HCV NS3/4A PROTEASE INHIBITORS [MOA]
C2605855|T121|N0000191970|NDFRT|SIMEPREVIR|SIMEPREVIR [CHEMICAL/INGREDIENT]
C3696072|T121||NDFRT|SIMEPREVIR SODIUM
C3696747|T121||NDFRT|SIMEPREVIR PILL
C3696511|T121||NDFRT|SIMEPREVIR 150 MG [OLYSIO]
C3696563|T121||NDFRT|SIMEPREVIR ORAL CAPSULE [OLYSIO]
C3696697|T121||NDFRT|SIMEPREVIR 150 MG
C3696720|T121||NDFRT|SIMEPREVIR ORAL CAPSULE
C3696748|T121||NDFRT|SIMEPREVIR ORAL PRODUCT
C3695381|T121||NDFRT|SIMEPREVIR 150 MG ORAL CAPSULE [OLYSIO]
C3695403|T121|N0000189930|NDFRT|SIMEPREVIR 150 MG ORAL CAPSULE|SIMEPREVIR 150MG CAP [VA PRODUCT]
C1738934|T121||NDFRT|BOCEPREVIR
C3209784|T121||NDFRT|BOCEPREVIR PILL
C3655064|T121||NDFRT|BOCEPREVIR:SUSC:PT:ISOLATE:ORDQN:GENOTYPING
C3154647|T121||NDFRT|BOCEPREVIR 200 MG
C3154648|T121||NDFRT|BOCEPREVIR ORAL CAPSULE
C3154649|T121|N0000182825|NDFRT|BOCEPREVIR 200 MG ORAL CAPSULE|BOCEPREVIR 200MG CAP [VA PRODUCT]
C3154651|T121||NDFRT|BOCEPREVIR 200 MG [VICTRELIS]
C3154652|T121||NDFRT|BOCEPREVIR ORAL CAPSULE [VICTRELIS]
C3209783|T121||NDFRT|BOCEPREVIR ORAL PRODUCT
C3154653|T121||NDFRT|BOCEPREVIR 200 MG ORAL CAPSULE [VICTRELIS]
C1876229|T121||NDFRT|TELAPREVIR
C3215243|T121||NDFRT|TELAPREVIR PILL
C3655063|T121||NDFRT|TELAPREVIR:SUSC:PT:ISOLATE:ORDQN:GENOTYPING
C3154700|T121||NDFRT|TELAPREVIR 375 MG
C3154702|T121||NDFRT|TELAPREVIR 375 MG [INCIVEK]
C3154710|T121||NDFRT|TELAPREVIR ORAL TABLET
C3154711|T121|N0000182827|NDFRT|TELAPREVIR 375 MG ORAL TABLET|TELAPREVIR 375MG TAB,28 [VA PRODUCT]
C3154712|T121||NDFRT|TELAPREVIR ORAL TABLET [INCIVEK]
C3215242|T121||NDFRT|TELAPREVIR ORAL PRODUCT
C3655696|T121||NDFRT|TELAPREVIR ISOLATE
C3154713|T121||NDFRT|TELAPREVIR 375 MG ORAL TABLET [INCIVEK]
C0717864|T121||NDFRT|RIBAVIRIN+INTERFERON ALPHA-2B
C0789390|T121|N0000164016|NDFRT|RIBAVIRIN 200 MG ORAL TABLET|RIBAVIRIN 200MG TAB [VA PRODUCT]
C0789393|T121|N0000165356|NDFRT|RIBAVIRIN 40 MG/ML ORAL SOLUTION|RIBAVIRIN 200MG/5ML SOLN,ORAL [VA PRODUCT]
C0979999|T121|N0000156300|NDFRT|RIBAVIRIN 20 MG/ML INHALANT SOLUTION|RIBAVIRIN 6GM/VIL INHL [VA PRODUCT]
C1128545|T121||NDFRT|RIBAVIRIN 200 MG
C1131183|T121||NDFRT|RIBAVIRIN 40 MG/ML
C0035525|T121|N0000005892|NDFRT|RIBAVIRIN|RIBAVIRIN [CHEMICAL/INGREDIENT]
C0073221|T121||NDFRT|RIBAVIRIN AMIDINE
C0627880|T121||NDFRT|TRIBUTYLRIBAVIRIN
C0935908|T121||NDFRT|PALIVIZUMAB/RIBAVIRIN
C1875630|T121|N0000022295|NDFRT|PEGINTERFERON/RIBAVIRIN|PEGINTERFERON/RIBAVIRIN
C3189667|T121||NDFRT|RIBAVIRIN POWDER
C3219702|T121||NDFRT|RIBAVIRIN PILL
C3547186|T121||NDFRT|RESPONSE TO RIBAVIRIN
C0979998|T121|N0000165984|NDFRT|RIBAVIRIN 200 MG ORAL CAPSULE|RIBAVIRIN 200MG CAP [VA PRODUCT]
C0361571|T121||NDFRT|RIBAVIRIN 100 MG ORAL CAPSULE
C0413496|T121||NDFRT|TRIBAVIRIN ADVERSE REACTION
C0717864|T121||NDFRT|RIBAVIRIN+INTERFERON ALPHA-2B
C0789390|T121|N0000164016|NDFRT|RIBAVIRIN 200 MG ORAL TABLET|RIBAVIRIN 200MG TAB [VA PRODUCT]
C0789393|T121|N0000165356|NDFRT|RIBAVIRIN 40 MG/ML ORAL SOLUTION|RIBAVIRIN 200MG/5ML SOLN,ORAL [VA PRODUCT]
C0979999|T121|N0000156300|NDFRT|RIBAVIRIN 20 MG/ML INHALANT SOLUTION|RIBAVIRIN 6GM/VIL INHL [VA PRODUCT]
C1128545|T121||NDFRT|RIBAVIRIN 200 MG
C1131183|T121||NDFRT|RIBAVIRIN 40 MG/ML
C1140523|T121||NDFRT|RIBAVIRIN 20 MG/ML
C1186936|T121||NDFRT|RIBAVIRIN 100 MG
C1240752|T121||NDFRT|RIBAVIRIN ORAL CAPSULE [REBETOL]
C1242547|T121||NDFRT|RIBAVIRIN ORAL TABLET [COPEGUS]
C1247842|T121||NDFRT|RIBAVIRIN ORAL CAPSULE
C1247843|T121||NDFRT|RIBAVIRIN ORAL SOLUTION
C1247844|T121||NDFRT|RIBAVIRIN ORAL TABLET
C1253016|T121||NDFRT|RIBAVIRIN INHALANT SOLUTION
C1382829|T121||NDFRT|RIBAVIRIN 400 MG
C1454123|T121||NDFRT|5-NOR CARBOCYCLIC RIBAVIRIN
C1589272|T121||NDFRT|RIBAVIRIN ORAL SOLUTION [REBETOL]
C1593466|T121||NDFRT|RIBAVIRIN 200 MG [REBETOL]
C1593727|T121||NDFRT|RIBAVIRIN 200 MG [COPEGUS]
C1601182|T121||NDFRT|RIBAVIRIN 200 MG [RIBASPHERE]
C1601183|T121||NDFRT|RIBAVIRIN ORAL CAPSULE [RIBASPHERE]
C1621221|T121||NDFRT|RIBAVIRIN INHALANT SOLUTION [VIRAZOLE]
C1626919|T121|N0000177127|NDFRT|RIBAVIRIN 400 MG ORAL TABLET|RIBAVIRIN 400MG TAB [VA PRODUCT]
C1641488|T121||NDFRT|RIBAVIRIN:MCNC:PT:SER/PLAS:QN
C1676705|T121|N0000177128|NDFRT|RIBAVIRIN 600 MG ORAL TABLET|RIBAVIRIN 600MG TAB [VA PRODUCT]
C1677789|T121||NDFRT|RIBAVIRIN 600 MG
C1694682|T121||NDFRT|RIBAVIRIN ORAL TABLET [RIBATAB]
C1702720|T121||NDFRT|RIBAVIRIN 400 MG [RIBASPHERE]
C1703270|T121||NDFRT|RIBAVIRIN 600 MG [RIBASPHERE]
C1704170|T121||NDFRT|RIBAVIRIN ORAL TABLET [RIBASPHERE]
C1878904|T121||NDFRT|RIBAVIRIN 400 MG [RIBATAB]
C1589271|T121||NDFRT|RIBAVIRIN 40 MG/ML [REBETOL]
C1616510|T121||NDFRT|RIBAVIRIN 20 MG/ML [VIRAZOLE]
C0733470|T121||NDFRT|HUMAN LEUKOCYTE INTERFERON
C3652465|T121||NDFRT|CONSDER REMOVING IF YOU GET TOO MANY FALSE POSITIVES AND ONLY INCLUDING INTERFERON AND RIBAVIRIN COMBINATIONS
C3653501|T121||NDFRT|DIRECT ACTING ANTIVIRALS
C3541967|T121||NDFRT|THIOSEMICARBAZONES, DIRECT ACTING ANTIVIRALS
C3653501|T121||NDFRT|DIRECT ACTING ANTIVIRALS
C3540755|T121||NDFRT|PROTEASE INHIBITORS, DIRECT ACTING ANTIVIRALS
C3541969|T121||NDFRT|NEURAMINIDASE INHIBITORS, DIRECT ACTING ANTIVIRALS
C3653443|T121||NDFRT|CYCLIC AMINES, DIRECT ACTING ANTIVIRALS
C3653392|T121||NDFRT|PHOSPHONIC ACID DERIVATIVES, DIRECT ACTING ANTIVIRALS
C0330845|T121||NDFRT|ASTRAGALUS PLANT
C1095897|T121|N0000022270|NDFRT|ASTRAGALUS PREPARATION|ASTRAGALUS
C3864824|T121||NDFRT|PARITAPREVIR
C3864824|T121||NDFRT|PARITAPREVIR
C3883274|T121||NDFRT|PARITAPREVIR DIHYDRATE
C3864967|T121||NDFRT|OMBITASVIR / PARITAPREVIR / RITONAVIR
C3865150|T121||NDFRT|PARITAPREVIR 75 MG
C3865210|T121||NDFRT|OMBITASVIR / PARITAPREVIR / RITONAVIR PILL
C3882783|T121||NDFRT|DASABUVIR / OMBITASVIR / PARITAPREVIR / RITONAVIR
C4075296|T121||NDFRT|PARITAPREVIR IN ORAL DOSAGE FORM
C4276327|T121||NDFRT|PARITAPREVIR 50 MG
C4298645|T121||NDFRT|PARITAPREVIR:SUSC:PT:ISOLATE:ORD:GENOTYPING
C3865188|T121||NDFRT|OMBITASVIR / PARITAPREVIR / RITONAVIR ORAL TABLET
C3865211|T121||NDFRT|OMBITASVIR / PARITAPREVIR / RITONAVIR ORAL PRODUCT
C4276383|T121||NDFRT|DASABUVIR / OMBITASVIR / PARITAPREVIR / RITONAVIR PILL
C3864964|T121|N0000191861|NDFRT|{2 (DASABUVIR 250 MG ORAL TABLET) / 2 (OMBITASVIR 12.5 MG / PARITAPREVIR 75 MG / RITONAVIR 50 MG ORAL TABLET) } PACK|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DOSE PACK,56 [VA PRODUCT]
C3871501|T121||NDFRT|DASABUVIR;OMBITASVIR, PARITAPREVIR, RITONAVIR ORAL TABLET
C3871617|T121||NDFRT|DASABUVIR;OMBITASVIR/PARITAPREVIR/RITONAVIR NA ORAL TABLET
C3882779|T121||NDFRT|DASABUVIR/OMBITASVIR/PARITAPREVIR/RITONAVIR ORAL KIT
C4047040|T121||NDFRT|OMBITASVIR / PARITAPREVIR / RITONAVIR ORAL TABLET [TECHNIVIE]
C4276384|T121||NDFRT|DASABUVIR / OMBITASVIR / PARITAPREVIR / RITONAVIR ORAL PRODUCT
C3854281|T121||NDFRT|{2 (DASABUVIR 250 MG ORAL TABLET) / 2 (OMBITASVIR 12.5 MG / PARITAPREVIR 75 MG / RITONAVIR 50 MG ORAL TABLET) } PACK [VIEKIRA PAK]
C3865125|T121|N0000192214|NDFRT|OMBITASVIR 12.5 MG / PARITAPREVIR 75 MG / RITONAVIR 50 MG ORAL TABLET|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DAILY PACK [VA PRODUCT]
C4046961|T121||NDFRT|OMBITASVIR 12.5 MG / PARITAPREVIR 75 MG / RITONAVIR 50 MG [TECHNIVIE]
C4276118|T121|N0000192787|NDFRT|DASABUVIR 200 MG / OMBITASVIR 8.33 MG / PARITAPREVIR 50 MG / RITONAVIR 33.33 MG EXTENDED RELEASE ORAL TABLET (3) 24HR PACK|DASABUVIR/OMBITASVIR/PARITAPREVIR/RITONAVIR TAB,SA DAILY PACK [VA PRODUCT]
C4276368|T121||NDFRT|DASABUVIR / OMBITASVIR / PARITAPREVIR / RITONAVIR EXTENDED RELEASE ORAL TABLET
C4046169|T121||NDFRT|OMBITASVIR 12.5 MG / PARITAPREVIR 75 MG / RITONAVIR 50 MG ORAL TABLET [TECHNIVIE]
C4275375|T121||NDFRT|24 HR DASABUVIR 200 MG / OMBITASVIR 8.33 MG / PARITAPREVIR 50 MG / RITONAVIR 33.33 MG EXTENDED RELEASE ORAL TABLET
C3696409|T121||NDFRT|OLYSIO
C3696630|T121||NDFRT|OLYSIO PILL
C3695381|T121||NDFRT|SIMEPREVIR 150 MG ORAL CAPSULE [OLYSIO]
C3696511|T121||NDFRT|SIMEPREVIR 150 MG [OLYSIO]
C3696563|T121||NDFRT|SIMEPREVIR ORAL CAPSULE [OLYSIO]
C3696631|T121||NDFRT|OLYSIO ORAL PRODUCT
C4080053|T121||NDFRT|GRAZOPREVIR
C4080453|T121||NDFRT|ELBASVIR / GRAZOPREVIR
C4255551|T121||NDFRT|GRAZOPREVIR ANHYDROUS
C4080449|T121||NDFRT|GRAZOPREVIR 100 MG
C4080450|T121||NDFRT|ELBASVIR / GRAZOPREVIR ORAL PRODUCT
C4080451|T121||NDFRT|ELBASVIR / GRAZOPREVIR PILL
C4080452|T121||NDFRT|ELBASVIR / GRAZOPREVIR ORAL TABLET
C4298643|T121||NDFRT|GRAZOPREVIR:SUSC:PT:ISOLATE:ORD:GENOTYPING
C4307658|T121||NDFRT|ELBASVIR-GRAZOPREVIR DRUG COMBINATION
C4080454|T121|N0000192438|NDFRT|ELBASVIR 50 MG / GRAZOPREVIR 100 MG ORAL TABLET|ELBASVIR 50MG/GRAZOPREVIR 100MG TAB [VA PRODUCT]
C4080457|T121||NDFRT|ELBASVIR / GRAZOPREVIR ORAL TABLET [ZEPATIER]
C4080456|T121||NDFRT|ELBASVIR 50 MG / GRAZOPREVIR 100 MG [ZEPATIER]
C4080460|T121||NDFRT|ELBASVIR 50 MG / GRAZOPREVIR 100 MG ORAL TABLET [ZEPATIER]
C3854280|T121||NDFRT|VIEKIRA PAK
C2976303|T121|N0000191981|NDFRT|SOFOSBUVIR|SOFOSBUVIR [CHEMICAL/INGREDIENT]
C3857383|T121||NDFRT|LEDIPASVIR
C3858025|T121||NDFRT|HARVONI
C3858199|T121||NDFRT|HARVONI PILL
C3858200|T121||NDFRT|HARVONI ORAL PRODUCT
C3852670|T121||NDFRT|OMBITASVIR
C3854280|T121||NDFRT|VIEKIRA PAK
C4080455|T121||NDFRT|ZEPATIER
C4080052|T121||NDFRT|ELBASVIR
C4299883|T121||NDFRT|ELBASVIR
C4080453|T121||NDFRT|ELBASVIR GRAZOPREVIR
C4080453|T121||NDFRT|GRAZOPREVIR
C3252090|T121||NDFRT|DACLATASVIR
C3892852|T121||NDFRT|DACLATASVIR DIHYDROCHLORIDE
C4047229|T121||NDFRT|DACLATASVIR PILL
C4298749|T121||NDFRT|DACLATASVIR
C4299898|T121||NDFRT|DACLATASVIR
C3851350|T121||NDFRT|LEDIPASVIR
C3858051|T121||NDFRT|LEDIPASVIR / SOFOSBUVIR
C3858262|T121||NDFRT|LEDIPASVIR 90 MG
C3858300|T121||NDFRT|LEDIPASVIR / SOFOSBUVIR ORAL TABLET
C3858321|T121||NDFRT|LEDIPASVIR / SOFOSBUVIR PILL
C3858322|T121||NDFRT|LEDIPASVIR / SOFOSBUVIR ORAL PRODUCT
C4075037|T121||NDFRT|LEDIPASVIR IN ORAL DOSAGE FORM
C4298751|T121||NDFRT|LEDIPASVIR:SUSC:PT:ISOLATE:ORD:GENOTYPING
C4299632|T121||NDFRT| ISOLATE
C3858080|T121|N0000191202|NDFRT|LEDIPASVIR 90 MG / SOFOSBUVIR 400 MG ORAL TABLET|LEDIPASVIR 90MG/SOFOSBUVIR 400MG TAB [VA PRODUCT]
C3858162|T121||NDFRT|LEDIPASVIR / SOFOSBUVIR ORAL TABLET [HARVONI]
C3858113|T121||NDFRT|LEDIPASVIR 90 MG / SOFOSBUVIR 400 MG [HARVONI]
C3857383|T121||NDFRT|LEDIPASVIR 90 MG / SOFOSBUVIR 400 MG ORAL TABLET [HARVONI]
C2605856|T121||NDFRT|435350, TMC
C2605856|T121||NDFRT|TMC435350
C2605856|T121||NDFRT|TMC-435350
C2605856|T121||NDFRT|TMC 435350
C2745868|T121||NDFRT|435, TMC
C2745868|T121||NDFRT|TMC435
C2745868|T121||NDFRT|TMC-435
C2745868|T121||NDFRT|TMC 435
C3696409|T121||NDFRT|OLYSIO
C2605855|T121|N0000191970|NDFRT|SIMEPREVIR|SIMEPREVIR [CHEMICAL/INGREDIENT]
C2605855|T121|N0000191970|NDFRT|SIMEPREVIR |SIMEPREVIR [CHEMICAL/INGREDIENT]
C2605855|T121|N0000191970|NDFRT|ANTIVIRAL SIMEPREVIR|SIMEPREVIR [CHEMICAL/INGREDIENT]
C2605855|T121|N0000191970|NDFRT|SIMEPREVIR |SIMEPREVIR [CHEMICAL/INGREDIENT]
C2605855|T121|N0000191970|NDFRT|N-(17-(2-(4-ISOPROPYLTHIAZOLE-2-YL)-7-METHOXY-8-METHYLQUINOLIN-4-YLOXY)-13-METHYL-2,14-DIOXO-3,13-DIAZATRICYCLO(13.3.0.04,6)OCTADEC-7-ENE-4-CARBONYL)(CYCLOPROPYL)SULFONAMIDE|SIMEPREVIR [CHEMICAL/INGREDIENT]
C2605855|T121|N0000191970|NDFRT|SIMEPREVIR [CHEMICAL/INGREDIENT]|SIMEPREVIR [CHEMICAL/INGREDIENT]
C2605855|T121|N0000191970|NDFRT|SIMEPREVIR |SIMEPREVIR [CHEMICAL/INGREDIENT]
C3696072|T121||NDFRT|SIMEPREVIR SODIUM
C3696072|T121||NDFRT|SIMEPREVIR (AS SODIUM)
C3696748|T121||NDFRT|SIMEPREVIR ORAL PRODUCT
C3696748|T121||NDFRT|ORAL FORM SIMEPREVIR 
C3696748|T121||NDFRT|ORAL FORM SIMEPREVIR
C4075528|T121||NDFRT|SIMEPREVIR + SOFOSBUVIR 
C4075528|T121||NDFRT|SIMEPREVIR + SOFOSBUVIR
C3696720|T121||NDFRT|SIMEPREVIR ORAL CAPSULE
C3696630|T121||NDFRT|OLYSIO PILL
C3695403|T121|N0000189930|NDFRT|SIMEPREVIR 150 MG ORAL CAPSULE|SIMEPREVIR 150MG CAP [VA PRODUCT]
C3695403|T121|N0000189930|NDFRT|SIMEPREVIR 150MG ORAL CAPSULE|SIMEPREVIR 150MG CAP [VA PRODUCT]
C3695403|T121|N0000189930|NDFRT|SIMEPREVIR SODIUM CAP 150 MG (BASE EQUIVALENT)|SIMEPREVIR 150MG CAP [VA PRODUCT]
C3695403|T121|N0000189930|NDFRT|SIMEPREVIR 150MG CAP|SIMEPREVIR 150MG CAP [VA PRODUCT]
C3695403|T121|N0000189930|NDFRT|SIMEPREVIR 150MG CAP [VA PRODUCT]|SIMEPREVIR 150MG CAP [VA PRODUCT]
C3695381|T121||NDFRT|SIMEPREVIR 150 MG ORAL CAPSULE [OLYSIO]
C3695381|T121||NDFRT|OLYSIO 150 MG ORAL CAPSULE
C3695381|T121||NDFRT|OLYSIO 150MG CAPSULE
C3695381|T121||NDFRT|SIMEPREVIR 150 MG (AS SIMEPREVIR SODIUM 154.4 MG ) ORAL CAPSULE [OLYSIO]
C3695381|T121||NDFRT|OLYSIO, 150 MG ORAL CAPSULE
C3696511|T121||NDFRT|SIMEPREVIR 150 MG [OLYSIO]
C3696563|T121||NDFRT|SIMEPREVIR ORAL CAPSULE [OLYSIO]
C3696631|T121||NDFRT|OLYSIO ORAL PRODUCT
C3154650|T121||NDFRT|VICTRELIS
C3154650|T121||NDFRT|VICRTELIS
C1738934|T121||NDFRT|N-(3-AMINO-1-(CYCLOBUTYLMETHYL)-2,3-DIOXOPROPYL)-3-(2-((((1,1-DIMETHYLETHYL)AMINO)CARBONYL)AMINO)-3,3-DIMETHYL-1-OXOBUTYL)-6,6-DIMETHYL-3-AZABICYCLO(3.1.0)HEXAN-2-CARBOXAMIDE
C1738934|T121||NDFRT|BOCEPREVIR
C1738934|T121||NDFRT|ANTIVIRALS BOCEPREVIR
C1738934|T121||NDFRT|ANTIVIRALS BOCEPREVIR 
C1738934|T121||NDFRT|BOCEPREVIR 
C1738934|T121||NDFRT|BOCEPREVIR 
C1738934|T121||NDFRT|3-AZABICYCLO(3.1.0)HEXANE-2-CARBOXAMIDE, N-(3-AMINO-1-(CYCLOBUTYLMETHYL)-2,3-DIOXOPROPYL)-3-((2S)-2-((((1,1- DIMETHYLETHYL)AMINO)CARBONYL)AMINO)-3,3-DIMETHYL-1-OXOBUTYL)-6,6- DIMETHYL-, (1R,2S,5S)-
C3154649|T121|N0000182825|NDFRT|BOCEPREVIR CAP 200 MG|BOCEPREVIR 200MG CAP [VA PRODUCT]
C3154649|T121|N0000182825|NDFRT|BOCEPREVIR 200MG CAP|BOCEPREVIR 200MG CAP [VA PRODUCT]
C3154649|T121|N0000182825|NDFRT|BOCEPREVIR 200 MG ORAL CAPSULE|BOCEPREVIR 200MG CAP [VA PRODUCT]
C3154649|T121|N0000182825|NDFRT|BOCEPREVIR 200MG CAP [VA PRODUCT]|BOCEPREVIR 200MG CAP [VA PRODUCT]
C3154649|T121|N0000182825|NDFRT|BOCEPREVIR 200MG ORAL CAPSULE|BOCEPREVIR 200MG CAP [VA PRODUCT]
C3154649|T121|N0000182825|NDFRT|BOCEPREVIR 200MG CAPSULE |BOCEPREVIR 200MG CAP [VA PRODUCT]
C3154649|T121|N0000182825|NDFRT|BOCEPREVIR 200MG CAPSULE|BOCEPREVIR 200MG CAP [VA PRODUCT]
C1741239|T121||NDFRT|SCH-503034
C1741239|T121||NDFRT|SCH 503034
C1741239|T121||NDFRT|SCH503034
C3896865|T121||NDFRT|EBP 520
C3240332|T121||NDFRT|VICTRELIS PILL
C3154648|T121||NDFRT|BOCEPREVIR ORAL CAPSULE
C3655064|T121||NDFRT|BOCEPREVIR:SUSC:PT:ISOLATE:ORDQN:GENOTYPING
C3655064|T121||NDFRT|BOCEPREVIR [SUSCEPTIBILITY] BY GENOTYPE METHOD
C3655064|T121||NDFRT|BOCEPREVIR ISLT GENOTYP
C3655064|T121||NDFRT|BOCEPREVIR:SUSCEPTIBILITY:POINT IN TIME:ISOLATE:QUANTITATIVE OR ORDINAL:GENOTYPING
C3154651|T121||NDFRT|BOCEPREVIR 200 MG [VICTRELIS]
C3154652|T121||NDFRT|BOCEPREVIR ORAL CAPSULE [VICTRELIS]
C3154653|T121||NDFRT|BOCEPREVIR 200 MG ORAL CAPSULE [VICTRELIS]
C3154653|T121||NDFRT|VICTRELIS 200 MG ORAL CAPSULE
C3154653|T121||NDFRT|VICTRELIS 200MG CAPSULE
C3154653|T121||NDFRT|VICTRELIS, 200 MG ORAL CAPSULE
C3240331|T121||NDFRT|VICTRELIS ORAL PRODUCT
C3154701|T121||NDFRT|INCIVEK
C1876229|T121||NDFRT|TELAPREVIR
C1876229|T121||NDFRT|ANTIVIRAL TELAPREVIR
C1876229|T121||NDFRT|ANTIVIRAL TELAPREVIR 
C1876229|T121||NDFRT|TELAPREVIR 
C1876229|T121||NDFRT|TELAPREVIR 
C3281323|T121||NDFRT|VRT-111950
C3281324|T121||NDFRT|MP-424
C3281325|T121||NDFRT|LY-570310
C1956374|T121||NDFRT|VX-950
C1956374|T121||NDFRT|VX 950
C1956374|T121||NDFRT|VX950 CPD
C3154711|T121|N0000182827|NDFRT|TELAPREVIR 375 MG ORAL TABLET|TELAPREVIR 375MG TAB,28 [VA PRODUCT]
C3154711|T121|N0000182827|NDFRT|TELAPREVIR TAB 375 MG|TELAPREVIR 375MG TAB,28 [VA PRODUCT]
C3154711|T121|N0000182827|NDFRT|TELAPREVIR 375MG TAB|TELAPREVIR 375MG TAB,28 [VA PRODUCT]
C3154711|T121|N0000182827|NDFRT|TELAPREVIR 375MG TAB,28 [VA PRODUCT]|TELAPREVIR 375MG TAB,28 [VA PRODUCT]
C3154711|T121|N0000182827|NDFRT|TELAPREVIR 375MG TAB,28|TELAPREVIR 375MG TAB,28 [VA PRODUCT]
C3154711|T121|N0000182827|NDFRT|TELAPREVIR 375MG TAB [VA PRODUCT]|TELAPREVIR 375MG TAB,28 [VA PRODUCT]
C3154711|T121|N0000182827|NDFRT|TELAPREVIR 375MG ORAL TABLET|TELAPREVIR 375MG TAB,28 [VA PRODUCT]
C3154711|T121|N0000182827|NDFRT|TELAPREVIR 375MG TAB,UD|TELAPREVIR 375MG TAB,28 [VA PRODUCT]
C3154711|T121|N0000182827|NDFRT|TELAPREVIR 375MG UD TAB|TELAPREVIR 375MG TAB,28 [VA PRODUCT]
C3154711|T121|N0000182827|NDFRT|TELAPREVIR 375MG TAB,UD [VA PRODUCT]|TELAPREVIR 375MG TAB,28 [VA PRODUCT]
C3154711|T121|N0000182827|NDFRT|TELAPREVIR 375MG TABLET|TELAPREVIR 375MG TAB,28 [VA PRODUCT]
C3154711|T121|N0000182827|NDFRT|TELAPREVIR 375MG TABLET |TELAPREVIR 375MG TAB,28 [VA PRODUCT]
C3226078|T121||NDFRT|INCIVEK PILL
C3154710|T121||NDFRT|TELAPREVIR ORAL TABLET
C3655063|T121||NDFRT|TELAPREVIR ISLT GENOTYP
C3655063|T121||NDFRT|TELAPREVIR [SUSCEPTIBILITY] BY GENOTYPE METHOD
C3655063|T121||NDFRT|TELAPREVIR:SUSC:PT:ISOLATE:ORDQN:GENOTYPING
C3655063|T121||NDFRT|TELAPREVIR:SUSCEPTIBILITY:POINT IN TIME:ISOLATE:QUANTITATIVE OR ORDINAL:GENOTYPING
C3154702|T121||NDFRT|TELAPREVIR 375 MG [INCIVEK]
C3154712|T121||NDFRT|TELAPREVIR ORAL TABLET [INCIVEK]
C3154713|T121||NDFRT|TELAPREVIR 375 MG ORAL TABLET [INCIVEK]
C3154713|T121||NDFRT|INCIVEK 375 MG ORAL TABLET
C3154713|T121||NDFRT|INCIVEK 375MG TABLET
C3154713|T121||NDFRT|INCIVEK, 375 MG ORAL TABLET
C3154713|T121||NDFRT|INCIVEK 375 MG ORAL TABLET, TWICE DAILY
C3226077|T121||NDFRT|INCIVEK ORAL PRODUCT
C0979954|T121|N0000165884|NDFRT|REBETRON, SINGLE DOSE 1000 MG/DAY ORAL AND INJECTABLE KIT|REBETRON 1000/PAK 3 PKT (1241-02) [VA PRODUCT]
C0979954|T121|N0000165884|NDFRT|REBETRON 1000/PAK 3 PKT (1241-02)|REBETRON 1000/PAK 3 PKT (1241-02) [VA PRODUCT]
C0979954|T121|N0000165884|NDFRT|REBETRON COMBINATION PACKAGE FOR PATIENTS < = 75 KG, INTRON A 6,000,000 UNT/ML SINGLE DOSE VIALS / 70 REBETOL CAPSULES|REBETRON 1000/PAK 3 PKT (1241-02) [VA PRODUCT]
C0979954|T121|N0000165884|NDFRT|REBETRON 1000/PAK 3 PKT (1241-02) [VA PRODUCT]|REBETRON 1000/PAK 3 PKT (1241-02) [VA PRODUCT]
C0979954|T121|N0000165884|NDFRT|{6 (0.5 ML) (INTERFERON ALFA-2B 6000000 UNT/ML INJECTABLE SOLUTION [INTRON A]) / 70 (RIBAVIRIN 200 MG ORAL CAPSULE [REBETOL]) } PACK [REBETRON COMBINATION PACKAGE FOR PATIENTS < = 75 KG, INTRON A 6,000,000 UNT/ML SINGLE DOSE VIALS / 70 REBETOL CAPSULES]|REBETRON 1000/PAK 3 PKT (1241-02) [VA PRODUCT]
C0979953|T121|N0000165885|NDFRT|REBETRON COMBINATION PACKAGE FOR PATIENTS < = 75 KG, INTRON A 6,000,000 UNT/ML MULTI-DOSE VIAL / 70 REBETOL CAPSULES|REBETRON 1000/MDV PKT (1236-02) [VA PRODUCT]
C0979953|T121|N0000165885|NDFRT|REBETRON 1000/MDV PKT (1236-02)|REBETRON 1000/MDV PKT (1236-02) [VA PRODUCT]
C0979953|T121|N0000165885|NDFRT|REBETRON 1000/MDV PKT (1236-02) [VA PRODUCT]|REBETRON 1000/MDV PKT (1236-02) [VA PRODUCT]
C0979953|T121|N0000165885|NDFRT|{1 (3 ML) (INTERFERON ALFA-2B 6000000 UNT/ML INJECTABLE SOLUTION [INTRON A]) / 70 (RIBAVIRIN 200 MG ORAL CAPSULE [REBETOL]) } PACK [REBETRON COMBINATION PACKAGE FOR PATIENTS < = 75 KG, INTRON A 6,000,000 UNT/ML MULTI-DOSE VIAL / 70 REBETOL CAPSULES]|REBETRON 1000/MDV PKT (1236-02) [VA PRODUCT]
C0979955|T121|N0000165886|NDFRT|REBETRON 1000/PEN PKT (1258-02)|REBETRON 1000/PEN PKT (1258-02) [VA PRODUCT]
C0979955|T121|N0000165886|NDFRT|REBETRON COMBINATION PACKAGE FOR PATIENTS < = 75 KG, INTRON A 15,000,000 UNT/ML MULTI-DOSE PEN / 70 REBETOL CAPSULES|REBETRON 1000/PEN PKT (1258-02) [VA PRODUCT]
C0979955|T121|N0000165886|NDFRT|REBETRON 1000/PEN PKT (1258-02) [VA PRODUCT]|REBETRON 1000/PEN PKT (1258-02) [VA PRODUCT]
C0979955|T121|N0000165886|NDFRT|{1 (1.2 ML) (INTERFERON ALFA-2B 15000000 UNT/ML INJECTABLE SOLUTION [INTRON A]) / 70 (RIBAVIRIN 200 MG ORAL CAPSULE [REBETOL]) } PACK [REBETRON COMBINATION PACKAGE FOR PATIENTS < = 75 KG, INTRON A 15,000,000 UNT/ML MULTI-DOSE PEN / 70 REBETOL CAPSULES]|REBETRON 1000/PEN PKT (1258-02) [VA PRODUCT]
C0979955|T121|N0000165886|NDFRT|INTERFERON ALFA-2B;RIBAVIRIN 3MILLION IU/0.2ML-200MG MULTIPLE ROUTES KIT [REBETRON 1000]|REBETRON 1000/PEN PKT (1258-02) [VA PRODUCT]
C0979957|T121|N0000165887|NDFRT|REBETRON, SINGLE DOSE 1200 MG/DAY ORAL AND INJECTABLE KIT|REBETRON 1200/PAK 3 PKT (1241-01) [VA PRODUCT]
C0979957|T121|N0000165887|NDFRT|REBETRON COMBINATION PACKAGE FOR PATIENTS > = 75 KG, INTRON A 6,000,000 UNT/ML SINGLE DOSE VIALS / 84 REBETOL CAPSULES|REBETRON 1200/PAK 3 PKT (1241-01) [VA PRODUCT]
C0979957|T121|N0000165887|NDFRT|REBETRON 1200/PAK 3 PKT (1241-01)|REBETRON 1200/PAK 3 PKT (1241-01) [VA PRODUCT]
C0979957|T121|N0000165887|NDFRT|REBETRON 1200/PAK 3 PKT (1241-01) [VA PRODUCT]|REBETRON 1200/PAK 3 PKT (1241-01) [VA PRODUCT]
C0979957|T121|N0000165887|NDFRT|{6 (0.5 ML) (INTERFERON ALFA-2B 6000000 UNT/ML INJECTABLE SOLUTION [INTRON A]) / 84 (RIBAVIRIN 200 MG ORAL CAPSULE [REBETOL]) } PACK [REBETRON COMBINATION PACKAGE FOR PATIENTS > = 75 KG, INTRON A 6,000,000 UNT/ML SINGLE DOSE VIALS / 84 REBETOL CAPSULES]|REBETRON 1200/PAK 3 PKT (1241-01) [VA PRODUCT]
C2342666|T121|N0000165889|NDFRT|REBETRON 1200/PEN PKT (1258-01)|REBETRON 1200/PEN PKT (1258-01) [VA PRODUCT]
C2342666|T121|N0000165889|NDFRT|REBETRON COMBINATION PACKAGE FOR PATIENTS > = 75 KG, INTRON A 15,000,000 UNT/ML MULTI-DOSE PEN / 84 REBETOL CAPSULES|REBETRON 1200/PEN PKT (1258-01) [VA PRODUCT]
C2342666|T121|N0000165889|NDFRT|{1 (1.2 ML INTERFERON ALFA-2B 15000000 UNT/ML INJECTABLE SOLUTION [INTRON A]) / 84 (RIBAVIRIN 200 MG ORAL CAPSULE [REBETOL]) } PACK [REBETRON COMBINATION PACKAGE FOR PATIENTS > = 75 KG, INTRON A 15,000,000 UNT/ML MULTI-DOSE PEN / 84 REBETOL CAPSULES]|REBETRON 1200/PEN PKT (1258-01) [VA PRODUCT]
C2342666|T121|N0000165889|NDFRT|REBETRON 1200/PEN PKT (1258-01) [VA PRODUCT]|REBETRON 1200/PEN PKT (1258-01) [VA PRODUCT]
C2342666|T121|N0000165889|NDFRT|{1 (1.2 ML) (INTERFERON ALFA-2B 15000000 UNT/ML INJECTABLE SOLUTION [INTRON A]) / 84 (RIBAVIRIN 200 MG ORAL CAPSULE [REBETOL]) } PACK [REBETRON COMBINATION PACKAGE FOR PATIENTS > = 75 KG, INTRON A 15,000,000 UNT/ML MULTI-DOSE PEN / 84 REBETOL CAPSULES]|REBETRON 1200/PEN PKT (1258-01) [VA PRODUCT]
C2342666|T121|N0000165889|NDFRT|INTERFERON ALFA-2B;RIBAVIRIN 3MILLION IU/0.2ML-200MG MULTIPLE ROUTES KIT [REBETRON 1200]|REBETRON 1200/PEN PKT (1258-01) [VA PRODUCT]
C0979959|T121|N0000165891|NDFRT|REBETRON, MULTIPLE DOSE 600 MG/DAY ORAL AND INJECTABLE KIT|REBETRON 600/MDV PKT (1236-03) [VA PRODUCT]
C0979959|T121|N0000165891|NDFRT|REBETRON COMBINATION PACKAGE FOR REBETOL DOSE REDUCTION, INTRON A 6,000,000 UNT/ML MULTI-DOSE VIAL / 42 REBETOL CAPSULES|REBETRON 600/MDV PKT (1236-03) [VA PRODUCT]
C0979959|T121|N0000165891|NDFRT|REBETRON 600/MDV PKT (1236-03)|REBETRON 600/MDV PKT (1236-03) [VA PRODUCT]
C0979959|T121|N0000165891|NDFRT|REBETRON 600/MDV PKT (1236-03) [VA PRODUCT]|REBETRON 600/MDV PKT (1236-03) [VA PRODUCT]
C0979959|T121|N0000165891|NDFRT|{1 (3 ML INTERFERON ALFA-2B 6000000 UNT/ML INJECTABLE SOLUTION [INTRON A]) / 42 (RIBAVIRIN 200 MG ORAL CAPSULE [REBETOL]) } PACK [REBETRON COMBINATION PACKAGE FOR REBETOL DOSE REDUCTION, INTRON A 6,000,000 UNT/ML MULTI-DOSE VIAL / 42 REBETOL CAPSULES]|REBETRON 600/MDV PKT (1236-03) [VA PRODUCT]
C0979959|T121|N0000165891|NDFRT|{1 (3 ML) (INTERFERON ALFA-2B 6000000 UNT/ML INJECTABLE SOLUTION [INTRON A]) / 42 (RIBAVIRIN 200 MG ORAL CAPSULE [REBETOL]) } PACK [REBETRON COMBINATION PACKAGE FOR REBETOL DOSE REDUCTION, INTRON A 6,000,000 UNT/ML MULTI-DOSE VIAL / 42 REBETOL CAPSULES]|REBETRON 600/MDV PKT (1236-03) [VA PRODUCT]
C0979959|T121|N0000165891|NDFRT|INTERFERON ALFA-2B;RIBAVIRIN 3MILLION IU/0.2ML-200MG MULTIPLE ROUTES KIT [REBETRON 600]|REBETRON 600/MDV PKT (1236-03) [VA PRODUCT]
C2342670|T121|N0000165892|NDFRT|REBETRON COMBINATION PACKAGE FOR REBETOL DOSE REDUCTION, INTRON A 15,000,000 UNT/ML MULTI-DOSE PEN / 42 REBETOL CAPSULES|REBETRON 600/PEN PKT (1258-03) [VA PRODUCT]
C2342670|T121|N0000165892|NDFRT|REBETRON 600/PEN PKT (1258-03)|REBETRON 600/PEN PKT (1258-03) [VA PRODUCT]
C2342670|T121|N0000165892|NDFRT|REBETRON 600/PEN PKT (1258-03) [VA PRODUCT]|REBETRON 600/PEN PKT (1258-03) [VA PRODUCT]
C2342670|T121|N0000165892|NDFRT|{1 (1.2 ML INTERFERON ALFA-2B 15000000 UNT/ML INJECTABLE SOLUTION [INTRON A]) / 42 (RIBAVIRIN 200 MG ORAL CAPSULE [REBETOL]) } PACK [REBETRON COMBINATION PACKAGE FOR REBETOL DOSE REDUCTION, INTRON A 15,000,000 UNT/ML MULTI-DOSE PEN / 42 REBETOL CAPSULES]|REBETRON 600/PEN PKT (1258-03) [VA PRODUCT]
C2342670|T121|N0000165892|NDFRT|{1 (1.2 ML) (INTERFERON ALFA-2B 15000000 UNT/ML INJECTABLE SOLUTION [INTRON A]) / 42 (RIBAVIRIN 200 MG ORAL CAPSULE [REBETOL]) } PACK [REBETRON COMBINATION PACKAGE FOR REBETOL DOSE REDUCTION, INTRON A 15,000,000 UNT/ML MULTI-DOSE PEN / 42 REBETOL CAPSULES]|REBETRON 600/PEN PKT (1258-03) [VA PRODUCT]
C1444872|T121||NDFRT|RIBAVIRIN 200MG CAPSULE+INTERFERON ALPHA-2B 3MILLION IU/VIAL INJECTION SOLUTION 
C1444872|T121||NDFRT|RIBAVIRIN 200MG CAPSULE+INTERFERON ALPHA-2B 3MILLION IU/VIAL INJECTION SOLUTION
C0705810|T121||NDFRT|INTERFERON ALFA-2B-RIBAVIRIN SINGLE DOSE 1000 MG/DAY ORAL AND INJECTABLE KIT
C0705812|T121||NDFRT|INTERFERON ALFA-2B-RIBAVIRIN SINGLE DOSE 600 MG/DAY ORAL AND INJECTABLE KIT
C0705811|T121||NDFRT|INTERFERON ALFA-2B-RIBAVIRIN SINGLE DOSE 1200 MG/DAY ORAL AND INJECTABLE KIT
C0789390|T121|N0000164016|NDFRT|RIBAVIRIN 200 MG ORAL TABLET|RIBAVIRIN 200MG TAB [VA PRODUCT]
C0789390|T121|N0000164016|NDFRT|RIBAVIRIN 200MG ORAL TABLET|RIBAVIRIN 200MG TAB [VA PRODUCT]
C0789390|T121|N0000164016|NDFRT|RIBAVIRIN 200MG TAB|RIBAVIRIN 200MG TAB [VA PRODUCT]
C0789390|T121|N0000164016|NDFRT|RIBAVIRIN TAB 200 MG|RIBAVIRIN 200MG TAB [VA PRODUCT]
C0789390|T121|N0000164016|NDFRT|RIBAVIRIN 200 MG ORAL TABLET, FILM COATED|RIBAVIRIN 200MG TAB [VA PRODUCT]
C0789390|T121|N0000164016|NDFRT|RIBAVIRIN 200MG TAB [VA PRODUCT]|RIBAVIRIN 200MG TAB [VA PRODUCT]
C0789390|T121|N0000164016|NDFRT|RIBAVIRIN 200 MG ORAL TABLET, FILM COATED [RIBAVIRIN]|RIBAVIRIN 200MG TAB [VA PRODUCT]
C0789390|T121|N0000164016|NDFRT|RIBAVIRIN 200MG TABLET |RIBAVIRIN 200MG TAB [VA PRODUCT]
C0789390|T121|N0000164016|NDFRT|RIBAVIRIN 200MG TABLET|RIBAVIRIN 200MG TAB [VA PRODUCT]
C0789390|T121|N0000164016|NDFRT|RIBAVIRIN, 200 MG ORAL TABLET|RIBAVIRIN 200MG TAB [VA PRODUCT]
C3473212|T121|N0000190073|NDFRT|RIBAVIRIN 200MG ORAL TABLET, RIBAVIRIN 400MG ORAL TABLET|RIBAVIRIN 200MG X 7/400MG X 7 TAB DOSEPACK,14 [VA PRODUCT]
C3473212|T121|N0000190073|NDFRT|RIBASPHERE RIBAPAK KIT|RIBAVIRIN 200MG X 7/400MG X 7 TAB DOSEPACK,14 [VA PRODUCT]
C3473212|T121|N0000190073|NDFRT|RIBAVIRIN TAB 200 MG & RIBAVIRIN TAB 400 MG DOSE PACK|RIBAVIRIN 200MG X 7/400MG X 7 TAB DOSEPACK,14 [VA PRODUCT]
C3473212|T121|N0000190073|NDFRT|{7 (RIBAVIRIN 200 MG ORAL TABLET) / 7 (RIBAVIRIN 400 MG ORAL TABLET) } PACK|RIBAVIRIN 200MG X 7/400MG X 7 TAB DOSEPACK,14 [VA PRODUCT]
C3473212|T121|N0000190073|NDFRT|RIBAPAK 600, 200 MG-400 MG ORAL TABLET|RIBAVIRIN 200MG X 7/400MG X 7 TAB DOSEPACK,14 [VA PRODUCT]
C3473212|T121|N0000190073|NDFRT|RIBAVIRIN 200MGX7/400MGX7 TAB DOSEPK 14|RIBAVIRIN 200MG X 7/400MG X 7 TAB DOSEPACK,14 [VA PRODUCT]
C3473212|T121|N0000190073|NDFRT|RIBAVIRIN 200MG X 7/400MG X 7 TAB DOSEPACK,14 [VA PRODUCT]|RIBAVIRIN 200MG X 7/400MG X 7 TAB DOSEPACK,14 [VA PRODUCT]
C3473212|T121|N0000190073|NDFRT|RIBAVIRIN 200MG X 7/400MG X 7 TAB DOSEPACK,14|RIBAVIRIN 200MG X 7/400MG X 7 TAB DOSEPACK,14 [VA PRODUCT]
C3473212|T121|N0000190073|NDFRT|RIBAVIRIN 200 MG (7) ORAL TABLET / RIBAVIRIN 400 MG (7) ORAL TABLET PACK|RIBAVIRIN 200MG X 7/400MG X 7 TAB DOSEPACK,14 [VA PRODUCT]
C3473212|T121|N0000190073|NDFRT|RIBAVIRIN;RIBAVIRIN 200 MG; 400 MG ORAL TABLET [RIBASPHERE RIBAPAK]|RIBAVIRIN 200MG X 7/400MG X 7 TAB DOSEPACK,14 [VA PRODUCT]
C3473212|T121|N0000190073|NDFRT|RIBASPHERE RIBAPAK 600MG/DAY DOSE PACK TABLET|RIBAVIRIN 200MG X 7/400MG X 7 TAB DOSEPACK,14 [VA PRODUCT]
C3700547|T121||NDFRT|RIBAVIRIN 200 MG ORAL TABLET, FILM COATED [MODERIBA]
C3700547|T121||NDFRT|MODERIBA 200 MG ORAL TABLET
C3700547|T121||NDFRT|RIBAVIRIN 200 MG ORAL TABLET [MODERIBA]
C3700547|T121||NDFRT|MODERIBA, 200 MG ORAL TABLET
C3700547|T121||NDFRT|MODERIBA 200MG TABLET
C1169961|T121||NDFRT|COPEGUS 200 MG ORAL TABLET
C1169961|T121||NDFRT|RIBAVIRIN 200 MG ORAL TABLET [COPEGUS]
C1169961|T121||NDFRT|COPEGUS 200MG TABLET
C1169961|T121||NDFRT|RIBAVIRIN 200 MG ORAL TABLET, FILM COATED [COPEGUS]
C1169961|T121||NDFRT|COPEGUS, 200 MG ORAL TABLET
C1694693|T121||NDFRT|RIBASPHERE, 200 MG ORAL TABLET
C1694693|T121||NDFRT|RIBASPHERE 200 MG ORAL TABLET
C1694693|T121||NDFRT|RIBAVIRIN 200 MG ORAL TABLET [RIBASPHERE]
C1694693|T121||NDFRT|RIBAVIRIN 200 MG ORAL TABLET, FILM COATED [RIBASPHERE]
C1694693|T121||NDFRT|RIBASPHERE 200MG TABLET
C0789393|T121|N0000165356|NDFRT|RIBAVIRIN 40 MG/ML ORAL SOLUTION|RIBAVIRIN 200MG/5ML SOLN,ORAL [VA PRODUCT]
C0789393|T121|N0000165356|NDFRT|RIBAVIRIN SOLN 40 MG/ML|RIBAVIRIN 200MG/5ML SOLN,ORAL [VA PRODUCT]
C0789393|T121|N0000165356|NDFRT|RIBAVIRIN 200MG/5ML SOLN,ORAL|RIBAVIRIN 200MG/5ML SOLN,ORAL [VA PRODUCT]
C0789393|T121|N0000165356|NDFRT|RIBAVIRIN 200MG/5ML ORAL SOLN|RIBAVIRIN 200MG/5ML SOLN,ORAL [VA PRODUCT]
C0789393|T121|N0000165356|NDFRT|RIBAVIRIN 200MG/5ML SOLN,ORAL [VA PRODUCT]|RIBAVIRIN 200MG/5ML SOLN,ORAL [VA PRODUCT]
C0789393|T121|N0000165356|NDFRT|RIBAVIRIN 40MG ORAL SOLUTION|RIBAVIRIN 200MG/5ML SOLN,ORAL [VA PRODUCT]
C0789393|T121|N0000165356|NDFRT|RIBAVIRIN 40MG/ML ORAL SOLUTION |RIBAVIRIN 200MG/5ML SOLN,ORAL [VA PRODUCT]
C0789393|T121|N0000165356|NDFRT|RIBAVIRIN 40MG/ML ORAL SOLUTION|RIBAVIRIN 200MG/5ML SOLN,ORAL [VA PRODUCT]
C1586219|T121||NDFRT|REBETOL 40 MG/ML ORAL SOLUTION
C1586219|T121||NDFRT|RIBAVIRIN 40 MG/ML ORAL SOLUTION [REBETOL]
C1586219|T121||NDFRT|REBETOL 40MG/ML SOLUTION
C1586219|T121||NDFRT|RIBAVIRIN 40 MG IN 1 ML ORAL LIQUID [REBETOL]
C1586219|T121||NDFRT|REBETOL, 40 MG/ML ORAL SOLUTION
C0350923|T121||NDFRT|RIBAVIRIN 20 MG/ML INHALANT SOLUTION [VIRAZID]
C0350923|T121||NDFRT|VIRAZID 20 MG/ML INHALANT SOLUTION
C0979999|T121|N0000156300|NDFRT|RIBAVIRIN 20 MG/ML INHALANT SOLUTION|RIBAVIRIN 6GM/VIL INHL [VA PRODUCT]
C0979999|T121|N0000156300|NDFRT|RIBAVIRIN 6GM/VI INHL SOLN|RIBAVIRIN 6GM/VIL INHL [VA PRODUCT]
C0979999|T121|N0000156300|NDFRT|RIBAVIRIN 6GM/VIL INHL [VA PRODUCT]|RIBAVIRIN 6GM/VIL INHL [VA PRODUCT]
C0979999|T121|N0000156300|NDFRT|RIBAVIRIN 6GM/VIL INHL|RIBAVIRIN 6GM/VIL INHL [VA PRODUCT]
C0979999|T121|N0000156300|NDFRT|RIBAVIRIN 6G POWDER FOR NEBULIZER SOLUTION|RIBAVIRIN 6GM/VIL INHL [VA PRODUCT]
C0979999|T121|N0000156300|NDFRT|RIBAVIRIN 6 GM INHALATION POWDER FOR SOLUTION|RIBAVIRIN 6GM/VIL INHL [VA PRODUCT]
C0979999|T121|N0000156300|NDFRT|RIBAVIRIN 6G/VIAL POWDER |RIBAVIRIN 6GM/VIL INHL [VA PRODUCT]
C0979999|T121|N0000156300|NDFRT|RIBAVIRIN 6G/VIAL POWDER|RIBAVIRIN 6GM/VIL INHL [VA PRODUCT]
C0979999|T121|N0000156300|NDFRT|RIBAVIRIN 6 GM POWDER FOR INHALANT SOLUTION|RIBAVIRIN 6GM/VIL INHL [VA PRODUCT]
C0979999|T121|N0000156300|NDFRT|RIBAVIRIN FOR INHAL SOLN 6 GM|RIBAVIRIN 6GM/VIL INHL [VA PRODUCT]
C0979999|T121|N0000156300|NDFRT|TRIBAVIRIN 6G INHALATION (PDR FOR RECON)|RIBAVIRIN 6GM/VIL INHL [VA PRODUCT]
C0979999|T121|N0000156300|NDFRT|TRIBAVIRIN 6G INHALATION (PDR FOR RECON) |RIBAVIRIN 6GM/VIL INHL [VA PRODUCT]
C0979999|T121|N0000156300|NDFRT|TRIBAVIRIN 6G INHALATION (PDR FOR RECON) |RIBAVIRIN 6GM/VIL INHL [VA PRODUCT]
C0979999|T121|N0000156300|NDFRT|RIBAVIRIN 6 G INHALATION POWDER FOR RECONSTITUTION|RIBAVIRIN 6GM/VIL INHL [VA PRODUCT]
C0708742|T121||NDFRT|RIBAVIRIN 20 MG/ML INHALANT SOLUTION [VIRAZOLE]
C0708742|T121||NDFRT|VIRAZOLE 20 MG/ML INHALANT SOLUTION
C0708742|T121||NDFRT|VIRAZOLE 6G POWDER FOR INHALATION SOLUTION
C0708742|T121||NDFRT|RIBAVIRIN 6 GM INHALATION POWDER FOR SOLUTION [VIRAZOLE]
C0708742|T121||NDFRT|RIBAVIRIN 6 G RESPIRATORY (INHALATION) POWDER, FOR SOLUTION [VIRAZOLE]
C0708742|T121||NDFRT|VIRAZOLE, 6 G INHALATION POWDER FOR RECONSTITUTION
C3701057|T121||NDFRT|RIBAVIRIN 200 MG [MODERIBA]
C1601182|T121||NDFRT|RIBAVIRIN 200 MG [RIBASPHERE]
C1593466|T121||NDFRT|RIBAVIRIN 200 MG [REBETOL]
C1593727|T121||NDFRT|RIBAVIRIN 200 MG [COPEGUS]
C1589271|T121||NDFRT|RIBAVIRIN 40 MG/ML [REBETOL]
C1622085|T121||NDFRT|VIRAZOLE
C1622085|T121||NDFRT|VILONA
C1622085|T121||NDFRT|ICN BRAND OF RIBAVIRIN
C0702025|T121||NDFRT|ICN-1229
C0702025|T121||NDFRT|ICN 1229
C0702025|T121||NDFRT|ICN1229
C0702024|T121||NDFRT|RIBAMIDE
C0702024|T121||NDFRT|RIBAMIDYL
C0702024|T121||NDFRT|RIBAMIDIL
C0035525|T121|N0000005892|NDFRT|RIBAVIRIN|RIBAVIRIN [CHEMICAL/INGREDIENT]
C0035525|T121|N0000005892|NDFRT|1H-1,2,4-TRIAZOLE-3-CARBOXAMIDE, 1-BETA-D-RIBOFURANOSYL-|RIBAVIRIN [CHEMICAL/INGREDIENT]
C0035525|T121|N0000005892|NDFRT|1-BETA-D-RIBOFURANOSYL-1,2,4-TRIAZOLO-3-CARBOXAMIDE|RIBAVIRIN [CHEMICAL/INGREDIENT]
C0035525|T121|N0000005892|NDFRT|1-BETA-D-RIBOFURANOSYL-1H-1,2,4-TRIAZOLE-3-CARBOXAMIDE|RIBAVIRIN [CHEMICAL/INGREDIENT]
C0035525|T121|N0000005892|NDFRT|RTCA|RIBAVIRIN [CHEMICAL/INGREDIENT]
C0035525|T121|N0000005892|NDFRT|RIBA|RIBAVIRIN [CHEMICAL/INGREDIENT]
C0035525|T121|N0000005892|NDFRT|RIBAVIRIN |RIBAVIRIN [CHEMICAL/INGREDIENT]
C0035525|T121|N0000005892|NDFRT|TRIBAVIRIN|RIBAVIRIN [CHEMICAL/INGREDIENT]
C0035525|T121|N0000005892|NDFRT|RIBAVIRIN [CHEMICAL/INGREDIENT]|RIBAVIRIN [CHEMICAL/INGREDIENT]
C0035525|T121|N0000005892|NDFRT|RIBOVIRIN|RIBAVIRIN [CHEMICAL/INGREDIENT]
C0035525|T121|N0000005892|NDFRT|TRIBAVIRIN |RIBAVIRIN [CHEMICAL/INGREDIENT]
C0035525|T121|N0000005892|NDFRT|1-.BETA.-D-RIBOFURANOSYL-1H-1,2, 4-TRIAZOLE-3-CARBOXAMIDE|RIBAVIRIN [CHEMICAL/INGREDIENT]
C0035525|T121|N0000005892|NDFRT|RIBAVIRIN |RIBAVIRIN [CHEMICAL/INGREDIENT]
C0035525|T121|N0000005892|NDFRT|RIBAVIRIN |RIBAVIRIN [CHEMICAL/INGREDIENT]
C2317046|T121||NDFRT|RESPIRATORY FORM RIBAVIRIN
C2317046|T121||NDFRT|RESPIRATORY FORM RIBAVIRIN 
C2315948|T121||NDFRT|ORAL FORM RIBAVIRIN 
C2315948|T121||NDFRT|ORAL FORM RIBAVIRIN
C2148525|T121||NDFRT|RIBAVIRIN 200MG CAPSULES GIVEN WITH INTERFERON ALFA-2B 
C2148525|T121||NDFRT|RIBAVIRIN 200MG CAPSULES GIVEN WITH INTERFERON ALFA-2B
C1626919|T121|N0000177127|NDFRT|RIBAVIRIN 400 MG ORAL TABLET|RIBAVIRIN 400MG TAB [VA PRODUCT]
C1626919|T121|N0000177127|NDFRT|RIBAVIRIN TAB 400 MG|RIBAVIRIN 400MG TAB [VA PRODUCT]
C1626919|T121|N0000177127|NDFRT|RIBAVIRIN 400MG ORAL TABLET|RIBAVIRIN 400MG TAB [VA PRODUCT]
C1626919|T121|N0000177127|NDFRT|RIBAVIRIN 400MG TAB|RIBAVIRIN 400MG TAB [VA PRODUCT]
C1626919|T121|N0000177127|NDFRT|RIBAVIRIN, 400 MG ORAL TABLET|RIBAVIRIN 400MG TAB [VA PRODUCT]
C1626919|T121|N0000177127|NDFRT|RIBAVIRIN 400MG TAB [VA PRODUCT]|RIBAVIRIN 400MG TAB [VA PRODUCT]
C1626919|T121|N0000177127|NDFRT|RIBAVIRIN 400 MG ORAL TABLET, FILM COATED|RIBAVIRIN 400MG TAB [VA PRODUCT]
C1626919|T121|N0000177127|NDFRT|RIBAVIRIN 400MG TABLET |RIBAVIRIN 400MG TAB [VA PRODUCT]
C1626919|T121|N0000177127|NDFRT|RIBAVIRIN 400MG TABLET|RIBAVIRIN 400MG TAB [VA PRODUCT]
C1676705|T121|N0000177128|NDFRT|RIBAVIRIN 600 MG ORAL TABLET|RIBAVIRIN 600MG TAB [VA PRODUCT]
C1676705|T121|N0000177128|NDFRT|RIBAVIRIN TAB 600 MG|RIBAVIRIN 600MG TAB [VA PRODUCT]
C1676705|T121|N0000177128|NDFRT|RIBAVIRIN 600MG TABLET |RIBAVIRIN 600MG TAB [VA PRODUCT]
C1676705|T121|N0000177128|NDFRT|RIBAVIRIN 600MG TABLET|RIBAVIRIN 600MG TAB [VA PRODUCT]
C1676705|T121|N0000177128|NDFRT|RIBAVIRIN, 600 MG ORAL TABLET|RIBAVIRIN 600MG TAB [VA PRODUCT]
C1676705|T121|N0000177128|NDFRT|RIBAVIRIN 600MG ORAL TABLET|RIBAVIRIN 600MG TAB [VA PRODUCT]
C1676705|T121|N0000177128|NDFRT|RIBAVIRIN 600MG TAB|RIBAVIRIN 600MG TAB [VA PRODUCT]
C1676705|T121|N0000177128|NDFRT|RIBAVIRIN 600MG TAB [VA PRODUCT]|RIBAVIRIN 600MG TAB [VA PRODUCT]
C1676705|T121|N0000177128|NDFRT|RIBAVIRIN 600 MG ORAL TABLET, FILM COATED|RIBAVIRIN 600MG TAB [VA PRODUCT]
C1170183|T121||NDFRT|COPEGUS
C1870873|T121||NDFRT|2-(3-AMINO-3-DEOXYXYLOFURANOSYL)THIAZOLE-4-CARBOXAMIDE
C3700973|T121||NDFRT|MODERIBA
C0637676|T121||NDFRT|METHYL 1-RIBOFURANOSYL-1,2,4-TRIAZOLE-3-CARBOXAMIDATE
C0637676|T121||NDFRT|MRTC
C0627880|T121||NDFRT|TB-RIBAVIRIN
C0627880|T121||NDFRT|TRIBUTYLRIBAVIRIN
C0640066|T121||NDFRT|3-RIBOFURANOSYL-1,2,4-TRIAZOLE-5-CARBOXAMIDE
C0076656|T121||NDFRT|2-RIBOFURANOSYLTHIAZOLE-4-CARBOXAMIDE
C0076656|T121||NDFRT|RIBOXAMIDE
C0076656|T121||NDFRT|TIAZOFURIN
C0076656|T121||NDFRT|TRANS CAROTID ARTERY REVASCULARIZATION
C0639452|T121||NDFRT|1-(5'-O-SULFAMOYL-BETA-D-RIBOFURANOSYL)(1,2,4)TRIAZOLE-3-CARBONITRILE
C0639452|T121||NDFRT|SRTCN
C1454123|T121||NDFRT|5'-NOR CARBOCYCLIC RIBAVIRIN
C0073218|T121||NDFRT|RIBAVIRIN 5'-DIPHOSPHATE
C0073218|T121||NDFRT|RIBAVIRIN-DP
C0637674|T121||NDFRT|ETHYL 1-RIBOFURANOSYL-1,2,4-TRIAZOLE-3-CARBOXIMIDATE
C0637674|T121||NDFRT|ERTC
C0764977|T121||NDFRT|4-FLUORO-1-RIBOFURANOSYL-1H-PYRAZOLE-3-CARBOXAMIDE
C0764977|T121||NDFRT|4-FRPC
C0605624|T121||NDFRT|1-(4-THIO-BETA-D-RIBOFURANOSYL)-1,2,4-TRIAZOLE-3-CARBOXAMIDE
C0632093|T121||NDFRT|5'-O-BETA-D-GLUCOPYRANOSYL RIBAVIRIN
C0632093|T121||NDFRT|5'-O-GLUCOPYRANOSYL RIBAVIRIN
C0647853|T121||NDFRT|2-(2',3'-DIDEOXYGLYCEROPENT-2-ENOFURANOSYL)THIAZOLE-4-CARBOXAMIDE
C0647853|T121||NDFRT|2',3'-DIDEHYDRO-2',3'-DIDEOXYTIAZOFURIN
C0640069|T121||NDFRT|2-RIBOFURANOSYL-1,2,3-TRIAZOLE-4,5-DICARBOXAMIDE
C1957632|T121||NDFRT|TIAZOFURIN MONOPHOSPHATE
C0632095|T121||NDFRT|5'-O-BETA-D-GALACTOPYRANOSYL RIBAVIRIN
C0632095|T121||NDFRT|5'-O-GALACTOPYRANOSYL RIBAVIRIN
C0073219|T121||NDFRT|1H-1,2,4-TRIAZOLE-3-CARBOXAMIDE, 1-(5-O-(AMINOSULFONYL)-BETA-D-RIBOFURANOSYL)-
C0073219|T121||NDFRT|5'-O-SULFAMOYL-1-RIBOFURANOSYL-1,2,4-TRIAZOLE-3-CARBOXAMIDE
C0073219|T121||NDFRT|RIBAVIRIN 5'-SULFAMATE
C0073219|T121||NDFRT|1-(5'-O-SULFAMOYL-BETA-RIBOFURANOSYL)-(1,2,4)TRIAZOLE-3-CARBOXAMIDE
C0140479|T121||NDFRT|RIBAVIRIN 2',3',5'-TRIACETATE
C0073221|T121||NDFRT|1-BETA-D-RIBOFURANOSYL-1,2,4-TRIAZOLE-3-CARBOXAMIDINE
C0073221|T121||NDFRT|RIBAMIDINE
C0073221|T121||NDFRT|RIBAVIRIN AMIDINE
C0073221|T121||NDFRT|TRAUMA CERTIFIED RN
C0073221|T121||NDFRT|TARIBAVIRIN
C0073221|T121||NDFRT|VIRAMIDINE
C0639450|T121||NDFRT|1-(5'-O-SULFAMOYL-BETA-RIBOFURANOSYL)(1,2,4)TRIAZOLE-3-THIOCARBOXAMIDE
C0639450|T121||NDFRT|SRTC
C0647851|T121||NDFRT|2-(2',3'-DIDEOXYGLYCEROPENTAFURANOSYL)THIAZOLE-4-CARBOXAMIDE
C0647851|T121||NDFRT|2',3'-DIDEOXYTIAZOFURIN
C0050823|T121||NDFRT|ADENYLYL-(3'-5')-VIRAZOLE
C0050823|T121||NDFRT|ADENYLYL-(3'-5')RIBAVIRIN
C0050823|T121||NDFRT|3'-ADENYLIC ACID, 3'-5'-ESTER WITH 1-BETA-D-RIBOFURANOSYL-1H-1,2,4-TRIAZOLE-3-CARBOXAMIDE
C2240463|T121|N0000190072|NDFRT|{7 (RIBAVIRIN 400 MG ORAL TABLET) / 7 (RIBAVIRIN 600 MG ORAL TABLET) } PACK|RIBAVIRIN 600MG X 7/400MG X 7 TAB DOSEPACK,14 [VA PRODUCT]
C2240463|T121|N0000190072|NDFRT|RIBAVIRIN 400MG ORAL TABLET, RIBAVIRIN 600MG ORAL TABLET|RIBAVIRIN 600MG X 7/400MG X 7 TAB DOSEPACK,14 [VA PRODUCT]
C2240463|T121|N0000190072|NDFRT|RIBAVIRIN 600MG X 7/400MG X 7 TAB DOSEPACK,14 [VA PRODUCT]|RIBAVIRIN 600MG X 7/400MG X 7 TAB DOSEPACK,14 [VA PRODUCT]
C2240463|T121|N0000190072|NDFRT|RIBAVIRIN 600MG X 7/400MG X 7 TAB DOSEPACK,14|RIBAVIRIN 600MG X 7/400MG X 7 TAB DOSEPACK,14 [VA PRODUCT]
C2240463|T121|N0000190072|NDFRT|RIBAVIRIN 600MGX7/400MGX7 TAB DOSEPK 14|RIBAVIRIN 600MG X 7/400MG X 7 TAB DOSEPACK,14 [VA PRODUCT]
C4075513|T121||NDFRT|RIBAVIRIN INJECTABLE PRODUCT
C4075513|T121||NDFRT|PARENTERAL FORM RIBAVIRIN 
C4075513|T121||NDFRT|PARENTERAL FORM RIBAVIRIN
C0361571|T121||NDFRT|RIBAVIRIN 100 MG ORAL CAPSULE
C0361571|T121||NDFRT|RIBAVIRIN 100MG CAPSULE
C0361571|T121||NDFRT|RIBAVIRIN 100MG CAPSULE 
C0361571|T121||NDFRT|RIBAVIRIN 100MG CAPSULE 
C0979998|T121|N0000165984|NDFRT|RIBAVIRIN 200 MG ORAL CAPSULE|RIBAVIRIN 200MG CAP [VA PRODUCT]
C0979998|T121|N0000165984|NDFRT|RIBAVIRIN 200MG ORAL CAPSULE|RIBAVIRIN 200MG CAP [VA PRODUCT]
C0979998|T121|N0000165984|NDFRT|RIBAVIRIN 200MG CAP|RIBAVIRIN 200MG CAP [VA PRODUCT]
C0979998|T121|N0000165984|NDFRT|RIBAVIRIN CAP 200 MG|RIBAVIRIN 200MG CAP [VA PRODUCT]
C0979998|T121|N0000165984|NDFRT|RIBAVIRIN 200MG CAP [VA PRODUCT]|RIBAVIRIN 200MG CAP [VA PRODUCT]
C0979998|T121|N0000165984|NDFRT|RIBAVIRIN 200 MG ORAL CAPSULE [RIBAVIRIN]|RIBAVIRIN 200MG CAP [VA PRODUCT]
C0979998|T121|N0000165984|NDFRT|RIBAVIRIN 200MG CAPSULE|RIBAVIRIN 200MG CAP [VA PRODUCT]
C0979998|T121|N0000165984|NDFRT|RIBAVIRIN 200MG CAPSULE |RIBAVIRIN 200MG CAP [VA PRODUCT]
C0979998|T121|N0000165984|NDFRT|RIBAVIRIN 200MG CAPSULE |RIBAVIRIN 200MG CAP [VA PRODUCT]
C0979998|T121|N0000165984|NDFRT|RIBAVIRIN, 200 MG ORAL CAPSULE|RIBAVIRIN 200MG CAP [VA PRODUCT]
C0717864|T121||NDFRT|INTERFERON ALFA-2B/RIBAVIRIN
C0717864|T121||NDFRT|INTERFERON ALFA-2B-RIBAVIRIN
C0717864|T121||NDFRT|RIBAVIRIN+INTERFERON ALPHA-2B 
C0717864|T121||NDFRT|RIBAVIRIN+INTERFERON ALPHA-2B
C0702029|T121||NDFRT|VIRAMIDE
C0731013|T121||NDFRT|VIRAZID
C1170576|T121||NDFRT|REBETOL
C1170576|T121||NDFRT|RIBAVIRIN MERCK BRAND
C1170576|T121||NDFRT|MERCK BRAND OF RIBAVIRIN
C1170576|T121||NDFRT|PFIZER BRAND OF RIBAVIRIN
C1170576|T121||NDFRT|ESSEX BRAND OF RIBAVIRIN
C1564036|T121||NDFRT|GROSSMAN BRAND OF RIBAVIRIN
C1564036|T121||NDFRT|VIRAZIDE
C1564036|T121||NDFRT|DERMATECH BRAND OF RIBAVIRIN
C1564336|T121||NDFRT|RIBASPHERE
C1564336|T121||NDFRT|THREE RIVERS PHARMACEUTICALS BRAND OF RIBAVIRIN
C0722990|T121||NDFRT|REBETRON
C1878903|T121||NDFRT|RIBATAB
C0935908|T121||NDFRT|PALIVIZUMAB/RIBAVIRIN
C0935908|T121||NDFRT|PALI/RIBA
C1339084|T121||NDFRT|RIBAVIRIN 400 MG ORAL CAPSULE
C2341626|T121||NDFRT|RIBAVIRIN 500MG ORAL TABLET
C2341626|T121||NDFRT|RIBAVIRIN 500 MG ORAL TABLET
C2341626|T121||NDFRT|RIBAVIRIN 500 MG ORAL TABLET, FILM COATED
C2341626|T121||NDFRT|RIBAVIRIN, 500 MG ORAL TABLET
C3222959|T121||NDFRT|COPEGUS PILL
C3232238|T121||NDFRT|REBETOL PILL
C3237959|T121||NDFRT|RIBATAB PILL
C3237961|T121||NDFRT|RIBASPHERE PILL
C1247842|T121||NDFRT|RIBAVIRIN ORAL CAPSULE
C1247844|T121||NDFRT|RIBAVIRIN ORAL TABLET
C3701173|T121||NDFRT|MODERIBA PILL
C1169620|T121||NDFRT|REBETOL 200 MG ORAL CAPSULE
C1169620|T121||NDFRT|RIBAVIRIN 200 MG ORAL CAPSULE [REBETOL]
C1169620|T121||NDFRT|REBETOL 200MG CAPSULE
C1169620|T121||NDFRT|REBETOL, 200 MG ORAL CAPSULE
C1584733|T121||NDFRT|RIBASPHERE 200 MG ORAL CAPSULE
C1584733|T121||NDFRT|RIBAVIRIN 200 MG ORAL CAPSULE [RIBASPHERE]
C1584733|T121||NDFRT|RIBASPHERE 200MG CAPSULE
C1584733|T121||NDFRT|RIBASPHERE, 200 MG ORAL CAPSULE
C2342580|T121||NDFRT|{6 (0.5 ML) (INTERFERON ALFA-2B 6000000 UNT/ML INJECTABLE SOLUTION) / 70 (RIBAVIRIN 200 MG ORAL CAPSULE) } PACK
C2342658|T121||NDFRT|{1 (3 ML) (INTERFERON ALFA-2B 6000000 UNT/ML INJECTABLE SOLUTION) / 70 (RIBAVIRIN 200 MG ORAL CAPSULE) } PACK
C2342661|T121||NDFRT|{1 (1.2 ML) (INTERFERON ALFA-2B 15000000 UNT/ML INJECTABLE SOLUTION) / 70 (RIBAVIRIN 200 MG ORAL CAPSULE) } PACK
C2342663|T121||NDFRT|{1 (3 ML) (INTERFERON ALFA-2B 6000000 UNT/ML INJECTABLE SOLUTION) / 84 (RIBAVIRIN 200 MG ORAL CAPSULE) } PACK
C2342664|T121||NDFRT|{6 (0.5 ML) (INTERFERON ALFA-2B 6000000 UNT/ML INJECTABLE SOLUTION) / 84 (RIBAVIRIN 200 MG ORAL CAPSULE) } PACK
C2342665|T121||NDFRT|{1 (1.2 ML) (INTERFERON ALFA-2B 15000000 UNT/ML INJECTABLE SOLUTION) / 84 (RIBAVIRIN 200 MG ORAL CAPSULE) } PACK
C2342667|T121||NDFRT|{1 (3 ML) (INTERFERON ALFA-2B 6000000 UNT/ML INJECTABLE SOLUTION) / 42 (RIBAVIRIN 200 MG ORAL CAPSULE) } PACK
C2342668|T121||NDFRT|{6 (0.5 ML) (INTERFERON ALFA-2B 6000000 UNT/ML INJECTABLE SOLUTION) / 42 (RIBAVIRIN 200 MG ORAL CAPSULE) } PACK
C2342669|T121||NDFRT|{1 (1.2 ML) (INTERFERON ALFA-2B 15000000 UNT/ML INJECTABLE SOLUTION) / 42 (RIBAVIRIN 200 MG ORAL CAPSULE) } PACK
C0413496|T121||NDFRT|ADVERSE REACTION TO TRIBAVIRIN
C0413496|T121||NDFRT|ADVERSE REACTION TO TRIBAVIRIN 
C0413496|T121||NDFRT|TRIBAVIRIN ADVERSE REACTION
C0413496|T121||NDFRT|TRIBAVIRIN ADVERSE REACTION 
C0413496|T121||NDFRT|RIBAVIRIN ADVERSE REACTION
C1595591|T121||NDFRT|RIBAVIRIN 20 MG/ML [VIRAZID]
C1616510|T121||NDFRT|RIBAVIRIN 20 MG/ML [VIRAZOLE]
C1240752|T121||NDFRT|RIBAVIRIN ORAL CAPSULE [REBETOL]
C1601183|T121||NDFRT|RIBAVIRIN ORAL CAPSULE [RIBASPHERE]
C0789392|T121||NDFRT|RIBAVIRIN 20 MG/ML ORAL SOLUTION
C1589272|T121||NDFRT|RIBAVIRIN ORAL SOLUTION [REBETOL]
C3701110|T121||NDFRT|RIBAVIRIN ORAL TABLET [MODERIBA]
C1242547|T121||NDFRT|RIBAVIRIN ORAL TABLET [COPEGUS]
C1704170|T121||NDFRT|RIBAVIRIN ORAL TABLET [RIBASPHERE]
C1694682|T121||NDFRT|RIBAVIRIN ORAL TABLET [RIBATAB]
C1621221|T121||NDFRT|RIBAVIRIN INHALANT SOLUTION [VIRAZOLE]
C1235816|T121||NDFRT|RIBAVIRIN INHALANT SOLUTION [VIRAZID]
C3701058|T121||NDFRT|RIBAVIRIN 400 MG [MODERIBA]
C1702720|T121||NDFRT|RIBAVIRIN 400 MG [RIBASPHERE]
C1878904|T121||NDFRT|RIBAVIRIN 400 MG [RIBATAB]
C3668937|T121||NDFRT|MODERIBA 400 MG ORAL TABLET
C3668937|T121||NDFRT|RIBAVIRIN 400 MG ORAL TABLET [MODERIBA]
C3668937|T121||NDFRT|RIBAVIRIN 400 MG ORAL TABLET, FILM COATED [MODERIBA]
C1694134|T121||NDFRT|RIBASPHERE, 400 MG ORAL TABLET
C1694134|T121||NDFRT|RIBASPHERE 400 MG ORAL TABLET
C1694134|T121||NDFRT|RIBAVIRIN 400 MG ORAL TABLET [RIBASPHERE]
C1694134|T121||NDFRT|RIBAVIRIN 400 MG ORAL TABLET, FILM COATED [RIBASPHERE]
C1694134|T121||NDFRT|RIBASPHERE 400MG TABLET
C1878399|T121||NDFRT|RIBATAB 400MG TABLET
C1878399|T121||NDFRT|RIBAVIRIN 400 MG ORAL TABLET [RIBATAB]
C1878399|T121||NDFRT|RIBATAB 400 MG ORAL TABLET
C1878399|T121||NDFRT|RIBATAB, 400 MG ORAL TABLET
C2240739|T121|N0000190071|NDFRT|{14 (RIBAVIRIN 400 MG ORAL TABLET) } PACK|RIBAVIRIN 400MG TAB DOSEPACK,14 [VA PRODUCT]
C2240739|T121|N0000190071|NDFRT|RIBAVIRIN 400MG TAB DOSEPACK 14|RIBAVIRIN 400MG TAB DOSEPACK,14 [VA PRODUCT]
C2240739|T121|N0000190071|NDFRT|RIBAVIRIN 400MG TAB DOSEPACK,14 [VA PRODUCT]|RIBAVIRIN 400MG TAB DOSEPACK,14 [VA PRODUCT]
C2240739|T121|N0000190071|NDFRT|RIBAVIRIN 400MG TAB DOSEPACK,14|RIBAVIRIN 400MG TAB DOSEPACK,14 [VA PRODUCT]
C1641488|T121||NDFRT|RIBAVIRIN:MCNC:PT:SER/PLAS:QN
C1641488|T121||NDFRT|RIBAVIRIN [MASS/VOLUME] IN SERUM OR PLASMA
C1641488|T121||NDFRT|RIBAVIRIN SERPL-MCNC
C1641488|T121||NDFRT|RIBAVIRIN:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE
C3668939|T121||NDFRT|RIBAVIRIN 600 MG ORAL TABLET [MODERIBA]
C3668939|T121||NDFRT|MODERIBA 600 MG ORAL TABLET
C3668939|T121||NDFRT|RIBAVIRIN 600 MG ORAL TABLET, FILM COATED [MODERIBA]
C1694694|T121||NDFRT|RIBASPHERE, 600 MG ORAL TABLET
C1694694|T121||NDFRT|RIBASPHERE 600 MG ORAL TABLET
C1694694|T121||NDFRT|RIBAVIRIN 600 MG ORAL TABLET [RIBASPHERE]
C1694694|T121||NDFRT|RIBAVIRIN 600 MG ORAL TABLET, FILM COATED [RIBASPHERE]
C1694694|T121||NDFRT|RIBASPHERE 600MG TABLET
C1878400|T121||NDFRT|RIBAVIRIN 600 MG ORAL TABLET [RIBATAB]
C1878400|T121||NDFRT|RIBATAB 600MG TABLET
C1878400|T121||NDFRT|RIBATAB 600 MG ORAL TABLET
C2240738|T121|N0000190070|NDFRT|{14 (RIBAVIRIN 600 MG ORAL TABLET) } PACK|RIBAVIRIN 600MG X 14 TAB DOSEPACK,14 [VA PRODUCT]
C2240738|T121|N0000190070|NDFRT|RIBAVIRIN 600 MG ORAL TABLET 7 DAY PACK|RIBAVIRIN 600MG X 14 TAB DOSEPACK,14 [VA PRODUCT]
C2240738|T121|N0000190070|NDFRT|RIBAVIRIN 600MG X 14 TAB DOSEPACK 14|RIBAVIRIN 600MG X 14 TAB DOSEPACK,14 [VA PRODUCT]
C2240738|T121|N0000190070|NDFRT|RIBAVIRIN 600MG X 14 TAB DOSEPACK,14 [VA PRODUCT]|RIBAVIRIN 600MG X 14 TAB DOSEPACK,14 [VA PRODUCT]
C2240738|T121|N0000190070|NDFRT|RIBAVIRIN 600MG X 14 TAB DOSEPACK,14|RIBAVIRIN 600MG X 14 TAB DOSEPACK,14 [VA PRODUCT]
C2240738|T121|N0000190070|NDFRT|RIBAVIRIN 600 MG ORAL TABLET 14 COUNT 7 DAY PACK|RIBAVIRIN 600MG X 14 TAB DOSEPACK,14 [VA PRODUCT]
C3701056|T121||NDFRT|RIBAVIRIN 600 MG [MODERIBA]
C1703270|T121||NDFRT|RIBAVIRIN 600 MG [RIBASPHERE]
C1878905|T121||NDFRT|RIBAVIRIN 600 MG [RIBATAB]
C0002199|T121|N0000006710|NDFRT|ALPHA INTERFERON|INTERFERON-ALPHA [CHEMICAL/INGREDIENT]
C0002199|T121|N0000006710|NDFRT|INTERFERON ALPHA|INTERFERON-ALPHA [CHEMICAL/INGREDIENT]
C0002199|T121|N0000006710|NDFRT|INTERFERON-ALPHA|INTERFERON-ALPHA [CHEMICAL/INGREDIENT]
C0002199|T121|N0000006710|NDFRT|INTERFERON ALFA|INTERFERON-ALPHA [CHEMICAL/INGREDIENT]
C0002199|T121|N0000006710|NDFRT|ALPHA-INTERFERON|INTERFERON-ALPHA [CHEMICAL/INGREDIENT]
C0002199|T121|N0000006710|NDFRT|INTERFERON, ALPHA|INTERFERON-ALPHA [CHEMICAL/INGREDIENT]
C0002199|T121|N0000006710|NDFRT|INTERFERON-ALPHA [CHEMICAL/INGREDIENT]|INTERFERON-ALPHA [CHEMICAL/INGREDIENT]
C0002199|T121|N0000006710|NDFRT|INTERFERON.ALPHA|INTERFERON-ALPHA [CHEMICAL/INGREDIENT]
C0002199|T121|N0000006710|NDFRT|IFNA|INTERFERON-ALPHA [CHEMICAL/INGREDIENT]
C0002199|T121|N0000006710|NDFRT|INTERFERON ALFA |INTERFERON-ALPHA [CHEMICAL/INGREDIENT]
C0002199|T121|N0000006710|NDFRT|INTERFERON ALFA |INTERFERON-ALPHA [CHEMICAL/INGREDIENT]
C0002199|T121|N0000006710|NDFRT|ALPHA INTERFERON |INTERFERON-ALPHA [CHEMICAL/INGREDIENT]
C0002199|T121|N0000006710|NDFRT|INTERFERON A|INTERFERON-ALPHA [CHEMICAL/INGREDIENT]
C0002199|T121|N0000006710|NDFRT|IFN-A|INTERFERON-ALPHA [CHEMICAL/INGREDIENT]
C0015980|T121|N0000007668|NDFRT|UNUSUAL BUT OCCASIONALLY USED|INTERFERON-BETA [CHEMICAL/INGREDIENT]
C0015980|T121|N0000007668|NDFRT|INTERFERON BETA|INTERFERON-BETA [CHEMICAL/INGREDIENT]
C0015980|T121|N0000007668|NDFRT|INTERFERON-BETA|INTERFERON-BETA [CHEMICAL/INGREDIENT]
C0015980|T121|N0000007668|NDFRT|INTERFERON BETA |INTERFERON-BETA [CHEMICAL/INGREDIENT]
C0015980|T121|N0000007668|NDFRT|INTERFERON, BETA|INTERFERON-BETA [CHEMICAL/INGREDIENT]
C0015980|T121|N0000007668|NDFRT|INTERFERON-BETA [CHEMICAL/INGREDIENT]|INTERFERON-BETA [CHEMICAL/INGREDIENT]
C0015980|T121|N0000007668|NDFRT|BETA-INTERFERON|INTERFERON-BETA [CHEMICAL/INGREDIENT]
C0015980|T121|N0000007668|NDFRT|INTERFERON.BETA|INTERFERON-BETA [CHEMICAL/INGREDIENT]
C0015980|T121|N0000007668|NDFRT|IFNB|INTERFERON-BETA [CHEMICAL/INGREDIENT]
C0015980|T121|N0000007668|NDFRT|INTERFERON BETA |INTERFERON-BETA [CHEMICAL/INGREDIENT]
C0015980|T121|N0000007668|NDFRT|BETA INTERFERON |INTERFERON-BETA [CHEMICAL/INGREDIENT]
C0015980|T121|N0000007668|NDFRT|IFN-B|INTERFERON-BETA [CHEMICAL/INGREDIENT]
C0015980|T121|N0000007668|NDFRT|ENDOGENOUS INTERFERON BETA|INTERFERON-BETA [CHEMICAL/INGREDIENT]
C0015980|T121|N0000007668|NDFRT|IFN-BETA|INTERFERON-BETA [CHEMICAL/INGREDIENT]
C0015980|T121|N0000007668|NDFRT|INTERFERON BETA, NATURAL|INTERFERON-BETA [CHEMICAL/INGREDIENT]
C0015980|T121|N0000007668|NDFRT|NATURAL HUMAN INTERFERON BETA|INTERFERON-BETA [CHEMICAL/INGREDIENT]
C0021747|T121|N0000008154|NDFRT|INTERFERON|INTERFERONS [CHEMICAL/INGREDIENT]
C0021747|T121|N0000008154|NDFRT|IFN|INTERFERONS [CHEMICAL/INGREDIENT]
C0021747|T121|N0000008154|NDFRT|INTERFERON |INTERFERONS [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|IFN-ALPHA CON 1|INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|CONSENSUS IFN-ALPHA|INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|RIFN-CON-1|INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|RECOMBINANT CONSENSUS INTERFERON ALPHA|INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|INTERFERON-ALPHA CON(1)|INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|INTERFERON ALFACON-1|INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|METHIONYL-INTERFERON-CONSENSUS|INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|METHIONYL INTERFERON CONSENSUS|INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|INTERFERON CONSENSUS, METHIONYL|INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|RECOMBINANT METHIONYL HUMAN CONSENSUS INTERFERON|INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|IFN ALFACON-1|INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|RECOMBINANT CONSENSUS INTERFERON|INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|R-METHUIFN-CON1|INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|CIFN|INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|INTERFERON ALFACON-1 AGENT|INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|CIFN (INTERFERON)|INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|INTERFERON ALFACON-1 |INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]|INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|INTERFERON ALFACON-1 AGENT |INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|INTERFERON ALFACON-1 PREPARATION|INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|CONSENSUS INTERFERON|INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0164613|T121|N0000004938|NDFRT|INTERFERON ALFACON-1 PREPARATION |INTERFERON ALFACON-1 [CHEMICAL/INGREDIENT]
C0021734|T121|N0000006291|NDFRT|INTERFERON ALFA-2A|INTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0021734|T121|N0000006291|NDFRT|RECOMBINANT INTERFERON ALPHA-2A|INTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0021734|T121|N0000006291|NDFRT|RECOMBINANT INTERFERON ALFA-2A|INTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0021734|T121|N0000006291|NDFRT|ALPHA 2 INTERFERON|INTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0021734|T121|N0000006291|NDFRT|IFN ALPHA-2A|INTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0021734|T121|N0000006291|NDFRT|RHUIFN-A 2A|INTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0021734|T121|N0000006291|NDFRT|IFN-ALPHA 2|INTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0021734|T121|N0000006291|NDFRT|INTERFERON ALFA 2A|INTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0021734|T121|N0000006291|NDFRT|INTERFERON ALFA|INTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0021734|T121|N0000006291|NDFRT|INTERFERON ALPHA-2A PREPARATION|INTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0021734|T121|N0000006291|NDFRT|INTERFERON ALFA-2A,RECOMBINANT|INTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0021734|T121|N0000006291|NDFRT|INTERFERON ALFA-2A [CHEMICAL/INGREDIENT]|INTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0021734|T121|N0000006291|NDFRT|INTERFERON ALFA-2A |INTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0021734|T121|N0000006291|NDFRT|INTERFERON ALPHA-2A |INTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0021734|T121|N0000006291|NDFRT|INTERFERON ALPHA-2A PREPARATION |INTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0021734|T121|N0000006291|NDFRT|INTERFERON ALPHA-2A|INTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0021734|T121|N0000006291|NDFRT|INTERFERON ALPHA-2A PREPARATION |INTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0021735|T121|N0000006294|NDFRT|INTERFERON ALFA-2B|INTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0021735|T121|N0000006294|NDFRT|IFN ALPHA-2B|INTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0021735|T121|N0000006294|NDFRT|RECOMBINANT INTERFERON ALFA-2B|INTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0021735|T121|N0000006294|NDFRT|INTERFERON ALPHA-2B|INTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0021735|T121|N0000006294|NDFRT|INTERFERON ALPHA-2B PREPARATION|INTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0021735|T121|N0000006294|NDFRT|INTERFERON ALFA 2-B|INTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0021735|T121|N0000006294|NDFRT|INTERFERON ALFA-2B,RECOMBINANT|INTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0021735|T121|N0000006294|NDFRT|RECOMBINANT INTERFERON ALPHA-2B|INTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0021735|T121|N0000006294|NDFRT|INTERFERON ALFA-2B [CHEMICAL/INGREDIENT]|INTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0021735|T121|N0000006294|NDFRT|INTERFERON ALPHA-2B, RECOMBINANT|INTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0021735|T121|N0000006294|NDFRT|IFNALPHA-2B, RECOMBINANT|INTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0021735|T121|N0000006294|NDFRT|INTERFERON ALFA-2B |INTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0021735|T121|N0000006294|NDFRT|INTERFERON ALPHA-2B |INTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0021735|T121|N0000006294|NDFRT|INTERFERON ALPHA-2B PREPARATION |INTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0021735|T121|N0000006294|NDFRT|INTERFERON ALPHA-2B PREPARATION |INTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0021735|T121|N0000006294|NDFRT|INTERFERON ALFA 2B|INTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0982233|T121|N0000147664|NDFRT|INTERFERON ALFA-3N,HUMAN LEUKOCYTE DERIVED|INTERFERON ALFA-3N,HUMAN LEUKOCYTE DERIVED
C0982234|T121||NDFRT|INTERFERON BETA-1A
C0982234|T121||NDFRT|INTERFERON BETA-1A 
C0982234|T121||NDFRT|INTERFERON BETA-1A,RECOMBINANT
C0982234|T121||NDFRT|RECOMBINANT INTERFERON BETA-1A
C0796545|T121|N0000178331|NDFRT|THIS IS THE ONLY IFNA VERSION I FEEL CONFIDENT SHOULD BE INCLUDED|PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|PEG INTERFERON ALFA-2B|PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|PEGYLATED INTERFERON ALFA-2B|PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|PEG-IFN-A 2B|PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|PEG-IFNA2B|PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|PEG-INTERFERON ALFA-2B|PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|PEG-IFNALPHA-2B|PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|PEG-IFN ALFA-2B|PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|PEGYLATED INTERFERON ALPHA-2B|PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|PEG INF ALPHA-2B|PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|PEG-INTERFERON ALPHA-2B|PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|PEGINTERFERON ALPHA-2B|PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|POLYETHYLENE GLYCOL-INTERFERON ALFA-2B|PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]|PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|POLYETHYLENE GLYCOL-INTERFERON ALPHA-2B|PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|PEG INF ALFA-2B|PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|PEG-IFN ALPHA-2B|PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|PEGINTERFERON ALFA-2B |PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|PEG-INTRON|PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|PEGINTERFERON ALFA-2B |PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|PEGINTERFERON ALFA-2B |PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|POLYETHYLENE GLYCOL INTERFERON ALFA-2B|PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0796545|T121|N0000178331|NDFRT|POLYETHYLENE GLYCOL IFN-A2B|PEGINTERFERON ALFA-2B [CHEMICAL/INGREDIENT]
C0391001|T121|N0000178330|NDFRT|PEG-IFN ALFA-2A|PEGINTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0391001|T121|N0000178330|NDFRT|PEG-IFN ALPHA-2A|PEGINTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0391001|T121|N0000178330|NDFRT|PEG-INTERFERON ALFA-2A|PEGINTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0391001|T121|N0000178330|NDFRT|PEGINTERFERON ALFA-2A|PEGINTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0391001|T121|N0000178330|NDFRT|PEGINTERFERON ALPHA-2A |PEGINTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0391001|T121|N0000178330|NDFRT|PEGINTERFERON ALPHA-2A|PEGINTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0391001|T121|N0000178330|NDFRT|PEGYLATED INTERFERON ALFA-2A|PEGINTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0391001|T121|N0000178330|NDFRT|POLYETHYLENE GLYCOL-INTERFERON ALFA-2A|PEGINTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0391001|T121|N0000178330|NDFRT|PEG-INTERFERON ALPHA-2A|PEGINTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0391001|T121|N0000178330|NDFRT|PEGYLATED INTERFERON ALPHA-2A|PEGINTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0391001|T121|N0000178330|NDFRT|POLYETHYLENE GLYCOL-INTERFERON ALPHA-2A|PEGINTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0391001|T121|N0000178330|NDFRT|PEGINTERFERON ALFA-2A [CHEMICAL/INGREDIENT]|PEGINTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0391001|T121|N0000178330|NDFRT|PEGINTERFERON ALFA-2A |PEGINTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0391001|T121|N0000178330|NDFRT|PEGINTERFERON ALFA-2A |PEGINTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C0391001|T121|N0000178330|NDFRT|PEG-IFNA2A|PEGINTERFERON ALFA-2A [CHEMICAL/INGREDIENT]
C3161968|T121||NDFRT|ANTIVIRAL ALPHA INTERFERONS
C3161968|T121||NDFRT|ANTIVIRAL ALPHA INTERFERONS 
C0301340|T121||NDFRT|INJECTABLE INTERFERON 
C0301340|T121||NDFRT|INJECTABLE INTERFERON
C0301340|T121||NDFRT|INJECTABLE INTERFERON 
C2969476|T121||NDFRT|INTERFERON DRUG &#X7C; PATIENT
C0733470|T121||NDFRT|HUMAN LEUKOCYTE INTERFERON
C0733470|T121||NDFRT|INTERFERON
C0733470|T121||NDFRT|IFN
C0063697|T121||NDFRT|ITF-ECP
C1522537|T121||NDFRT|RECOMBINANT INTERFERON
C1522537|T121||NDFRT|IFN
C1522537|T121||NDFRT|HUMAN LEUKOCYTE INTERFERON
C1621234|T121|N0000021274|NDFRT|INTERFERON ALFA-N3|INTERFERON ALFA-3N
C1621234|T121|N0000021274|NDFRT|INTERFERON ALFA-3N|INTERFERON ALFA-3N
C1621234|T121|N0000021274|NDFRT|INTERFERON ALPHA-N3 AGENT|INTERFERON ALFA-3N
C1621234|T121|N0000021274|NDFRT|INTERFERON ALFA-N3 AGENT|INTERFERON ALFA-3N
C1621234|T121|N0000021274|NDFRT|INTERFERON ALFA-N3 |INTERFERON ALFA-3N
C1621234|T121|N0000021274|NDFRT|INTERFERON ALPHA-N3 AGENT |INTERFERON ALFA-3N
C1621234|T121|N0000021274|NDFRT|INTERFERON ALPHA-N3 PREPARATION|INTERFERON ALFA-3N
C1621234|T121|N0000021274|NDFRT|INTERFERON ALPHA-N3 PREPARATION |INTERFERON ALFA-3N
C1621234|T121|N0000021274|NDFRT|ALFA-N3 INTERFERON|INTERFERON ALFA-3N
C0876233|T121||NDFRT|INTERFERON ALFA-N1 LYMPHOBLASTOID
C0876233|T121||NDFRT|INTERFERON ALFA-N1, LYMPHOBLASTOID
C0876233|T121||NDFRT|INTERFERON ALFA-N1 LYMPHOBLASTOID 
C1610033|T121||NDFRT|HUMAN LEUKOCYTE INTERFERON
C1610033|T121||NDFRT|ALPHA INTERFERON
C1610033|T121||NDFRT|LEUKOCYTE INTERFERON
C1610033|T121||NDFRT|IFN ALPHA
C1610033|T121||NDFRT|INTERFERON ALFA-N3
C1610033|T121||NDFRT|INTERFERON ALPHA
C1610033|T121||NDFRT|ALFA-N3 INTERFERON
C1610033|T121||NDFRT|LYMPHOBLAST INTERFERON
C1610033|T121||NDFRT|LYMPHOBLASTOID INTERFERON
C1610033|T121||NDFRT|INTERFERON ALPHA, HUMAN
C0949830|T121||NDFRT|ASTRAGALUS GUMMIFER
C0949830|T121||NDFRT|ASTRAGALUS GUMMIFERS
C0949830|T121||NDFRT|GUMMIFER, ASTRAGALUS
C0949830|T121||NDFRT|GUMMIFERS, ASTRAGALUS
C0949830|T121||NDFRT|ASTRAGALUS GUMMIFER LABILL.
C0330845|T121||NDFRT|ASTRAGALUS
C0330845|T121||NDFRT|ASTRAGALUS PLANTS
C0330845|T121||NDFRT|PLANT, ASTRAGALUS
C0330845|T121||NDFRT|PLANTS, ASTRAGALUS
C0330845|T121||NDFRT|ASTRAGALUS PLANT
C0330845|T121||NDFRT|ASTRAGALUS L., 1753
C0330845|T121||NDFRT|ASTRAGALUS (PLANTS)
C0330845|T121||NDFRT|ASTRAGALUS SPECIES
C0330845|T121||NDFRT|ASTRAGALUS SPECIES 
C0330845|T121||NDFRT|LOCOWEEDS
C0330845|T121||NDFRT|ASTRAGALUS 
C0330845|T121||NDFRT|ASTRAGALUS, NOS
C0330845|T121||NDFRT|LOCOWEEDS, NOS
C0949831|T121||NDFRT|MEMBRANACEUS, ASTRAGALUS
C0949831|T121||NDFRT|ASTRAGALUS MEMBRANACEUS
C0949831|T121||NDFRT|ASTRAGALUS MEMBRANACEUS MOENCH
C1135771|T121||NDFRT|LOCOWEEDS, WOOLY
C1135771|T121||NDFRT|WOOLY LOCOWEEDS
C1135771|T121||NDFRT|WOOLY LOCOWEED
C1135771|T121||NDFRT|LOCOWEED, WOOLY
C0949829|T121||NDFRT|MILK VETCH
C0949829|T121||NDFRT|MILKVETCH
C0949829|T121||NDFRT|MILK VETCHS
C0949829|T121||NDFRT|VETCHS, MILK
C0949829|T121||NDFRT|VETCH, MILK
C2757825|T121||NDFRT|ASTRAGALUS MEMBRANACEUS VAR. MONGHOLICUS (BUNGE) P.K.HSIAO
C2757825|T121||NDFRT|ASTRAGALUS PENDULIFLORUS SUBSP. MONGHOLICUS
C2757825|T121||NDFRT|ASTRAGALUS PENDULIFLORUS VAR. MONGHOLICUS
C2757825|T121||NDFRT|ASTRAGALUS PENDULIFLORUS VAR. MONGHOLICUS (BUNGE) X.Y.ZHU
C2757825|T121||NDFRT|ASTRAGALUS MONGHOLICUS BUNGE
C2757825|T121||NDFRT|ASTRAGALUS PENDULIFLORUS SUBSP. MONGHOLICUS VAR. MONGHOLICUS
C2757825|T121||NDFRT|ASTRAGALUS PENDULIFLORUS SUBSP. MONGHOLICUS (BUNGE) X.Y.ZHU
C2757825|T121||NDFRT|ASTRAGALUS MONGHOLICUS
C2757825|T121||NDFRT|ASTRAGALUS MEMBRANACEUS VAR. MONGHOLICUS
C1075624|T121||NDFRT|ASTRAGALUS MEMBRANACEUS F. PROPINQUUS
C1075624|T121||NDFRT|ASTRAGALUS MEMBRANACEUS F. PROPINQUUS (SCHISCHKIN) KITAG.
C1095897|T121|N0000022270|NDFRT|ASTRAGALUS PREPARATION|ASTRAGALUS
C1095897|T121|N0000022270|NDFRT|ASTRAGALUS|ASTRAGALUS
C1095897|T121|N0000022270|NDFRT|ASTRAGALUS |ASTRAGALUS
C1095897|T121|N0000022270|NDFRT|ASTRAGALUS EXTRACT|ASTRAGALUS
C1177063|T121|N0000163694|NDFRT|ASTRAGALUS EXTRACT PWDR|ASTRAGALUS EXTRACT PWDR [VA PRODUCT]
C1177063|T121|N0000163694|NDFRT|ASTRAGALUS EXTRACT PWDR [VA PRODUCT]|ASTRAGALUS EXTRACT PWDR [VA PRODUCT]
C3864824|T121||NDFRT|PARITAPREVIR
C3864824|T121||NDFRT|PARITAPREVIR 
C3864824|T121||NDFRT|PARITAPREVIR 
C3883274|T121||NDFRT|PARITAPREVIR DIHYDRATE
C4046856|T121||NDFRT|TECHNIVIE
C3864967|T121||NDFRT|OMBITASVIR / PARITAPREVIR / RITONAVIR
C3864967|T121||NDFRT|OMBITASVIR/PARITAPREVIR/RITONAVIR
C3864967|T121||NDFRT|OMBITASVIR + PARITAPREVIR + RITONAVIR
C3864967|T121||NDFRT|OMBITASVIR + PARITAPREVIR + RITONAVIR 
C3864967|T121||NDFRT|OMBITASVIR + PARITAPREVIR + RITONAVIR 
C4075296|T121||NDFRT|ORAL FORM PARITAPREVIR 
C4075296|T121||NDFRT|ORAL FORM PARITAPREVIR
C3865211|T121||NDFRT|OMBITASVIR / PARITAPREVIR / RITONAVIR ORAL PRODUCT
C3865211|T121||NDFRT|ORAL FORM OMBITASVIR + PARITAPREVIR + RITONAVIR
C3865211|T121||NDFRT|ORAL FORM OMBITASVIR + PARITAPREVIR + RITONAVIR 
C4046961|T121||NDFRT|OMBITASVIR 12.5 MG / PARITAPREVIR 75 MG / RITONAVIR 50 MG [TECHNIVIE]
C3865125|T121|N0000192214|NDFRT|OMBITASVIR 12.5 MG / PARITAPREVIR 75 MG / RITONAVIR 50 MG ORAL TABLET|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DAILY PACK [VA PRODUCT]
C3865125|T121|N0000192214|NDFRT|OMBITASVIR/PARITAPREVIR/RITONAVIR 12.5 MG-75 MG-50 MG ORAL TABLET|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DAILY PACK [VA PRODUCT]
C3865125|T121|N0000192214|NDFRT|OMBITASVIR, PARITAPREVIR, RITONAVIR 12.5-75-50MG ORAL TABLET|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DAILY PACK [VA PRODUCT]
C3865125|T121|N0000192214|NDFRT|OMBITASVIR-PARITAPREVIR-RITONAVIR TAB 12.5-75-50 MG|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DAILY PACK [VA PRODUCT]
C3865188|T121||NDFRT|OMBITASVIR / PARITAPREVIR / RITONAVIR ORAL TABLET
C4047089|T121||NDFRT|TECHNIVIE PILL
C4047040|T121||NDFRT|OMBITASVIR / PARITAPREVIR / RITONAVIR ORAL TABLET [TECHNIVIE]
C4047090|T121||NDFRT|TECHNIVIE ORAL PRODUCT
C3854281|T121||NDFRT|{2 (DASABUVIR 250 MG ORAL TABLET) / 2 (OMBITASVIR 12.5 MG / PARITAPREVIR 75 MG / RITONAVIR 50 MG ORAL TABLET) } PACK [VIEKIRA PAK]
C3854281|T121||NDFRT|VIEKIRA PAK
C3854281|T121||NDFRT|VIEKIRA PAK KIT
C3854281|T121||NDFRT|VIEKIRA PAK, ORAL KIT
C3854281|T121||NDFRT|DASABUVIR;OMBITASVIR/PARITAPREVIR/RITONAVIR NA ORAL TABLET [VIEKIRA PAK]
C3864964|T121|N0000191861|NDFRT|{2 (DASABUVIR 250 MG ORAL TABLET) / 2 (OMBITASVIR 12.5 MG / PARITAPREVIR 75 MG / RITONAVIR 50 MG ORAL TABLET) } PACK|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DOSE PACK,56 [VA PRODUCT]
C3864964|T121|N0000191861|NDFRT|OMBITAS-PARITAPRE-RITON & DASAB TAB PAK 12.5-75-50 & 250 MG|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DOSE PACK,56 [VA PRODUCT]
C3864964|T121|N0000191861|NDFRT|DASABUVIR/OMBITASVIR/PARITAPREVIR/RITONAVIR DAILY DOSE PACK [VA PRODUCT]|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DOSE PACK,56 [VA PRODUCT]
C3864964|T121|N0000191861|NDFRT|VIEKIRA DAILY PAK|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DOSE PACK,56 [VA PRODUCT]
C3864964|T121|N0000191861|NDFRT|DASABUVIR/OMBITASVIR/PARITAPREVIR/RITONAVIR DAILY DOSE PACK|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DOSE PACK,56 [VA PRODUCT]
C3864964|T121|N0000191861|NDFRT|TECHNIVIE DOSE PACK,56|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DOSE PACK,56 [VA PRODUCT]
C3864964|T121|N0000191861|NDFRT|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DOSE PACK,56|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DOSE PACK,56 [VA PRODUCT]
C3864964|T121|N0000191861|NDFRT|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DOSE PACK,56 [VA PRODUCT]|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DOSE PACK,56 [VA PRODUCT]
C3864964|T121|N0000191861|NDFRT|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DAILY PACK [VA PRODUCT]|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DOSE PACK,56 [VA PRODUCT]
C3864964|T121|N0000191861|NDFRT|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DAILY PACK|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DOSE PACK,56 [VA PRODUCT]
C3864964|T121|N0000191861|NDFRT|TECHNIVIE DAILY PACK|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DOSE PACK,56 [VA PRODUCT]
C4046169|T121||NDFRT|TECHNIVIE 12.5 MG / 75 MG / 50 MG ORAL TABLET
C4046169|T121||NDFRT|TECHNIVIE KIT
C4046169|T121||NDFRT|RITONAVIR 50 MG / OMBITASVIR HEMINONAHYDRATE 12.5 MG / PARITAPREVIR DIHYDRATE 75 MG ORAL TABLET, FILM COATED [TECHNIVIE]
C4046169|T121||NDFRT|TECHNIVIE 12.5MG-75MG-50MG TABLET
C4046169|T121||NDFRT|OMBITASVIR/PARITAPREVIR/RITONAVIR 12.5 MG-75 MG-50 MG ORAL TABLET [TECHNIVIE]
C4046169|T121||NDFRT|OMBITASVIR 12.5 MG / PARITAPREVIR 75 MG / RITONAVIR 50 MG ORAL TABLET [TECHNIVIE]
C4046169|T121||NDFRT|TECHNIVIE, 12.5 MG-75 MG-50 MG ORAL TABLET
C4080053|T121||NDFRT|GRAZOPREVIR
C4080455|T121||NDFRT|ZEPATIER
C4080456|T121||NDFRT|ELBASVIR 50 MG / GRAZOPREVIR 100 MG [ZEPATIER]
C4080458|T121||NDFRT|ZEPATIER ORAL PRODUCT
C4080452|T121||NDFRT|ELBASVIR / GRAZOPREVIR ORAL TABLET
C4080454|T121|N0000192438|NDFRT|ELBASVIR, GRAZOPREVIR 50-100MG ORAL TABLET|ELBASVIR 50MG/GRAZOPREVIR 100MG TAB [VA PRODUCT]
C4080454|T121|N0000192438|NDFRT|ELBASVIR/GRAZOPREVIR 50 MG-100 MG ORAL TABLET|ELBASVIR 50MG/GRAZOPREVIR 100MG TAB [VA PRODUCT]
C4080454|T121|N0000192438|NDFRT|ELBASVIR 50 MG / GRAZOPREVIR 100 MG ORAL TABLET|ELBASVIR 50MG/GRAZOPREVIR 100MG TAB [VA PRODUCT]
C4080459|T121||NDFRT|ZEPATIER PILL
C4080457|T121||NDFRT|ELBASVIR / GRAZOPREVIR ORAL TABLET [ZEPATIER]
C4080460|T121||NDFRT|ZEPATIER 50MG-100MG TABLET
C4080460|T121||NDFRT|ZEPATIER 50 MG / 100 MG ORAL TABLET
C4080460|T121||NDFRT|ZEPATIER (ELBASVIR 50 MG / GRAZOPREVIR 100 MG) ORAL TABLET
C4080460|T121||NDFRT|ELBASVIR 50 MG / GRAZOPREVIR 100 MG ORAL TABLET, FILM COATED [ZEPATIER]
C4080460|T121||NDFRT|ELBASVIR/GRAZOPREVIR 50 MG-100 MG ORAL TABLET [ZEPATIER]
C4080460|T121||NDFRT|ELBASVIR 50 MG / GRAZOPREVIR 100 MG ORAL TABLET [ZEPATIER]
C2976304|T121||NDFRT|PSI-7977
C2976304|T121||NDFRT|7977, PSI
C2976304|T121||NDFRT|PSI7977
C2976304|T121||NDFRT|PSI 7977
C3530149|T121||NDFRT|GS-7977
C3530149|T121||NDFRT|GS7977
C3530149|T121||NDFRT|GS 7977
C2976303|T121|N0000191981|NDFRT|L-ALANINE, N-[[P(S),2'R]-2'-DEOXY-2'-FLUORO-2'-METHYL-P-PHENYL-5'-URIDYLYL]-, 1-METHYLETHYL ESTER|SOFOSBUVIR [CHEMICAL/INGREDIENT]
C2976303|T121|N0000191981|NDFRT|SOFOSBUVIR|SOFOSBUVIR [CHEMICAL/INGREDIENT]
C2976303|T121|N0000191981|NDFRT|ANTIVIRALS SOFOSBUVIR|SOFOSBUVIR [CHEMICAL/INGREDIENT]
C2976303|T121|N0000191981|NDFRT|SOFOSBUVIR |SOFOSBUVIR [CHEMICAL/INGREDIENT]
C2976303|T121|N0000191981|NDFRT|SOFOSBUVIR |SOFOSBUVIR [CHEMICAL/INGREDIENT]
C2976303|T121|N0000191981|NDFRT|2-((5-(2,4-DIOXO-3,4-DIHYDRO-2H-PYRIMIDIN-1-YL)-4-FLUORO-3-HYDROXY-4-METHYLTETRAHYDROFURAN-2-YLMETHOXY)PHENOXYPHOSPHORYLAMINO)PROPIONIC ACID ISOPROPYL ESTER|SOFOSBUVIR [CHEMICAL/INGREDIENT]
C2976303|T121|N0000191981|NDFRT|SOFOSBUVIR [CHEMICAL/INGREDIENT]|SOFOSBUVIR [CHEMICAL/INGREDIENT]
C2976303|T121|N0000191981|NDFRT|SOFOSBUVIR |SOFOSBUVIR [CHEMICAL/INGREDIENT]
C3700471|T121||NDFRT|SOVALDI
C3858025|T121||NDFRT|HARVONI
C3858051|T121||NDFRT|LEDIPASVIR / SOFOSBUVIR
C3858051|T121||NDFRT|LEDIPASVIR-SOFOSBUVIR
C3858051|T121||NDFRT|LEDIPASVIR/SOFOSBUVIR
C3858051|T121||NDFRT|LEDIPASVIR + SOFOSBUVIR
C3858051|T121||NDFRT|ANTIVIRAL LEDIPASVIR + SOFOSBUVIR
C3858051|T121||NDFRT|LEDIPASVIR + SOFOSBUVIR 
C3858051|T121||NDFRT|LEDIPASVIR, SOFOSBUVIR DRUG COMBINATION
C3858051|T121||NDFRT|LEDIPASVIR - SOFOSBUVIR
C3858051|T121||NDFRT|LEDIPASVIR + SOFOSBUVIR 
C3696724|T121||NDFRT|SOFOSBUVIR ORAL PRODUCT
C3696724|T121||NDFRT|ORAL FORM SOFOSBUVIR
C3696724|T121||NDFRT|ORAL FORM SOFOSBUVIR 
C3857383|T121||NDFRT|LEDIPASVIR 90 MG / SOFOSBUVIR 400 MG ORAL TABLET [HARVONI]
C3857383|T121||NDFRT|LEDIPASVIR 90 MG / SOFOSBUVIR 400 MG ORAL TABLET, FILM COATED [HARVONI]
C3857383|T121||NDFRT|HARVONI 90 MG / 400 MG ORAL TABLET
C3857383|T121||NDFRT|HARVONI (LEDIPASVIR 90 MG / SOFOSBUVIR 400 MG) ORAL TABLET
C3857383|T121||NDFRT|HARVONI 90MG-400MG TABLET
C3857383|T121||NDFRT|LEDIPASVIR/SOFOSBUVIR 90 MG-400 MG ORAL TABLET [HARVONI]
C3857383|T121||NDFRT|HARVONI, 90 MG-400 MG ORAL TABLET
C3857383|T121||NDFRT|LEDIPASVIR 90 MG / SOFOSBUVIR 400 MG ORAL TABLET, FILM COATED [HARVONI ACCESS]
C3858162|T121||NDFRT|LEDIPASVIR / SOFOSBUVIR ORAL TABLET [HARVONI]
C3852670|T121||NDFRT|OMBITASVIR
C3852670|T121||NDFRT|OMBITASVIR 
C3852670|T121||NDFRT|OMBITASVIR 
C3883273|T121||NDFRT|OMBITASVIR HEMINONAHYDRATE
C4075325|T121||NDFRT|ORAL FORM OMBITASVIR
C4075325|T121||NDFRT|ORAL FORM OMBITASVIR 
C4080052|T121||NDFRT|ELBASVIR
C3252090|T121||NDFRT|DACLATASVIR
C3252090|T121||NDFRT|DACLATASVIR 
C3252090|T121||NDFRT|DACLATASVIR 
C3252090|T121||NDFRT|ANTIVIRAL DACLATASVIR
C3252090|T121||NDFRT|DACLATASVIR 
C3892852|T121||NDFRT|DACLATASVIR DIHYDROCHLORIDE
C3892852|T121||NDFRT|DACLATASVIR (AS DIHYDROCHLORIDE)
C4046850|T121||NDFRT|DAKLINZA
C4047230|T121||NDFRT|DACLATASVIR ORAL PRODUCT
C4047230|T121||NDFRT|ORAL FORM DACLATASVIR
C4047230|T121||NDFRT|ORAL FORM DACLATASVIR 
C4047078|T121||NDFRT|DAKLINZA PILL
C3857361|T121|N0000191806|NDFRT|DACLATASVIR 30 MG ORAL TABLET|DACLATASVIR 30MG TAB [VA PRODUCT]
C3857361|T121|N0000191806|NDFRT|DACLATASVIR DIHYDROCHLORIDE 30 MG ORAL TABLET|DACLATASVIR 30MG TAB [VA PRODUCT]
C3857361|T121|N0000191806|NDFRT|DACLATASVIR (AS DACLATASVIR DIHYDROCHLORIDE 33 MG) 30 MG ORAL TABLET|DACLATASVIR 30MG TAB [VA PRODUCT]
C3857361|T121|N0000191806|NDFRT|DACLATASVIR 30MG ORAL TABLET|DACLATASVIR 30MG TAB [VA PRODUCT]
C3857361|T121|N0000191806|NDFRT|DACLATASVIR 30MG TAB|DACLATASVIR 30MG TAB [VA PRODUCT]
C3857361|T121|N0000191806|NDFRT|DACLATASVIR DIHYDROCHLORIDE TAB 30 MG (BASE EQUIVALENT)|DACLATASVIR 30MG TAB [VA PRODUCT]
C3857361|T121|N0000191806|NDFRT|DACLATASVIR 30MG TAB [VA PRODUCT]|DACLATASVIR 30MG TAB [VA PRODUCT]
C4047197|T121||NDFRT|DACLATASVIR ORAL TABLET
C3892515|T121|N0000191807|NDFRT|DACLATASVIR DIHYDROCHLORIDE 60 MG ORAL TABLET|DACLATASVIR 60MG TAB [VA PRODUCT]
C3892515|T121|N0000191807|NDFRT|DACLATASVIR 60 MG ORAL TABLET|DACLATASVIR 60MG TAB [VA PRODUCT]
C3892515|T121|N0000191807|NDFRT|DACLATASVIR 60MG ORAL TABLET|DACLATASVIR 60MG TAB [VA PRODUCT]
C3892515|T121|N0000191807|NDFRT|DACLATASVIR (AS DACLATASVIR DIHYDROCHLORIDE 66 MG) 60 MG ORAL TABLET|DACLATASVIR 60MG TAB [VA PRODUCT]
C3892515|T121|N0000191807|NDFRT|DACLATASVIR 60MG TAB|DACLATASVIR 60MG TAB [VA PRODUCT]
C3892515|T121|N0000191807|NDFRT|DACLATASVIR DIHYDROCHLORIDE TAB 60 MG (BASE EQUIVALENT)|DACLATASVIR 60MG TAB [VA PRODUCT]
C3892515|T121|N0000191807|NDFRT|DACLATASVIR 60MG TAB [VA PRODUCT]|DACLATASVIR 60MG TAB [VA PRODUCT]
C3852655|T121||NDFRT|GS-5885
C3851350|T121||NDFRT|LEDIPASVIR
C3851350|T121||NDFRT|LEDIPASVIR 
C3851350|T121||NDFRT|LEDIPASVIR 
C4075037|T121||NDFRT|ORAL FORM LEDIPASVIR 
C4075037|T121||NDFRT|ORAL FORM LEDIPASVIR
C3858322|T121||NDFRT|LEDIPASVIR / SOFOSBUVIR ORAL PRODUCT
C3858322|T121||NDFRT|ORAL FORM LEDIPASVIR + SOFOSBUVIR
C3858322|T121||NDFRT|ORAL FORM LEDIPASVIR + SOFOSBUVIR 
C3858113|T121||NDFRT|LEDIPASVIR 90 MG / SOFOSBUVIR 400 MG [HARVONI]
C3858080|T121|N0000191202|NDFRT|LEDIPASVIR 90 MG / SOFOSBUVIR 400 MG ORAL TABLET|LEDIPASVIR 90MG/SOFOSBUVIR 400MG TAB [VA PRODUCT]
C3858080|T121|N0000191202|NDFRT|LEDIPASVIR, SOFOSBUVIR 90-400MG ORAL TABLET|LEDIPASVIR 90MG/SOFOSBUVIR 400MG TAB [VA PRODUCT]
C3858080|T121|N0000191202|NDFRT|LEDIPASVIR-SOFOSBUVIR TAB 90-400 MG|LEDIPASVIR 90MG/SOFOSBUVIR 400MG TAB [VA PRODUCT]
C3858080|T121|N0000191202|NDFRT|LEDIPASVIR-SOFOSBUVIR 90 MG-400 MG ORAL TABLET|LEDIPASVIR 90MG/SOFOSBUVIR 400MG TAB [VA PRODUCT]
C3858080|T121|N0000191202|NDFRT|LEDIPASVIR/SOFOSBUVIR 90 MG-400 MG ORAL TABLET|LEDIPASVIR 90MG/SOFOSBUVIR 400MG TAB [VA PRODUCT]
C3858080|T121|N0000191202|NDFRT|LEDIPASVIR 90MG/SOFOSBUVIR 400MG TAB|LEDIPASVIR 90MG/SOFOSBUVIR 400MG TAB [VA PRODUCT]
C3858080|T121|N0000191202|NDFRT|LEDIPASVIR 90MG/SOFOSBUVIR 400MG TAB [VA PRODUCT]|LEDIPASVIR 90MG/SOFOSBUVIR 400MG TAB [VA PRODUCT]
C3858300|T121||NDFRT|LEDIPASVIR / SOFOSBUVIR ORAL TABLET
C3858199|T121||NDFRT|HARVONI PILL
C3858200|T121||NDFRT|HARVONI ORAL PRODUCT
