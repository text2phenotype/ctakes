C0019029|T034||LNC|HEMOGLOBIN CONCENTRATION RESULT
C0019046|T034|LP32067-8|LNC|HEMOGLOBIN|HEMOGLOBIN
C0518015|T034||LNC|HEMOGLOBIN MEASUREMENT
C0019047|T034||LNC|ABNORMAL HAEMOGLOBIN
C0019047|T034||LNC|ABNORMAL HEMOGLOBIN
C0019047|T034||LNC|ABNORMAL HEMOGLOBIN 
C0019047|T034||LNC|ABNORMAL HEMOGLOBIN, NOS
C0019046|T034|LP32067-8|LNC|HEMOGLOBIN|HEMOGLOBIN
C0019046|T034|LP32067-8|LNC|HGB|HEMOGLOBIN
C0019046|T034|LP32067-8|LNC|HB|HEMOGLOBIN
C0019046|T034|LP32067-8|LNC|HAEMOGLOBIN|HEMOGLOBIN
C0019046|T034|LP32067-8|LNC|HB - HAEMOGLOBIN|HEMOGLOBIN
C0019046|T034|LP32067-8|LNC|HB - HEMOGLOBIN|HEMOGLOBIN
C0019046|T034|LP32067-8|LNC|HGB - HAEMOGLOBIN|HEMOGLOBIN
C0019046|T034|LP32067-8|LNC|HGB - HEMOGLOBIN|HEMOGLOBIN
C0019046|T034|LP32067-8|LNC|HEMOGLOBIN |HEMOGLOBIN
C0019046|T034|LP32067-8|LNC|HEMOGLOBIN, NOS|HEMOGLOBIN
C0019046|T034|LP32067-8|LNC|HAEMOGLOBIN, NOS|HEMOGLOBIN
C1988917|T034|LP49432-5|LNC|HEMOGLOBIN &#X7C; BLOOD VENOUS|HEMOGLOBIN &#X7C; BLOOD VENOUS
C1988910|T034|LP43135-0|LNC|HEMOGLOBIN &#X7C; BLD-SER-PLAS|HEMOGLOBIN &#X7C; BLD-SER-PLAS
C1988911|T034|LP43637-5|LNC|HEMOGLOBIN &#X7C; BLOOD ARTERIAL|HEMOGLOBIN &#X7C; BLOOD ARTERIAL
C1988916|T034|LP49433-3|LNC|HEMOGLOBIN &#X7C; BLOOD MIXED VENOUS|HEMOGLOBIN &#X7C; BLOOD MIXED VENOUS
C1988912|T034|LP49434-1|LNC|HEMOGLOBIN &#X7C; BLOOD CAPILLARY|HEMOGLOBIN &#X7C; BLOOD CAPILLARY
C0518015|T034||LNC|HAEMOGLOBIN
C0518015|T034||LNC|HAEM
C0518015|T034||LNC|HEMOGLOBIN MEASUREMENT
C0518015|T034||LNC|HEMOGLOBIN
C0518015|T034||LNC|HEMOGLOBIN MEASUREMENT 
C0518015|T034||LNC|TEST;HAEMOGLOBIN
C0518015|T034||LNC|BLOOD COUNT HEMOGLOBIN
C0518015|T034||LNC|HEMOGLOBIN LEVEL
C0518015|T034||LNC|MEASUREMENT OF HEMOGLOBIN (HGB)
C0518015|T034||LNC|HEMOGLOBIN DETERMINATION 
C0518015|T034||LNC|HEMOGLOBIN DETERMINATION
C0518015|T034||LNC|HAEMOGLOBIN DETERMINATION
C0518015|T034||LNC|HGB
C0518015|T034||LNC|BLOOD COUNT; HEMOGLOBIN (HGB)
C0518015|T034||LNC|FHGB
C0518015|T034||LNC|HEMOGLOBIN DETERMINATION, NOS
C0518015|T034||LNC|HAEMOGLOBIN DETERMINATION, NOS
C0518015|T034||LNC|TEST;HEMOGLOBIN
C0518015|T034||LNC|HAEMOGLOBIN TEST
C0518015|T034||LNC|HEMOGLOBIN TEST
C0587341|T034||LNC|HB ESTIMATION
C0587341|T034||LNC|HAEMOGLOBIN ESTIMATION
C0587341|T034||LNC|HEMOGLOBIN ESTIMATION
C0587341|T034||LNC|HEMOGLOBIN ESTIMATION NOS
C0587341|T034||LNC|HAEMOGLOBIN ESTIMATION NOS
C0587341|T034||LNC|HEMOGLOBIN ESTIMATION (& LEVEL)
C0587341|T034||LNC|HAEMOGLOBIN ESTIMATION (& LEVEL) 
C0587341|T034||LNC|HEMOGLOBIN ESTIMATION NOS 
C0587341|T034||LNC|HAEMOGLOBIN ESTIMATION NOS 
C0587341|T034||LNC|HAEMOGLOBIN ESTIMATION (& LEVEL)
C0587341|T034||LNC|HAEMOGLOBIN ESTIMATION LEVEL
C0587341|T034||LNC|HEMOGLOBIN ESTIMATION LEVEL
C0587341|T034||LNC|HAEMOGLOBIN LEVEL ESTIMATION
C0587341|T034||LNC|HB ESTIMATION 
C0587341|T034||LNC|HEMOGLOBIN LEVEL ESTIMATION 
C0587341|T034||LNC|HEMOGLOBIN LEVEL ESTIMATION
C0474563|T034||LNC|HEMOGLOBIN; PLASMA
C0474563|T034||LNC|MEASUREMENT OF TOTAL HEMOGLOBIN CONCENTRATION IN PLASMA SPECIMEN
C0474563|T034||LNC|MEASUREMENT OF TOTAL HAEMOGLOBIN CONCENTRATION IN PLASMA SPECIMEN
C0474563|T034||LNC|HAEMOGLOBIN DETERMINATION, PLASMA
C0474563|T034||LNC|HEMOGLOBIN DETERMINATION, PLASMA 
C0474563|T034||LNC|MEASUREMENT OF TOTAL HEMOGLOBIN CONCENTRATION IN PLASMA SPECIMEN 
C0474563|T034||LNC|HEMOGLOBIN DETERMINATION, PLASMA
C0474563|T034||LNC|PLASMA HEMOGLOBIN MEASUREMENT 
C0474563|T034||LNC|PLASMA HEMOGLOBIN MEASUREMENT
C0474563|T034||LNC|MEASUREMENT OF HEMOGLOBIN IN PLASMA
C0474563|T034||LNC|PLASMA HEMOGLOBIN LEVEL
C0474563|T034||LNC|ASSAY OF HEMOGLOBIN PLASMA
C0474563|T034||LNC|PLASMA HEMOGLOBINS TEST
C0474563|T034||LNC|PLASMA HAEMOGLOBIN LEVEL
C0474563|T034||LNC|ASSAY OF PLASMA HEMOGLOBIN
C4066087|T034||LNC|CALCULATED HEMOGLOBIN LEVEL
C4066087|T034||LNC|HEMOGLOBIN CALCULATED
C4066087|T034||LNC|CALCULATED HEMOGLOBIN LEVEL 
C0200694|T034||LNC|MEASUREMENT OF TOTAL HEMOGLOBIN CONCENTRATION AND HEMATOCRIT 
C0200694|T034||LNC|HEMOGLOBIN AND HEMATOCRIT DETERMINATION
C0200694|T034||LNC|MEASUREMENT OF TOTAL HEMOGLOBIN CONCENTRATION AND HEMATOCRIT
C0200694|T034||LNC|MEASUREMENT OF TOTAL HAEMOGLOBIN CONCENTRATION AND HAEMATOCRIT
C0200694|T034||LNC|HEMOGLOBIN AND HEMATOCRIT DETERMINATION 
C0200694|T034||LNC|HAEMOGLOBIN AND HAEMATOCRIT DETERMINATION
C0200694|T034||LNC|H & H DETERMINATION
C0200694|T034||LNC|TOTAL HEMOGLOBIN CONCENTRATION AND HEMATOCRIT
C0200694|T034||LNC|TOTAL HEMOGLOBIN CONCENTRATION AND HEMATOCRIT 
C0200694|T034||LNC|HAEMOGLOBIN AND HEMATOCRIT DETERMINATION
C0523149|T034||LNC|SEMI-QUANTITATIVE MEASUREMENT OF TOTAL HAEMOGLOBIN IN BLOOD SPECIMEN
C0523149|T034||LNC|SEMI-QUANTITATIVE MEASUREMENT OF TOTAL HEMOGLOBIN IN BLOOD SPECIMEN
C0523149|T034||LNC|HAEMOGLOBIN DETERMINATION, BLOOD, SEMI-QUANTITATIVE
C0523149|T034||LNC|SEMI-QUANTITATIVE MEASUREMENT OF TOTAL HEMOGLOBIN IN BLOOD SPECIMEN 
C0523149|T034||LNC|HEMOGLOBIN DETERMINATION, BLOOD, SEMI-QUANTITATIVE 
C0523149|T034||LNC|HEMOGLOBIN DETERMINATION, BLOOD, SEMI-QUANTITATIVE
C1314664|T034||LNC|HAEMOGLOBIN CONCENTRATION
C1314664|T034||LNC|HEMOGLOBIN LEVEL
C1314664|T034||LNC|HAEMOGLOBIN LEVEL
C1314664|T034||LNC|HB - HAEMOGLOBIN LEVEL
C1314664|T034||LNC|HB - HEMOGLOBIN CONCENTRATION
C1314664|T034||LNC|HB - HEMOGLOBIN LEVEL
C1314664|T034||LNC|HB - HAEMOGLOBIN CONCENTRATION
C1314664|T034||LNC|HEMOGLOBIN CONCENTRATION
