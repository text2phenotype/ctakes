C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE AIRWAY DISEASE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0034067|T047|155573002|SNOMEDCT_US|EMPHYSEMA|EMPHYSEMA (DISORDER)
C0034067|T047|155573002|SNOMEDCT_US|PULMONARY EMPHYSEMA|EMPHYSEMA (DISORDER)
C0034067|T047|155573002|SNOMEDCT_US|EMPHYSEMA, UNSPECIFIED|EMPHYSEMA (DISORDER)
C0034067|T047|155573002|SNOMEDCT_US|EMPHYSEMAS PULM|EMPHYSEMA (DISORDER)
C0034067|T047|155573002|SNOMEDCT_US|EMPHYSEMA PULM|EMPHYSEMA (DISORDER)
C0034067|T047|155573002|SNOMEDCT_US|PULM EMPHYSEMAS|EMPHYSEMA (DISORDER)
C0034067|T047|155573002|SNOMEDCT_US|PULM EMPHYSEMA|EMPHYSEMA (DISORDER)
C0034067|T047|155573002|SNOMEDCT_US|EMPHYSEMA |EMPHYSEMA (DISORDER)
C0034067|T047|155573002|SNOMEDCT_US|EMPHYSEMA (LUNG)(PULMONARY) NOS|EMPHYSEMA (DISORDER)
C0034067|T047|155573002|SNOMEDCT_US|EMPHYSEMAS, PULMONARY|EMPHYSEMA (DISORDER)
C0034067|T047|155573002|SNOMEDCT_US|PULMONARY EMPHYSEMAS|EMPHYSEMA (DISORDER)
C0034067|T047|155573002|SNOMEDCT_US|PULMONARY EMPHYSEMA [DISEASE/FINDING]|EMPHYSEMA (DISORDER)
C0034067|T047|155573002|SNOMEDCT_US|EMPHYSEMA, PULMONARY|EMPHYSEMA (DISORDER)
C0034067|T047|155573002|SNOMEDCT_US|EMPHYSEMA |EMPHYSEMA (DISORDER)
C0034067|T047|155573002|SNOMEDCT_US|EMPHYSEMA PULMONARY|EMPHYSEMA (DISORDER)
C0034067|T047|155573002|SNOMEDCT_US|EMPHYSEMA OF LUNG|EMPHYSEMA (DISORDER)
C0034067|T047|155573002|SNOMEDCT_US|PULMONARY EMPHYSEMA |EMPHYSEMA (DISORDER)
C0034067|T047|155573002|SNOMEDCT_US|EMPHYSEMA OF LUNG, NOS|EMPHYSEMA (DISORDER)
C0034067|T047|155573002|SNOMEDCT_US|PULMONARY EMPHYSEMA, NOS|EMPHYSEMA (DISORDER)
C0034067|T047|155573002|SNOMEDCT_US|EMPHYSEMA (PULMONARY)|EMPHYSEMA (DISORDER)
C0008677|T047|63480004|SNOMEDCT_US|UNSPECIFIED CHRONIC BRONCHITIS|CHRONIC BRONCHITIS (DISORDER)
C0008677|T047|63480004|SNOMEDCT_US|CHRONIC BRONCHITIS|CHRONIC BRONCHITIS (DISORDER)
C0008677|T047|63480004|SNOMEDCT_US|CHRONIC BRONCHITIS |CHRONIC BRONCHITIS (DISORDER)
C0008677|T047|63480004|SNOMEDCT_US|CHRONIC BRONCHITIS NOS|CHRONIC BRONCHITIS (DISORDER)
C0008677|T047|63480004|SNOMEDCT_US|BRONCHITIS, CHRONIC|CHRONIC BRONCHITIS (DISORDER)
C0008677|T047|63480004|SNOMEDCT_US|BRONCHITIS, CHRONIC [DISEASE/FINDING]|CHRONIC BRONCHITIS (DISORDER)
C0008677|T047|63480004|SNOMEDCT_US|BRONCHITIS;CHRONIC|CHRONIC BRONCHITIS (DISORDER)
C0008677|T047|63480004|SNOMEDCT_US|CHRONIC BRONCHITIS |CHRONIC BRONCHITIS (DISORDER)
C0008677|T047|63480004|SNOMEDCT_US|CHRONIC BRONCHITIS NOS |CHRONIC BRONCHITIS (DISORDER)
C0008677|T047|63480004|SNOMEDCT_US|-- CHRONIC BRONCHITIS|CHRONIC BRONCHITIS (DISORDER)
C0008677|T047|63480004|SNOMEDCT_US|CHRONIC BRONCHITIS, UNSPECIFIED|CHRONIC BRONCHITIS (DISORDER)
C0008677|T047|63480004|SNOMEDCT_US|BRONCHITIS CHRONIC|CHRONIC BRONCHITIS (DISORDER)
C0008677|T047|63480004|SNOMEDCT_US|BRONCHITIS CHRONIC NOS|CHRONIC BRONCHITIS (DISORDER)
C0008677|T047|63480004|SNOMEDCT_US|BRONCHITIS; CHRONIC|CHRONIC BRONCHITIS (DISORDER)
C0008677|T047|63480004|SNOMEDCT_US|CHRONIC; BRONCHITIS|CHRONIC BRONCHITIS (DISORDER)
C0008677|T047|63480004|SNOMEDCT_US|CHRONIC BRONCHITIS, NOS|CHRONIC BRONCHITIS (DISORDER)
C0024117|T047|413846005|SNOMEDCT_US|COPD|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|PULMONARY DISEASE, CHRONIC OBSTRUCTIVE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMONARY DISEASE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE AIRWAY DISEASE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMONARY DISEASE, UNSPECIFIED|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE LUNG DISEASE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE AIRWAYS DISEASE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE LUNG DIS|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|PULM DIS CHRONIC OBSTRUCTIVE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULM DIS|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE AIRWAY DIS|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|COLD (CHRONIC OBSTRUCTIVE LUNG DISEASE)|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMONARY DISEASE |CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMONARY DISEASE (COPD)|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE AIRWAY DISEASE NOS|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE LUNG DISEASE NOS|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|PULMONARY DISEASE, CHRONIC OBSTRUCTIVE [DISEASE/FINDING]|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|LESS PREFERRED TERM|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC AIRWAYS DISEASE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE AIRWAYS DISEASE NOS |CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE LUNG DISEASE |CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE AIRWAYS DISEASE NOS|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMONARY DISEASE NOS|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|-- COPD|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|OBSTRUCTIVE PULMONARY DISEASE (COPD), CHRONIC|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|COPD, CHRONIC OBSTRUCTIVE PULMONARY DISEASE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|PULMONARY DISEASE (COPD), CHRONIC OBSTRUCTIVE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMONARY DISEASE, (COPD)|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|DISEASE (COPD), CHRONIC OBSTRUCTIVE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING |CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCT AIRWAYS DISEASE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE BRONCHOPNEUMOPATHY|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|OBSTRUCTIVE AIRWAYS DISEASE (CHRONIC)|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC AIRFLOW LIMITATION|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC AIRWAY OBSTRUCTION|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|COAD - CHRONIC OBSTRUCTIVE AIRWAYS DISEASE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|COLD - CHRONIC OBSTRUCTIVE LUNG DISEASE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|COPD - CHRONIC OBSTRUCTIVE PULMONARY DISEASE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC AIRWAY DISEASE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC IRREVERSIBLE AIRWAY OBSTRUCTION|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CAFL - CHRONIC AIRFLOW LIMITATION|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CAL - CHRONIC AIRFLOW LIMITATION|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|DISEASE (OR DISORDER); RESPIRATORY TRACT, CHRONIC, OBSTRUCTIVE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|DISEASE (OR DISORDER); RESPIRATORY TRACT, OBSTRUCTIVE, CHRONIC|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|LUNG; DISEASE, OBSTRUCTIVE (CHRONIC)|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|LUNG; OBSTRUCTION, DISEASE, CHRONIC|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|OBSTRUCTION; AIRWAY, CHRONIC|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|OBSTRUCTION; LUNG, DISEASE, CHRONIC|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|AIRWAY; OBSTRUCTION, CHRONIC|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|RESPIRATORY TRACT; DISORDER, CHRONIC, OBSTRUCTIVE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|RESPIRATORY TRACT; DISORDER, OBSTRUCTIVE, CHRONIC|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE LUNG DISEASE, NOS|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTRUCTIVE LUNG DISEASE [AMBIGUOUS]|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC AIRWAY OBSTRUCTION; NOT OTHERWISE SPECIFIED|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|COPD NOS|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTR AIRWAYS DISEASE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTR LUNG DISEASE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0024117|T047|413846005|SNOMEDCT_US|CHRONIC OBSTR PULMON DISEASE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE FINDING
C0375334|T047||SNOMEDCT_US|CHRONIC OBSTRUCTIVE ASTHMA WITH STATUS ASTHMATICUS
C0375334|T047||SNOMEDCT_US|CHRONIC OBSTRUCTIVE ASTHMA WITH STATUS ASTHMATICUS 
C0375334|T047||SNOMEDCT_US|CH OB ASTHMA W STAT ASTH
C0348818|T047|196001008|SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMONARY DISEASE WITH ACUTE LOWER RESPIRATORY INFECTION|CHRONIC OBSTRUCTIVE PULMONARY DISEASE WITH ACUTE LOWER RESPIRATORY INFECTION (DISORDER)
C0348818|T047|196001008|SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMON DISEASE W ACUTE LOWER RESP INFCT|CHRONIC OBSTRUCTIVE PULMONARY DISEASE WITH ACUTE LOWER RESPIRATORY INFECTION (DISORDER)
C0348818|T047|196001008|SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMONARY DISEASE WITH ACUTE LOWER RESPIRATORY INFECTION |CHRONIC OBSTRUCTIVE PULMONARY DISEASE WITH ACUTE LOWER RESPIRATORY INFECTION (DISORDER)
C0348818|T047|196001008|SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMONARY DISEASE WITH ACUTE LOWER RESPIRATORY INFECTION |CHRONIC OBSTRUCTIVE PULMONARY DISEASE WITH ACUTE LOWER RESPIRATORY INFECTION (DISORDER)
C3508933|T047||SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMONARY DISEASE WITH EXACERBATION 
C3508933|T047||SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMONARY DISEASE WITH EXACERBATION
C1527303|T047|13645005|SNOMEDCT_US|AIRFLOW OBSTRUCTIONS, CHRONIC|CAO - CHRONIC AIRFLOW OBSTRUCTION
C1527303|T047|13645005|SNOMEDCT_US|CHRONIC AIRFLOW OBSTRUCTIONS|CAO - CHRONIC AIRFLOW OBSTRUCTION
C1527303|T047|13645005|SNOMEDCT_US|CHRONIC AIRFLOW OBSTRUCTION|CAO - CHRONIC AIRFLOW OBSTRUCTION
C1527303|T047|13645005|SNOMEDCT_US|CAO - CHRONIC AIRFLOW OBSTRUCTION|CAO - CHRONIC AIRFLOW OBSTRUCTION
C1527303|T047|13645005|SNOMEDCT_US|AIRFLOW OBSTRUCTION, CHRONIC|CAO - CHRONIC AIRFLOW OBSTRUCTION
C3714496|T047|10169006|SNOMEDCT_US|CHRONIC AIRWAY DISEASE|CHRONIC OBSTRUCTIVE PULMONARY DISEASE OF HORSES
C3714496|T047|10169006|SNOMEDCT_US|COPD|CHRONIC OBSTRUCTIVE PULMONARY DISEASE OF HORSES
C0348693|T047|196231009|SNOMEDCT_US|OTHER SPECIFIED CHRONIC OBSTRUCTIVE PULMONARY DISEASE|[X]OTHER SPECIFIED CHRONIC OBSTRUCTIVE PULMONARY DISEASE (DISORDER)
C0348693|T047|196231009|SNOMEDCT_US|OTHER SPECIFIED CHRONIC OBSTRUCTIVE AIRWAYS DISEASE|[X]OTHER SPECIFIED CHRONIC OBSTRUCTIVE PULMONARY DISEASE (DISORDER)
C0348693|T047|196231009|SNOMEDCT_US|[X]OTHER SPECIFIED CHRONIC OBSTRUCTIVE PULMONARY DISEASE |[X]OTHER SPECIFIED CHRONIC OBSTRUCTIVE PULMONARY DISEASE (DISORDER)
C0348693|T047|196231009|SNOMEDCT_US|OTHER SPECIFIED CHRONIC OBSTRUCTIVE AIRWAYS DISEASE |[X]OTHER SPECIFIED CHRONIC OBSTRUCTIVE PULMONARY DISEASE (DISORDER)
C0348693|T047|196231009|SNOMEDCT_US|[X]OTHER SPECIFIED CHRONIC OBSTRUCTIVE PULMONARY DISEASE|[X]OTHER SPECIFIED CHRONIC OBSTRUCTIVE PULMONARY DISEASE (DISORDER)
C0155874|T047|195950008|SNOMEDCT_US|OBSTRUCTIVE CHRONIC BRONCHITIS|EMPHYSEMATOUS BRONCHITIS (DISORDER)
C0155874|T047|195950008|SNOMEDCT_US|CHRONIC OBSTRUCTIVE BRONCHITIS|EMPHYSEMATOUS BRONCHITIS (DISORDER)
C0155874|T047|195950008|SNOMEDCT_US|CHRONIC BRONCHITIS WITH EMPHYSEMA|EMPHYSEMATOUS BRONCHITIS (DISORDER)
C0155874|T047|195950008|SNOMEDCT_US|EMPHYSEMATOUS BRONCHITIS|EMPHYSEMATOUS BRONCHITIS (DISORDER)
C0155874|T047|195950008|SNOMEDCT_US|CHRONIC OBSTRUCTIVE BRONCHITIS |EMPHYSEMATOUS BRONCHITIS (DISORDER)
C0155874|T047|195950008|SNOMEDCT_US|OBSTRUCTIVE CHRONIC BRONCHITIS NOS |EMPHYSEMATOUS BRONCHITIS (DISORDER)
C0155874|T047|195950008|SNOMEDCT_US|EMPHYSEMATOUS BRONCHITIS |EMPHYSEMATOUS BRONCHITIS (DISORDER)
C0155874|T047|195950008|SNOMEDCT_US|OBSTRUCTIVE CHRONIC BRONCHITIS NOS|EMPHYSEMATOUS BRONCHITIS (DISORDER)
C0155874|T047|195950008|SNOMEDCT_US|BRONCHITIS WITH AIRWAY OBSTRUCTION|EMPHYSEMATOUS BRONCHITIS (DISORDER)
C0155874|T047|195950008|SNOMEDCT_US|COB - CHRONIC OBSTRUCTIVE BRONCHITIS|EMPHYSEMATOUS BRONCHITIS (DISORDER)
C0155874|T047|195950008|SNOMEDCT_US|BRONCHITIS; CHRONIC, OBSTRUCTIVE|EMPHYSEMATOUS BRONCHITIS (DISORDER)
C0155874|T047|195950008|SNOMEDCT_US|BRONCHITIS; EMPHYSEMATOUS|EMPHYSEMATOUS BRONCHITIS (DISORDER)
C0155874|T047|195950008|SNOMEDCT_US|CHRONIC; BRONCHITIS, OBSTRUCTIVE|EMPHYSEMATOUS BRONCHITIS (DISORDER)
C0155874|T047|195950008|SNOMEDCT_US|EMPHYSEMATOUS; BRONCHITIS|EMPHYSEMATOUS BRONCHITIS (DISORDER)
C0155874|T047|195950008|SNOMEDCT_US|CHRONIC OBSTRUCTIVE BRONCHITIS  [AMBIGUOUS]|EMPHYSEMATOUS BRONCHITIS (DISORDER)
C0155874|T047|195950008|SNOMEDCT_US|CHRONIC BRONCHITIS & EMPHYSEMA|EMPHYSEMATOUS BRONCHITIS (DISORDER)
C0155874|T047|195950008|SNOMEDCT_US|EMPHYSEMA WITH CHRONIC BRONCHITIS|EMPHYSEMATOUS BRONCHITIS (DISORDER)
C0155874|T047|195950008|SNOMEDCT_US|CHRONIC BRONCHITIS, OBSTRUCTIVE|EMPHYSEMATOUS BRONCHITIS (DISORDER)
C0155874|T047|195950008|SNOMEDCT_US|BRONCHITIS WITH EMPHYSEMA|EMPHYSEMATOUS BRONCHITIS (DISORDER)
C0155874|T047|195950008|SNOMEDCT_US|BRONCHITIS, EMPHYSEMATOUS|EMPHYSEMATOUS BRONCHITIS (DISORDER)
C0730607|T047|313299006|SNOMEDCT_US|SEVERE CHRONIC OBSTRUCTIVE PULMONARY DISEASE|SEVERE CHRONIC OBSTRUCTIVE PULMONARY DISEASE (DISORDER)
C0730607|T047|313299006|SNOMEDCT_US|SEVERE CHRONIC OBSTRUCTIVE PULMONARY DISEASE |SEVERE CHRONIC OBSTRUCTIVE PULMONARY DISEASE (DISORDER)
C0730607|T047|313299006|SNOMEDCT_US|SEVERE CHRONIC OBSTRUCTIVE PULMONARY DISEASE |SEVERE CHRONIC OBSTRUCTIVE PULMONARY DISEASE (DISORDER)
C0730607|T047|313299006|SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMONARY DISEASE SEVERE|SEVERE CHRONIC OBSTRUCTIVE PULMONARY DISEASE (DISORDER)
C0730604|T047|313296004|SNOMEDCT_US|MILD CHRONIC OBSTRUCTIVE PULMONARY DISEASE|MILD CHRONIC OBSTRUCTIVE PULMONARY DISEASE (DISORDER)
C0730604|T047|313296004|SNOMEDCT_US|MILD CHRONIC OBSTRUCTIVE PULMONARY DISEASE |MILD CHRONIC OBSTRUCTIVE PULMONARY DISEASE (DISORDER)
C0730604|T047|313296004|SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMONARY DISEASE MILD|MILD CHRONIC OBSTRUCTIVE PULMONARY DISEASE (DISORDER)
C0730604|T047|313296004|SNOMEDCT_US|MILD CHRONIC OBSTRUCTIVE PULMONARY DISEASE |MILD CHRONIC OBSTRUCTIVE PULMONARY DISEASE (DISORDER)
C0730605|T047|313297008|SNOMEDCT_US|MODERATE CHRONIC OBSTRUCTIVE PULMONARY DISEASE |MODERATE CHRONIC OBSTRUCTIVE PULMONARY DISEASE (DISORDER)
C0730605|T047|313297008|SNOMEDCT_US|MODERATE CHRONIC OBSTRUCTIVE PULMONARY DISEASE|MODERATE CHRONIC OBSTRUCTIVE PULMONARY DISEASE (DISORDER)
C0730605|T047|313297008|SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMONARY DISEASE MODERATE|MODERATE CHRONIC OBSTRUCTIVE PULMONARY DISEASE (DISORDER)
C0730605|T047|313297008|SNOMEDCT_US|MODERATE CHRONIC OBSTRUCTIVE PULMONARY DISEASE |MODERATE CHRONIC OBSTRUCTIVE PULMONARY DISEASE (DISORDER)
C3662842|T047|1761000119103|SNOMEDCT_US|CHRONIC OBSTRUCTIVE AIRWAY DISEASE WITH ASTHMA |CHRONIC OBSTRUCTIVE AIRWAY DISEASE WITH ASTHMA (DISORDER)
C3662842|T047|1761000119103|SNOMEDCT_US|CHRONIC OBSTRUCTIVE AIRWAY DISEASE WITH ASTHMA|CHRONIC OBSTRUCTIVE AIRWAY DISEASE WITH ASTHMA (DISORDER)
C1847014|T047||SNOMEDCT_US|PULMONARY DISEASE, CHRONIC OBSTRUCTIVE, SEVERE EARLY-ONSET
C0494659|T047||SNOMEDCT_US|OTHER CHRONIC OBSTRUCTIVE PULMONARY DISEASE
C0029607|T047|196230005|SNOMEDCT_US|OTHER EMPHYSEMA|[X]OTHER EMPHYSEMA (MORPHOLOGIC ABNORMALITY)
C0029607|T047|196230005|SNOMEDCT_US|EMPHYSEMA NEC|[X]OTHER EMPHYSEMA (MORPHOLOGIC ABNORMALITY)
C0029607|T047|196230005|SNOMEDCT_US|OTHER EMPHYSEMA (MORPHOLOGIC ABNORMALITY)|[X]OTHER EMPHYSEMA (MORPHOLOGIC ABNORMALITY)
C0029607|T047|196230005|SNOMEDCT_US|OTHER EMPHYSEMA NOS|[X]OTHER EMPHYSEMA (MORPHOLOGIC ABNORMALITY)
C0029607|T047|196230005|SNOMEDCT_US|[X]OTHER EMPHYSEMA|[X]OTHER EMPHYSEMA (MORPHOLOGIC ABNORMALITY)
C0029607|T047|196230005|SNOMEDCT_US|[X]OTHER EMPHYSEMA (MORPHOLOGIC ABNORMALITY)|[X]OTHER EMPHYSEMA (MORPHOLOGIC ABNORMALITY)
C0029607|T047|196230005|SNOMEDCT_US|OTHER EMPHYSEMA NOS (MORPHOLOGIC ABNORMALITY)|[X]OTHER EMPHYSEMA (MORPHOLOGIC ABNORMALITY)
C0849659|T047||SNOMEDCT_US|CHRONIC AIRWAYS LIMITATION
C0348817|T047|196002001|SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMONARY DISEASE WITH ACUTE EXACERBATION, UNSPECIFIED|CHRONIC OBSTRUCTIVE PULMONARY DISEASE WITH ACUTE EXACERBATION, UNSPECIFIED (DISORDER)
C0348817|T047|196002001|SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMONARY DISEASE WITH ACUTE EXACERBATION, UNSPECIFIED |CHRONIC OBSTRUCTIVE PULMONARY DISEASE WITH ACUTE EXACERBATION, UNSPECIFIED (DISORDER)
C0221227|T047|68328006|SNOMEDCT_US|CENTRILOBULAR EMPHYSEMA|CENTRIACINAR EMPHYSEMA (DISORDER)
C0221227|T047|68328006|SNOMEDCT_US|CENTRIACINAR EMPHYSEMA |CENTRIACINAR EMPHYSEMA (DISORDER)
C0221227|T047|68328006|SNOMEDCT_US|CENTRIACINAR EMPHYSEMA|CENTRIACINAR EMPHYSEMA (DISORDER)
C0221227|T047|68328006|SNOMEDCT_US|EMPHYSEMA, CENTRILOBULAR|CENTRIACINAR EMPHYSEMA (DISORDER)
C0221227|T047|68328006|SNOMEDCT_US|EMPHYSEMAS, CENTRIACINAR|CENTRIACINAR EMPHYSEMA (DISORDER)
C0221227|T047|68328006|SNOMEDCT_US|CENTRIACINAR EMPHYSEMAS|CENTRIACINAR EMPHYSEMA (DISORDER)
C0221227|T047|68328006|SNOMEDCT_US|EMPHYSEMA, CENTRIACINAR|CENTRIACINAR EMPHYSEMA (DISORDER)
C0221227|T047|68328006|SNOMEDCT_US|CENTRILOBULAR EMPHYSEMAS|CENTRIACINAR EMPHYSEMA (DISORDER)
C0221227|T047|68328006|SNOMEDCT_US|EMPHYSEMAS, CENTRILOBULAR|CENTRIACINAR EMPHYSEMA (DISORDER)
C0221227|T047|68328006|SNOMEDCT_US|CENTRIACINAR EMPHYSEMA |CENTRIACINAR EMPHYSEMA (DISORDER)
C0221227|T047|68328006|SNOMEDCT_US|CENTRILOBULAR; EMPHYSEMA|CENTRIACINAR EMPHYSEMA (DISORDER)
C0221227|T047|68328006|SNOMEDCT_US|EMPHYSEMA; CENTRILOBULAR|CENTRIACINAR EMPHYSEMA (DISORDER)
C0221227|T047|68328006|SNOMEDCT_US|LUNG OR PULMONARY EMPHYSEMA, CENTRIACINAR|CENTRIACINAR EMPHYSEMA (DISORDER)
C0221227|T047|68328006|SNOMEDCT_US|LUNG OR PULMONARY EMPHYSEMA, CENTRILOBULAR|CENTRIACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|PANLOBULAR EMPHYSEMA|PANACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|PANACINAR EMPHYSEMA|PANACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|PANACINAR EMPHYSEMA |PANACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|PANLOBULAR EMPHYSEMAS|PANACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|PANACINAR EMPHYSEMAS|PANACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|EMPHYSEMAS, PANLOBULAR|PANACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|EMPHYSEMA, PANACINAR|PANACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|EMPHYSEMAS, PANACINAR|PANACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|EMPHYSEMA, PANLOBULAR|PANACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|ALVEOLAR EMPHYSEMA OF LUNG|PANACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|VESICULAR EMPHYSEMA|PANACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|PANACINAR EMPHYSEMA |PANACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|EMPHYSEMA; PANACINAR|PANACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|EMPHYSEMA; PANLOBULAR|PANACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|EMPHYSEMA; VESICULAR|PANACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|PANACINAR; EMPHYSEMA|PANACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|PANLOBULAR; EMPHYSEMA|PANACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|VESICULAR; EMPHYSEMA|PANACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|EMPHYSEMA, VESICULAR|PANACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|LUNG OR PULMONARY EMPHYSEMA, PANACINAR|PANACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|LUNG OR PULMONARY EMPHYSEMA, PANLOBULAR|PANACINAR EMPHYSEMA (DISORDER)
C0264393|T047|4981000|SNOMEDCT_US|LUNG OR PULMONARY EMPHYSEMA, VESICULAR|PANACINAR EMPHYSEMA (DISORDER)
C1277261|T047|135836000|SNOMEDCT_US|END STAGE CHRONIC OBSTRUCTIVE PULMONARY DISEASE|END STAGE CHRONIC OBSTRUCTIVE AIRWAYS DISEASE (DISORDER)
C1277261|T047|135836000|SNOMEDCT_US|END STAGE CHRONIC OBSTRUCTIVE PULMONARY DISEASE |END STAGE CHRONIC OBSTRUCTIVE AIRWAYS DISEASE (DISORDER)
C1277261|T047|135836000|SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMONARY DISEASE END STAGE|END STAGE CHRONIC OBSTRUCTIVE AIRWAYS DISEASE (DISORDER)
C1277261|T047|135836000|SNOMEDCT_US|END STAGE CHRONIC OBSTRUCTIVE AIRWAYS DISEASE |END STAGE CHRONIC OBSTRUCTIVE AIRWAYS DISEASE (DISORDER)
C1277261|T047|135836000|SNOMEDCT_US|END STAGE CHRONIC OBSTRUCTIVE AIRWAYS DISEASE|END STAGE CHRONIC OBSTRUCTIVE AIRWAYS DISEASE (DISORDER)
C1969833|T047||SNOMEDCT_US|COPD, SEVERE EARLY-ONSET
C4040148|T047|106001000119101|SNOMEDCT_US|CHRONIC OBSTRUCTIVE LUNG DISEASE CO-OCCURRENT WITH ACUTE BRONCHITIS |CHRONIC OBSTRUCTIVE LUNG DISEASE CO-OCCURRENT WITH ACUTE BRONCHITIS (DISORDER)
C4040148|T047|106001000119101|SNOMEDCT_US|CHRONIC OBSTRUCTIVE LUNG DISEASE CO-OCCURRENT WITH ACUTE BRONCHITIS|CHRONIC OBSTRUCTIVE LUNG DISEASE CO-OCCURRENT WITH ACUTE BRONCHITIS (DISORDER)
C0340044|T047|195951007|SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMONARY DISEASE WITH (ACUTE) EXACERBATION|ACUTE EXACERBATION OF CHRONIC OBSTRUCTIVE PULMONARY DISEASE
C0340044|T047|195951007|SNOMEDCT_US|CHRONIC OBSTRUCTIVE PULMONARY DISEASE W (ACUTE) EXACERBATION|ACUTE EXACERBATION OF CHRONIC OBSTRUCTIVE PULMONARY DISEASE
C0340044|T047|195951007|SNOMEDCT_US|ACUTE EXACERBATION OF CHRONIC OBSTRUCTIVE AIRWAYS DISEASE |ACUTE EXACERBATION OF CHRONIC OBSTRUCTIVE PULMONARY DISEASE
C0340044|T047|195951007|SNOMEDCT_US|ACUTE EXACERBATION OF CHRONIC OBSTRUCTIVE AIRWAYS DISEASE|ACUTE EXACERBATION OF CHRONIC OBSTRUCTIVE PULMONARY DISEASE
C0340044|T047|195951007|SNOMEDCT_US|ACUTE EXACERBATION OF COPD|ACUTE EXACERBATION OF CHRONIC OBSTRUCTIVE PULMONARY DISEASE
C0340044|T047|195951007|SNOMEDCT_US|ACUTE EXACERBATION OF CHRONIC OBSTRUCTIVE PULMONARY DISEASE|ACUTE EXACERBATION OF CHRONIC OBSTRUCTIVE PULMONARY DISEASE
C1385064|T047||SNOMEDCT_US|DISEASE (OR DISORDER); LUNG, OBSTRUCTIVE (CHRONIC)
C0155883|T047||SNOMEDCT_US|CHRONIC OBSTRUCTIVE ASTHMA
C0155883|T047||SNOMEDCT_US|CHRONIC OBSTRUCTIVE ASTHMA 
C0155883|T047||SNOMEDCT_US|CHRONIC OBSTRUCTIVE ASTHMA (WITH OBSTRUCTIVE PULMONARY DISEASE)
