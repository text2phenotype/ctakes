C0010076|T005|DE|0000016152|AOD|Coronaviridae|Coronaviridae
C0010076|T005|PT|3108-0765|CSP|Coronaviridae|Coronaviridae
C0010076|T005|MH|D003332|MSH|Coronaviridae|Coronaviridae
C0010076|T005|PT|X73lD|RCD|Coronaviridae|Coronaviridae
C0010076|T005|PT|C113205|NCI|Coronaviridae|Coronaviridae
C0010076|T005|SY|243607003|SNOMEDCT_US|Coronaviridae|Coronaviridae
C0010076|T005|PN|U001830|MTH|Coronaviridae|Coronaviridae
C0010076|T005|PT|0000003373|CHV|coronaviridae|coronaviridae
C0010076|T005|PT|C113205|NCI_CDISC|CORONAVIRIDAE|CORONAVIRIDAE
C0010076|T005|OF|243607003|SNOMEDCT_US|Coronaviridae (organism)|Coronaviridae (organism)
C0010076|T005|IS|88711001|SNOMEDCT_US|Coronavirus group|Coronavirus group
C0010076|T005|SY|243607003|SNOMEDCT_US|Coronavirus group|Coronavirus group
C0010076|T005|IS|88711001|SNOMEDCT_US|Coronavirus group, NOS|Coronavirus group, NOS
C0010076|T005|PT|243607003|SNOMEDCT_US|Family Coronaviridae|Family Coronaviridae
C0010076|T005|FN|243607003|SNOMEDCT_US|Family Coronaviridae (organism)|Family Coronaviridae (organism)
C0010076|T005|IS|243607003|SNOMEDCT_US|Family: Coronavirus group|Family: Coronavirus group
C0010076|T005|SY|X73lD|RCD|Family: Coronavirus group|Family: Coronavirus group
C0010077|T116|PEP|D014759|MSH|Coronavirus gpE1|Coronavirus gpE1
C0010077|T123|PEP|D014759|MSH|Coronavirus gpE1|Coronavirus gpE1
C0010079|T116|PEP|D014759|MSH|Coronavirus Peplomer Protein E1|Coronavirus Peplomer Protein E1
C0010079|T123|PEP|D014759|MSH|Coronavirus Peplomer Protein E1|Coronavirus Peplomer Protein E1
C0010080|T116|PEP|D014759|MSH|Coronavirus Peplomer Protein E2 JHM|Coronavirus Peplomer Protein E2 JHM
C0010080|T123|PEP|D014759|MSH|Coronavirus Peplomer Protein E2 JHM|Coronavirus Peplomer Protein E2 JHM
C0014338|T005|OAS|51225001|SNOMEDCT_US|Bluecomb disease virus|Bluecomb disease virus
C0014338|T005|SY|422912001|SNOMEDCT_US|Bluecomb disease virus|Bluecomb disease virus
C0014338|T005|ET|D004752|MSH|Bluecomb Virus|Bluecomb Virus
C0014338|T005|PM|D004752|MSH|Bluecomb Viruses|Bluecomb Viruses
C0014338|T005|MH|D004752|MSH|Coronavirus, Turkey|Coronavirus, Turkey
C0014338|T005|PM|D004752|MSH|Coronaviruses, Turkey|Coronaviruses, Turkey
C0014338|T005|OAP|51225001|SNOMEDCT_US|Enteritis of turkeys coronavirus|Enteritis of turkeys coronavirus
C0014338|T005|SY|422912001|SNOMEDCT_US|Enteritis of turkeys coronavirus|Enteritis of turkeys coronavirus
C0014338|T005|OAF|51225001|SNOMEDCT_US|Enteritis of turkeys coronavirus (organism)|Enteritis of turkeys coronavirus (organism)
C0014338|T005|ET|D004752|MSH|Enteritis Virus, Turkey|Enteritis Virus, Turkey
C0014338|T005|PM|D004752|MSH|Enteritis Viruses, Turkey|Enteritis Viruses, Turkey
C0014338|T005|DEV|D004752|MSH|TRANSM ENTERITIS VIRUS OF TURKEYS|TRANSM ENTERITIS VIRUS OF TURKEYS
C0014338|T005|DEV|D004752|MSH|TRANSM ENTERITIS VIRUS TURKEYS|TRANSM ENTERITIS VIRUS TURKEYS
C0014338|T005|ET|D004752|MSH|Transmissible Enteritis Virus of Turkeys|Transmissible Enteritis Virus of Turkeys
C0014338|T005|ET|D004752|MSH|Transmissible Enteritis Virus, Turkeys|Transmissible Enteritis Virus, Turkeys
C0014338|T005|OAS|51225001|SNOMEDCT_US|Turkey coronavirus|Turkey coronavirus
C0014338|T005|PT|422912001|SNOMEDCT_US|Turkey coronavirus|Turkey coronavirus
C0014338|T005|ET|D004752|MSH|Turkey Coronavirus|Turkey Coronavirus
C0014338|T005|FN|422912001|SNOMEDCT_US|Turkey coronavirus (organism)|Turkey coronavirus (organism)
C0014338|T005|PM|D004752|MSH|Turkey Coronaviruses|Turkey Coronaviruses
C0014338|T005|LPN|LP19955-1|LNC|Turkey enteritis coronavirus|Turkey enteritis coronavirus
C0014338|T005|CN|MTHU011313|LNC|Turkey enteritis coronavirus|Turkey enteritis coronavirus
C0014338|T005|PM|D004752|MSH|Turkey Enteritis Virus|Turkey Enteritis Virus
C0014338|T005|PM|D004752|MSH|Turkey Enteritis Viruses|Turkey Enteritis Viruses
C0017161|T005|SY|80073003|SNOMEDCT_US|Coronavirus 777|Coronavirus 777
C0017161|T005|DEV|D005760|MSH|GASTEROENTERITIS VIRUS PORCINE TRANSM|GASTEROENTERITIS VIRUS PORCINE TRANSM
C0017161|T005|ET|D005760|MSH|Gastroenteritis Virus of Swine|Gastroenteritis Virus of Swine
C0017161|T005|ET|D005760|MSH|Gastroenteritis Virus, Porcine Transmissible|Gastroenteritis Virus, Porcine Transmissible
C0017161|T005|DEV|D005760|MSH|PORCINE TRANSM GASTROENTERITIS VIRUS|PORCINE TRANSM GASTROENTERITIS VIRUS
C0017161|T005|PT|80073003|SNOMEDCT_US|Porcine transmissible gastroenteritis virus|Porcine transmissible gastroenteritis virus
C0017161|T005|ET|D005760|MSH|Porcine Transmissible Gastroenteritis Virus|Porcine Transmissible Gastroenteritis Virus
C0017161|T005|ET|3108-0765|CSP|porcine transmissible gastroenteritis virus|porcine transmissible gastroenteritis virus
C0017161|T005|FN|80073003|SNOMEDCT_US|Porcine transmissible gastroenteritis virus (organism)|Porcine transmissible gastroenteritis virus (organism)
C0017161|T005|PM|D005760|MSH|Swine Gastroenteritis Virus|Swine Gastroenteritis Virus
C0017161|T005|PM|D005760|MSH|Swine Gastroenteritis Viruses|Swine Gastroenteritis Viruses
C0017161|T005|ET|D005760|MSH|TGE Virus|TGE Virus
C0017161|T005|PM|D005760|MSH|TGE Viruses|TGE Viruses
C0017161|T005|DEV|D005760|MSH|TRANSM GASTROENTERITIS VIRUS|TRANSM GASTROENTERITIS VIRUS
C0017161|T005|DEV|D005760|MSH|TRANSM GASTROENTERITIS VIRUS SWINE|TRANSM GASTROENTERITIS VIRUS SWINE
C0017161|T005|LPN|LP19950-2|LNC|Transmissible gastroenteritis virus|Transmissible gastroenteritis virus
C0017161|T005|MH|D005760|MSH|Transmissible gastroenteritis virus|Transmissible gastroenteritis virus
C0017161|T005|SY|80073003|SNOMEDCT_US|Transmissible gastroenteritis virus|Transmissible gastroenteritis virus
C0017161|T005|ET|D005760|MSH|Transmissible Gastroenteritis Virus, Swine|Transmissible Gastroenteritis Virus, Swine
C0019185|T005|ET|D006517|MSH|Gastroenteritis Virus, Murine|Gastroenteritis Virus, Murine
C0019185|T005|PM|D006517|MSH|Gastroenteritis Viruses, Murine|Gastroenteritis Viruses, Murine
C0019185|T005|ET|D006517|MSH|Hepatitis Virus, Mouse|Hepatitis Virus, Mouse
C0019185|T005|PM|D006517|MSH|Hepatitis Viruses, Mouse|Hepatitis Viruses, Mouse
C0019185|T005|DE|0000016153|AOD|mouse hepatitis virus|mouse hepatitis virus
C0019185|T005|ET|3108-0815|CSP|mouse hepatitis virus|mouse hepatitis virus
C0019185|T005|ET|D006517|MSH|Mouse Hepatitis Virus|Mouse Hepatitis Virus
C0019185|T005|PM|D006517|MSH|Mouse Hepatitis Viruses|Mouse Hepatitis Viruses
C0019185|T005|ET|D006517|MSH|Murine coronavirus|Murine coronavirus
C0019185|T005|PT|697943002|SNOMEDCT_US|Murine coronavirus|Murine coronavirus
C0019185|T005|FN|697943002|SNOMEDCT_US|Murine coronavirus (organism)|Murine coronavirus (organism)
C0019185|T005|PM|D006517|MSH|Murine coronaviruses|Murine coronaviruses
C0019185|T005|ET|D006517|MSH|Murine Gastroenteritis Virus|Murine Gastroenteritis Virus
C0019185|T005|PM|D006517|MSH|Murine Gastroenteritis Viruses|Murine Gastroenteritis Viruses
C0019185|T005|MH|D006517|MSH|Murine hepatitis virus|Murine hepatitis virus
C0019185|T005|PT|80129000|SNOMEDCT_US|Murine hepatitis virus|Murine hepatitis virus
C0019185|T005|PT|3108-0815|CSP|murine hepatitis virus|murine hepatitis virus
C0019185|T005|FN|80129000|SNOMEDCT_US|Murine hepatitis virus (organism)|Murine hepatitis virus (organism)
C0019185|T005|PM|D006517|MSH|Murine hepatitis viruses|Murine hepatitis viruses
C0027610|T005|LPN|LP19603-7|LNC|Bovine coronavirus|Bovine coronavirus
C0027610|T005|PT|407372004|SNOMEDCT_US|Bovine coronavirus|Bovine coronavirus
C0027610|T005|PN|NOCODE|MTH|Bovine coronavirus|Bovine coronavirus
C0027610|T005|ET|D017938|MSH|Bovine Coronavirus|Bovine Coronavirus
C0027610|T005|ET|3108-0765|CSP|bovine coronavirus|bovine coronavirus
C0027610|T005|FN|407372004|SNOMEDCT_US|Bovine coronavirus (organism)|Bovine coronavirus (organism)
C0027610|T005|PM|D017938|MSH|Bovine Coronaviruses|Bovine Coronaviruses
C0027610|T005|MH|D017938|MSH|Coronavirus, Bovine|Coronavirus, Bovine
C0027610|T005|PM|D017938|MSH|Coronaviruses, Bovine|Coronaviruses, Bovine
C0126544|T116|CE|C067997|MSH|M protein, BECV F15|M protein, BECV F15
C0126544|T116|PCE|C067997|MSH|M protein, Bovine enteric coronavirus F15|M protein, Bovine enteric coronavirus F15
C0126544|T116|CE|C067997|MSH|matrix protein, BECV F15|matrix protein, BECV F15
C0174990|T116|NM|C078034|MSH|coronavirus receptor|coronavirus receptor
C0174990|T192|NM|C078034|MSH|coronavirus receptor|coronavirus receptor
C0174990|T116|CE|C078034|MSH|coronavirus receptors|coronavirus receptors
C0174990|T192|CE|C078034|MSH|coronavirus receptors|coronavirus receptors
C0174990|T116|CE|C078034|MSH|receptor, coronavirus|receptor, coronavirus
C0174990|T192|CE|C078034|MSH|receptor, coronavirus|receptor, coronavirus
C0199848|T061|PT|90640007|SNOMEDCT_US|Coronavirus vaccination|Coronavirus vaccination
C0199848|T061|FN|90640007|SNOMEDCT_US|Coronavirus vaccination (procedure)|Coronavirus vaccination (procedure)
C0206419|T005|ET|3108-0765|CSP|Coronavirus|Coronavirus
C0206419|T005|PT|X73lE|RCD|Coronavirus|Coronavirus
C0206419|T005|LPN|LP16680-8|LNC|Coronavirus|Coronavirus
C0206419|T005|OAP|88711001|SNOMEDCT_US|Coronavirus|Coronavirus
C0206419|T005|OAP|243608008|SNOMEDCT_US|Coronavirus|Coronavirus
C0206419|T005|PT|C26431|NCI|Coronavirus|Coronavirus
C0206419|T005|MH|D017934|MSH|Coronavirus|Coronavirus
C0206419|T005|PT|0000020927|CHV|coronavirus|coronavirus
C0206419|T005|OAF|88711001|SNOMEDCT_US|Coronavirus (living organism) (organism)|Coronavirus (living organism) (organism)
C0206419|T005|OF|88711001|SNOMEDCT_US|Coronavirus (living organism) [Ambiguous]|Coronavirus (living organism) [Ambiguous]
C0206419|T005|OF|243608008|SNOMEDCT_US|Coronavirus (organism)|Coronavirus (organism)
C0206419|T005|IS|88711001|SNOMEDCT_US|Coronavirus, NOS|Coronavirus, NOS
C0206419|T005|PT|U005409|LCH|Coronaviruses|Coronaviruses
C0206419|T005|PM|D017934|MSH|Coronaviruses|Coronaviruses
C0206419|T005|PT|sh85032882|LCH_NW|Coronaviruses|Coronaviruses
C0206419|T005|SY|0000020927|CHV|coronaviruses|coronaviruses
C0206419|T005|OAS|243608008|SNOMEDCT_US|Genus Coronavirus|Genus Coronavirus
C0206419|T005|OAF|243608008|SNOMEDCT_US|Genus Coronavirus (organism)|Genus Coronavirus (organism)
C0206419|T005|SY|X73lE|RCD|Genus: Coronavirus|Genus: Coronavirus
C0206419|T005|OAS|243608008|SNOMEDCT_US|Genus: Coronavirus|Genus: Coronavirus
C0206419|T005|PN|U002406|MTH|Genus: Coronavirus|Genus: Coronavirus
C0206421|T005|LPN|LP14096-9|LNC|Canine coronavirus|Canine coronavirus
C0206421|T005|PT|16365004|SNOMEDCT_US|Canine coronavirus|Canine coronavirus
C0206421|T005|ET|D017939|MSH|Canine Coronavirus|Canine Coronavirus
C0206421|T005|ET|3108-0765|CSP|canine coronavirus|canine coronavirus
C0206421|T005|FN|16365004|SNOMEDCT_US|Canine coronavirus (organism)|Canine coronavirus (organism)
C0206421|T005|PM|D017939|MSH|Canine Coronaviruses|Canine Coronaviruses
C0206421|T005|ET|D017939|MSH|Canine respiratory coronavirus|Canine respiratory coronavirus
C0206421|T005|PM|D017939|MSH|Canine respiratory coronaviruses|Canine respiratory coronaviruses
C0206421|T005|MH|D017939|MSH|Coronavirus, Canine|Coronavirus, Canine
C0206421|T005|PM|D017939|MSH|Coronaviruses, Canine|Coronaviruses, Canine
C0206422|T005|SY|0000020928|CHV|coronavirus human|coronavirus human
C0206422|T005|AB|X73lF|RCD|Enveloped ssRNA no DNA: 1 neg|Enveloped ssRNA no DNA: 1 neg
C0206422|T005|AB|X73lF|RCD|Enveloped ssRNA virus no DNA step with one neg-sense genome|Enveloped ssRNA virus no DNA step with one neg-sense genome
C0206422|T005|IS|84101006|SNOMEDCT_US|Enveloped ssRNA virus without a DNA step with single-stranded negative-sense genome|Enveloped ssRNA virus without a DNA step with single-stranded negative-sense genome
C0206422|T005|SY|X73lF|RCD|Enveloped ssRNA virus without a DNA step with single-stranded negative-sense genome|Enveloped ssRNA virus without a DNA step with single-stranded negative-sense genome
C0206422|T005|IS|84101006|SNOMEDCT_US|Enveloped ssRNA virus without a DNA step with single-stranded negative-sense genome (organism)|Enveloped ssRNA virus without a DNA step with single-stranded negative-sense genome (organism)
C0206422|T005|SY|X73lF|RCD|HCV - Human coronavirus|HCV - Human coronavirus
C0206422|T005|SY|84101006|SNOMEDCT_US|HCV - Human coronavirus|HCV - Human coronavirus
C0206422|T005|PT|X73lF|RCD|Human coronavirus|Human coronavirus
C0206422|T005|LPN|LP35707-6|LNC|Human coronavirus|Human coronavirus
C0206422|T005|LG|LG32771-4|LNC|Human coronavirus|Human coronavirus
C0206422|T005|PT|84101006|SNOMEDCT_US|Human coronavirus|Human coronavirus
C0206422|T005|ET|3108-0765|CSP|human coronavirus|human coronavirus
C0206422|T005|PT|0000020928|CHV|human coronavirus|human coronavirus
C0206422|T005|FN|84101006|SNOMEDCT_US|Human coronavirus (organism)|Human coronavirus (organism)
C0206423|T005|MH|D017941|MSH|Coronavirus, Rat|Coronavirus, Rat
C0206423|T005|PT|12231001|SNOMEDCT_US|Rat coronavirus|Rat coronavirus
C0206423|T005|ET|D017941|MSH|Rat Coronavirus|Rat Coronavirus
C0206423|T005|FN|12231001|SNOMEDCT_US|Rat coronavirus (organism)|Rat coronavirus (organism)
C0206750|T047|OAP|187467005|SNOMEDCT_US|[X]Coronavirus infection, unspecified|[X]Coronavirus infection, unspecified
C0206750|T047|OP|AyuDC|RCD|[X]Coronavirus infection, unspecified|[X]Coronavirus infection, unspecified
C0206750|T047|OAF|187467005|SNOMEDCT_US|[X]Coronavirus infection, unspecified (disorder)|[X]Coronavirus infection, unspecified (disorder)
C0206750|T047|OA|AyuDC|RCD|[X]Coronavirus infection,unspc|[X]Coronavirus infection,unspc
C0206750|T047|SY|0000021065|CHV|corona infection virus|corona infection virus
C0206750|T047|SY|0000021065|CHV|corona infections virus|corona infections virus
C0206750|T047|LLT|10053983|MDR|Corona virus infection|Corona virus infection
C0206750|T047|PT|10053983|MDR|Corona virus infection|Corona virus infection
C0206750|T047|SY|318393|MEDCIN|coronavirus|coronavirus
C0206750|T047|DEV|D018352|MSH|CORONAVIRUS INFECT|CORONAVIRUS INFECT
C0206750|T047|PM|D018352|MSH|Coronavirus Infection|Coronavirus Infection
C0206750|T047|PT|A795.|RCD|Coronavirus infection|Coronavirus infection
C0206750|T047|PT|318393|MEDCIN|Coronavirus infection|Coronavirus infection
C0206750|T047|LLT|10051905|MDR|Coronavirus infection|Coronavirus infection
C0206750|T047|PT|186747009|SNOMEDCT_US|Coronavirus infection|Coronavirus infection
C0206750|T047|PT|0000021065|CHV|coronavirus infection|coronavirus infection
C0206750|T047|FN|318393|MEDCIN|Coronavirus infection (diagnosis)|Coronavirus infection (diagnosis)
C0206750|T047|FN|186747009|SNOMEDCT_US|Coronavirus infection (disorder)|Coronavirus infection (disorder)
C0206750|T047|OP|AyuDC|RCDSY|Coronavirus infection, unspecified|Coronavirus infection, unspecified
C0206750|T047|PT|B34.2|ICD10CM|Coronavirus infection, unspecified|Coronavirus infection, unspecified
C0206750|T047|AB|B34.2|ICD10CM|Coronavirus infection, unspecified|Coronavirus infection, unspecified
C0206750|T047|PT|B34.2|ICD10|Coronavirus infection, unspecified|Coronavirus infection, unspecified
C0206750|T047|OA|AyuDC|RCDSY|Coronavirus infection,unspc|Coronavirus infection,unspc
C0206750|T047|MH|D018352|MSH|Coronavirus Infections|Coronavirus Infections
C0206750|T047|PN|NOCODE|MTH|Coronavirus Infections|Coronavirus Infections
C0206750|T047|PT|sh90004313|LCH_NW|Coronavirus infections|Coronavirus infections
C0206750|T047|DEV|D018352|MSH|INFECT CORONAVIRUS|INFECT CORONAVIRUS
C0206750|T047|PM|D018352|MSH|Infection, Coronavirus|Infection, Coronavirus
C0206750|T047|PT|MTHU038700|ICPC2ICD10ENG|infection; viral, coronavirus|infection; viral, coronavirus
C0206750|T047|ET|D018352|MSH|Infections, Coronavirus|Infections, Coronavirus
C0246449|T116|NM|C067997|MSH|M protein, Coronavirus|M protein, Coronavirus
C0255554|T116|CE|C087632|MSH|6b protein, coronavirus|6b protein, coronavirus
C0255554|T116|NM|C087632|MSH|glycoprotein 6b, coronavirus|glycoprotein 6b, coronavirus
C0255556|T116|PCE|C087633|MSH|NS2 protein, bovine coronavirus (BCV)|NS2 protein, bovine coronavirus (BCV)
C0255557|T116|PCE|C087633|MSH|NS2 protein, human coronavirus (HCV)|NS2 protein, human coronavirus (HCV)
C0255558|T116|NM|C087633|MSH|nonstructural protein, coronavirus|nonstructural protein, coronavirus
C0255558|T116|CE|C087633|MSH|NS protein, coronavirus|NS protein, coronavirus
C0255568|T116|PCE|C087637|MSH|gene 1 protein, Human coronavirus (HCV)|gene 1 protein, Human coronavirus (HCV)
C0255568|T123|PCE|C087637|MSH|gene 1 protein, Human coronavirus (HCV)|gene 1 protein, Human coronavirus (HCV)
C0255573|T116|NM|C087637|MSH|gene 1 protein, Coronavirus|gene 1 protein, Coronavirus
C0255573|T123|NM|C087637|MSH|gene 1 protein, Coronavirus|gene 1 protein, Coronavirus
C0310685|T116|OAP|78742002|SNOMEDCT_US|Bovine rota - coronavirus vaccine|Bovine rota - coronavirus vaccine
C0310685|T121|OAP|78742002|SNOMEDCT_US|Bovine rota - coronavirus vaccine|Bovine rota - coronavirus vaccine
C0310685|T129|OAP|78742002|SNOMEDCT_US|Bovine rota - coronavirus vaccine|Bovine rota - coronavirus vaccine
C0310685|T116|OAF|78742002|SNOMEDCT_US|Bovine rota - coronavirus vaccine (product)|Bovine rota - coronavirus vaccine (product)
C0310685|T121|OAF|78742002|SNOMEDCT_US|Bovine rota - coronavirus vaccine (product)|Bovine rota - coronavirus vaccine (product)
C0310685|T129|OAF|78742002|SNOMEDCT_US|Bovine rota - coronavirus vaccine (product)|Bovine rota - coronavirus vaccine (product)
C0310685|T116|OF|78742002|SNOMEDCT_US|Bovine rota - coronavirus vaccine (substance)|Bovine rota - coronavirus vaccine (substance)
C0310685|T121|OF|78742002|SNOMEDCT_US|Bovine rota - coronavirus vaccine (substance)|Bovine rota - coronavirus vaccine (substance)
C0310685|T129|OF|78742002|SNOMEDCT_US|Bovine rota - coronavirus vaccine (substance)|Bovine rota - coronavirus vaccine (substance)
C0310701|T116|OAP|72390003|SNOMEDCT_US|Canine coronavirus vaccine|Canine coronavirus vaccine
C0310701|T121|OAP|72390003|SNOMEDCT_US|Canine coronavirus vaccine|Canine coronavirus vaccine
C0310701|T129|OAP|72390003|SNOMEDCT_US|Canine coronavirus vaccine|Canine coronavirus vaccine
C0310701|T116|OAP|449238002|SNOMEDCT_US|Canine coronavirus vaccine|Canine coronavirus vaccine
C0310701|T121|OAP|449238002|SNOMEDCT_US|Canine coronavirus vaccine|Canine coronavirus vaccine
C0310701|T129|OAP|449238002|SNOMEDCT_US|Canine coronavirus vaccine|Canine coronavirus vaccine
C0310701|T116|OAF|72390003|SNOMEDCT_US|Canine coronavirus vaccine (product)|Canine coronavirus vaccine (product)
C0310701|T121|OAF|72390003|SNOMEDCT_US|Canine coronavirus vaccine (product)|Canine coronavirus vaccine (product)
C0310701|T129|OAF|72390003|SNOMEDCT_US|Canine coronavirus vaccine (product)|Canine coronavirus vaccine (product)
C0310701|T116|OF|72390003|SNOMEDCT_US|Canine coronavirus vaccine (substance)|Canine coronavirus vaccine (substance)
C0310701|T121|OF|72390003|SNOMEDCT_US|Canine coronavirus vaccine (substance)|Canine coronavirus vaccine (substance)
C0310701|T129|OF|72390003|SNOMEDCT_US|Canine coronavirus vaccine (substance)|Canine coronavirus vaccine (substance)
C0310701|T116|OAF|449238002|SNOMEDCT_US|Canine coronavirus vaccine (substance)|Canine coronavirus vaccine (substance)
C0310701|T121|OAF|449238002|SNOMEDCT_US|Canine coronavirus vaccine (substance)|Canine coronavirus vaccine (substance)
C0310701|T129|OAF|449238002|SNOMEDCT_US|Canine coronavirus vaccine (substance)|Canine coronavirus vaccine (substance)
C0310702|T116|OAP|61898000|SNOMEDCT_US|Canine coronavirus - parvovirus vaccine|Canine coronavirus - parvovirus vaccine
C0310702|T121|OAP|61898000|SNOMEDCT_US|Canine coronavirus - parvovirus vaccine|Canine coronavirus - parvovirus vaccine
C0310702|T129|OAP|61898000|SNOMEDCT_US|Canine coronavirus - parvovirus vaccine|Canine coronavirus - parvovirus vaccine
C0310702|T116|OAF|61898000|SNOMEDCT_US|Canine coronavirus - parvovirus vaccine (product)|Canine coronavirus - parvovirus vaccine (product)
C0310702|T121|OAF|61898000|SNOMEDCT_US|Canine coronavirus - parvovirus vaccine (product)|Canine coronavirus - parvovirus vaccine (product)
C0310702|T129|OAF|61898000|SNOMEDCT_US|Canine coronavirus - parvovirus vaccine (product)|Canine coronavirus - parvovirus vaccine (product)
C0310702|T116|OF|61898000|SNOMEDCT_US|Canine coronavirus - parvovirus vaccine (substance)|Canine coronavirus - parvovirus vaccine (substance)
C0310702|T121|OF|61898000|SNOMEDCT_US|Canine coronavirus - parvovirus vaccine (substance)|Canine coronavirus - parvovirus vaccine (substance)
C0310702|T129|OF|61898000|SNOMEDCT_US|Canine coronavirus - parvovirus vaccine (substance)|Canine coronavirus - parvovirus vaccine (substance)
C0310705|T116|OAP|44765006|SNOMEDCT_US|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine
C0310705|T121|OAP|44765006|SNOMEDCT_US|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine
C0310705|T129|OAP|44765006|SNOMEDCT_US|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine
C0310705|T116|OAF|44765006|SNOMEDCT_US|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine (product)|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine (product)
C0310705|T121|OAF|44765006|SNOMEDCT_US|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine (product)|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine (product)
C0310705|T129|OAF|44765006|SNOMEDCT_US|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine (product)|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine (product)
C0310705|T116|OF|44765006|SNOMEDCT_US|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine (substance)|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine (substance)
C0310705|T121|OF|44765006|SNOMEDCT_US|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine (substance)|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine (substance)
C0310705|T129|OF|44765006|SNOMEDCT_US|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine (substance)|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine (substance)
C0310907|T116|OAP|14254009|SNOMEDCT_US|Bovine rota - coronavirus vaccine - clostridium perfringens type C - escherichia coli bacterin - toxoid|Bovine rota - coronavirus vaccine - clostridium perfringens type C - escherichia coli bacterin - toxoid
C0310907|T121|OAP|14254009|SNOMEDCT_US|Bovine rota - coronavirus vaccine - clostridium perfringens type C - escherichia coli bacterin - toxoid|Bovine rota - coronavirus vaccine - clostridium perfringens type C - escherichia coli bacterin - toxoid
C0310907|T129|OAP|14254009|SNOMEDCT_US|Bovine rota - coronavirus vaccine - clostridium perfringens type C - escherichia coli bacterin - toxoid|Bovine rota - coronavirus vaccine - clostridium perfringens type C - escherichia coli bacterin - toxoid
C0310907|T116|OAF|14254009|SNOMEDCT_US|Bovine rota - coronavirus vaccine - clostridium perfringens type C - escherichia coli bacterin - toxoid (product)|Bovine rota - coronavirus vaccine - clostridium perfringens type C - escherichia coli bacterin - toxoid (product)
C0310907|T121|OAF|14254009|SNOMEDCT_US|Bovine rota - coronavirus vaccine - clostridium perfringens type C - escherichia coli bacterin - toxoid (product)|Bovine rota - coronavirus vaccine - clostridium perfringens type C - escherichia coli bacterin - toxoid (product)
C0310907|T129|OAF|14254009|SNOMEDCT_US|Bovine rota - coronavirus vaccine - clostridium perfringens type C - escherichia coli bacterin - toxoid (product)|Bovine rota - coronavirus vaccine - clostridium perfringens type C - escherichia coli bacterin - toxoid (product)
C0310907|T116|OF|14254009|SNOMEDCT_US|Bovine rota - coronavirus vaccine - clostridium perfringens type C - escherichia coli bacterin - toxoid (substance)|Bovine rota - coronavirus vaccine - clostridium perfringens type C - escherichia coli bacterin - toxoid (substance)
C0310907|T121|OF|14254009|SNOMEDCT_US|Bovine rota - coronavirus vaccine - clostridium perfringens type C - escherichia coli bacterin - toxoid (substance)|Bovine rota - coronavirus vaccine - clostridium perfringens type C - escherichia coli bacterin - toxoid (substance)
C0310907|T129|OF|14254009|SNOMEDCT_US|Bovine rota - coronavirus vaccine - clostridium perfringens type C - escherichia coli bacterin - toxoid (substance)|Bovine rota - coronavirus vaccine - clostridium perfringens type C - escherichia coli bacterin - toxoid (substance)
C0310908|T116|OAP|9819008|SNOMEDCT_US|Bovine rota - coronavirus vaccine - escherichia coli bacterin|Bovine rota - coronavirus vaccine - escherichia coli bacterin
C0310908|T121|OAP|9819008|SNOMEDCT_US|Bovine rota - coronavirus vaccine - escherichia coli bacterin|Bovine rota - coronavirus vaccine - escherichia coli bacterin
C0310908|T129|OAP|9819008|SNOMEDCT_US|Bovine rota - coronavirus vaccine - escherichia coli bacterin|Bovine rota - coronavirus vaccine - escherichia coli bacterin
C0310908|T116|OAF|9819008|SNOMEDCT_US|Bovine rota - coronavirus vaccine - escherichia coli bacterin (product)|Bovine rota - coronavirus vaccine - escherichia coli bacterin (product)
C0310908|T121|OAF|9819008|SNOMEDCT_US|Bovine rota - coronavirus vaccine - escherichia coli bacterin (product)|Bovine rota - coronavirus vaccine - escherichia coli bacterin (product)
C0310908|T129|OAF|9819008|SNOMEDCT_US|Bovine rota - coronavirus vaccine - escherichia coli bacterin (product)|Bovine rota - coronavirus vaccine - escherichia coli bacterin (product)
C0310908|T116|OF|9819008|SNOMEDCT_US|Bovine rota - coronavirus vaccine - escherichia coli bacterin (substance)|Bovine rota - coronavirus vaccine - escherichia coli bacterin (substance)
C0310908|T121|OF|9819008|SNOMEDCT_US|Bovine rota - coronavirus vaccine - escherichia coli bacterin (substance)|Bovine rota - coronavirus vaccine - escherichia coli bacterin (substance)
C0310908|T129|OF|9819008|SNOMEDCT_US|Bovine rota - coronavirus vaccine - escherichia coli bacterin (substance)|Bovine rota - coronavirus vaccine - escherichia coli bacterin (substance)
C0310914|T116|OAP|67519008|SNOMEDCT_US|Canine coronavirus vaccine - leptospira bacterin|Canine coronavirus vaccine - leptospira bacterin
C0310914|T121|OAP|67519008|SNOMEDCT_US|Canine coronavirus vaccine - leptospira bacterin|Canine coronavirus vaccine - leptospira bacterin
C0310914|T129|OAP|67519008|SNOMEDCT_US|Canine coronavirus vaccine - leptospira bacterin|Canine coronavirus vaccine - leptospira bacterin
C0310914|T116|OAF|67519008|SNOMEDCT_US|Canine coronavirus vaccine - leptospira bacterin (product)|Canine coronavirus vaccine - leptospira bacterin (product)
C0310914|T121|OAF|67519008|SNOMEDCT_US|Canine coronavirus vaccine - leptospira bacterin (product)|Canine coronavirus vaccine - leptospira bacterin (product)
C0310914|T129|OAF|67519008|SNOMEDCT_US|Canine coronavirus vaccine - leptospira bacterin (product)|Canine coronavirus vaccine - leptospira bacterin (product)
C0310914|T116|OF|67519008|SNOMEDCT_US|Canine coronavirus vaccine - leptospira bacterin (substance)|Canine coronavirus vaccine - leptospira bacterin (substance)
C0310914|T121|OF|67519008|SNOMEDCT_US|Canine coronavirus vaccine - leptospira bacterin (substance)|Canine coronavirus vaccine - leptospira bacterin (substance)
C0310914|T129|OF|67519008|SNOMEDCT_US|Canine coronavirus vaccine - leptospira bacterin (substance)|Canine coronavirus vaccine - leptospira bacterin (substance)
C0310915|T116|OAP|9079002|SNOMEDCT_US|Canine coronavirus - parvovirus vaccine - leptospira bacterin|Canine coronavirus - parvovirus vaccine - leptospira bacterin
C0310915|T121|OAP|9079002|SNOMEDCT_US|Canine coronavirus - parvovirus vaccine - leptospira bacterin|Canine coronavirus - parvovirus vaccine - leptospira bacterin
C0310915|T129|OAP|9079002|SNOMEDCT_US|Canine coronavirus - parvovirus vaccine - leptospira bacterin|Canine coronavirus - parvovirus vaccine - leptospira bacterin
C0310915|T116|OAF|9079002|SNOMEDCT_US|Canine coronavirus - parvovirus vaccine - leptospira bacterin (product)|Canine coronavirus - parvovirus vaccine - leptospira bacterin (product)
C0310915|T121|OAF|9079002|SNOMEDCT_US|Canine coronavirus - parvovirus vaccine - leptospira bacterin (product)|Canine coronavirus - parvovirus vaccine - leptospira bacterin (product)
C0310915|T129|OAF|9079002|SNOMEDCT_US|Canine coronavirus - parvovirus vaccine - leptospira bacterin (product)|Canine coronavirus - parvovirus vaccine - leptospira bacterin (product)
C0310915|T116|OF|9079002|SNOMEDCT_US|Canine coronavirus - parvovirus vaccine - leptospira bacterin (substance)|Canine coronavirus - parvovirus vaccine - leptospira bacterin (substance)
C0310915|T121|OF|9079002|SNOMEDCT_US|Canine coronavirus - parvovirus vaccine - leptospira bacterin (substance)|Canine coronavirus - parvovirus vaccine - leptospira bacterin (substance)
C0310915|T129|OF|9079002|SNOMEDCT_US|Canine coronavirus - parvovirus vaccine - leptospira bacterin (substance)|Canine coronavirus - parvovirus vaccine - leptospira bacterin (substance)
C0310916|T116|OAP|30777008|SNOMEDCT_US|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine - leptospira bacterin|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine - leptospira bacterin
C0310916|T121|OAP|30777008|SNOMEDCT_US|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine - leptospira bacterin|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine - leptospira bacterin
C0310916|T129|OAP|30777008|SNOMEDCT_US|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine - leptospira bacterin|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine - leptospira bacterin
C0310916|T116|OAF|30777008|SNOMEDCT_US|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine - leptospira bacterin (product)|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine - leptospira bacterin (product)
C0310916|T121|OAF|30777008|SNOMEDCT_US|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine - leptospira bacterin (product)|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine - leptospira bacterin (product)
C0310916|T129|OAF|30777008|SNOMEDCT_US|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine - leptospira bacterin (product)|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine - leptospira bacterin (product)
C0310916|T116|OF|30777008|SNOMEDCT_US|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine - leptospira bacterin (substance)|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine - leptospira bacterin (substance)
C0310916|T121|OF|30777008|SNOMEDCT_US|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine - leptospira bacterin (substance)|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine - leptospira bacterin (substance)
C0310916|T129|OF|30777008|SNOMEDCT_US|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine - leptospira bacterin (substance)|Canine distemper - adenovirus type 2 - coronavirus - parainfluenza - parvovirus vaccine - leptospira bacterin (substance)
C0311097|T074|OAP|64592008|SNOMEDCT_US|Mycoplasma pulmonis - rodent coronavirus - sendai virus antibody test kit|Mycoplasma pulmonis - rodent coronavirus - sendai virus antibody test kit
C0311097|T074|OAF|64592008|SNOMEDCT_US|Mycoplasma pulmonis - rodent coronavirus - sendai virus antibody test kit (substance)|Mycoplasma pulmonis - rodent coronavirus - sendai virus antibody test kit (substance)
C0311110|T074|OAP|49159001|SNOMEDCT_US|Rat coronavirus sialodacryoadenitis virus antibody test kit|Rat coronavirus sialodacryoadenitis virus antibody test kit
C0311110|T074|OAF|49159001|SNOMEDCT_US|Rat coronavirus sialodacryoadenitis virus antibody test kit (substance)|Rat coronavirus sialodacryoadenitis virus antibody test kit (substance)
C0318856|T005|PM|D045722|MSH|Coronavirus, Porcine Respiratory|Coronavirus, Porcine Respiratory
C0318856|T005|LPN|LP19934-6|LNC|Porcine respiratory coronavirus|Porcine respiratory coronavirus
C0318856|T005|PT|15226006|SNOMEDCT_US|Porcine respiratory coronavirus|Porcine respiratory coronavirus
C0318856|T005|MH|D045722|MSH|Porcine Respiratory Coronavirus|Porcine Respiratory Coronavirus
C0318856|T005|FN|15226006|SNOMEDCT_US|Porcine respiratory coronavirus (organism)|Porcine respiratory coronavirus (organism)
C0318856|T005|PM|D045722|MSH|Respiratory Coronavirus, Porcine|Respiratory Coronavirus, Porcine
C0318858|T005|OAP|81773004|SNOMEDCT_US|Neonatal calf diarrhea coronavirus|Neonatal calf diarrhea coronavirus
C0318858|T005|OAF|81773004|SNOMEDCT_US|Neonatal calf diarrhea coronavirus (organism)|Neonatal calf diarrhea coronavirus (organism)
C0318858|T005|OAP|81773004|SNOMEDCT_US|Neonatal calf diarrhoea coronavirus|Neonatal calf diarrhoea coronavirus
C0318859|T005|OAP|64219004|SNOMEDCT_US|Winter dysentery bovine coronavirus|Winter dysentery bovine coronavirus
C0318859|T005|OAF|64219004|SNOMEDCT_US|Winter dysentery bovine coronavirus (organism)|Winter dysentery bovine coronavirus (organism)
C0318861|T005|PEP|D000073641|MSH|Human enteric coronavirus|Human enteric coronavirus
C0318861|T005|PT|70986004|SNOMEDCT_US|Human enteric coronavirus|Human enteric coronavirus
C0318861|T005|FN|70986004|SNOMEDCT_US|Human enteric coronavirus (organism)|Human enteric coronavirus (organism)
C0318861|T005|PM|D000073641|MSH|Human enteric coronaviruses|Human enteric coronaviruses
C0348984|T047|OA|A7y00|RCD|Coronavir caus dis clas oth ch|Coronavir caus dis clas oth ch
C0348984|T047|OA|A7y00|RCD|Coronavirus as cause of dis classified to other chapters|Coronavirus as cause of dis classified to other chapters
C0348984|T047|OP|A7y00|RCD|Coronavirus as the cause of diseases classified to other chapters|Coronavirus as the cause of diseases classified to other chapters
C0348984|T047|OAP|186758000|SNOMEDCT_US|Coronavirus as the cause of diseases classified to other chapters|Coronavirus as the cause of diseases classified to other chapters
C0348984|T047|OAP|187587009|SNOMEDCT_US|Coronavirus as the cause of diseases classified to other chapters|Coronavirus as the cause of diseases classified to other chapters
C0348984|T047|OF|187587009|SNOMEDCT_US|Coronavirus as the cause of diseases classified to other chapters|Coronavirus as the cause of diseases classified to other chapters
C0348984|T047|PT|B97.2|ICD10|Coronavirus as the cause of diseases classified to other chapters|Coronavirus as the cause of diseases classified to other chapters
C0348984|T047|OAF|187587009|SNOMEDCT_US|Coronavirus as the cause of diseases classified to other chapters (disorder)|Coronavirus as the cause of diseases classified to other chapters (disorder)
C0348984|T047|OAF|186758000|SNOMEDCT_US|Coronavirus as the cause of diseases classified to other chapters (disorder)|Coronavirus as the cause of diseases classified to other chapters (disorder)
C0368227|T201|LC|5099-7|LNC|Coronavirus Ab [Units/volume] in Serum|Coronavirus Ab [Units/volume] in Serum
C0368227|T201|DN|5099-7|LNC|Coronavirus Ab Qn (S)|Coronavirus Ab Qn (S)
C0368227|T201|OSN|5099-7|LNC|Coronavirus Ab Ser-aCnc|Coronavirus Ab Ser-aCnc
C0368227|T201|LN|5099-7|LNC|Coronavirus Ab:ACnc:Pt:Ser:Qn|Coronavirus Ab:ACnc:Pt:Ser:Qn
C0368227|T201|MTH_LN|5099-7|LNC|Coronavirus Antibody:Arbitrary Concentration:Point in time:Serum:Quantitative|Coronavirus Antibody:Arbitrary Concentration:Point in time:Serum:Quantitative
C0369034|T116|LPN|LP37778-5|LNC|Coronavirus Ab|Coronavirus Ab
C0369034|T129|LPN|LP37778-5|LNC|Coronavirus Ab|Coronavirus Ab
C0369034|T116|CN|MTHU022123|LNC|Coronavirus Ab|Coronavirus Ab
C0369034|T129|CN|MTHU022123|LNC|Coronavirus Ab|Coronavirus Ab
C0369034|T116|PT|120814005|SNOMEDCT_US|Coronavirus antibody|Coronavirus antibody
C0369034|T129|PT|120814005|SNOMEDCT_US|Coronavirus antibody|Coronavirus antibody
C0369034|T116|MTH_CN|MTHU022123|LNC|Coronavirus Antibody|Coronavirus Antibody
C0369034|T129|MTH_CN|MTHU022123|LNC|Coronavirus Antibody|Coronavirus Antibody
C0369034|T116|FN|120814005|SNOMEDCT_US|Coronavirus antibody (substance)|Coronavirus antibody (substance)
C0369034|T129|FN|120814005|SNOMEDCT_US|Coronavirus antibody (substance)|Coronavirus antibody (substance)
C0389916|T114|CE|C099602|MSH|N protein, Coronavirus|N protein, Coronavirus
C0389916|T116|CE|C099602|MSH|N protein, Coronavirus|N protein, Coronavirus
C0389916|T114|NM|C099602|MSH|nucleocapsid protein, Coronavirus|nucleocapsid protein, Coronavirus
C0389916|T116|NM|C099602|MSH|nucleocapsid protein, Coronavirus|nucleocapsid protein, Coronavirus
C0528529|T116|NM|C099456|MSH|3C-like proteinase, Coronavirus|3C-like proteinase, Coronavirus
C0528529|T126|NM|C099456|MSH|3C-like proteinase, Coronavirus|3C-like proteinase, Coronavirus
C0528529|T116|CE|C099456|MSH|M(pro) protein, Coronavirus|M(pro) protein, Coronavirus
C0528529|T126|CE|C099456|MSH|M(pro) protein, Coronavirus|M(pro) protein, Coronavirus
C0528529|T116|CE|C099456|MSH|main proteinase, Coronavirus|main proteinase, Coronavirus
C0528529|T126|CE|C099456|MSH|main proteinase, Coronavirus|main proteinase, Coronavirus
C0528529|T116|CE|C099456|MSH|Mpro protein, Coronavirus|Mpro protein, Coronavirus
C0528529|T126|CE|C099456|MSH|Mpro protein, Coronavirus|Mpro protein, Coronavirus
C0653195|T116|CE|C076115|MSH|I protein, BCV|I protein, BCV
C0653195|T116|CE|C076115|MSH|I protein, bovine coronavirus|I protein, bovine coronavirus
C0653195|T116|NM|C076115|MSH|internal ORF protein, bovine coronavirus|internal ORF protein, bovine coronavirus
C0753268|T116|PCE|C060814|MSH|HE protein, Coronavirus|HE protein, Coronavirus
C0766211|T116|CE|C118611|MSH|3b protein, coronavirus|3b protein, coronavirus
C0766211|T116|NM|C118611|MSH|glycoprotein 3b, coronavirus|glycoprotein 3b, coronavirus
C0803579|T201|OSN|20779-5|LNC|BCV Ag Tiss Ql IF|BCV Ag Tiss Ql IF
C0803579|T201|LC|20779-5|LNC|Bovine coronavirus Ag [Presence] in Tissue by Immunofluorescence|Bovine coronavirus Ag [Presence] in Tissue by Immunofluorescence
C0803579|T201|DN|20779-5|LNC|Bovine coronavirus Ag IF Ql (Tiss)|Bovine coronavirus Ag IF Ql (Tiss)
C0803579|T201|LN|20779-5|LNC|Bovine coronavirus Ag:PrThr:Pt:Tiss:Ord:IF|Bovine coronavirus Ag:PrThr:Pt:Tiss:Ord:IF
C0803579|T201|MTH_LN|20779-5|LNC|Bovine coronavirus Antigen:Presence or Threshold:Point in time:Tissue, unspecified:Ordinal:Immune Fluorescence|Bovine coronavirus Antigen:Presence or Threshold:Point in time:Tissue, unspecified:Ordinal:Immune Fluorescence
C0805362|T129|OAS|709225000|SNOMEDCT_US|Antigen of Bovine coronavirus|Antigen of Bovine coronavirus
C0805362|T129|OAF|709225000|SNOMEDCT_US|Antigen of Bovine coronavirus (substance)|Antigen of Bovine coronavirus (substance)
C0805362|T129|LPN|LP37387-5|LNC|Bovine coronavirus Ag|Bovine coronavirus Ag
C0805362|T129|OAP|709225000|SNOMEDCT_US|Bovine coronavirus Ag|Bovine coronavirus Ag
C0805362|T129|CN|MTHU009322|LNC|Bovine coronavirus Ag|Bovine coronavirus Ag
C0805362|T129|MTH_CN|MTHU009322|LNC|Bovine coronavirus Antigen|Bovine coronavirus Antigen
C0805362|T129|OAS|709225000|SNOMEDCT_US|Bovine coronavirus antigen|Bovine coronavirus antigen
C0880795|T201|LC|23372-6|LNC|Porcine respiratory coronavirus Ab [Presence] in Serum|Porcine respiratory coronavirus Ab [Presence] in Serum
C0880795|T201|DN|23372-6|LNC|Porcine respiratory coronavirus Ab Ql (S)|Porcine respiratory coronavirus Ab Ql (S)
C0880795|T201|LN|23372-6|LNC|Porcine respiratory coronavirus Ab:PrThr:Pt:Ser:Ord|Porcine respiratory coronavirus Ab:PrThr:Pt:Ser:Ord
C0880795|T201|PN|NOCODE|MTH|Porcine respiratory coronavirus Antibody:Arbitrary Concentration:Point in time:Serum:Ordinal|Porcine respiratory coronavirus Antibody:Arbitrary Concentration:Point in time:Serum:Ordinal
C0880795|T201|MTH_LN|23372-6|LNC|Porcine respiratory coronavirus Antibody:Presence or Threshold:Point in time:Serum:Ordinal|Porcine respiratory coronavirus Antibody:Presence or Threshold:Point in time:Serum:Ordinal
C0880795|T201|OSN|23372-6|LNC|PRCoV Ab Ser Ql|PRCoV Ab Ser Ql
C0880796|T201|LC|23374-2|LNC|Porcine respiratory coronavirus Ab [Presence] in Serum by Immunoassay|Porcine respiratory coronavirus Ab [Presence] in Serum by Immunoassay
C0880796|T201|DN|23374-2|LNC|Porcine respiratory coronavirus Ab IA Ql (S)|Porcine respiratory coronavirus Ab IA Ql (S)
C0880796|T201|LN|23374-2|LNC|Porcine respiratory coronavirus Ab:PrThr:Pt:Ser:Ord:IA|Porcine respiratory coronavirus Ab:PrThr:Pt:Ser:Ord:IA
C0880796|T201|MTH_LN|23374-2|LNC|Porcine respiratory coronavirus Antibody:Presence or Threshold:Point in time:Serum:Ordinal:Enzyme Immunoassay|Porcine respiratory coronavirus Antibody:Presence or Threshold:Point in time:Serum:Ordinal:Enzyme Immunoassay
C0880796|T201|OSN|23374-2|LNC|PRCoV Ab Ser Ql IA|PRCoV Ab Ser Ql IA
C0880797|T201|LC|23376-7|LNC|Porcine respiratory coronavirus Ag [Presence] in Unspecified specimen by Immune stain|Porcine respiratory coronavirus Ag [Presence] in Unspecified specimen by Immune stain
C0880797|T201|DN|23376-7|LNC|Porcine respiratory coronavirus Ag Immune stain Ql (Unsp spec)|Porcine respiratory coronavirus Ag Immune stain Ql (Unsp spec)
C0880797|T201|LN|23376-7|LNC|Porcine respiratory coronavirus Ag:PrThr:Pt:XXX:Ord:Immune stain|Porcine respiratory coronavirus Ag:PrThr:Pt:XXX:Ord:Immune stain
C0880797|T201|MTH_LN|23376-7|LNC|Porcine respiratory coronavirus Antigen:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:Immune stain|Porcine respiratory coronavirus Antigen:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:Immune stain
C0880797|T201|OSN|23376-7|LNC|PRCoV Ag XXX Ql ImStn|PRCoV Ag XXX Ql ImStn
C0880798|T201|LC|23377-5|LNC|Porcine respiratory coronavirus Ag [Presence] in Small intestine Tissue by Immune stain|Porcine respiratory coronavirus Ag [Presence] in Small intestine Tissue by Immune stain
C0880798|T201|DN|23377-5|LNC|Porcine respiratory coronavirus Ag Immune stain Ql (Small intestine Tissue)|Porcine respiratory coronavirus Ag Immune stain Ql (Small intestine Tissue)
C0880798|T201|LN|23377-5|LNC|Porcine respiratory coronavirus Ag:PrThr:Pt:Tsmi:Ord:Immune stain|Porcine respiratory coronavirus Ag:PrThr:Pt:Tsmi:Ord:Immune stain
C0880798|T201|MTH_LN|23377-5|LNC|Porcine respiratory coronavirus Antigen:Presence or Threshold:Point in time:Tissue small intestine:Ordinal:Immune stain|Porcine respiratory coronavirus Antigen:Presence or Threshold:Point in time:Tissue small intestine:Ordinal:Immune stain
C0880798|T201|OSN|23377-5|LNC|PRCoV Ag TSMI Ql ImStn|PRCoV Ag TSMI Ql ImStn
C0880799|T201|MTH_LN|23378-3|LNC|Porcine respiratory coronavirus ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe|Porcine respiratory coronavirus ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe
C0880799|T201|LC|23378-3|LNC|Porcine respiratory coronavirus RNA [Presence] in Unspecified specimen by Probe|Porcine respiratory coronavirus RNA [Presence] in Unspecified specimen by Probe
C0880799|T201|DN|23378-3|LNC|Porcine respiratory coronavirus RNA Probe Ql (Unsp spec)|Porcine respiratory coronavirus RNA Probe Ql (Unsp spec)
C0880799|T201|LN|23378-3|LNC|Porcine respiratory coronavirus RNA:PrThr:Pt:XXX:Ord:Probe|Porcine respiratory coronavirus RNA:PrThr:Pt:XXX:Ord:Probe
C0880799|T201|OSN|23378-3|LNC|PRCoV RNA XXX Ql Probe|PRCoV RNA XXX Ql Probe
C0880934|T201|OSN|23540-8|LNC|TCoV Ser Ql IF|TCoV Ser Ql IF
C0880934|T201|LC|23540-8|LNC|Turkey enteritis coronavirus [Presence] in Serum by Immunofluorescence|Turkey enteritis coronavirus [Presence] in Serum by Immunofluorescence
C0880934|T201|DN|23540-8|LNC|Turkey enteritis coronavirus IF Ql (S)|Turkey enteritis coronavirus IF Ql (S)
C0880934|T201|MTH_LN|23540-8|LNC|Turkey enteritis coronavirus:Presence or Threshold:Point in time:Serum:Ordinal:Immune Fluorescence|Turkey enteritis coronavirus:Presence or Threshold:Point in time:Serum:Ordinal:Immune Fluorescence
C0880934|T201|LN|23540-8|LNC|Turkey enteritis coronavirus:PrThr:Pt:Ser:Ord:IF|Turkey enteritis coronavirus:PrThr:Pt:Ser:Ord:IF
C0881088|T201|OSN|23716-4|LNC|FCoV Ab Ser Ql IA|FCoV Ab Ser Ql IA
C0881088|T201|LC|23716-4|LNC|Feline coronavirus Ab [Presence] in Serum by Immunoassay|Feline coronavirus Ab [Presence] in Serum by Immunoassay
C0881088|T201|DN|23716-4|LNC|Feline coronavirus Ab IA Ql (S)|Feline coronavirus Ab IA Ql (S)
C0881088|T201|LN|23716-4|LNC|Feline coronavirus Ab:PrThr:Pt:Ser:Ord:IA|Feline coronavirus Ab:PrThr:Pt:Ser:Ord:IA
C0881088|T201|MTH_LN|23716-4|LNC|Feline coronavirus Antibody:Presence or Threshold:Point in time:Serum:Ordinal:Enzyme Immunoassay|Feline coronavirus Antibody:Presence or Threshold:Point in time:Serum:Ordinal:Enzyme Immunoassay
C0881089|T201|OSN|23717-2|LNC|FCoV Ab Ser Ql|FCoV Ab Ser Ql
C0881089|T201|LC|23717-2|LNC|Feline coronavirus Ab [Presence] in Serum|Feline coronavirus Ab [Presence] in Serum
C0881089|T201|DN|23717-2|LNC|Feline coronavirus Ab Ql (S)|Feline coronavirus Ab Ql (S)
C0881089|T201|LN|23717-2|LNC|Feline coronavirus Ab:PrThr:Pt:Ser:Ord|Feline coronavirus Ab:PrThr:Pt:Ser:Ord
C0881089|T201|MTH_LN|23717-2|LNC|Feline coronavirus Antibody:Presence or Threshold:Point in time:Serum:Ordinal|Feline coronavirus Antibody:Presence or Threshold:Point in time:Serum:Ordinal
C0881090|T201|OSN|23718-0|LNC|FCoV Ab Titr Ser|FCoV Ab Titr Ser
C0881090|T201|DN|23718-0|LNC|Feline coronavirus Ab (S) [Titer]|Feline coronavirus Ab (S) [Titer]
C0881090|T201|LC|23718-0|LNC|Feline coronavirus Ab [Titer] in Serum|Feline coronavirus Ab [Titer] in Serum
C0881090|T201|LN|23718-0|LNC|Feline coronavirus Ab:Titr:Pt:Ser:Qn|Feline coronavirus Ab:Titr:Pt:Ser:Qn
C0881090|T201|MTH_LN|23718-0|LNC|Feline coronavirus Antibody:Dilution Factor (Titer):Point in time:Serum:Quantitative|Feline coronavirus Antibody:Dilution Factor (Titer):Point in time:Serum:Quantitative
C0882387|T201|LC|23373-4|LNC|Porcine respiratory coronavirus Ab [Presence] in Serum by Neutralization test|Porcine respiratory coronavirus Ab [Presence] in Serum by Neutralization test
C0882387|T201|DN|23373-4|LNC|Porcine respiratory coronavirus Ab Neut test Ql (S)|Porcine respiratory coronavirus Ab Neut test Ql (S)
C0882387|T201|LN|23373-4|LNC|Porcine respiratory coronavirus Ab:PrThr:Pt:Ser:Ord:Neut|Porcine respiratory coronavirus Ab:PrThr:Pt:Ser:Ord:Neut
C0882387|T201|MTH_LN|23373-4|LNC|Porcine respiratory coronavirus Antibody:Presence or Threshold:Point in time:Serum:Ordinal:Neutralization|Porcine respiratory coronavirus Antibody:Presence or Threshold:Point in time:Serum:Ordinal:Neutralization
C0882387|T201|OSN|23373-4|LNC|PRCoV Ab Ser Ql Nt|PRCoV Ab Ser Ql Nt
C0882422|T201|LC|23687-7|LNC|Canine coronavirus Ab [Presence] in Serum by Immunofluorescence|Canine coronavirus Ab [Presence] in Serum by Immunofluorescence
C0882422|T201|DN|23687-7|LNC|Canine coronavirus Ab IF Ql (S)|Canine coronavirus Ab IF Ql (S)
C0882422|T201|LN|23687-7|LNC|Canine coronavirus Ab:PrThr:Pt:Ser:Ord:IF|Canine coronavirus Ab:PrThr:Pt:Ser:Ord:IF
C0882422|T201|MTH_LN|23687-7|LNC|Canine coronavirus Antibody:Presence or Threshold:Point in time:Serum:Ordinal:Immune Fluorescence|Canine coronavirus Antibody:Presence or Threshold:Point in time:Serum:Ordinal:Immune Fluorescence
C0882422|T201|OSN|23687-7|LNC|CCV Ab Ser Ql IF|CCV Ab Ser Ql IF
C0882423|T201|LC|23688-5|LNC|Canine coronavirus Ag [Presence] in Tissue by Immunofluorescence|Canine coronavirus Ag [Presence] in Tissue by Immunofluorescence
C0882423|T201|DN|23688-5|LNC|Canine coronavirus Ag IF Ql (Tiss)|Canine coronavirus Ag IF Ql (Tiss)
C0882423|T201|LN|23688-5|LNC|Canine coronavirus Ag:PrThr:Pt:Tiss:Ord:IF|Canine coronavirus Ag:PrThr:Pt:Tiss:Ord:IF
C0882423|T201|MTH_LN|23688-5|LNC|Canine coronavirus Antigen:Presence or Threshold:Point in time:Tissue, unspecified:Ordinal:Immune Fluorescence|Canine coronavirus Antigen:Presence or Threshold:Point in time:Tissue, unspecified:Ordinal:Immune Fluorescence
C0882423|T201|OSN|23688-5|LNC|CCV Ag Tiss Ql IF|CCV Ag Tiss Ql IF
C0882751|T116|LPN|LP37510-2|LNC|Canine coronavirus Ab|Canine coronavirus Ab
C0882751|T129|LPN|LP37510-2|LNC|Canine coronavirus Ab|Canine coronavirus Ab
C0882751|T116|CN|MTHU011428|LNC|Canine coronavirus Ab|Canine coronavirus Ab
C0882751|T129|CN|MTHU011428|LNC|Canine coronavirus Ab|Canine coronavirus Ab
C0882751|T116|MTH_CN|MTHU011428|LNC|Canine coronavirus Antibody|Canine coronavirus Antibody
C0882751|T129|MTH_CN|MTHU011428|LNC|Canine coronavirus Antibody|Canine coronavirus Antibody
C0883053|T116|LPN|LP38135-7|LNC|Feline coronavirus Ab|Feline coronavirus Ab
C0883053|T129|LPN|LP38135-7|LNC|Feline coronavirus Ab|Feline coronavirus Ab
C0883053|T116|CN|MTHU011458|LNC|Feline coronavirus Ab|Feline coronavirus Ab
C0883053|T129|CN|MTHU011458|LNC|Feline coronavirus Ab|Feline coronavirus Ab
C0883053|T116|MTH_CN|MTHU011458|LNC|Feline coronavirus Antibody|Feline coronavirus Antibody
C0883053|T129|MTH_CN|MTHU011458|LNC|Feline coronavirus Antibody|Feline coronavirus Antibody
C0883320|T116|SY|709962005|SNOMEDCT_US|Anti-Porcine respiratory coronavirus antibody|Anti-Porcine respiratory coronavirus antibody
C0883320|T129|SY|709962005|SNOMEDCT_US|Anti-Porcine respiratory coronavirus antibody|Anti-Porcine respiratory coronavirus antibody
C0883320|T116|SY|709962005|SNOMEDCT_US|Antibody to Porcine respiratory coronavirus|Antibody to Porcine respiratory coronavirus
C0883320|T129|SY|709962005|SNOMEDCT_US|Antibody to Porcine respiratory coronavirus|Antibody to Porcine respiratory coronavirus
C0883320|T116|FN|709962005|SNOMEDCT_US|Antibody to Porcine respiratory coronavirus (substance)|Antibody to Porcine respiratory coronavirus (substance)
C0883320|T129|FN|709962005|SNOMEDCT_US|Antibody to Porcine respiratory coronavirus (substance)|Antibody to Porcine respiratory coronavirus (substance)
C0883320|T116|LPN|LP39469-9|LNC|Porcine respiratory coronavirus Ab|Porcine respiratory coronavirus Ab
C0883320|T129|LPN|LP39469-9|LNC|Porcine respiratory coronavirus Ab|Porcine respiratory coronavirus Ab
C0883320|T116|CN|MTHU011210|LNC|Porcine respiratory coronavirus Ab|Porcine respiratory coronavirus Ab
C0883320|T129|CN|MTHU011210|LNC|Porcine respiratory coronavirus Ab|Porcine respiratory coronavirus Ab
C0883320|T116|PT|709962005|SNOMEDCT_US|Porcine respiratory coronavirus Ab|Porcine respiratory coronavirus Ab
C0883320|T129|PT|709962005|SNOMEDCT_US|Porcine respiratory coronavirus Ab|Porcine respiratory coronavirus Ab
C0883320|T116|SY|709962005|SNOMEDCT_US|Porcine respiratory coronavirus antibody|Porcine respiratory coronavirus antibody
C0883320|T129|SY|709962005|SNOMEDCT_US|Porcine respiratory coronavirus antibody|Porcine respiratory coronavirus antibody
C0883320|T116|MTH_CN|MTHU011210|LNC|Porcine respiratory coronavirus Antibody|Porcine respiratory coronavirus Antibody
C0883320|T129|MTH_CN|MTHU011210|LNC|Porcine respiratory coronavirus Antibody|Porcine respiratory coronavirus Antibody
C0883321|T116|LPN|LP39470-7|LNC|Porcine respiratory coronavirus Ag|Porcine respiratory coronavirus Ag
C0883321|T129|LPN|LP39470-7|LNC|Porcine respiratory coronavirus Ag|Porcine respiratory coronavirus Ag
C0883321|T116|CN|MTHU011212|LNC|Porcine respiratory coronavirus Ag|Porcine respiratory coronavirus Ag
C0883321|T129|CN|MTHU011212|LNC|Porcine respiratory coronavirus Ag|Porcine respiratory coronavirus Ag
C0883321|T116|MTH_CN|MTHU011212|LNC|Porcine respiratory coronavirus Antigen|Porcine respiratory coronavirus Antigen
C0883321|T129|MTH_CN|MTHU011212|LNC|Porcine respiratory coronavirus Antigen|Porcine respiratory coronavirus Antigen
C0883322|T114|MTH_CN|MTHU011214|LNC|Porcine respiratory coronavirus ribonucleic acid|Porcine respiratory coronavirus ribonucleic acid
C0883322|T114|LPN|LP39471-5|LNC|Porcine respiratory coronavirus RNA|Porcine respiratory coronavirus RNA
C0883322|T114|CN|MTHU011214|LNC|Porcine respiratory coronavirus RNA|Porcine respiratory coronavirus RNA
C0883322|T114|PT|707945006|SNOMEDCT_US|Porcine respiratory coronavirus RNA|Porcine respiratory coronavirus RNA
C0883322|T114|SY|707945006|SNOMEDCT_US|Ribonucleic acid of Porcine respiratory coronavirus|Ribonucleic acid of Porcine respiratory coronavirus
C0883322|T114|FN|707945006|SNOMEDCT_US|Ribonucleic acid of Porcine respiratory coronavirus (substance)|Ribonucleic acid of Porcine respiratory coronavirus (substance)
C0883460|T116|OAS|709320007|SNOMEDCT_US|Antigen of Canine coronavirus|Antigen of Canine coronavirus
C0883460|T129|OAS|709320007|SNOMEDCT_US|Antigen of Canine coronavirus|Antigen of Canine coronavirus
C0883460|T116|OAF|709320007|SNOMEDCT_US|Antigen of Canine coronavirus (substance)|Antigen of Canine coronavirus (substance)
C0883460|T129|OAF|709320007|SNOMEDCT_US|Antigen of Canine coronavirus (substance)|Antigen of Canine coronavirus (substance)
C0883460|T116|LPN|LP37511-0|LNC|Canine coronavirus Ag|Canine coronavirus Ag
C0883460|T129|LPN|LP37511-0|LNC|Canine coronavirus Ag|Canine coronavirus Ag
C0883460|T116|OAP|709320007|SNOMEDCT_US|Canine coronavirus Ag|Canine coronavirus Ag
C0883460|T129|OAP|709320007|SNOMEDCT_US|Canine coronavirus Ag|Canine coronavirus Ag
C0883460|T116|CN|MTHU011430|LNC|Canine coronavirus Ag|Canine coronavirus Ag
C0883460|T129|CN|MTHU011430|LNC|Canine coronavirus Ag|Canine coronavirus Ag
C0883460|T116|MTH_CN|MTHU011430|LNC|Canine coronavirus Antigen|Canine coronavirus Antigen
C0883460|T129|MTH_CN|MTHU011430|LNC|Canine coronavirus Antigen|Canine coronavirus Antigen
C0883460|T116|OAS|709320007|SNOMEDCT_US|Canine coronavirus antigen|Canine coronavirus antigen
C0883460|T129|OAS|709320007|SNOMEDCT_US|Canine coronavirus antigen|Canine coronavirus antigen
C0936087|T005|MH|D016765|MSH|Coronavirus, Feline|Coronavirus, Feline
C0936087|T005|ET|D016765|MSH|Coronavirus, Feline Enteric|Coronavirus, Feline Enteric
C0936087|T005|PM|D016765|MSH|Coronaviruses, Feline|Coronaviruses, Feline
C0936087|T005|PM|D016765|MSH|Coronaviruses, Feline Enteric|Coronaviruses, Feline Enteric
C0936087|T005|PM|D016765|MSH|Enteric Coronavirus, Feline|Enteric Coronavirus, Feline
C0936087|T005|PM|D016765|MSH|Enteric Coronaviruses, Feline|Enteric Coronaviruses, Feline
C0936087|T005|ET|D016765|MSH|FECV|FECV
C0936087|T005|LPN|LP14108-2|LNC|Feline coronavirus|Feline coronavirus
C0936087|T005|PT|407366004|SNOMEDCT_US|Feline coronavirus|Feline coronavirus
C0936087|T005|PM|D016765|MSH|Feline Coronavirus|Feline Coronavirus
C0936087|T005|PT|0000052845|CHV|feline coronavirus|feline coronavirus
C0936087|T005|FN|407366004|SNOMEDCT_US|Feline coronavirus (organism)|Feline coronavirus (organism)
C0936087|T005|PM|D016765|MSH|Feline Coronaviruses|Feline Coronaviruses
C0936087|T005|OAS|49835008|SNOMEDCT_US|Feline enteric coronavirus|Feline enteric coronavirus
C0936087|T005|SY|407366004|SNOMEDCT_US|Feline enteric coronavirus|Feline enteric coronavirus
C0936087|T005|ET|D016765|MSH|Feline Enteric Coronavirus|Feline Enteric Coronavirus
C0936087|T005|PM|D016765|MSH|Feline Enteric Coronaviruses|Feline Enteric Coronaviruses
C0949525|T005|PEP|D017934|MSH|Coronavirus, Rabbit|Coronavirus, Rabbit
C0949525|T005|PM|D017934|MSH|Coronaviruses, Rabbit|Coronaviruses, Rabbit
C0949525|T005|ET|D017934|MSH|Rabbit Coronavirus|Rabbit Coronavirus
C0949525|T005|PM|D017934|MSH|Rabbit Coronaviruses|Rabbit Coronaviruses
C0949880|T005|OAP|418746002|SNOMEDCT_US|Coronavirus 229E|Coronavirus 229E
C0949880|T005|LA|LA26147-1|LNC|Coronavirus 229E|Coronavirus 229E
C0949880|T005|OAF|418746002|SNOMEDCT_US|Coronavirus 229E (organism)|Coronavirus 229E (organism)
C0949880|T005|MH|D028941|MSH|Coronavirus 229E, Human|Coronavirus 229E, Human
C0949880|T005|DSV|D028941|MSH|CORONAVIRUS HUMAN A 229 E|CORONAVIRUS HUMAN A 229 E
C0949880|T005|ET|D028941|MSH|HCoV-229E|HCoV-229E
C0949880|T005|LPN|LP35708-4|LNC|Human coronavirus 229E|Human coronavirus 229E
C0949880|T005|PT|407370007|SNOMEDCT_US|Human coronavirus 229E|Human coronavirus 229E
C0949880|T005|PN|NOCODE|MTH|Human coronavirus 229E|Human coronavirus 229E
C0949880|T005|ET|D028941|MSH|Human Coronavirus 229E|Human Coronavirus 229E
C0949880|T005|FN|407370007|SNOMEDCT_US|Human coronavirus 229E (organism)|Human coronavirus 229E (organism)
C0949880|T005|IS|407370007|SNOMEDCT_US|Human coronavirus 299E|Human coronavirus 299E
C0949880|T005|OF|407370007|SNOMEDCT_US|Human coronavirus 299E (organism)|Human coronavirus 299E (organism)
C0949880|T005|DSV|D028941|MSH|HUMAN CORONAVIRUS A 229 E|HUMAN CORONAVIRUS A 229 E
C0949881|T005|DSV|D028962|MSH|CORONAVIRUS HUMAN OC 043|CORONAVIRUS HUMAN OC 043
C0949881|T005|MH|D028962|MSH|Coronavirus OC43, Human|Coronavirus OC43, Human
C0949881|T005|ET|D028962|MSH|HCoV-OC43|HCoV-OC43
C0949881|T005|DSV|D028962|MSH|HUMAN CORONAVIRUS OC 043|HUMAN CORONAVIRUS OC 043
C0949881|T005|LPN|LP35710-0|LNC|Human coronavirus OC43|Human coronavirus OC43
C0949881|T005|PT|407371006|SNOMEDCT_US|Human coronavirus OC43|Human coronavirus OC43
C0949881|T005|ET|D028962|MSH|Human Coronavirus OC43|Human Coronavirus OC43
C0949881|T005|FN|407371006|SNOMEDCT_US|Human coronavirus OC43 (organism)|Human coronavirus OC43 (organism)
C1146968|T201|LC|31283-5|LNC|Canine coronavirus Ab [Presence] in Serum|Canine coronavirus Ab [Presence] in Serum
C1146968|T201|DN|31283-5|LNC|Canine coronavirus Ab Ql (S)|Canine coronavirus Ab Ql (S)
C1146968|T201|LN|31283-5|LNC|Canine coronavirus Ab:PrThr:Pt:Ser:Ord|Canine coronavirus Ab:PrThr:Pt:Ser:Ord
C1146968|T201|MTH_LN|31283-5|LNC|Canine coronavirus Antibody:Presence or Threshold:Point in time:Serum:Ordinal|Canine coronavirus Antibody:Presence or Threshold:Point in time:Serum:Ordinal
C1146968|T201|OSN|31283-5|LNC|CCV Ab Ser Ql|CCV Ab Ser Ql
C1147070|T201|OSN|31385-8|LNC|FCoV Ab Ser-aCnc|FCoV Ab Ser-aCnc
C1147070|T201|LC|31385-8|LNC|Feline coronavirus Ab [Units/volume] in Serum|Feline coronavirus Ab [Units/volume] in Serum
C1147070|T201|DN|31385-8|LNC|Feline coronavirus Ab Qn (S)|Feline coronavirus Ab Qn (S)
C1147070|T201|LN|31385-8|LNC|Feline coronavirus Ab:ACnc:Pt:Ser:Qn|Feline coronavirus Ab:ACnc:Pt:Ser:Qn
C1147070|T201|MTH_LN|31385-8|LNC|Feline coronavirus Antibody:Arbitrary Concentration:Point in time:Serum:Quantitative|Feline coronavirus Antibody:Arbitrary Concentration:Point in time:Serum:Quantitative
C1175175|T047|PT|3181|MEDLINEPLUS|Coronavirus Infections|Coronavirus Infections
C1175175|T047|SY|330007|MEDCIN|coronavirus sars-associated|coronavirus sars-associated
C1175175|T047|ET|D045169|MSH|Respiratory Syndrome, Acute, Severe|Respiratory Syndrome, Acute, Severe
C1175175|T047|ET|D045169|MSH|Respiratory Syndrome, Severe Acute|Respiratory Syndrome, Severe Acute
C1175175|T047|SY|272816|MEDCIN|SARS|SARS
C1175175|T047|AB|C85064|NCI|SARS|SARS
C1175175|T047|LPN|LP71047-2|LNC|SARS|SARS
C1175175|T047|SY|0000055815|CHV|SARS|SARS
C1175175|T047|ET|3181|MEDLINEPLUS|SARS|SARS
C1175175|T047|LA|LA10504-1|LNC|SARS|SARS
C1175175|T047|LLT|10061986|MDR|SARS|SARS
C1175175|T047|SY|C85064|NCI_NICHD|SARS|SARS
C1175175|T047|ET|5004-0074|CSP|SARS|SARS
C1175175|T047|SY|398447004|SNOMEDCT_US|SARS|SARS
C1175175|T047|ET|D045169|MSH|SARS (Severe Acute Respiratory Syndrome)|SARS (Severe Acute Respiratory Syndrome)
C1175175|T047|AB|079.82|ICD9CM|SARS assoc coronavirus|SARS assoc coronavirus
C1175175|T047|PT|079.82|ICD9CM|SARS-associated coronavirus|SARS-associated coronavirus
C1175175|T047|PT|330007|MEDCIN|SARS-associated coronavirus|SARS-associated coronavirus
C1175175|T047|FN|330007|MEDCIN|SARS-associated coronavirus (diagnosis)|SARS-associated coronavirus (diagnosis)
C1175175|T047|SY|398447004|SNOMEDCT_US|SARS-CoV infection|SARS-CoV infection
C1175175|T047|PT|C85064|NCI|Severe Acute Respiratory Syndrome|Severe Acute Respiratory Syndrome
C1175175|T047|ET|3181|MEDLINEPLUS|Severe Acute Respiratory Syndrome|Severe Acute Respiratory Syndrome
C1175175|T047|MH|D045169|MSH|Severe Acute Respiratory Syndrome|Severe Acute Respiratory Syndrome
C1175175|T047|PT|C85064|NCI_NICHD|Severe Acute Respiratory Syndrome|Severe Acute Respiratory Syndrome
C1175175|T047|PN|NOCODE|MTH|Severe Acute Respiratory Syndrome|Severe Acute Respiratory Syndrome
C1175175|T047|LLT|10061982|MDR|Severe acute respiratory syndrome|Severe acute respiratory syndrome
C1175175|T047|PT|10061982|MDR|Severe acute respiratory syndrome|Severe acute respiratory syndrome
C1175175|T047|PT|398447004|SNOMEDCT_US|Severe acute respiratory syndrome|Severe acute respiratory syndrome
C1175175|T047|PT|5004-0074|CSP|severe acute respiratory syndrome|severe acute respiratory syndrome
C1175175|T047|FN|398447004|SNOMEDCT_US|Severe acute respiratory syndrome (disorder)|Severe acute respiratory syndrome (disorder)
C1175175|T047|PT|0000055815|CHV|severe acute respiratory syndrome (SARS)|severe acute respiratory syndrome (SARS)
C1175175|T047|PT|272816|MEDCIN|severe acute respiratory syndrome (SARS)|severe acute respiratory syndrome (SARS)
C1175175|T047|FN|272816|MEDCIN|severe acute respiratory syndrome (SARS) (diagnosis)|severe acute respiratory syndrome (SARS) (diagnosis)
C1175175|T047|ET|J12.81|ICD10CM|Severe acute respiratory syndrome NOS|Severe acute respiratory syndrome NOS
C1175743|T005|SY|0000055818|CHV|coronavirus SARS|coronavirus SARS
C1175743|T005|PM|D045473|MSH|Coronavirus, SARS|Coronavirus, SARS
C1175743|T005|PM|D045473|MSH|Coronavirus, SARS-Associated|Coronavirus, SARS-Associated
C1175743|T005|PM|D045473|MSH|Coronavirus, SARS-Related|Coronavirus, SARS-Related
C1175743|T005|PM|D045473|MSH|Coronavirus, Urbani SARS-Associated|Coronavirus, Urbani SARS-Associated
C1175743|T005|SY|C112432|NCI_CDISC|HCoV-SARS|HCoV-SARS
C1175743|T005|SY|C112432|NCI_CDISC|SARS|SARS
C1175743|T005|SY|415360003|SNOMEDCT_US|SARS|SARS
C1175743|T005|DEV|D045473|MSH|SARS ASSOC CORONAVIRUS|SARS ASSOC CORONAVIRUS
C1175743|T005|PM|D045473|MSH|SARS Associated Coronavirus|SARS Associated Coronavirus
C1175743|T005|LPN|LP35807-4|LNC|SARS coronavirus|SARS coronavirus
C1175743|T005|SY|0000055818|CHV|SARS coronavirus|SARS coronavirus
C1175743|T005|CN|MTHU044721|LNC|SARS coronavirus|SARS coronavirus
C1175743|T005|PT|415360003|SNOMEDCT_US|SARS coronavirus|SARS coronavirus
C1175743|T005|PN|NOCODE|MTH|SARS coronavirus|SARS coronavirus
C1175743|T005|PT|C112432|NCI|SARS Coronavirus|SARS Coronavirus
C1175743|T005|ET|D045473|MSH|SARS Coronavirus|SARS Coronavirus
C1175743|T005|PT|C112432|NCI_CDISC|SARS CORONAVIRUS|SARS CORONAVIRUS
C1175743|T005|OF|415360003|SNOMEDCT_US|SARS coronavirus (organism)|SARS coronavirus (organism)
C1175743|T005|DEV|D045473|MSH|SARS RELAT CORONAVIRUS|SARS RELAT CORONAVIRUS
C1175743|T005|PM|D045473|MSH|SARS Related Coronavirus|SARS Related Coronavirus
C1175743|T005|PT|0000055818|CHV|SARS virus|SARS virus
C1175743|T005|PT|5004-0073|CSP|SARS virus|SARS virus
C1175743|T005|SY|415360003|SNOMEDCT_US|SARS virus|SARS virus
C1175743|T005|MH|D045473|MSH|SARS Virus|SARS Virus
C1175743|T005|ET|D045473|MSH|SARS-Associated Coronavirus|SARS-Associated Coronavirus
C1175743|T005|PM|D045473|MSH|SARS-Associated Coronavirus, Urbani|SARS-Associated Coronavirus, Urbani
C1175743|T005|ET|D045473|MSH|SARS-CoV|SARS-CoV
C1175743|T005|SY|C112432|NCI|SARS-CoV|SARS-CoV
C1175743|T005|SY|415360003|SNOMEDCT_US|SARS-CoV|SARS-CoV
C1175743|T005|SY|0000055818|CHV|sars-cov|sars-cov
C1175743|T005|ET|D045473|MSH|SARS-Related Coronavirus|SARS-Related Coronavirus
C1175743|T005|SY|415360003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus|Severe acute respiratory syndrome (SARS) coronavirus
C1175743|T005|OF|415360003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus (organism)|Severe acute respiratory syndrome (SARS) coronavirus (organism)
C1175743|T005|SY|415360003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus|Severe acute respiratory syndrome coronavirus
C1175743|T005|SY|C112432|NCI_CDISC|Severe Acute Respiratory Syndrome Coronavirus|Severe Acute Respiratory Syndrome Coronavirus
C1175743|T005|OF|415360003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus (organism)|Severe acute respiratory syndrome coronavirus (organism)
C1175743|T005|PM|D045473|MSH|Severe acute respiratory syndrome related coronavirus|Severe acute respiratory syndrome related coronavirus
C1175743|T005|ET|D045473|MSH|Severe Acute Respiratory Syndrome Virus|Severe Acute Respiratory Syndrome Virus
C1175743|T005|ET|D045473|MSH|Severe acute respiratory syndrome-related coronavirus|Severe acute respiratory syndrome-related coronavirus
C1175743|T005|SY|415360003|SNOMEDCT_US|Severe acute respiratory syndrome-related coronavirus|Severe acute respiratory syndrome-related coronavirus
C1175743|T005|FN|415360003|SNOMEDCT_US|Severe acute respiratory syndrome-related coronavirus (organism)|Severe acute respiratory syndrome-related coronavirus (organism)
C1175743|T005|DEV|D045473|MSH|URBANI SARS ASSOC CORONAVIRUS|URBANI SARS ASSOC CORONAVIRUS
C1175743|T005|PM|D045473|MSH|Urbani SARS Associated Coronavirus|Urbani SARS Associated Coronavirus
C1175743|T005|ET|D045473|MSH|Urbani SARS-Associated Coronavirus|Urbani SARS-Associated Coronavirus
C1175743|T005|SY|0000055818|CHV|virus SARS|virus SARS
C1258835|T116|CE|C099602|MSH|N protein, SARS virus|N protein, SARS virus
C1258835|T123|CE|C099602|MSH|N protein, SARS virus|N protein, SARS virus
C1258835|T116|CE|C099602|MSH|N protein, SARS-CoV|N protein, SARS-CoV
C1258835|T123|CE|C099602|MSH|N protein, SARS-CoV|N protein, SARS-CoV
C1258835|T116|PCE|C099602|MSH|N protein, Severe acute respiratory syndrome virus|N protein, Severe acute respiratory syndrome virus
C1258835|T123|PCE|C099602|MSH|N protein, Severe acute respiratory syndrome virus|N protein, Severe acute respiratory syndrome virus
C1258836|T116|CE|C067997|MSH|M protein, SARS virus|M protein, SARS virus
C1258836|T123|CE|C067997|MSH|M protein, SARS virus|M protein, SARS virus
C1258836|T116|CE|C067997|MSH|M protein, SARS-CoV|M protein, SARS-CoV
C1258836|T123|CE|C067997|MSH|M protein, SARS-CoV|M protein, SARS-CoV
C1258836|T116|PCE|C067997|MSH|M protein, Severe acute respiratory syndrome virus|M protein, Severe acute respiratory syndrome virus
C1258836|T123|PCE|C067997|MSH|M protein, Severe acute respiratory syndrome virus|M protein, Severe acute respiratory syndrome virus
C1258836|T116|CE|C067997|MSH|SARS-CoV M protein|SARS-CoV M protein
C1258836|T123|CE|C067997|MSH|SARS-CoV M protein|SARS-CoV M protein
C1258836|T116|CE|C067997|MSH|SARS-CoV membrane structural protein|SARS-CoV membrane structural protein
C1258836|T123|CE|C067997|MSH|SARS-CoV membrane structural protein|SARS-CoV membrane structural protein
C1260415|T047|SY|441590008|SNOMEDCT_US|Pneumonia caused by Severe acute respiratory syndrome coronavirus|Pneumonia caused by Severe acute respiratory syndrome coronavirus
C1260415|T047|FN|441590008|SNOMEDCT_US|Pneumonia caused by Severe acute respiratory syndrome coronavirus (disorder)|Pneumonia caused by Severe acute respiratory syndrome coronavirus (disorder)
C1260415|T047|AB|480.3|ICD9CM|Pneumonia due to SARS|Pneumonia due to SARS
C1260415|T047|AB|J12.81|ICD10CM|Pneumonia due to SARS-associated coronavirus|Pneumonia due to SARS-associated coronavirus
C1260415|T047|PT|480.3|ICD9CM|Pneumonia due to SARS-associated coronavirus|Pneumonia due to SARS-associated coronavirus
C1260415|T047|PT|J12.81|ICD10CM|Pneumonia due to SARS-associated coronavirus|Pneumonia due to SARS-associated coronavirus
C1260415|T047|PT|441590008|SNOMEDCT_US|Pneumonia due to Severe acute respiratory syndrome coronavirus|Pneumonia due to Severe acute respiratory syndrome coronavirus
C1260415|T047|OF|441590008|SNOMEDCT_US|Pneumonia due to Severe acute respiratory syndrome coronavirus (disorder)|Pneumonia due to Severe acute respiratory syndrome coronavirus (disorder)
C1260451|T033|PT|123661|MEDCIN|exposure to SARS|exposure to SARS
C1260451|T033|AB|V01.82|ICD9CM|Exposure to SARS|Exposure to SARS
C1260451|T033|FN|123661|MEDCIN|exposure to SARS (history)|exposure to SARS (history)
C1260451|T033|PT|V01.82|ICD9CM|Exposure to SARS-associated coronavirus|Exposure to SARS-associated coronavirus
C1275826|T059|PT|399150003|SNOMEDCT_US|PCR test for SARS|PCR test for SARS
C1275826|T059|SY|399150003|SNOMEDCT_US|Polymerase chain reaction test for SARS|Polymerase chain reaction test for SARS
C1275826|T059|OF|399150003|SNOMEDCT_US|Polymerase chain reaction test for SARS (procedure)|Polymerase chain reaction test for SARS (procedure)
C1275826|T059|SY|399150003|SNOMEDCT_US|Polymerase chain reaction test for severe acute respiratory syndrome|Polymerase chain reaction test for severe acute respiratory syndrome
C1275826|T059|FN|399150003|SNOMEDCT_US|Polymerase chain reaction test for severe acute respiratory syndrome (procedure)|Polymerase chain reaction test for severe acute respiratory syndrome (procedure)
C1275826|T059|SY|399150003|SNOMEDCT_US|SARS-CoV PCR|SARS-CoV PCR
C1294675|T059|SY|121973000|SNOMEDCT_US|Coronavirus antibody assay|Coronavirus antibody assay
C1294675|T059|OF|121973000|SNOMEDCT_US|Coronavirus antibody assay (procedure)|Coronavirus antibody assay (procedure)
C1294675|T059|PT|121973000|SNOMEDCT_US|Measurement of coronavirus antibody|Measurement of coronavirus antibody
C1294675|T059|FN|121973000|SNOMEDCT_US|Measurement of coronavirus antibody (procedure)|Measurement of coronavirus antibody (procedure)
C1294866|T059|PT|117945005|SNOMEDCT_US|Bovine coronavirus antigen assay|Bovine coronavirus antigen assay
C1294866|T059|FN|117945005|SNOMEDCT_US|Bovine coronavirus antigen assay (procedure)|Bovine coronavirus antigen assay (procedure)
C1312200|T116|NM|C477905|MSH|papain-like proteinase 2|papain-like proteinase 2
C1312200|T126|NM|C477905|MSH|papain-like proteinase 2|papain-like proteinase 2
C1312200|T116|CE|C477905|MSH|PLP-2, coronavirus|PLP-2, coronavirus
C1312200|T126|CE|C477905|MSH|PLP-2, coronavirus|PLP-2, coronavirus
C1316427|T201|MTH_LN|33964-8|LNC|SARS coronavirus Urbani ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar|SARS coronavirus Urbani ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar
C1316427|T201|LC|33964-8|LNC|SARS coronavirus Urbani RNA [Presence] in Unspecified specimen by NAA with probe detection|SARS coronavirus Urbani RNA [Presence] in Unspecified specimen by NAA with probe detection
C1316427|T201|DN|33964-8|LNC|SARS coronavirus Urbani RNA NAA+probe Ql (Unsp spec)|SARS coronavirus Urbani RNA NAA+probe Ql (Unsp spec)
C1316427|T201|LN|33964-8|LNC|SARS coronavirus Urbani RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar|SARS coronavirus Urbani RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar
C1316427|T201|OSN|33964-8|LNC|SARS-CoV Urb RNA XXX Ql NAA+probe|SARS-CoV Urb RNA XXX Ql NAA+probe
C1316428|T201|MTH_LN|33965-5|LNC|SARS coronavirus Urbani ribonucleic acid:Presence or Threshold:Point in time:Stool = Fecal:Ordinal:DNA Nucleic Acid Probe.amp.tar|SARS coronavirus Urbani ribonucleic acid:Presence or Threshold:Point in time:Stool = Fecal:Ordinal:DNA Nucleic Acid Probe.amp.tar
C1316428|T201|LC|33965-5|LNC|SARS coronavirus Urbani RNA [Presence] in Stool by NAA with probe detection|SARS coronavirus Urbani RNA [Presence] in Stool by NAA with probe detection
C1316428|T201|DN|33965-5|LNC|SARS coronavirus Urbani RNA NAA+probe Ql (Stl)|SARS coronavirus Urbani RNA NAA+probe Ql (Stl)
C1316428|T201|LN|33965-5|LNC|SARS coronavirus Urbani RNA:PrThr:Pt:Stool:Ord:Probe.amp.tar|SARS coronavirus Urbani RNA:PrThr:Pt:Stool:Ord:Probe.amp.tar
C1316428|T201|OSN|33965-5|LNC|SARS-CoV Urb RNA Stl Ql NAA+probe|SARS-CoV Urb RNA Stl Ql NAA+probe
C1316429|T201|MTH_LN|33966-3|LNC|SARS coronavirus Urbani ribonucleic acid:Presence or Threshold:Point in time:Nose (nasal passage):Ordinal:DNA Nucleic Acid Probe.amp.tar|SARS coronavirus Urbani ribonucleic acid:Presence or Threshold:Point in time:Nose (nasal passage):Ordinal:DNA Nucleic Acid Probe.amp.tar
C1316429|T201|LC|33966-3|LNC|SARS coronavirus Urbani RNA [Presence] in Nose by NAA with probe detection|SARS coronavirus Urbani RNA [Presence] in Nose by NAA with probe detection
C1316429|T201|DN|33966-3|LNC|SARS coronavirus Urbani RNA NAA+probe Ql (Nose)|SARS coronavirus Urbani RNA NAA+probe Ql (Nose)
C1316429|T201|LN|33966-3|LNC|SARS coronavirus Urbani RNA:PrThr:Pt:Nose:Ord:Probe.amp.tar|SARS coronavirus Urbani RNA:PrThr:Pt:Nose:Ord:Probe.amp.tar
C1316429|T201|OSN|33966-3|LNC|SARS-CoV Urb RNA Nose Ql NAA+probe|SARS-CoV Urb RNA Nose Ql NAA+probe
C1316430|T201|MTH_LN|33967-1|LNC|SARS coronavirus Urbani ribonucleic acid:Presence or Threshold:Point in time:Serum/Plasma:Ordinal:DNA Nucleic Acid Probe.amp.tar|SARS coronavirus Urbani ribonucleic acid:Presence or Threshold:Point in time:Serum/Plasma:Ordinal:DNA Nucleic Acid Probe.amp.tar
C1316430|T201|LC|33967-1|LNC|SARS coronavirus Urbani RNA [Presence] in Serum or Plasma by NAA with probe detection|SARS coronavirus Urbani RNA [Presence] in Serum or Plasma by NAA with probe detection
C1316430|T201|DN|33967-1|LNC|SARS coronavirus Urbani RNA NAA+probe Ql|SARS coronavirus Urbani RNA NAA+probe Ql
C1316430|T201|LN|33967-1|LNC|SARS coronavirus Urbani RNA:PrThr:Pt:Ser/Plas:Ord:Probe.amp.tar|SARS coronavirus Urbani RNA:PrThr:Pt:Ser/Plas:Ord:Probe.amp.tar
C1316430|T201|OSN|33967-1|LNC|SARS-CoV Urb RNA SerPl Ql NAA+probe|SARS-CoV Urb RNA SerPl Ql NAA+probe
C1316431|T201|LC|33968-9|LNC|SARS coronavirus Urbani Ab [Presence] in Serum by Immunoassay|SARS coronavirus Urbani Ab [Presence] in Serum by Immunoassay
C1316431|T201|DN|33968-9|LNC|SARS coronavirus Urbani Ab IA Ql (S)|SARS coronavirus Urbani Ab IA Ql (S)
C1316431|T201|LN|33968-9|LNC|SARS coronavirus Urbani Ab:PrThr:Pt:Ser:Ord:IA|SARS coronavirus Urbani Ab:PrThr:Pt:Ser:Ord:IA
C1316431|T201|MTH_LN|33968-9|LNC|SARS coronavirus Urbani Antibody:Presence or Threshold:Point in time:Serum:Ordinal:Enzyme Immunoassay|SARS coronavirus Urbani Antibody:Presence or Threshold:Point in time:Serum:Ordinal:Enzyme Immunoassay
C1316431|T201|OSN|33968-9|LNC|SARS-CoV Urb Ab Ser Ql IA|SARS-CoV Urb Ab Ser Ql IA
C1316432|T201|LC|33969-7|LNC|SARS coronavirus Urbani Ab [Units/volume] in Serum by Immunoassay|SARS coronavirus Urbani Ab [Units/volume] in Serum by Immunoassay
C1316432|T201|DN|33969-7|LNC|SARS coronavirus Urbani Ab IA Qn (S)|SARS coronavirus Urbani Ab IA Qn (S)
C1316432|T201|LN|33969-7|LNC|SARS coronavirus Urbani Ab:ACnc:Pt:Ser:Qn:IA|SARS coronavirus Urbani Ab:ACnc:Pt:Ser:Qn:IA
C1316432|T201|MTH_LN|33969-7|LNC|SARS coronavirus Urbani Antibody:Arbitrary Concentration:Point in time:Serum:Quantitative:Enzyme Immunoassay|SARS coronavirus Urbani Antibody:Arbitrary Concentration:Point in time:Serum:Quantitative:Enzyme Immunoassay
C1316432|T201|OSN|33969-7|LNC|SARS-CoV Urb Ab Ser IA-aCnc|SARS-CoV Urb Ab Ser IA-aCnc
C1316433|T201|LC|33970-5|LNC|SARS coronavirus Urbani Ab [Presence] in Serum by Immunofluorescence|SARS coronavirus Urbani Ab [Presence] in Serum by Immunofluorescence
C1316433|T201|DN|33970-5|LNC|SARS coronavirus Urbani Ab IF Ql (S)|SARS coronavirus Urbani Ab IF Ql (S)
C1316433|T201|LN|33970-5|LNC|SARS coronavirus Urbani Ab:PrThr:Pt:Ser:Ord:IF|SARS coronavirus Urbani Ab:PrThr:Pt:Ser:Ord:IF
C1316433|T201|MTH_LN|33970-5|LNC|SARS coronavirus Urbani Antibody:Presence or Threshold:Point in time:Serum:Ordinal:Immune Fluorescence|SARS coronavirus Urbani Antibody:Presence or Threshold:Point in time:Serum:Ordinal:Immune Fluorescence
C1316433|T201|OSN|33970-5|LNC|SARS-CoV Urb Ab Ser Ql IF|SARS-CoV Urb Ab Ser Ql IF
C1316434|T201|LC|33971-3|LNC|SARS coronavirus Urbani Ab [Titer] in Serum by Immunofluorescence|SARS coronavirus Urbani Ab [Titer] in Serum by Immunofluorescence
C1316434|T201|DN|33971-3|LNC|SARS coronavirus Urbani Ab IF (S) [Titer]|SARS coronavirus Urbani Ab IF (S) [Titer]
C1316434|T201|LN|33971-3|LNC|SARS coronavirus Urbani Ab:Titr:Pt:Ser:Qn:IF|SARS coronavirus Urbani Ab:Titr:Pt:Ser:Qn:IF
C1316434|T201|MTH_LN|33971-3|LNC|SARS coronavirus Urbani Antibody:Dilution Factor (Titer):Point in time:Serum:Quantitative:Immune Fluorescence|SARS coronavirus Urbani Antibody:Dilution Factor (Titer):Point in time:Serum:Quantitative:Immune Fluorescence
C1316434|T201|OSN|33971-3|LNC|SARS-CoV Urb Ab Titr Ser IF|SARS-CoV Urb Ab Titr Ser IF
C1316435|T201|LC|33972-1|LNC|SARS coronavirus Urbani Ab [Presence] in Serum|SARS coronavirus Urbani Ab [Presence] in Serum
C1316435|T201|DN|33972-1|LNC|SARS coronavirus Urbani Ab Ql (S)|SARS coronavirus Urbani Ab Ql (S)
C1316435|T201|LN|33972-1|LNC|SARS coronavirus Urbani Ab:PrThr:Pt:Ser:Ord|SARS coronavirus Urbani Ab:PrThr:Pt:Ser:Ord
C1316435|T201|MTH_LN|33972-1|LNC|SARS coronavirus Urbani Antibody:Presence or Threshold:Point in time:Serum:Ordinal|SARS coronavirus Urbani Antibody:Presence or Threshold:Point in time:Serum:Ordinal
C1316435|T201|OSN|33972-1|LNC|SARS-CoV Urb Ab Ser Ql|SARS-CoV Urb Ab Ser Ql
C1316436|T201|LC|33973-9|LNC|SARS coronavirus Urbani Ab [Units/volume] in Serum|SARS coronavirus Urbani Ab [Units/volume] in Serum
C1316436|T201|DN|33973-9|LNC|SARS coronavirus Urbani Ab Qn (S)|SARS coronavirus Urbani Ab Qn (S)
C1316436|T201|LN|33973-9|LNC|SARS coronavirus Urbani Ab:ACnc:Pt:Ser:Qn|SARS coronavirus Urbani Ab:ACnc:Pt:Ser:Qn
C1316436|T201|MTH_LN|33973-9|LNC|SARS coronavirus Urbani Antibody:Arbitrary Concentration:Point in time:Serum:Quantitative|SARS coronavirus Urbani Antibody:Arbitrary Concentration:Point in time:Serum:Quantitative
C1316436|T201|OSN|33973-9|LNC|SARS-CoV Urb Ab Ser-aCnc|SARS-CoV Urb Ab Ser-aCnc
C1316437|T201|DN|33974-7|LNC|SARS coronavirus Urbani Ab (S) [Titer]|SARS coronavirus Urbani Ab (S) [Titer]
C1316437|T201|LC|33974-7|LNC|SARS coronavirus Urbani Ab [Titer] in Serum|SARS coronavirus Urbani Ab [Titer] in Serum
C1316437|T201|LN|33974-7|LNC|SARS coronavirus Urbani Ab:Titr:Pt:Ser:Qn|SARS coronavirus Urbani Ab:Titr:Pt:Ser:Qn
C1316437|T201|MTH_LN|33974-7|LNC|SARS coronavirus Urbani Antibody:Dilution Factor (Titer):Point in time:Serum:Quantitative|SARS coronavirus Urbani Antibody:Dilution Factor (Titer):Point in time:Serum:Quantitative
C1316437|T201|OSN|33974-7|LNC|SARS-CoV Urb Ab Titr Ser|SARS-CoV Urb Ab Titr Ser
C1316438|T201|MTH_LN|33975-4|LNC|SARS coronavirus Urbani ribonucleic acid:Presence or Threshold:Point in time:Sputum:Ordinal:DNA Nucleic Acid Probe.amp.tar|SARS coronavirus Urbani ribonucleic acid:Presence or Threshold:Point in time:Sputum:Ordinal:DNA Nucleic Acid Probe.amp.tar
C1316438|T201|LC|33975-4|LNC|SARS coronavirus Urbani RNA [Presence] in Sputum by NAA with probe detection|SARS coronavirus Urbani RNA [Presence] in Sputum by NAA with probe detection
C1316438|T201|DN|33975-4|LNC|SARS coronavirus Urbani RNA NAA+probe Ql (Sput)|SARS coronavirus Urbani RNA NAA+probe Ql (Sput)
C1316438|T201|LN|33975-4|LNC|SARS coronavirus Urbani RNA:PrThr:Pt:Sputum:Ord:Probe.amp.tar|SARS coronavirus Urbani RNA:PrThr:Pt:Sputum:Ord:Probe.amp.tar
C1316438|T201|OSN|33975-4|LNC|SARS-CoV Urb RNA Spt Ql NAA+probe|SARS-CoV Urb RNA Spt Ql NAA+probe
C1317705|T116|SY|709905009|SNOMEDCT_US|Anti-Severe acute respiratory syndrome coronavirus urbani antibody|Anti-Severe acute respiratory syndrome coronavirus urbani antibody
C1317705|T129|SY|709905009|SNOMEDCT_US|Anti-Severe acute respiratory syndrome coronavirus urbani antibody|Anti-Severe acute respiratory syndrome coronavirus urbani antibody
C1317705|T116|SY|709905009|SNOMEDCT_US|Antibody to Severe acute respiratory syndrome coronavirus urbani|Antibody to Severe acute respiratory syndrome coronavirus urbani
C1317705|T129|SY|709905009|SNOMEDCT_US|Antibody to Severe acute respiratory syndrome coronavirus urbani|Antibody to Severe acute respiratory syndrome coronavirus urbani
C1317705|T116|FN|709905009|SNOMEDCT_US|Antibody to Severe acute respiratory syndrome coronavirus urbani (substance)|Antibody to Severe acute respiratory syndrome coronavirus urbani (substance)
C1317705|T129|FN|709905009|SNOMEDCT_US|Antibody to Severe acute respiratory syndrome coronavirus urbani (substance)|Antibody to Severe acute respiratory syndrome coronavirus urbani (substance)
C1317705|T116|LPN|LP39712-2|LNC|SARS coronavirus Urbani Ab|SARS coronavirus Urbani Ab
C1317705|T129|LPN|LP39712-2|LNC|SARS coronavirus Urbani Ab|SARS coronavirus Urbani Ab
C1317705|T116|CN|MTHU015801|LNC|SARS coronavirus Urbani Ab|SARS coronavirus Urbani Ab
C1317705|T129|CN|MTHU015801|LNC|SARS coronavirus Urbani Ab|SARS coronavirus Urbani Ab
C1317705|T116|SY|709905009|SNOMEDCT_US|SARS coronavirus Urbani Ab|SARS coronavirus Urbani Ab
C1317705|T129|SY|709905009|SNOMEDCT_US|SARS coronavirus Urbani Ab|SARS coronavirus Urbani Ab
C1317705|T116|MTH_CN|MTHU015801|LNC|SARS coronavirus Urbani Antibody|SARS coronavirus Urbani Antibody
C1317705|T129|MTH_CN|MTHU015801|LNC|SARS coronavirus Urbani Antibody|SARS coronavirus Urbani Antibody
C1317705|T116|PT|709905009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus urbani Ab|Severe acute respiratory syndrome coronavirus urbani Ab
C1317705|T129|PT|709905009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus urbani Ab|Severe acute respiratory syndrome coronavirus urbani Ab
C1317705|T116|SY|709905009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus urbani antibody|Severe acute respiratory syndrome coronavirus urbani antibody
C1317705|T129|SY|709905009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus urbani antibody|Severe acute respiratory syndrome coronavirus urbani antibody
C1317706|T114|MTH_CN|MTHU015799|LNC|SARS coronavirus Urbani ribonucleic acid|SARS coronavirus Urbani ribonucleic acid
C1317706|T123|MTH_CN|MTHU015799|LNC|SARS coronavirus Urbani ribonucleic acid|SARS coronavirus Urbani ribonucleic acid
C1317706|T114|PN|NOCODE|MTH|SARS coronavirus Urbani ribonucleic acid|SARS coronavirus Urbani ribonucleic acid
C1317706|T123|PN|NOCODE|MTH|SARS coronavirus Urbani ribonucleic acid|SARS coronavirus Urbani ribonucleic acid
C1317706|T114|LPN|LP39713-0|LNC|SARS coronavirus Urbani RNA|SARS coronavirus Urbani RNA
C1317706|T123|LPN|LP39713-0|LNC|SARS coronavirus Urbani RNA|SARS coronavirus Urbani RNA
C1317706|T114|CN|MTHU015799|LNC|SARS coronavirus Urbani RNA|SARS coronavirus Urbani RNA
C1317706|T123|CN|MTHU015799|LNC|SARS coronavirus Urbani RNA|SARS coronavirus Urbani RNA
C1394032|T047|PT|330006|MEDCIN|coronavirus as cause of disease classified elsewhere|coronavirus as cause of disease classified elsewhere
C1394032|T047|FN|330006|MEDCIN|coronavirus as cause of disease classified elsewhere (diagnosis)|coronavirus as cause of disease classified elsewhere (diagnosis)
C1394032|T047|AB|B97.2|ICD10CM|Coronavirus as the cause of diseases classified elsewhere|Coronavirus as the cause of diseases classified elsewhere
C1394032|T047|HT|B97.2|ICD10CM|Coronavirus as the cause of diseases classified elsewhere|Coronavirus as the cause of diseases classified elsewhere
C1394032|T047|PT|MTHU019530|ICPC2ICD10ENG|coronavirus; as cause of disease classified elsewhere|coronavirus; as cause of disease classified elsewhere
C1400736|T047|PT|MTHU038701|ICPC2ICD10ENG|infection; viral, coronavirus, as cause of disease classified elsewhere|infection; viral, coronavirus, as cause of disease classified elsewhere
C1400736|T047|PT|MTHU080923|ICPC2ICD10ENG|viral; infection, coronavirus, as cause of disease classified elsewhere|viral; infection, coronavirus, as cause of disease classified elsewhere
C1430045|T116|PCE|C087637|MSH|gene 1a protein, Coronavirus|gene 1a protein, Coronavirus
C1430045|T123|PCE|C087637|MSH|gene 1a protein, Coronavirus|gene 1a protein, Coronavirus
C1430046|T116|PCE|C087637|MSH|gene 1b protein, Coronavirus|gene 1b protein, Coronavirus
C1430046|T123|PCE|C087637|MSH|gene 1b protein, Coronavirus|gene 1b protein, Coronavirus
C1433062|T116|NM|C479931|MSH|3C-like protease, SARS coronavirus|3C-like protease, SARS coronavirus
C1433062|T126|NM|C479931|MSH|3C-like protease, SARS coronavirus|3C-like protease, SARS coronavirus
C1433062|T116|CE|C479931|MSH|3C-like protease, severe acute respiratory syndrome coronavirus|3C-like protease, severe acute respiratory syndrome coronavirus
C1433062|T126|CE|C479931|MSH|3C-like protease, severe acute respiratory syndrome coronavirus|3C-like protease, severe acute respiratory syndrome coronavirus
C1433062|T116|CE|C479931|MSH|3CL(pro) protein, SARS-CoV|3CL(pro) protein, SARS-CoV
C1433062|T126|CE|C479931|MSH|3CL(pro) protein, SARS-CoV|3CL(pro) protein, SARS-CoV
C1433062|T116|CE|C479931|MSH|M(pro) protein, SARS-CoV|M(pro) protein, SARS-CoV
C1433062|T126|CE|C479931|MSH|M(pro) protein, SARS-CoV|M(pro) protein, SARS-CoV
C1433062|T116|CE|C479931|MSH|papain-like protease, SARS coronavirus|papain-like protease, SARS coronavirus
C1433062|T126|CE|C479931|MSH|papain-like protease, SARS coronavirus|papain-like protease, SARS coronavirus
C1433062|T116|CE|C479931|MSH|PLpro, SARS-CoV|PLpro, SARS-CoV
C1433062|T126|CE|C479931|MSH|PLpro, SARS-CoV|PLpro, SARS-CoV
C1433062|T116|CE|C479931|MSH|SARS coronavirus main protease|SARS coronavirus main protease
C1433062|T126|CE|C479931|MSH|SARS coronavirus main protease|SARS coronavirus main protease
C1433062|T116|CE|C479931|MSH|SARS-CoV main protease|SARS-CoV main protease
C1433062|T126|CE|C479931|MSH|SARS-CoV main protease|SARS-CoV main protease
C1439114|T116|CE|C412015|MSH|HCoV helicase protein, Human coronavirus 229E|HCoV helicase protein, Human coronavirus 229E
C1439114|T126|CE|C412015|MSH|HCoV helicase protein, Human coronavirus 229E|HCoV helicase protein, Human coronavirus 229E
C1439114|T116|CE|C412015|MSH|HCoV SF1 RNA helicase protein, Human coronavirus 229E|HCoV SF1 RNA helicase protein, Human coronavirus 229E
C1439114|T126|CE|C412015|MSH|HCoV SF1 RNA helicase protein, Human coronavirus 229E|HCoV SF1 RNA helicase protein, Human coronavirus 229E
C1439114|T116|CE|C412015|MSH|p66(HEL) protein, Human coronavirus 229E|p66(HEL) protein, Human coronavirus 229E
C1439114|T126|CE|C412015|MSH|p66(HEL) protein, Human coronavirus 229E|p66(HEL) protein, Human coronavirus 229E
C1439114|T116|NM|C412015|MSH|p66HEL protein, Human coronavirus 229E|p66HEL protein, Human coronavirus 229E
C1439114|T126|NM|C412015|MSH|p66HEL protein, Human coronavirus 229E|p66HEL protein, Human coronavirus 229E
C1443246|T047|SY|408688009|SNOMEDCT_US|Healthcare associated SARS|Healthcare associated SARS
C1443246|T047|PT|408688009|SNOMEDCT_US|Healthcare associated severe acute respiratory syndrome|Healthcare associated severe acute respiratory syndrome
C1443246|T047|FN|408688009|SNOMEDCT_US|Healthcare associated severe acute respiratory syndrome (disorder)|Healthcare associated severe acute respiratory syndrome (disorder)
C1447200|T116|PCE|C078034|MSH|mmCGM1 protein, Coronavirus|mmCGM1 protein, Coronavirus
C1447200|T192|PCE|C078034|MSH|mmCGM1 protein, Coronavirus|mmCGM1 protein, Coronavirus
C1447201|T116|PCE|C078034|MSH|mmCGM2 protein, Coronavirus|mmCGM2 protein, Coronavirus
C1447201|T192|PCE|C078034|MSH|mmCGM2 protein, Coronavirus|mmCGM2 protein, Coronavirus
C1450568|T116|CE|C483945|MSH|nonstructural protein 9, SARS-CoV|nonstructural protein 9, SARS-CoV
C1450568|T123|CE|C483945|MSH|nonstructural protein 9, SARS-CoV|nonstructural protein 9, SARS-CoV
C1450568|T116|NM|C483945|MSH|nsp9 protein, SARS virus|nsp9 protein, SARS virus
C1450568|T123|NM|C483945|MSH|nsp9 protein, SARS virus|nsp9 protein, SARS virus
C1452735|T116|CE|C487105|MSH|3a protein, SARS-CoV|3a protein, SARS-CoV
C1452735|T123|CE|C487105|MSH|3a protein, SARS-CoV|3a protein, SARS-CoV
C1452735|T116|NM|C487105|MSH|3a protein, severe acute respiratory syndrome coronavirus|3a protein, severe acute respiratory syndrome coronavirus
C1452735|T123|NM|C487105|MSH|3a protein, severe acute respiratory syndrome coronavirus|3a protein, severe acute respiratory syndrome coronavirus
C1454704|T116|CE|C488151|MSH|7a protein, SARS virus|7a protein, SARS virus
C1454704|T123|CE|C488151|MSH|7a protein, SARS virus|7a protein, SARS virus
C1454704|T116|CE|C488151|MSH|7a protein, severe acute respiratory syndrome coronavirus|7a protein, severe acute respiratory syndrome coronavirus
C1454704|T123|CE|C488151|MSH|7a protein, severe acute respiratory syndrome coronavirus|7a protein, severe acute respiratory syndrome coronavirus
C1454704|T116|CE|C488151|MSH|accessory protein 7a, SARS virus|accessory protein 7a, SARS virus
C1454704|T123|CE|C488151|MSH|accessory protein 7a, SARS virus|accessory protein 7a, SARS virus
C1454704|T116|CE|C488151|MSH|ORF7a protein, SARS virus|ORF7a protein, SARS virus
C1454704|T123|CE|C488151|MSH|ORF7a protein, SARS virus|ORF7a protein, SARS virus
C1454704|T116|CE|C488151|MSH|ORF8 protein, SARS virus|ORF8 protein, SARS virus
C1454704|T123|CE|C488151|MSH|ORF8 protein, SARS virus|ORF8 protein, SARS virus
C1454704|T116|NM|C488151|MSH|sars7a protein, SARS virus|sars7a protein, SARS virus
C1454704|T123|NM|C488151|MSH|sars7a protein, SARS virus|sars7a protein, SARS virus
C1454704|T116|CE|C488151|MSH|U122 protein, SARS virus|U122 protein, SARS virus
C1454704|T123|CE|C488151|MSH|U122 protein, SARS virus|U122 protein, SARS virus
C1454704|T116|CE|C488151|MSH|X4 protein, SARS virus|X4 protein, SARS virus
C1454704|T123|CE|C488151|MSH|X4 protein, SARS virus|X4 protein, SARS virus
C1478824|T005|LA|LA26149-7|LNC|Coronavirus NL63|Coronavirus NL63
C1478824|T005|MH|D058957|MSH|Coronavirus NL63, Human|Coronavirus NL63, Human
C1478824|T005|ET|D058957|MSH|HCoV-NL63|HCoV-NL63
C1478824|T005|LPN|LP35709-2|LNC|Human coronavirus NL63|Human coronavirus NL63
C1478824|T005|PT|417818007|SNOMEDCT_US|Human coronavirus NL63|Human coronavirus NL63
C1478824|T005|PN|NOCODE|MTH|Human coronavirus NL63|Human coronavirus NL63
C1478824|T005|ET|D058957|MSH|Human Coronavirus NL63|Human Coronavirus NL63
C1478824|T005|FN|417818007|SNOMEDCT_US|Human coronavirus NL63 (organism)|Human coronavirus NL63 (organism)
C1478824|T005|PM|D058957|MSH|NL63, Human Coronavirus|NL63, Human Coronavirus
C1499881|T005|PT|415493006|SNOMEDCT_US|SARS coronavirus TWS|SARS coronavirus TWS
C1499881|T005|OF|415493006|SNOMEDCT_US|SARS coronavirus TWS (organism)|SARS coronavirus TWS (organism)
C1499881|T005|SY|415493006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TWS|Severe acute respiratory syndrome (SARS) coronavirus TWS
C1499881|T005|OF|415493006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TWS (organism)|Severe acute respiratory syndrome (SARS) coronavirus TWS (organism)
C1499881|T005|SY|415493006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TWS|Severe acute respiratory syndrome coronavirus TWS
C1499881|T005|FN|415493006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TWS (organism)|Severe acute respiratory syndrome coronavirus TWS (organism)
C1499882|T005|PT|415467004|SNOMEDCT_US|SARS coronavirus TW-HP1|SARS coronavirus TW-HP1
C1499882|T005|OF|415467004|SNOMEDCT_US|SARS coronavirus TW-HP1 (organism)|SARS coronavirus TW-HP1 (organism)
C1499882|T005|SY|415467004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-HP1|Severe acute respiratory syndrome (SARS) coronavirus TW-HP1
C1499882|T005|OF|415467004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-HP1 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW-HP1 (organism)
C1499882|T005|SY|415467004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-HP1|Severe acute respiratory syndrome coronavirus TW-HP1
C1499882|T005|FN|415467004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-HP1 (organism)|Severe acute respiratory syndrome coronavirus TW-HP1 (organism)
C1499883|T005|PT|415468009|SNOMEDCT_US|SARS coronavirus TW-HP2|SARS coronavirus TW-HP2
C1499883|T005|OF|415468009|SNOMEDCT_US|SARS coronavirus TW-HP2 (organism)|SARS coronavirus TW-HP2 (organism)
C1499883|T005|SY|415468009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-HP2|Severe acute respiratory syndrome (SARS) coronavirus TW-HP2
C1499883|T005|OF|415468009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-HP2 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW-HP2 (organism)
C1499883|T005|SY|415468009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-HP2|Severe acute respiratory syndrome coronavirus TW-HP2
C1499883|T005|FN|415468009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-HP2 (organism)|Severe acute respiratory syndrome coronavirus TW-HP2 (organism)
C1499884|T005|PT|415469001|SNOMEDCT_US|SARS coronavirus TW-HP3|SARS coronavirus TW-HP3
C1499884|T005|OF|415469001|SNOMEDCT_US|SARS coronavirus TW-HP3 (organism)|SARS coronavirus TW-HP3 (organism)
C1499884|T005|SY|415469001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-HP3|Severe acute respiratory syndrome (SARS) coronavirus TW-HP3
C1499884|T005|OF|415469001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-HP3 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW-HP3 (organism)
C1499884|T005|SY|415469001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-HP3|Severe acute respiratory syndrome coronavirus TW-HP3
C1499884|T005|FN|415469001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-HP3 (organism)|Severe acute respiratory syndrome coronavirus TW-HP3 (organism)
C1499885|T005|PT|415470000|SNOMEDCT_US|SARS coronavirus TW-HP4|SARS coronavirus TW-HP4
C1499885|T005|OF|415470000|SNOMEDCT_US|SARS coronavirus TW-HP4 (organism)|SARS coronavirus TW-HP4 (organism)
C1499885|T005|SY|415470000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-HP4|Severe acute respiratory syndrome (SARS) coronavirus TW-HP4
C1499885|T005|OF|415470000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-HP4 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW-HP4 (organism)
C1499885|T005|SY|415470000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-HP4|Severe acute respiratory syndrome coronavirus TW-HP4
C1499885|T005|FN|415470000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-HP4 (organism)|Severe acute respiratory syndrome coronavirus TW-HP4 (organism)
C1499886|T005|PT|415471001|SNOMEDCT_US|SARS coronavirus TW-JC2|SARS coronavirus TW-JC2
C1499886|T005|OF|415471001|SNOMEDCT_US|SARS coronavirus TW-JC2 (organism)|SARS coronavirus TW-JC2 (organism)
C1499886|T005|SY|415471001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-JC2|Severe acute respiratory syndrome (SARS) coronavirus TW-JC2
C1499886|T005|OF|415471001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-JC2 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW-JC2 (organism)
C1499886|T005|SY|415471001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-JC2|Severe acute respiratory syndrome coronavirus TW-JC2
C1499886|T005|FN|415471001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-JC2 (organism)|Severe acute respiratory syndrome coronavirus TW-JC2 (organism)
C1499887|T005|PT|415472008|SNOMEDCT_US|SARS coronavirus TW-KC1|SARS coronavirus TW-KC1
C1499887|T005|PN|NOCODE|MTH|SARS coronavirus TW-KC1|SARS coronavirus TW-KC1
C1499887|T005|OF|415472008|SNOMEDCT_US|SARS coronavirus TW-KC1 (organism)|SARS coronavirus TW-KC1 (organism)
C1499887|T005|SY|415472008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-KC1|Severe acute respiratory syndrome (SARS) coronavirus TW-KC1
C1499887|T005|OF|415472008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-KC1 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW-KC1 (organism)
C1499887|T005|SY|415472008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-KC1|Severe acute respiratory syndrome coronavirus TW-KC1
C1499887|T005|FN|415472008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-KC1 (organism)|Severe acute respiratory syndrome coronavirus TW-KC1 (organism)
C1499889|T005|PT|415463000|SNOMEDCT_US|SARS coronavirus TW-GD1|SARS coronavirus TW-GD1
C1499889|T005|OF|415463000|SNOMEDCT_US|SARS coronavirus TW-GD1 (organism)|SARS coronavirus TW-GD1 (organism)
C1499889|T005|SY|415463000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-GD1|Severe acute respiratory syndrome (SARS) coronavirus TW-GD1
C1499889|T005|OF|415463000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-GD1 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW-GD1 (organism)
C1499889|T005|SY|415463000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-GD1|Severe acute respiratory syndrome coronavirus TW-GD1
C1499889|T005|FN|415463000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-GD1 (organism)|Severe acute respiratory syndrome coronavirus TW-GD1 (organism)
C1499890|T005|PT|415464006|SNOMEDCT_US|SARS coronavirus TW-GD2|SARS coronavirus TW-GD2
C1499890|T005|OF|415464006|SNOMEDCT_US|SARS coronavirus TW-GD2 (organism)|SARS coronavirus TW-GD2 (organism)
C1499890|T005|SY|415464006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-GD2|Severe acute respiratory syndrome (SARS) coronavirus TW-GD2
C1499890|T005|OF|415464006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-GD2 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW-GD2 (organism)
C1499890|T005|SY|415464006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-GD2|Severe acute respiratory syndrome coronavirus TW-GD2
C1499890|T005|FN|415464006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-GD2 (organism)|Severe acute respiratory syndrome coronavirus TW-GD2 (organism)
C1499891|T005|PT|415465007|SNOMEDCT_US|SARS coronavirus TW-GD3|SARS coronavirus TW-GD3
C1499891|T005|OF|415465007|SNOMEDCT_US|SARS coronavirus TW-GD3 (organism)|SARS coronavirus TW-GD3 (organism)
C1499891|T005|SY|415465007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-GD3|Severe acute respiratory syndrome (SARS) coronavirus TW-GD3
C1499891|T005|OF|415465007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-GD3 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW-GD3 (organism)
C1499891|T005|SY|415465007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-GD3|Severe acute respiratory syndrome coronavirus TW-GD3
C1499891|T005|FN|415465007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-GD3 (organism)|Severe acute respiratory syndrome coronavirus TW-GD3 (organism)
C1499893|T005|PT|415466008|SNOMEDCT_US|SARS coronavirus TW-GD5|SARS coronavirus TW-GD5
C1499893|T005|OF|415466008|SNOMEDCT_US|SARS coronavirus TW-GD5 (organism)|SARS coronavirus TW-GD5 (organism)
C1499893|T005|SY|415466008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-GD5|Severe acute respiratory syndrome (SARS) coronavirus TW-GD5
C1499893|T005|OF|415466008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-GD5 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW-GD5 (organism)
C1499893|T005|SY|415466008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-GD5|Severe acute respiratory syndrome coronavirus TW-GD5
C1499893|T005|FN|415466008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-GD5 (organism)|Severe acute respiratory syndrome coronavirus TW-GD5 (organism)
C1499897|T005|PT|415475005|SNOMEDCT_US|SARS coronavirus TW-YM4|SARS coronavirus TW-YM4
C1499897|T005|OF|415475005|SNOMEDCT_US|SARS coronavirus TW-YM4 (organism)|SARS coronavirus TW-YM4 (organism)
C1499897|T005|SY|415475005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-YM4|Severe acute respiratory syndrome (SARS) coronavirus TW-YM4
C1499897|T005|OF|415475005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-YM4 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW-YM4 (organism)
C1499897|T005|SY|415475005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-YM4|Severe acute respiratory syndrome coronavirus TW-YM4
C1499897|T005|FN|415475005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-YM4 (organism)|Severe acute respiratory syndrome coronavirus TW-YM4 (organism)
C1499898|T005|PT|415474009|SNOMEDCT_US|SARS coronavirus TW-PH1|SARS coronavirus TW-PH1
C1499898|T005|OF|415474009|SNOMEDCT_US|SARS coronavirus TW-PH1 (organism)|SARS coronavirus TW-PH1 (organism)
C1499898|T005|SY|415474009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-PH1|Severe acute respiratory syndrome (SARS) coronavirus TW-PH1
C1499898|T005|OF|415474009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-PH1 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW-PH1 (organism)
C1499898|T005|SY|415474009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-PH1|Severe acute respiratory syndrome coronavirus TW-PH1
C1499898|T005|FN|415474009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-PH1 (organism)|Severe acute respiratory syndrome coronavirus TW-PH1 (organism)
C1519126|T044|PT|C39229|NCI_BioC|SARS Coronavirus Protease|SARS Coronavirus Protease
C1519126|T044|PT|C39229|NCI|SARS Coronavirus Protease Pathway|SARS Coronavirus Protease Pathway
C1531863|T005|PT|415444001|SNOMEDCT_US|SARS coronavirus Sin850|SARS coronavirus Sin850
C1531863|T005|OF|415444001|SNOMEDCT_US|SARS coronavirus Sin850 (organism)|SARS coronavirus Sin850 (organism)
C1531863|T005|SY|415444001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin850|Severe acute respiratory syndrome (SARS) coronavirus Sin850
C1531863|T005|OF|415444001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin850 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Sin850 (organism)
C1531863|T005|SY|415444001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin850|Severe acute respiratory syndrome coronavirus Sin850
C1531863|T005|FN|415444001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin850 (organism)|Severe acute respiratory syndrome coronavirus Sin850 (organism)
C1531864|T005|PT|415445000|SNOMEDCT_US|SARS coronavirus Sin852|SARS coronavirus Sin852
C1531864|T005|OF|415445000|SNOMEDCT_US|SARS coronavirus Sin852 (organism)|SARS coronavirus Sin852 (organism)
C1531864|T005|SY|415445000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin852|Severe acute respiratory syndrome (SARS) coronavirus Sin852
C1531864|T005|OF|415445000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin852 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Sin852 (organism)
C1531864|T005|SY|415445000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin852|Severe acute respiratory syndrome coronavirus Sin852
C1531864|T005|FN|415445000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin852 (organism)|Severe acute respiratory syndrome coronavirus Sin852 (organism)
C1531865|T005|PT|415446004|SNOMEDCT_US|SARS coronavirus Sin_WNV|SARS coronavirus Sin_WNV
C1531865|T005|OF|415446004|SNOMEDCT_US|SARS coronavirus Sin_WNV (organism)|SARS coronavirus Sin_WNV (organism)
C1531865|T005|SY|415446004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin_WNV|Severe acute respiratory syndrome (SARS) coronavirus Sin_WNV
C1531865|T005|OF|415446004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin_WNV (organism)|Severe acute respiratory syndrome (SARS) coronavirus Sin_WNV (organism)
C1531865|T005|SY|415446004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin_WNV|Severe acute respiratory syndrome coronavirus Sin_WNV
C1531865|T005|FN|415446004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin_WNV (organism)|Severe acute respiratory syndrome coronavirus Sin_WNV (organism)
C1531866|T005|PT|415447008|SNOMEDCT_US|SARS coronavirus SinP1|SARS coronavirus SinP1
C1531866|T005|OF|415447008|SNOMEDCT_US|SARS coronavirus SinP1 (organism)|SARS coronavirus SinP1 (organism)
C1531866|T005|SY|415447008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus SinP1|Severe acute respiratory syndrome (SARS) coronavirus SinP1
C1531866|T005|OF|415447008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus SinP1 (organism)|Severe acute respiratory syndrome (SARS) coronavirus SinP1 (organism)
C1531866|T005|SY|415447008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus SinP1|Severe acute respiratory syndrome coronavirus SinP1
C1531866|T005|FN|415447008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus SinP1 (organism)|Severe acute respiratory syndrome coronavirus SinP1 (organism)
C1531867|T005|PT|415448003|SNOMEDCT_US|SARS coronavirus SinP2|SARS coronavirus SinP2
C1531867|T005|OF|415448003|SNOMEDCT_US|SARS coronavirus SinP2 (organism)|SARS coronavirus SinP2 (organism)
C1531867|T005|SY|415448003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus SinP2|Severe acute respiratory syndrome (SARS) coronavirus SinP2
C1531867|T005|OF|415448003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus SinP2 (organism)|Severe acute respiratory syndrome (SARS) coronavirus SinP2 (organism)
C1531867|T005|SY|415448003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus SinP2|Severe acute respiratory syndrome coronavirus SinP2
C1531867|T005|FN|415448003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus SinP2 (organism)|Severe acute respiratory syndrome coronavirus SinP2 (organism)
C1531868|T005|PT|415449006|SNOMEDCT_US|SARS coronavirus SinP3|SARS coronavirus SinP3
C1531868|T005|OF|415449006|SNOMEDCT_US|SARS coronavirus SinP3 (organism)|SARS coronavirus SinP3 (organism)
C1531868|T005|SY|415449006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus SinP3|Severe acute respiratory syndrome (SARS) coronavirus SinP3
C1531868|T005|OF|415449006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus SinP3 (organism)|Severe acute respiratory syndrome (SARS) coronavirus SinP3 (organism)
C1531868|T005|SY|415449006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus SinP3|Severe acute respiratory syndrome coronavirus SinP3
C1531868|T005|FN|415449006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus SinP3 (organism)|Severe acute respiratory syndrome coronavirus SinP3 (organism)
C1531869|T005|PT|415450006|SNOMEDCT_US|SARS coronavirus SinP4|SARS coronavirus SinP4
C1531869|T005|OF|415450006|SNOMEDCT_US|SARS coronavirus SinP4 (organism)|SARS coronavirus SinP4 (organism)
C1531869|T005|SY|415450006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus SinP4|Severe acute respiratory syndrome (SARS) coronavirus SinP4
C1531869|T005|OF|415450006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus SinP4 (organism)|Severe acute respiratory syndrome (SARS) coronavirus SinP4 (organism)
C1531869|T005|SY|415450006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus SinP4|Severe acute respiratory syndrome coronavirus SinP4
C1531869|T005|FN|415450006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus SinP4 (organism)|Severe acute respiratory syndrome coronavirus SinP4 (organism)
C1531870|T005|PT|415451005|SNOMEDCT_US|SARS coronavirus SinP5|SARS coronavirus SinP5
C1531870|T005|OF|415451005|SNOMEDCT_US|SARS coronavirus SinP5 (organism)|SARS coronavirus SinP5 (organism)
C1531870|T005|SY|415451005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus SinP5|Severe acute respiratory syndrome (SARS) coronavirus SinP5
C1531870|T005|OF|415451005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus SinP5 (organism)|Severe acute respiratory syndrome (SARS) coronavirus SinP5 (organism)
C1531870|T005|SY|415451005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus SinP5|Severe acute respiratory syndrome coronavirus SinP5
C1531870|T005|FN|415451005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus SinP5 (organism)|Severe acute respiratory syndrome coronavirus SinP5 (organism)
C1531946|T005|PT|415499005|SNOMEDCT_US|SARS coronavirus ZS-C|SARS coronavirus ZS-C
C1531946|T005|OF|415499005|SNOMEDCT_US|SARS coronavirus ZS-C (organism)|SARS coronavirus ZS-C (organism)
C1531946|T005|SY|415499005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus ZS-C|Severe acute respiratory syndrome (SARS) coronavirus ZS-C
C1531946|T005|OF|415499005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus ZS-C (organism)|Severe acute respiratory syndrome (SARS) coronavirus ZS-C (organism)
C1531946|T005|SY|415499005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus ZS-C|Severe acute respiratory syndrome coronavirus ZS-C
C1531946|T005|FN|415499005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus ZS-C (organism)|Severe acute respiratory syndrome coronavirus ZS-C (organism)
C1532052|T005|PT|415452003|SNOMEDCT_US|SARS coronavirus SoD|SARS coronavirus SoD
C1532052|T005|OF|415452003|SNOMEDCT_US|SARS coronavirus SoD (organism)|SARS coronavirus SoD (organism)
C1532052|T005|SY|415452003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus SoD|Severe acute respiratory syndrome (SARS) coronavirus SoD
C1532052|T005|OF|415452003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus SoD (organism)|Severe acute respiratory syndrome (SARS) coronavirus SoD (organism)
C1532052|T005|SY|415452003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus SoD|Severe acute respiratory syndrome coronavirus SoD
C1532052|T005|FN|415452003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus SoD (organism)|Severe acute respiratory syndrome coronavirus SoD (organism)
C1532053|T005|PT|415453008|SNOMEDCT_US|SARS coronavirus SZ1|SARS coronavirus SZ1
C1532053|T005|OF|415453008|SNOMEDCT_US|SARS coronavirus SZ1 (organism)|SARS coronavirus SZ1 (organism)
C1532053|T005|SY|415453008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus SZ1|Severe acute respiratory syndrome (SARS) coronavirus SZ1
C1532053|T005|OF|415453008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus SZ1 (organism)|Severe acute respiratory syndrome (SARS) coronavirus SZ1 (organism)
C1532053|T005|SY|415453008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus SZ1|Severe acute respiratory syndrome coronavirus SZ1
C1532053|T005|FN|415453008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus SZ1 (organism)|Severe acute respiratory syndrome coronavirus SZ1 (organism)
C1532054|T005|PT|415454002|SNOMEDCT_US|SARS coronavirus SZ13|SARS coronavirus SZ13
C1532054|T005|OF|415454002|SNOMEDCT_US|SARS coronavirus SZ13 (organism)|SARS coronavirus SZ13 (organism)
C1532054|T005|SY|415454002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus SZ13|Severe acute respiratory syndrome (SARS) coronavirus SZ13
C1532054|T005|OF|415454002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus SZ13 (organism)|Severe acute respiratory syndrome (SARS) coronavirus SZ13 (organism)
C1532054|T005|SY|415454002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus SZ13|Severe acute respiratory syndrome coronavirus SZ13
C1532054|T005|FN|415454002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus SZ13 (organism)|Severe acute respiratory syndrome coronavirus SZ13 (organism)
C1532055|T005|PT|415455001|SNOMEDCT_US|SARS coronavirus SZ16|SARS coronavirus SZ16
C1532055|T005|OF|415455001|SNOMEDCT_US|SARS coronavirus SZ16 (organism)|SARS coronavirus SZ16 (organism)
C1532055|T005|SY|415455001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus SZ16|Severe acute respiratory syndrome (SARS) coronavirus SZ16
C1532055|T005|OF|415455001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus SZ16 (organism)|Severe acute respiratory syndrome (SARS) coronavirus SZ16 (organism)
C1532055|T005|SY|415455001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus SZ16|Severe acute respiratory syndrome coronavirus SZ16
C1532055|T005|FN|415455001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus SZ16 (organism)|Severe acute respiratory syndrome coronavirus SZ16 (organism)
C1532056|T005|PT|415456000|SNOMEDCT_US|SARS coronavirus SZ3|SARS coronavirus SZ3
C1532056|T005|OF|415456000|SNOMEDCT_US|SARS coronavirus SZ3 (organism)|SARS coronavirus SZ3 (organism)
C1532056|T005|SY|415456000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus SZ3|Severe acute respiratory syndrome (SARS) coronavirus SZ3
C1532056|T005|OF|415456000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus SZ3 (organism)|Severe acute respiratory syndrome (SARS) coronavirus SZ3 (organism)
C1532056|T005|SY|415456000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus SZ3|Severe acute respiratory syndrome coronavirus SZ3
C1532056|T005|FN|415456000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus SZ3 (organism)|Severe acute respiratory syndrome coronavirus SZ3 (organism)
C1532057|T005|PT|415457009|SNOMEDCT_US|SARS coronavirus Taiwan|SARS coronavirus Taiwan
C1532057|T005|OF|415457009|SNOMEDCT_US|SARS coronavirus Taiwan (organism)|SARS coronavirus Taiwan (organism)
C1532057|T005|SY|415457009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Taiwan|Severe acute respiratory syndrome (SARS) coronavirus Taiwan
C1532057|T005|OF|415457009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Taiwan (organism)|Severe acute respiratory syndrome (SARS) coronavirus Taiwan (organism)
C1532057|T005|SY|415457009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Taiwan|Severe acute respiratory syndrome coronavirus Taiwan
C1532057|T005|FN|415457009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Taiwan (organism)|Severe acute respiratory syndrome coronavirus Taiwan (organism)
C1532058|T005|PT|415458004|SNOMEDCT_US|SARS coronavirus Taiwan TC1|SARS coronavirus Taiwan TC1
C1532058|T005|OF|415458004|SNOMEDCT_US|SARS coronavirus Taiwan TC1 (organism)|SARS coronavirus Taiwan TC1 (organism)
C1532058|T005|SY|415458004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Taiwan TC1|Severe acute respiratory syndrome (SARS) coronavirus Taiwan TC1
C1532058|T005|OF|415458004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Taiwan TC1 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Taiwan TC1 (organism)
C1532058|T005|SY|415458004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Taiwan TC1|Severe acute respiratory syndrome coronavirus Taiwan TC1
C1532058|T005|FN|415458004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Taiwan TC1 (organism)|Severe acute respiratory syndrome coronavirus Taiwan TC1 (organism)
C1532059|T005|PT|415459007|SNOMEDCT_US|SARS coronavirus Taiwan TC2|SARS coronavirus Taiwan TC2
C1532059|T005|OF|415459007|SNOMEDCT_US|SARS coronavirus Taiwan TC2 (organism)|SARS coronavirus Taiwan TC2 (organism)
C1532059|T005|SY|415459007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Taiwan TC2|Severe acute respiratory syndrome (SARS) coronavirus Taiwan TC2
C1532059|T005|OF|415459007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Taiwan TC2 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Taiwan TC2 (organism)
C1532059|T005|SY|415459007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Taiwan TC2|Severe acute respiratory syndrome coronavirus Taiwan TC2
C1532059|T005|FN|415459007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Taiwan TC2 (organism)|Severe acute respiratory syndrome coronavirus Taiwan TC2 (organism)
C1532060|T005|PT|415460002|SNOMEDCT_US|SARS coronavirus Taiwan TC3|SARS coronavirus Taiwan TC3
C1532060|T005|OF|415460002|SNOMEDCT_US|SARS coronavirus Taiwan TC3 (organism)|SARS coronavirus Taiwan TC3 (organism)
C1532060|T005|SY|415460002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Taiwan TC3|Severe acute respiratory syndrome (SARS) coronavirus Taiwan TC3
C1532060|T005|OF|415460002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Taiwan TC3 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Taiwan TC3 (organism)
C1532060|T005|SY|415460002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Taiwan TC3|Severe acute respiratory syndrome coronavirus Taiwan TC3
C1532060|T005|FN|415460002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Taiwan TC3 (organism)|Severe acute respiratory syndrome coronavirus Taiwan TC3 (organism)
C1532061|T005|PT|415461003|SNOMEDCT_US|SARS coronavirus Tor2|SARS coronavirus Tor2
C1532061|T005|OF|415461003|SNOMEDCT_US|SARS coronavirus Tor2 (organism)|SARS coronavirus Tor2 (organism)
C1532061|T005|SY|415461003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Tor2|Severe acute respiratory syndrome (SARS) coronavirus Tor2
C1532061|T005|OF|415461003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Tor2 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Tor2 (organism)
C1532061|T005|SY|415461003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Tor2|Severe acute respiratory syndrome coronavirus Tor2
C1532061|T005|FN|415461003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Tor2 (organism)|Severe acute respiratory syndrome coronavirus Tor2 (organism)
C1532062|T005|PT|415473003|SNOMEDCT_US|SARS coronavirus TW-KC2|SARS coronavirus TW-KC2
C1532062|T005|PN|NOCODE|MTH|SARS coronavirus TW-KC2|SARS coronavirus TW-KC2
C1532062|T005|OF|415473003|SNOMEDCT_US|SARS coronavirus TW-KC2 (organism)|SARS coronavirus TW-KC2 (organism)
C1532062|T005|SY|415473003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-KC2|Severe acute respiratory syndrome (SARS) coronavirus TW-KC2
C1532062|T005|OF|415473003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW-KC2 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW-KC2 (organism)
C1532062|T005|SY|415473003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-KC2|Severe acute respiratory syndrome coronavirus TW-KC2
C1532062|T005|FN|415473003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW-KC2 (organism)|Severe acute respiratory syndrome coronavirus TW-KC2 (organism)
C1532063|T005|PT|415476006|SNOMEDCT_US|SARS coronavirus TW1|SARS coronavirus TW1
C1532063|T005|OF|415476006|SNOMEDCT_US|SARS coronavirus TW1 (organism)|SARS coronavirus TW1 (organism)
C1532063|T005|SY|415476006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW1|Severe acute respiratory syndrome (SARS) coronavirus TW1
C1532063|T005|OF|415476006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW1 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW1 (organism)
C1532063|T005|SY|415476006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW1|Severe acute respiratory syndrome coronavirus TW1
C1532063|T005|FN|415476006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW1 (organism)|Severe acute respiratory syndrome coronavirus TW1 (organism)
C1532064|T005|PT|415477002|SNOMEDCT_US|SARS coronavirus TW10|SARS coronavirus TW10
C1532064|T005|OF|415477002|SNOMEDCT_US|SARS coronavirus TW10 (organism)|SARS coronavirus TW10 (organism)
C1532064|T005|SY|415477002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW10|Severe acute respiratory syndrome (SARS) coronavirus TW10
C1532064|T005|OF|415477002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW10 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW10 (organism)
C1532064|T005|SY|415477002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW10|Severe acute respiratory syndrome coronavirus TW10
C1532064|T005|FN|415477002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW10 (organism)|Severe acute respiratory syndrome coronavirus TW10 (organism)
C1532065|T005|PT|415478007|SNOMEDCT_US|SARS coronavirus TW11|SARS coronavirus TW11
C1532065|T005|OF|415478007|SNOMEDCT_US|SARS coronavirus TW11 (organism)|SARS coronavirus TW11 (organism)
C1532065|T005|SY|415478007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW11|Severe acute respiratory syndrome (SARS) coronavirus TW11
C1532065|T005|OF|415478007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW11 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW11 (organism)
C1532065|T005|SY|415478007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW11|Severe acute respiratory syndrome coronavirus TW11
C1532065|T005|FN|415478007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW11 (organism)|Severe acute respiratory syndrome coronavirus TW11 (organism)
C1532066|T005|PT|415479004|SNOMEDCT_US|SARS coronavirus TW2|SARS coronavirus TW2
C1532066|T005|OF|415479004|SNOMEDCT_US|SARS coronavirus TW2 (organism)|SARS coronavirus TW2 (organism)
C1532066|T005|SY|415479004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW2|Severe acute respiratory syndrome (SARS) coronavirus TW2
C1532066|T005|OF|415479004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW2 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW2 (organism)
C1532066|T005|SY|415479004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW2|Severe acute respiratory syndrome coronavirus TW2
C1532066|T005|FN|415479004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW2 (organism)|Severe acute respiratory syndrome coronavirus TW2 (organism)
C1532067|T005|PT|415480001|SNOMEDCT_US|SARS coronavirus TW3|SARS coronavirus TW3
C1532067|T005|OF|415480001|SNOMEDCT_US|SARS coronavirus TW3 (organism)|SARS coronavirus TW3 (organism)
C1532067|T005|SY|415480001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW3|Severe acute respiratory syndrome (SARS) coronavirus TW3
C1532067|T005|OF|415480001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW3 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW3 (organism)
C1532067|T005|SY|415480001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW3|Severe acute respiratory syndrome coronavirus TW3
C1532067|T005|FN|415480001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW3 (organism)|Severe acute respiratory syndrome coronavirus TW3 (organism)
C1532068|T005|PT|415481002|SNOMEDCT_US|SARS coronavirus TW4|SARS coronavirus TW4
C1532068|T005|OF|415481002|SNOMEDCT_US|SARS coronavirus TW4 (organism)|SARS coronavirus TW4 (organism)
C1532068|T005|SY|415481002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW4|Severe acute respiratory syndrome (SARS) coronavirus TW4
C1532068|T005|OF|415481002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW4 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW4 (organism)
C1532068|T005|SY|415481002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW4|Severe acute respiratory syndrome coronavirus TW4
C1532068|T005|FN|415481002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW4 (organism)|Severe acute respiratory syndrome coronavirus TW4 (organism)
C1532069|T005|PT|415482009|SNOMEDCT_US|SARS coronavirus TW5|SARS coronavirus TW5
C1532069|T005|OF|415482009|SNOMEDCT_US|SARS coronavirus TW5 (organism)|SARS coronavirus TW5 (organism)
C1532069|T005|SY|415482009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW5|Severe acute respiratory syndrome (SARS) coronavirus TW5
C1532069|T005|OF|415482009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW5 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW5 (organism)
C1532069|T005|SY|415482009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW5|Severe acute respiratory syndrome coronavirus TW5
C1532069|T005|FN|415482009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW5 (organism)|Severe acute respiratory syndrome coronavirus TW5 (organism)
C1532070|T005|PT|415483004|SNOMEDCT_US|SARS coronavirus TW6|SARS coronavirus TW6
C1532070|T005|OF|415483004|SNOMEDCT_US|SARS coronavirus TW6 (organism)|SARS coronavirus TW6 (organism)
C1532070|T005|SY|415483004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW6|Severe acute respiratory syndrome (SARS) coronavirus TW6
C1532070|T005|OF|415483004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW6 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW6 (organism)
C1532070|T005|SY|415483004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW6|Severe acute respiratory syndrome coronavirus TW6
C1532070|T005|FN|415483004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW6 (organism)|Severe acute respiratory syndrome coronavirus TW6 (organism)
C1532071|T005|PT|415484005|SNOMEDCT_US|SARS coronavirus TW7|SARS coronavirus TW7
C1532071|T005|OF|415484005|SNOMEDCT_US|SARS coronavirus TW7 (organism)|SARS coronavirus TW7 (organism)
C1532071|T005|SY|415484005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW7|Severe acute respiratory syndrome (SARS) coronavirus TW7
C1532071|T005|OF|415484005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW7 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW7 (organism)
C1532071|T005|SY|415484005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW7|Severe acute respiratory syndrome coronavirus TW7
C1532071|T005|FN|415484005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW7 (organism)|Severe acute respiratory syndrome coronavirus TW7 (organism)
C1532072|T005|PT|415485006|SNOMEDCT_US|SARS coronavirus TW8|SARS coronavirus TW8
C1532072|T005|OF|415485006|SNOMEDCT_US|SARS coronavirus TW8 (organism)|SARS coronavirus TW8 (organism)
C1532072|T005|SY|415485006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW8|Severe acute respiratory syndrome (SARS) coronavirus TW8
C1532072|T005|OF|415485006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW8 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW8 (organism)
C1532072|T005|SY|415485006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW8|Severe acute respiratory syndrome coronavirus TW8
C1532072|T005|FN|415485006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW8 (organism)|Severe acute respiratory syndrome coronavirus TW8 (organism)
C1532073|T005|PT|415486007|SNOMEDCT_US|SARS coronavirus TW9|SARS coronavirus TW9
C1532073|T005|OF|415486007|SNOMEDCT_US|SARS coronavirus TW9 (organism)|SARS coronavirus TW9 (organism)
C1532073|T005|SY|415486007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW9|Severe acute respiratory syndrome (SARS) coronavirus TW9
C1532073|T005|OF|415486007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW9 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW9 (organism)
C1532073|T005|SY|415486007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW9|Severe acute respiratory syndrome coronavirus TW9
C1532073|T005|FN|415486007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW9 (organism)|Severe acute respiratory syndrome coronavirus TW9 (organism)
C1532074|T005|PT|415487003|SNOMEDCT_US|SARS coronavirus TWC|SARS coronavirus TWC
C1532074|T005|OF|415487003|SNOMEDCT_US|SARS coronavirus TWC (organism)|SARS coronavirus TWC (organism)
C1532074|T005|SY|415487003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TWC|Severe acute respiratory syndrome (SARS) coronavirus TWC
C1532074|T005|OF|415487003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TWC (organism)|Severe acute respiratory syndrome (SARS) coronavirus TWC (organism)
C1532074|T005|SY|415487003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TWC|Severe acute respiratory syndrome coronavirus TWC
C1532074|T005|FN|415487003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TWC (organism)|Severe acute respiratory syndrome coronavirus TWC (organism)
C1532075|T005|PT|415488008|SNOMEDCT_US|SARS coronavirus TWC2|SARS coronavirus TWC2
C1532075|T005|OF|415488008|SNOMEDCT_US|SARS coronavirus TWC2 (organism)|SARS coronavirus TWC2 (organism)
C1532075|T005|SY|415488008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TWC2|Severe acute respiratory syndrome (SARS) coronavirus TWC2
C1532075|T005|OF|415488008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TWC2 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TWC2 (organism)
C1532075|T005|SY|415488008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TWC2|Severe acute respiratory syndrome coronavirus TWC2
C1532075|T005|FN|415488008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TWC2 (organism)|Severe acute respiratory syndrome coronavirus TWC2 (organism)
C1532076|T005|PT|415489000|SNOMEDCT_US|SARS coronavirus TWC3|SARS coronavirus TWC3
C1532076|T005|OF|415489000|SNOMEDCT_US|SARS coronavirus TWC3 (organism)|SARS coronavirus TWC3 (organism)
C1532076|T005|SY|415489000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TWC3|Severe acute respiratory syndrome (SARS) coronavirus TWC3
C1532076|T005|OF|415489000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TWC3 (organism)|Severe acute respiratory syndrome (SARS) coronavirus TWC3 (organism)
C1532076|T005|SY|415489000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TWC3|Severe acute respiratory syndrome coronavirus TWC3
C1532076|T005|FN|415489000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TWC3 (organism)|Severe acute respiratory syndrome coronavirus TWC3 (organism)
C1532077|T005|PT|415490009|SNOMEDCT_US|SARS coronavirus TWH|SARS coronavirus TWH
C1532077|T005|OF|415490009|SNOMEDCT_US|SARS coronavirus TWH (organism)|SARS coronavirus TWH (organism)
C1532077|T005|SY|415490009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TWH|Severe acute respiratory syndrome (SARS) coronavirus TWH
C1532077|T005|OF|415490009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TWH (organism)|Severe acute respiratory syndrome (SARS) coronavirus TWH (organism)
C1532077|T005|SY|415490009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TWH|Severe acute respiratory syndrome coronavirus TWH
C1532077|T005|FN|415490009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TWH (organism)|Severe acute respiratory syndrome coronavirus TWH (organism)
C1532078|T005|PT|415491008|SNOMEDCT_US|SARS coronavirus TWJ|SARS coronavirus TWJ
C1532078|T005|OF|415491008|SNOMEDCT_US|SARS coronavirus TWJ (organism)|SARS coronavirus TWJ (organism)
C1532078|T005|SY|415491008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TWJ|Severe acute respiratory syndrome (SARS) coronavirus TWJ
C1532078|T005|OF|415491008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TWJ (organism)|Severe acute respiratory syndrome (SARS) coronavirus TWJ (organism)
C1532078|T005|SY|415491008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TWJ|Severe acute respiratory syndrome coronavirus TWJ
C1532078|T005|FN|415491008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TWJ (organism)|Severe acute respiratory syndrome coronavirus TWJ (organism)
C1532079|T005|PT|415492001|SNOMEDCT_US|SARS coronavirus TWK|SARS coronavirus TWK
C1532079|T005|OF|415492001|SNOMEDCT_US|SARS coronavirus TWK (organism)|SARS coronavirus TWK (organism)
C1532079|T005|SY|415492001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TWK|Severe acute respiratory syndrome (SARS) coronavirus TWK
C1532079|T005|OF|415492001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TWK (organism)|Severe acute respiratory syndrome (SARS) coronavirus TWK (organism)
C1532079|T005|SY|415492001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TWK|Severe acute respiratory syndrome coronavirus TWK
C1532079|T005|FN|415492001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TWK (organism)|Severe acute respiratory syndrome coronavirus TWK (organism)
C1532080|T005|PT|415494000|SNOMEDCT_US|SARS coronavirus TWY|SARS coronavirus TWY
C1532080|T005|OF|415494000|SNOMEDCT_US|SARS coronavirus TWY (organism)|SARS coronavirus TWY (organism)
C1532080|T005|SY|415494000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TWY|Severe acute respiratory syndrome (SARS) coronavirus TWY
C1532080|T005|OF|415494000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TWY (organism)|Severe acute respiratory syndrome (SARS) coronavirus TWY (organism)
C1532080|T005|SY|415494000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TWY|Severe acute respiratory syndrome coronavirus TWY
C1532080|T005|FN|415494000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TWY (organism)|Severe acute respiratory syndrome coronavirus TWY (organism)
C1532081|T005|PT|415496003|SNOMEDCT_US|SARS coronavirus Vietnam|SARS coronavirus Vietnam
C1532081|T005|OF|415496003|SNOMEDCT_US|SARS coronavirus Vietnam (organism)|SARS coronavirus Vietnam (organism)
C1532081|T005|SY|415496003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Vietnam|Severe acute respiratory syndrome (SARS) coronavirus Vietnam
C1532081|T005|OF|415496003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Vietnam (organism)|Severe acute respiratory syndrome (SARS) coronavirus Vietnam (organism)
C1532081|T005|SY|415496003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Vietnam|Severe acute respiratory syndrome coronavirus Vietnam
C1532081|T005|FN|415496003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Vietnam (organism)|Severe acute respiratory syndrome coronavirus Vietnam (organism)
C1532082|T005|PT|415497007|SNOMEDCT_US|SARS coronavirus WHU|SARS coronavirus WHU
C1532082|T005|OF|415497007|SNOMEDCT_US|SARS coronavirus WHU (organism)|SARS coronavirus WHU (organism)
C1532082|T005|SY|415497007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus WHU|Severe acute respiratory syndrome (SARS) coronavirus WHU
C1532082|T005|OF|415497007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus WHU (organism)|Severe acute respiratory syndrome (SARS) coronavirus WHU (organism)
C1532082|T005|SY|415497007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus WHU|Severe acute respiratory syndrome coronavirus WHU
C1532082|T005|FN|415497007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus WHU (organism)|Severe acute respiratory syndrome coronavirus WHU (organism)
C1532083|T005|PT|415498002|SNOMEDCT_US|SARS coronavirus ZS-B|SARS coronavirus ZS-B
C1532083|T005|OF|415498002|SNOMEDCT_US|SARS coronavirus ZS-B (organism)|SARS coronavirus ZS-B (organism)
C1532083|T005|SY|415498002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus ZS-B|Severe acute respiratory syndrome (SARS) coronavirus ZS-B
C1532083|T005|OF|415498002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus ZS-B (organism)|Severe acute respiratory syndrome (SARS) coronavirus ZS-B (organism)
C1532083|T005|SY|415498002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus ZS-B|Severe acute respiratory syndrome coronavirus ZS-B
C1532083|T005|FN|415498002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus ZS-B (organism)|Severe acute respiratory syndrome coronavirus ZS-B (organism)
C1532720|T005|PT|415391009|SNOMEDCT_US|SARS coronavirus HGZ8L1-B|SARS coronavirus HGZ8L1-B
C1532720|T005|OF|415391009|SNOMEDCT_US|SARS coronavirus HGZ8L1-B (organism)|SARS coronavirus HGZ8L1-B (organism)
C1532720|T005|SY|415391009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HGZ8L1-B|Severe acute respiratory syndrome (SARS) coronavirus HGZ8L1-B
C1532720|T005|OF|415391009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HGZ8L1-B (organism)|Severe acute respiratory syndrome (SARS) coronavirus HGZ8L1-B (organism)
C1532720|T005|SY|415391009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HGZ8L1-B|Severe acute respiratory syndrome coronavirus HGZ8L1-B
C1532720|T005|FN|415391009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HGZ8L1-B (organism)|Severe acute respiratory syndrome coronavirus HGZ8L1-B (organism)
C1532721|T005|PT|415392002|SNOMEDCT_US|SARS coronavirus HGZ8L2|SARS coronavirus HGZ8L2
C1532721|T005|OF|415392002|SNOMEDCT_US|SARS coronavirus HGZ8L2 (organism)|SARS coronavirus HGZ8L2 (organism)
C1532721|T005|SY|415392002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HGZ8L2|Severe acute respiratory syndrome (SARS) coronavirus HGZ8L2
C1532721|T005|OF|415392002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HGZ8L2 (organism)|Severe acute respiratory syndrome (SARS) coronavirus HGZ8L2 (organism)
C1532721|T005|SY|415392002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HGZ8L2|Severe acute respiratory syndrome coronavirus HGZ8L2
C1532721|T005|FN|415392002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HGZ8L2 (organism)|Severe acute respiratory syndrome coronavirus HGZ8L2 (organism)
C1532722|T005|PT|415393007|SNOMEDCT_US|SARS coronavirus HKU-36871|SARS coronavirus HKU-36871
C1532722|T005|OF|415393007|SNOMEDCT_US|SARS coronavirus HKU-36871 (organism)|SARS coronavirus HKU-36871 (organism)
C1532722|T005|SY|415393007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HKU-36871|Severe acute respiratory syndrome (SARS) coronavirus HKU-36871
C1532722|T005|OF|415393007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HKU-36871 (organism)|Severe acute respiratory syndrome (SARS) coronavirus HKU-36871 (organism)
C1532722|T005|SY|415393007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HKU-36871|Severe acute respiratory syndrome coronavirus HKU-36871
C1532722|T005|FN|415393007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HKU-36871 (organism)|Severe acute respiratory syndrome coronavirus HKU-36871 (organism)
C1532723|T005|PT|415394001|SNOMEDCT_US|SARS coronavirus HKU-39849|SARS coronavirus HKU-39849
C1532723|T005|OF|415394001|SNOMEDCT_US|SARS coronavirus HKU-39849 (organism)|SARS coronavirus HKU-39849 (organism)
C1532723|T005|SY|415394001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HKU-39849|Severe acute respiratory syndrome (SARS) coronavirus HKU-39849
C1532723|T005|OF|415394001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HKU-39849 (organism)|Severe acute respiratory syndrome (SARS) coronavirus HKU-39849 (organism)
C1532723|T005|SY|415394001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HKU-39849|Severe acute respiratory syndrome coronavirus HKU-39849
C1532723|T005|FN|415394001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HKU-39849 (organism)|Severe acute respiratory syndrome coronavirus HKU-39849 (organism)
C1532724|T005|PT|415395000|SNOMEDCT_US|SARS coronavirus HKU-65806|SARS coronavirus HKU-65806
C1532724|T005|OF|415395000|SNOMEDCT_US|SARS coronavirus HKU-65806 (organism)|SARS coronavirus HKU-65806 (organism)
C1532724|T005|SY|415395000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HKU-65806|Severe acute respiratory syndrome (SARS) coronavirus HKU-65806
C1532724|T005|OF|415395000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HKU-65806 (organism)|Severe acute respiratory syndrome (SARS) coronavirus HKU-65806 (organism)
C1532724|T005|SY|415395000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HKU-65806|Severe acute respiratory syndrome coronavirus HKU-65806
C1532724|T005|FN|415395000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HKU-65806 (organism)|Severe acute respiratory syndrome coronavirus HKU-65806 (organism)
C1532791|T005|PT|415361004|SNOMEDCT_US|SARS coronavirus AS|SARS coronavirus AS
C1532791|T005|OF|415361004|SNOMEDCT_US|SARS coronavirus AS (organism)|SARS coronavirus AS (organism)
C1532791|T005|SY|415361004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus AS|Severe acute respiratory syndrome (SARS) coronavirus AS
C1532791|T005|OF|415361004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus AS (organism)|Severe acute respiratory syndrome (SARS) coronavirus AS (organism)
C1532791|T005|SY|415361004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus AS|Severe acute respiratory syndrome coronavirus AS
C1532791|T005|FN|415361004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus AS (organism)|Severe acute respiratory syndrome coronavirus AS (organism)
C1532792|T005|PT|415362006|SNOMEDCT_US|SARS coronavirus BJ01|SARS coronavirus BJ01
C1532792|T005|OF|415362006|SNOMEDCT_US|SARS coronavirus BJ01 (organism)|SARS coronavirus BJ01 (organism)
C1532792|T005|SY|415362006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus BJ01|Severe acute respiratory syndrome (SARS) coronavirus BJ01
C1532792|T005|OF|415362006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus BJ01 (organism)|Severe acute respiratory syndrome (SARS) coronavirus BJ01 (organism)
C1532792|T005|SY|415362006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus BJ01|Severe acute respiratory syndrome coronavirus BJ01
C1532792|T005|FN|415362006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus BJ01 (organism)|Severe acute respiratory syndrome coronavirus BJ01 (organism)
C1532793|T005|PT|415363001|SNOMEDCT_US|SARS coronavirus BJ02|SARS coronavirus BJ02
C1532793|T005|OF|415363001|SNOMEDCT_US|SARS coronavirus BJ02 (organism)|SARS coronavirus BJ02 (organism)
C1532793|T005|SY|415363001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus BJ02|Severe acute respiratory syndrome (SARS) coronavirus BJ02
C1532793|T005|OF|415363001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus BJ02 (organism)|Severe acute respiratory syndrome (SARS) coronavirus BJ02 (organism)
C1532793|T005|SY|415363001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus BJ02|Severe acute respiratory syndrome coronavirus BJ02
C1532793|T005|FN|415363001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus BJ02 (organism)|Severe acute respiratory syndrome coronavirus BJ02 (organism)
C1532794|T005|PT|415364007|SNOMEDCT_US|SARS coronavirus BJ03|SARS coronavirus BJ03
C1532794|T005|OF|415364007|SNOMEDCT_US|SARS coronavirus BJ03 (organism)|SARS coronavirus BJ03 (organism)
C1532794|T005|SY|415364007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus BJ03|Severe acute respiratory syndrome (SARS) coronavirus BJ03
C1532794|T005|OF|415364007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus BJ03 (organism)|Severe acute respiratory syndrome (SARS) coronavirus BJ03 (organism)
C1532794|T005|SY|415364007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus BJ03|Severe acute respiratory syndrome coronavirus BJ03
C1532794|T005|FN|415364007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus BJ03 (organism)|Severe acute respiratory syndrome coronavirus BJ03 (organism)
C1532795|T005|PT|415365008|SNOMEDCT_US|SARS coronavirus BJ04|SARS coronavirus BJ04
C1532795|T005|OF|415365008|SNOMEDCT_US|SARS coronavirus BJ04 (organism)|SARS coronavirus BJ04 (organism)
C1532795|T005|SY|415365008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus BJ04|Severe acute respiratory syndrome (SARS) coronavirus BJ04
C1532795|T005|OF|415365008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus BJ04 (organism)|Severe acute respiratory syndrome (SARS) coronavirus BJ04 (organism)
C1532795|T005|SY|415365008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus BJ04|Severe acute respiratory syndrome coronavirus BJ04
C1532795|T005|FN|415365008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus BJ04 (organism)|Severe acute respiratory syndrome coronavirus BJ04 (organism)
C1532796|T005|PT|415366009|SNOMEDCT_US|SARS coronavirus BJ2232|SARS coronavirus BJ2232
C1532796|T005|OF|415366009|SNOMEDCT_US|SARS coronavirus BJ2232 (organism)|SARS coronavirus BJ2232 (organism)
C1532796|T005|SY|415366009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus BJ2232|Severe acute respiratory syndrome (SARS) coronavirus BJ2232
C1532796|T005|OF|415366009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus BJ2232 (organism)|Severe acute respiratory syndrome (SARS) coronavirus BJ2232 (organism)
C1532796|T005|SY|415366009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus BJ2232|Severe acute respiratory syndrome coronavirus BJ2232
C1532796|T005|FN|415366009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus BJ2232 (organism)|Severe acute respiratory syndrome coronavirus BJ2232 (organism)
C1532797|T005|PT|415367000|SNOMEDCT_US|SARS coronavirus BJ302|SARS coronavirus BJ302
C1532797|T005|OF|415367000|SNOMEDCT_US|SARS coronavirus BJ302 (organism)|SARS coronavirus BJ302 (organism)
C1532797|T005|SY|415367000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus BJ302|Severe acute respiratory syndrome (SARS) coronavirus BJ302
C1532797|T005|OF|415367000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus BJ302 (organism)|Severe acute respiratory syndrome (SARS) coronavirus BJ302 (organism)
C1532797|T005|SY|415367000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus BJ302|Severe acute respiratory syndrome coronavirus BJ302
C1532797|T005|FN|415367000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus BJ302 (organism)|Severe acute respiratory syndrome coronavirus BJ302 (organism)
C1532798|T005|PT|415368005|SNOMEDCT_US|SARS coronavirus CUHK-AG01|SARS coronavirus CUHK-AG01
C1532798|T005|OF|415368005|SNOMEDCT_US|SARS coronavirus CUHK-AG01 (organism)|SARS coronavirus CUHK-AG01 (organism)
C1532798|T005|SY|415368005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus CUHK-AG01|Severe acute respiratory syndrome (SARS) coronavirus CUHK-AG01
C1532798|T005|OF|415368005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus CUHK-AG01 (organism)|Severe acute respiratory syndrome (SARS) coronavirus CUHK-AG01 (organism)
C1532798|T005|SY|415368005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus CUHK-AG01|Severe acute respiratory syndrome coronavirus CUHK-AG01
C1532798|T005|FN|415368005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus CUHK-AG01 (organism)|Severe acute respiratory syndrome coronavirus CUHK-AG01 (organism)
C1532799|T005|PT|415369002|SNOMEDCT_US|SARS coronavirus CUHK-AG02|SARS coronavirus CUHK-AG02
C1532799|T005|OF|415369002|SNOMEDCT_US|SARS coronavirus CUHK-AG02 (organism)|SARS coronavirus CUHK-AG02 (organism)
C1532799|T005|SY|415369002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus CUHK-AG02|Severe acute respiratory syndrome (SARS) coronavirus CUHK-AG02
C1532799|T005|OF|415369002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus CUHK-AG02 (organism)|Severe acute respiratory syndrome (SARS) coronavirus CUHK-AG02 (organism)
C1532799|T005|SY|415369002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus CUHK-AG02|Severe acute respiratory syndrome coronavirus CUHK-AG02
C1532799|T005|FN|415369002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus CUHK-AG02 (organism)|Severe acute respiratory syndrome coronavirus CUHK-AG02 (organism)
C1532800|T005|PT|415370001|SNOMEDCT_US|SARS coronavirus CUHK-AG03|SARS coronavirus CUHK-AG03
C1532800|T005|OF|415370001|SNOMEDCT_US|SARS coronavirus CUHK-AG03 (organism)|SARS coronavirus CUHK-AG03 (organism)
C1532800|T005|SY|415370001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus CUHK-AG03|Severe acute respiratory syndrome (SARS) coronavirus CUHK-AG03
C1532800|T005|OF|415370001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus CUHK-AG03 (organism)|Severe acute respiratory syndrome (SARS) coronavirus CUHK-AG03 (organism)
C1532800|T005|SY|415370001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus CUHK-AG03|Severe acute respiratory syndrome coronavirus CUHK-AG03
C1532800|T005|FN|415370001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus CUHK-AG03 (organism)|Severe acute respiratory syndrome coronavirus CUHK-AG03 (organism)
C1532801|T005|PT|415371002|SNOMEDCT_US|SARS coronavirus CUHK-L2|SARS coronavirus CUHK-L2
C1532801|T005|OF|415371002|SNOMEDCT_US|SARS coronavirus CUHK-L2 (organism)|SARS coronavirus CUHK-L2 (organism)
C1532801|T005|SY|415371002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus CUHK-L2|Severe acute respiratory syndrome (SARS) coronavirus CUHK-L2
C1532801|T005|OF|415371002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus CUHK-L2 (organism)|Severe acute respiratory syndrome (SARS) coronavirus CUHK-L2 (organism)
C1532801|T005|SY|415371002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus CUHK-L2|Severe acute respiratory syndrome coronavirus CUHK-L2
C1532801|T005|FN|415371002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus CUHK-L2 (organism)|Severe acute respiratory syndrome coronavirus CUHK-L2 (organism)
C1532802|T005|PT|415372009|SNOMEDCT_US|SARS coronavirus CUHK-Su10|SARS coronavirus CUHK-Su10
C1532802|T005|OF|415372009|SNOMEDCT_US|SARS coronavirus CUHK-Su10 (organism)|SARS coronavirus CUHK-Su10 (organism)
C1532802|T005|SY|415372009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus CUHK-Su10|Severe acute respiratory syndrome (SARS) coronavirus CUHK-Su10
C1532802|T005|OF|415372009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus CUHK-Su10 (organism)|Severe acute respiratory syndrome (SARS) coronavirus CUHK-Su10 (organism)
C1532802|T005|SY|415372009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus CUHK-Su10|Severe acute respiratory syndrome coronavirus CUHK-Su10
C1532802|T005|FN|415372009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus CUHK-Su10 (organism)|Severe acute respiratory syndrome coronavirus CUHK-Su10 (organism)
C1532803|T005|PT|415373004|SNOMEDCT_US|SARS coronavirus CUHK-W1|SARS coronavirus CUHK-W1
C1532803|T005|OF|415373004|SNOMEDCT_US|SARS coronavirus CUHK-W1 (organism)|SARS coronavirus CUHK-W1 (organism)
C1532803|T005|SY|415373004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus CUHK-W1|Severe acute respiratory syndrome (SARS) coronavirus CUHK-W1
C1532803|T005|OF|415373004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus CUHK-W1 (organism)|Severe acute respiratory syndrome (SARS) coronavirus CUHK-W1 (organism)
C1532803|T005|SY|415373004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus CUHK-W1|Severe acute respiratory syndrome coronavirus CUHK-W1
C1532803|T005|FN|415373004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus CUHK-W1 (organism)|Severe acute respiratory syndrome coronavirus CUHK-W1 (organism)
C1532804|T005|PT|415374005|SNOMEDCT_US|SARS coronavirus cw037|SARS coronavirus cw037
C1532804|T005|OF|415374005|SNOMEDCT_US|SARS coronavirus cw037 (organism)|SARS coronavirus cw037 (organism)
C1532804|T005|SY|415374005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus cw037|Severe acute respiratory syndrome (SARS) coronavirus cw037
C1532804|T005|OF|415374005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus cw037 (organism)|Severe acute respiratory syndrome (SARS) coronavirus cw037 (organism)
C1532804|T005|SY|415374005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus cw037|Severe acute respiratory syndrome coronavirus cw037
C1532804|T005|FN|415374005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus cw037 (organism)|Severe acute respiratory syndrome coronavirus cw037 (organism)
C1532805|T005|PT|415375006|SNOMEDCT_US|SARS coronavirus cw049|SARS coronavirus cw049
C1532805|T005|OF|415375006|SNOMEDCT_US|SARS coronavirus cw049 (organism)|SARS coronavirus cw049 (organism)
C1532805|T005|SY|415375006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus cw049|Severe acute respiratory syndrome (SARS) coronavirus cw049
C1532805|T005|OF|415375006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus cw049 (organism)|Severe acute respiratory syndrome (SARS) coronavirus cw049 (organism)
C1532805|T005|SY|415375006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus cw049|Severe acute respiratory syndrome coronavirus cw049
C1532805|T005|FN|415375006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus cw049 (organism)|Severe acute respiratory syndrome coronavirus cw049 (organism)
C1532806|T005|PT|415376007|SNOMEDCT_US|SARS coronavirus FRA|SARS coronavirus FRA
C1532806|T005|OF|415376007|SNOMEDCT_US|SARS coronavirus FRA (organism)|SARS coronavirus FRA (organism)
C1532806|T005|SY|415376007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus FRA|Severe acute respiratory syndrome (SARS) coronavirus FRA
C1532806|T005|OF|415376007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus FRA (organism)|Severe acute respiratory syndrome (SARS) coronavirus FRA (organism)
C1532806|T005|SY|415376007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus FRA|Severe acute respiratory syndrome coronavirus FRA
C1532806|T005|FN|415376007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus FRA (organism)|Severe acute respiratory syndrome coronavirus FRA (organism)
C1532807|T005|PT|415377003|SNOMEDCT_US|SARS coronavirus Frankfurt 1|SARS coronavirus Frankfurt 1
C1532807|T005|OF|415377003|SNOMEDCT_US|SARS coronavirus Frankfurt 1 (organism)|SARS coronavirus Frankfurt 1 (organism)
C1532807|T005|SY|415377003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Frankfurt 1|Severe acute respiratory syndrome (SARS) coronavirus Frankfurt 1
C1532807|T005|OF|415377003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Frankfurt 1 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Frankfurt 1 (organism)
C1532807|T005|SY|415377003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Frankfurt 1|Severe acute respiratory syndrome coronavirus Frankfurt 1
C1532807|T005|FN|415377003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Frankfurt 1 (organism)|Severe acute respiratory syndrome coronavirus Frankfurt 1 (organism)
C1532808|T005|PT|415378008|SNOMEDCT_US|SARS coronavirus GD01|SARS coronavirus GD01
C1532808|T005|OF|415378008|SNOMEDCT_US|SARS coronavirus GD01 (organism)|SARS coronavirus GD01 (organism)
C1532808|T005|SY|415378008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GD01|Severe acute respiratory syndrome (SARS) coronavirus GD01
C1532808|T005|OF|415378008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GD01 (organism)|Severe acute respiratory syndrome (SARS) coronavirus GD01 (organism)
C1532808|T005|SY|415378008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GD01|Severe acute respiratory syndrome coronavirus GD01
C1532808|T005|FN|415378008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GD01 (organism)|Severe acute respiratory syndrome coronavirus GD01 (organism)
C1532809|T005|PT|415379000|SNOMEDCT_US|SARS coronavirus GD03T0013|SARS coronavirus GD03T0013
C1532809|T005|OF|415379000|SNOMEDCT_US|SARS coronavirus GD03T0013 (organism)|SARS coronavirus GD03T0013 (organism)
C1532809|T005|SY|415379000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GD03T0013|Severe acute respiratory syndrome (SARS) coronavirus GD03T0013
C1532809|T005|OF|415379000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GD03T0013 (organism)|Severe acute respiratory syndrome (SARS) coronavirus GD03T0013 (organism)
C1532809|T005|SY|415379000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GD03T0013|Severe acute respiratory syndrome coronavirus GD03T0013
C1532809|T005|FN|415379000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GD03T0013 (organism)|Severe acute respiratory syndrome coronavirus GD03T0013 (organism)
C1532810|T005|PT|415380002|SNOMEDCT_US|SARS coronavirus GD69|SARS coronavirus GD69
C1532810|T005|OF|415380002|SNOMEDCT_US|SARS coronavirus GD69 (organism)|SARS coronavirus GD69 (organism)
C1532810|T005|SY|415380002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GD69|Severe acute respiratory syndrome (SARS) coronavirus GD69
C1532810|T005|OF|415380002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GD69 (organism)|Severe acute respiratory syndrome (SARS) coronavirus GD69 (organism)
C1532810|T005|SY|415380002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GD69|Severe acute respiratory syndrome coronavirus GD69
C1532810|T005|FN|415380002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GD69 (organism)|Severe acute respiratory syndrome coronavirus GD69 (organism)
C1532811|T005|PT|415381003|SNOMEDCT_US|SARS coronavirus GZ-A|SARS coronavirus GZ-A
C1532811|T005|OF|415381003|SNOMEDCT_US|SARS coronavirus GZ-A (organism)|SARS coronavirus GZ-A (organism)
C1532811|T005|SY|415381003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GZ-A|Severe acute respiratory syndrome (SARS) coronavirus GZ-A
C1532811|T005|OF|415381003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GZ-A (organism)|Severe acute respiratory syndrome (SARS) coronavirus GZ-A (organism)
C1532811|T005|SY|415381003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GZ-A|Severe acute respiratory syndrome coronavirus GZ-A
C1532811|T005|FN|415381003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GZ-A (organism)|Severe acute respiratory syndrome coronavirus GZ-A (organism)
C1532812|T005|PT|415382005|SNOMEDCT_US|SARS coronavirus GZ-B|SARS coronavirus GZ-B
C1532812|T005|OF|415382005|SNOMEDCT_US|SARS coronavirus GZ-B (organism)|SARS coronavirus GZ-B (organism)
C1532812|T005|SY|415382005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GZ-B|Severe acute respiratory syndrome (SARS) coronavirus GZ-B
C1532812|T005|OF|415382005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GZ-B (organism)|Severe acute respiratory syndrome (SARS) coronavirus GZ-B (organism)
C1532812|T005|SY|415382005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GZ-B|Severe acute respiratory syndrome coronavirus GZ-B
C1532812|T005|FN|415382005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GZ-B (organism)|Severe acute respiratory syndrome coronavirus GZ-B (organism)
C1532813|T005|PT|415383000|SNOMEDCT_US|SARS coronavirus GZ-C|SARS coronavirus GZ-C
C1532813|T005|OF|415383000|SNOMEDCT_US|SARS coronavirus GZ-C (organism)|SARS coronavirus GZ-C (organism)
C1532813|T005|SY|415383000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GZ-C|Severe acute respiratory syndrome (SARS) coronavirus GZ-C
C1532813|T005|OF|415383000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GZ-C (organism)|Severe acute respiratory syndrome (SARS) coronavirus GZ-C (organism)
C1532813|T005|SY|415383000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GZ-C|Severe acute respiratory syndrome coronavirus GZ-C
C1532813|T005|FN|415383000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GZ-C (organism)|Severe acute respiratory syndrome coronavirus GZ-C (organism)
C1532814|T005|PT|415384006|SNOMEDCT_US|SARS coronavirus GZ-D|SARS coronavirus GZ-D
C1532814|T005|OF|415384006|SNOMEDCT_US|SARS coronavirus GZ-D (organism)|SARS coronavirus GZ-D (organism)
C1532814|T005|SY|415384006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GZ-D|Severe acute respiratory syndrome (SARS) coronavirus GZ-D
C1532814|T005|OF|415384006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GZ-D (organism)|Severe acute respiratory syndrome (SARS) coronavirus GZ-D (organism)
C1532814|T005|SY|415384006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GZ-D|Severe acute respiratory syndrome coronavirus GZ-D
C1532814|T005|FN|415384006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GZ-D (organism)|Severe acute respiratory syndrome coronavirus GZ-D (organism)
C1532815|T005|PT|415385007|SNOMEDCT_US|SARS coronavirus GZ02|SARS coronavirus GZ02
C1532815|T005|OF|415385007|SNOMEDCT_US|SARS coronavirus GZ02 (organism)|SARS coronavirus GZ02 (organism)
C1532815|T005|SY|415385007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GZ02|Severe acute respiratory syndrome (SARS) coronavirus GZ02
C1532815|T005|OF|415385007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GZ02 (organism)|Severe acute respiratory syndrome (SARS) coronavirus GZ02 (organism)
C1532815|T005|SY|415385007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GZ02|Severe acute respiratory syndrome coronavirus GZ02
C1532815|T005|FN|415385007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GZ02 (organism)|Severe acute respiratory syndrome coronavirus GZ02 (organism)
C1532816|T005|PT|415386008|SNOMEDCT_US|SARS coronavirus GZ43|SARS coronavirus GZ43
C1532816|T005|OF|415386008|SNOMEDCT_US|SARS coronavirus GZ43 (organism)|SARS coronavirus GZ43 (organism)
C1532816|T005|SY|415386008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GZ43|Severe acute respiratory syndrome (SARS) coronavirus GZ43
C1532816|T005|OF|415386008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GZ43 (organism)|Severe acute respiratory syndrome (SARS) coronavirus GZ43 (organism)
C1532816|T005|SY|415386008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GZ43|Severe acute respiratory syndrome coronavirus GZ43
C1532816|T005|FN|415386008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GZ43 (organism)|Severe acute respiratory syndrome coronavirus GZ43 (organism)
C1532817|T005|PT|415387004|SNOMEDCT_US|SARS coronavirus GZ50|SARS coronavirus GZ50
C1532817|T005|OF|415387004|SNOMEDCT_US|SARS coronavirus GZ50 (organism)|SARS coronavirus GZ50 (organism)
C1532817|T005|SY|415387004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GZ50|Severe acute respiratory syndrome (SARS) coronavirus GZ50
C1532817|T005|OF|415387004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GZ50 (organism)|Severe acute respiratory syndrome (SARS) coronavirus GZ50 (organism)
C1532817|T005|SY|415387004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GZ50|Severe acute respiratory syndrome coronavirus GZ50
C1532817|T005|FN|415387004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GZ50 (organism)|Severe acute respiratory syndrome coronavirus GZ50 (organism)
C1532818|T005|PT|415388009|SNOMEDCT_US|SARS coronavirus GZ60|SARS coronavirus GZ60
C1532818|T005|OF|415388009|SNOMEDCT_US|SARS coronavirus GZ60 (organism)|SARS coronavirus GZ60 (organism)
C1532818|T005|SY|415388009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GZ60|Severe acute respiratory syndrome (SARS) coronavirus GZ60
C1532818|T005|OF|415388009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus GZ60 (organism)|Severe acute respiratory syndrome (SARS) coronavirus GZ60 (organism)
C1532818|T005|SY|415388009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GZ60|Severe acute respiratory syndrome coronavirus GZ60
C1532818|T005|FN|415388009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus GZ60 (organism)|Severe acute respiratory syndrome coronavirus GZ60 (organism)
C1532819|T005|PT|415389001|SNOMEDCT_US|SARS coronavirus HB|SARS coronavirus HB
C1532819|T005|OF|415389001|SNOMEDCT_US|SARS coronavirus HB (organism)|SARS coronavirus HB (organism)
C1532819|T005|SY|415389001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HB|Severe acute respiratory syndrome (SARS) coronavirus HB
C1532819|T005|OF|415389001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HB (organism)|Severe acute respiratory syndrome (SARS) coronavirus HB (organism)
C1532819|T005|SY|415389001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HB|Severe acute respiratory syndrome coronavirus HB
C1532819|T005|FN|415389001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HB (organism)|Severe acute respiratory syndrome coronavirus HB (organism)
C1532820|T005|PT|415390005|SNOMEDCT_US|SARS coronavirus HGZ8L1-A|SARS coronavirus HGZ8L1-A
C1532820|T005|OF|415390005|SNOMEDCT_US|SARS coronavirus HGZ8L1-A (organism)|SARS coronavirus HGZ8L1-A (organism)
C1532820|T005|SY|415390005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HGZ8L1-A|Severe acute respiratory syndrome (SARS) coronavirus HGZ8L1-A
C1532820|T005|OF|415390005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HGZ8L1-A (organism)|Severe acute respiratory syndrome (SARS) coronavirus HGZ8L1-A (organism)
C1532820|T005|SY|415390005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HGZ8L1-A|Severe acute respiratory syndrome coronavirus HGZ8L1-A
C1532820|T005|FN|415390005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HGZ8L1-A (organism)|Severe acute respiratory syndrome coronavirus HGZ8L1-A (organism)
C1532878|T005|PT|415396004|SNOMEDCT_US|SARS coronavirus HKU-66078|SARS coronavirus HKU-66078
C1532878|T005|OF|415396004|SNOMEDCT_US|SARS coronavirus HKU-66078 (organism)|SARS coronavirus HKU-66078 (organism)
C1532878|T005|SY|415396004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HKU-66078|Severe acute respiratory syndrome (SARS) coronavirus HKU-66078
C1532878|T005|OF|415396004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HKU-66078 (organism)|Severe acute respiratory syndrome (SARS) coronavirus HKU-66078 (organism)
C1532878|T005|SY|415396004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HKU-66078|Severe acute respiratory syndrome coronavirus HKU-66078
C1532878|T005|FN|415396004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HKU-66078 (organism)|Severe acute respiratory syndrome coronavirus HKU-66078 (organism)
C1532879|T005|PT|415397008|SNOMEDCT_US|SARS coronavirus Hong Kong/03/2003|SARS coronavirus Hong Kong/03/2003
C1532879|T005|OF|415397008|SNOMEDCT_US|SARS coronavirus Hong Kong/03/2003 (organism)|SARS coronavirus Hong Kong/03/2003 (organism)
C1532879|T005|SY|415397008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Hong Kong/03/2003|Severe acute respiratory syndrome (SARS) coronavirus Hong Kong/03/2003
C1532879|T005|OF|415397008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Hong Kong/03/2003 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Hong Kong/03/2003 (organism)
C1532879|T005|SY|415397008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Hong Kong/03/2003|Severe acute respiratory syndrome coronavirus Hong Kong/03/2003
C1532879|T005|FN|415397008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Hong Kong/03/2003 (organism)|Severe acute respiratory syndrome coronavirus Hong Kong/03/2003 (organism)
C1532880|T005|PT|415398003|SNOMEDCT_US|SARS coronavirus HPZ-2003|SARS coronavirus HPZ-2003
C1532880|T005|OF|415398003|SNOMEDCT_US|SARS coronavirus HPZ-2003 (organism)|SARS coronavirus HPZ-2003 (organism)
C1532880|T005|SY|415398003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HPZ-2003|Severe acute respiratory syndrome (SARS) coronavirus HPZ-2003
C1532880|T005|OF|415398003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HPZ-2003 (organism)|Severe acute respiratory syndrome (SARS) coronavirus HPZ-2003 (organism)
C1532880|T005|SY|415398003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HPZ-2003|Severe acute respiratory syndrome coronavirus HPZ-2003
C1532880|T005|FN|415398003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HPZ-2003 (organism)|Severe acute respiratory syndrome coronavirus HPZ-2003 (organism)
C1532881|T005|PT|415399006|SNOMEDCT_US|SARS coronavirus HSR 1|SARS coronavirus HSR 1
C1532881|T005|OF|415399006|SNOMEDCT_US|SARS coronavirus HSR 1 (organism)|SARS coronavirus HSR 1 (organism)
C1532881|T005|SY|415399006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HSR 1|Severe acute respiratory syndrome (SARS) coronavirus HSR 1
C1532881|T005|OF|415399006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HSR 1 (organism)|Severe acute respiratory syndrome (SARS) coronavirus HSR 1 (organism)
C1532881|T005|SY|415399006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HSR 1|Severe acute respiratory syndrome coronavirus HSR 1
C1532881|T005|FN|415399006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HSR 1 (organism)|Severe acute respiratory syndrome coronavirus HSR 1 (organism)
C1532882|T005|PT|415400004|SNOMEDCT_US|SARS coronavirus HSZ-A|SARS coronavirus HSZ-A
C1532882|T005|OF|415400004|SNOMEDCT_US|SARS coronavirus HSZ-A (organism)|SARS coronavirus HSZ-A (organism)
C1532882|T005|SY|415400004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HSZ-A|Severe acute respiratory syndrome (SARS) coronavirus HSZ-A
C1532882|T005|OF|415400004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HSZ-A (organism)|Severe acute respiratory syndrome (SARS) coronavirus HSZ-A (organism)
C1532882|T005|SY|415400004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HSZ-A|Severe acute respiratory syndrome coronavirus HSZ-A
C1532882|T005|FN|415400004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HSZ-A (organism)|Severe acute respiratory syndrome coronavirus HSZ-A (organism)
C1532883|T005|PT|415401000|SNOMEDCT_US|SARS coronavirus HSZ-Bb|SARS coronavirus HSZ-Bb
C1532883|T005|OF|415401000|SNOMEDCT_US|SARS coronavirus HSZ-Bb (organism)|SARS coronavirus HSZ-Bb (organism)
C1532883|T005|SY|415401000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HSZ-Bb|Severe acute respiratory syndrome (SARS) coronavirus HSZ-Bb
C1532883|T005|OF|415401000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HSZ-Bb (organism)|Severe acute respiratory syndrome (SARS) coronavirus HSZ-Bb (organism)
C1532883|T005|SY|415401000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HSZ-Bb|Severe acute respiratory syndrome coronavirus HSZ-Bb
C1532883|T005|FN|415401000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HSZ-Bb (organism)|Severe acute respiratory syndrome coronavirus HSZ-Bb (organism)
C1532884|T005|PT|415402007|SNOMEDCT_US|SARS coronavirus HSZ-Bc|SARS coronavirus HSZ-Bc
C1532884|T005|OF|415402007|SNOMEDCT_US|SARS coronavirus HSZ-Bc (organism)|SARS coronavirus HSZ-Bc (organism)
C1532884|T005|SY|415402007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HSZ-Bc|Severe acute respiratory syndrome (SARS) coronavirus HSZ-Bc
C1532884|T005|OF|415402007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HSZ-Bc (organism)|Severe acute respiratory syndrome (SARS) coronavirus HSZ-Bc (organism)
C1532884|T005|SY|415402007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HSZ-Bc|Severe acute respiratory syndrome coronavirus HSZ-Bc
C1532884|T005|FN|415402007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HSZ-Bc (organism)|Severe acute respiratory syndrome coronavirus HSZ-Bc (organism)
C1532885|T005|PT|415403002|SNOMEDCT_US|SARS coronavirus HSZ-Cb|SARS coronavirus HSZ-Cb
C1532885|T005|OF|415403002|SNOMEDCT_US|SARS coronavirus HSZ-Cb (organism)|SARS coronavirus HSZ-Cb (organism)
C1532885|T005|SY|415403002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HSZ-Cb|Severe acute respiratory syndrome (SARS) coronavirus HSZ-Cb
C1532885|T005|OF|415403002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HSZ-Cb (organism)|Severe acute respiratory syndrome (SARS) coronavirus HSZ-Cb (organism)
C1532885|T005|SY|415403002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HSZ-Cb|Severe acute respiratory syndrome coronavirus HSZ-Cb
C1532885|T005|FN|415403002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HSZ-Cb (organism)|Severe acute respiratory syndrome coronavirus HSZ-Cb (organism)
C1532886|T005|PT|415404008|SNOMEDCT_US|SARS coronavirus HSZ-Cc|SARS coronavirus HSZ-Cc
C1532886|T005|OF|415404008|SNOMEDCT_US|SARS coronavirus HSZ-Cc (organism)|SARS coronavirus HSZ-Cc (organism)
C1532886|T005|SY|415404008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HSZ-Cc|Severe acute respiratory syndrome (SARS) coronavirus HSZ-Cc
C1532886|T005|OF|415404008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HSZ-Cc (organism)|Severe acute respiratory syndrome (SARS) coronavirus HSZ-Cc (organism)
C1532886|T005|SY|415404008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HSZ-Cc|Severe acute respiratory syndrome coronavirus HSZ-Cc
C1532886|T005|FN|415404008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HSZ-Cc (organism)|Severe acute respiratory syndrome coronavirus HSZ-Cc (organism)
C1532887|T005|PT|415405009|SNOMEDCT_US|SARS coronavirus HSZ2-A|SARS coronavirus HSZ2-A
C1532887|T005|OF|415405009|SNOMEDCT_US|SARS coronavirus HSZ2-A (organism)|SARS coronavirus HSZ2-A (organism)
C1532887|T005|SY|415405009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HSZ2-A|Severe acute respiratory syndrome (SARS) coronavirus HSZ2-A
C1532887|T005|OF|415405009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HSZ2-A (organism)|Severe acute respiratory syndrome (SARS) coronavirus HSZ2-A (organism)
C1532887|T005|SY|415405009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HSZ2-A|Severe acute respiratory syndrome coronavirus HSZ2-A
C1532887|T005|FN|415405009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HSZ2-A (organism)|Severe acute respiratory syndrome coronavirus HSZ2-A (organism)
C1532888|T005|PT|415406005|SNOMEDCT_US|SARS coronavirus HZS2-Bb|SARS coronavirus HZS2-Bb
C1532888|T005|OF|415406005|SNOMEDCT_US|SARS coronavirus HZS2-Bb (organism)|SARS coronavirus HZS2-Bb (organism)
C1532888|T005|SY|415406005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HSZ2-Bb|Severe acute respiratory syndrome (SARS) coronavirus HSZ2-Bb
C1532888|T005|OF|415406005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HSZ2-Bb (organism)|Severe acute respiratory syndrome (SARS) coronavirus HSZ2-Bb (organism)
C1532888|T005|SY|415406005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HSZ2-Bb|Severe acute respiratory syndrome coronavirus HSZ2-Bb
C1532888|T005|FN|415406005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HSZ2-Bb (organism)|Severe acute respiratory syndrome coronavirus HSZ2-Bb (organism)
C1532889|T005|PT|415407001|SNOMEDCT_US|SARS coronavirus HZS2-C|SARS coronavirus HZS2-C
C1532889|T005|OF|415407001|SNOMEDCT_US|SARS coronavirus HZS2-C (organism)|SARS coronavirus HZS2-C (organism)
C1532889|T005|SY|415407001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HZS2-C|Severe acute respiratory syndrome (SARS) coronavirus HZS2-C
C1532889|T005|OF|415407001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HZS2-C (organism)|Severe acute respiratory syndrome (SARS) coronavirus HZS2-C (organism)
C1532889|T005|SY|415407001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HZS2-C|Severe acute respiratory syndrome coronavirus HZS2-C
C1532889|T005|FN|415407001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HZS2-C (organism)|Severe acute respiratory syndrome coronavirus HZS2-C (organism)
C1532890|T005|PT|415408006|SNOMEDCT_US|SARS coronavirus HZS2-D|SARS coronavirus HZS2-D
C1532890|T005|OF|415408006|SNOMEDCT_US|SARS coronavirus HZS2-D (organism)|SARS coronavirus HZS2-D (organism)
C1532890|T005|SY|415408006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HZS2-D|Severe acute respiratory syndrome (SARS) coronavirus HZS2-D
C1532890|T005|OF|415408006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HZS2-D (organism)|Severe acute respiratory syndrome (SARS) coronavirus HZS2-D (organism)
C1532890|T005|SY|415408006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HZS2-D|Severe acute respiratory syndrome coronavirus HZS2-D
C1532890|T005|FN|415408006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HZS2-D (organism)|Severe acute respiratory syndrome coronavirus HZS2-D (organism)
C1532891|T005|PT|415409003|SNOMEDCT_US|SARS coronavirus HZS2-E|SARS coronavirus HZS2-E
C1532891|T005|OF|415409003|SNOMEDCT_US|SARS coronavirus HZS2-E (organism)|SARS coronavirus HZS2-E (organism)
C1532891|T005|SY|415409003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HZS2-E|Severe acute respiratory syndrome (SARS) coronavirus HZS2-E
C1532891|T005|OF|415409003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HZS2-E (organism)|Severe acute respiratory syndrome (SARS) coronavirus HZS2-E (organism)
C1532891|T005|SY|415409003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HZS2-E|Severe acute respiratory syndrome coronavirus HZS2-E
C1532891|T005|FN|415409003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HZS2-E (organism)|Severe acute respiratory syndrome coronavirus HZS2-E (organism)
C1532892|T005|PT|415410008|SNOMEDCT_US|SARS coronavirus HZS2-Fb|SARS coronavirus HZS2-Fb
C1532892|T005|OF|415410008|SNOMEDCT_US|SARS coronavirus HZS2-Fb (organism)|SARS coronavirus HZS2-Fb (organism)
C1532892|T005|SY|415410008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HZS2-Fb|Severe acute respiratory syndrome (SARS) coronavirus HZS2-Fb
C1532892|T005|OF|415410008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HZS2-Fb (organism)|Severe acute respiratory syndrome (SARS) coronavirus HZS2-Fb (organism)
C1532892|T005|SY|415410008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HZS2-Fb|Severe acute respiratory syndrome coronavirus HZS2-Fb
C1532892|T005|FN|415410008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HZS2-Fb (organism)|Severe acute respiratory syndrome coronavirus HZS2-Fb (organism)
C1532893|T005|PT|415411007|SNOMEDCT_US|SARS coronavirus HZS2-Fc|SARS coronavirus HZS2-Fc
C1532893|T005|OF|415411007|SNOMEDCT_US|SARS coronavirus HZS2-Fc (organism)|SARS coronavirus HZS2-Fc (organism)
C1532893|T005|SY|415411007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HZS2-Fc|Severe acute respiratory syndrome (SARS) coronavirus HZS2-Fc
C1532893|T005|OF|415411007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HZS2-Fc (organism)|Severe acute respiratory syndrome (SARS) coronavirus HZS2-Fc (organism)
C1532893|T005|SY|415411007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HZS2-Fc|Severe acute respiratory syndrome coronavirus HZS2-Fc
C1532893|T005|FN|415411007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HZS2-Fc (organism)|Severe acute respiratory syndrome coronavirus HZS2-Fc (organism)
C1532894|T005|PT|415412000|SNOMEDCT_US|SARS coronavirus JMD|SARS coronavirus JMD
C1532894|T005|OF|415412000|SNOMEDCT_US|SARS coronavirus JMD (organism)|SARS coronavirus JMD (organism)
C1532894|T005|SY|415412000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HZS2-JMD|Severe acute respiratory syndrome (SARS) coronavirus HZS2-JMD
C1532894|T005|OF|415412000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HZS2-JMD (organism)|Severe acute respiratory syndrome (SARS) coronavirus HZS2-JMD (organism)
C1532894|T005|SY|415412000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HZS2-JMD|Severe acute respiratory syndrome coronavirus HZS2-JMD
C1532894|T005|FN|415412000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HZS2-JMD (organism)|Severe acute respiratory syndrome coronavirus HZS2-JMD (organism)
C1532895|T005|PT|415413005|SNOMEDCT_US|SARS coronavirus LC1|SARS coronavirus LC1
C1532895|T005|OF|415413005|SNOMEDCT_US|SARS coronavirus LC1 (organism)|SARS coronavirus LC1 (organism)
C1532895|T005|SY|415413005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus LC1|Severe acute respiratory syndrome (SARS) coronavirus LC1
C1532895|T005|OF|415413005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus LC1 (organism)|Severe acute respiratory syndrome (SARS) coronavirus LC1 (organism)
C1532895|T005|SY|415413005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus LC1|Severe acute respiratory syndrome coronavirus LC1
C1532895|T005|FN|415413005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus LC1 (organism)|Severe acute respiratory syndrome coronavirus LC1 (organism)
C1532896|T005|PT|415414004|SNOMEDCT_US|SARS coronavirus LC2|SARS coronavirus LC2
C1532896|T005|OF|415414004|SNOMEDCT_US|SARS coronavirus LC2 (organism)|SARS coronavirus LC2 (organism)
C1532896|T005|SY|415414004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus LC2|Severe acute respiratory syndrome (SARS) coronavirus LC2
C1532896|T005|OF|415414004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus LC2 (organism)|Severe acute respiratory syndrome (SARS) coronavirus LC2 (organism)
C1532896|T005|SY|415414004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus LC2|Severe acute respiratory syndrome coronavirus LC2
C1532896|T005|FN|415414004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus LC2 (organism)|Severe acute respiratory syndrome coronavirus LC2 (organism)
C1532897|T005|PT|415415003|SNOMEDCT_US|SARS coronavirus LC3|SARS coronavirus LC3
C1532897|T005|OF|415415003|SNOMEDCT_US|SARS coronavirus LC3 (organism)|SARS coronavirus LC3 (organism)
C1532897|T005|SY|415415003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus LC3|Severe acute respiratory syndrome (SARS) coronavirus LC3
C1532897|T005|OF|415415003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus LC3 (organism)|Severe acute respiratory syndrome (SARS) coronavirus LC3 (organism)
C1532897|T005|SY|415415003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus LC3|Severe acute respiratory syndrome coronavirus LC3
C1532897|T005|FN|415415003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus LC3 (organism)|Severe acute respiratory syndrome coronavirus LC3 (organism)
C1532898|T005|PT|415416002|SNOMEDCT_US|SARS coronavirus LC4|SARS coronavirus LC4
C1532898|T005|OF|415416002|SNOMEDCT_US|SARS coronavirus LC4 (organism)|SARS coronavirus LC4 (organism)
C1532898|T005|SY|415416002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus LC4|Severe acute respiratory syndrome (SARS) coronavirus LC4
C1532898|T005|OF|415416002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus LC4 (organism)|Severe acute respiratory syndrome (SARS) coronavirus LC4 (organism)
C1532898|T005|SY|415416002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus LC4|Severe acute respiratory syndrome coronavirus LC4
C1532898|T005|FN|415416002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus LC4 (organism)|Severe acute respiratory syndrome coronavirus LC4 (organism)
C1532899|T005|PT|415417006|SNOMEDCT_US|SARS coronavirus LC5|SARS coronavirus LC5
C1532899|T005|OF|415417006|SNOMEDCT_US|SARS coronavirus LC5 (organism)|SARS coronavirus LC5 (organism)
C1532899|T005|SY|415417006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus LC5|Severe acute respiratory syndrome (SARS) coronavirus LC5
C1532899|T005|OF|415417006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus LC5 (organism)|Severe acute respiratory syndrome (SARS) coronavirus LC5 (organism)
C1532899|T005|SY|415417006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus LC5|Severe acute respiratory syndrome coronavirus LC5
C1532899|T005|FN|415417006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus LC5 (organism)|Severe acute respiratory syndrome coronavirus LC5 (organism)
C1532900|T005|PT|415418001|SNOMEDCT_US|SARS coronavirus NS-1|SARS coronavirus NS-1
C1532900|T005|OF|415418001|SNOMEDCT_US|SARS coronavirus NS-1 (organism)|SARS coronavirus NS-1 (organism)
C1532900|T005|SY|415418001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus NS-1|Severe acute respiratory syndrome (SARS) coronavirus NS-1
C1532900|T005|OF|415418001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus NS-1 (organism)|Severe acute respiratory syndrome (SARS) coronavirus NS-1 (organism)
C1532900|T005|SY|415418001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus NS-1|Severe acute respiratory syndrome coronavirus NS-1
C1532900|T005|FN|415418001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus NS-1 (organism)|Severe acute respiratory syndrome coronavirus NS-1 (organism)
C1532901|T005|PT|415419009|SNOMEDCT_US|SARS coronavirus PUMC01|SARS coronavirus PUMC01
C1532901|T005|OF|415419009|SNOMEDCT_US|SARS coronavirus PUMC01 (organism)|SARS coronavirus PUMC01 (organism)
C1532901|T005|SY|415419009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus PUMC01|Severe acute respiratory syndrome (SARS) coronavirus PUMC01
C1532901|T005|OF|415419009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus PUMC01 (organism)|Severe acute respiratory syndrome (SARS) coronavirus PUMC01 (organism)
C1532901|T005|SY|415419009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus PUMC01|Severe acute respiratory syndrome coronavirus PUMC01
C1532901|T005|FN|415419009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus PUMC01 (organism)|Severe acute respiratory syndrome coronavirus PUMC01 (organism)
C1532902|T005|PT|415420003|SNOMEDCT_US|SARS coronavirus PUMC02|SARS coronavirus PUMC02
C1532902|T005|OF|415420003|SNOMEDCT_US|SARS coronavirus PUMC02 (organism)|SARS coronavirus PUMC02 (organism)
C1532902|T005|SY|415420003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus PUMC02|Severe acute respiratory syndrome (SARS) coronavirus PUMC02
C1532902|T005|OF|415420003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus PUMC02 (organism)|Severe acute respiratory syndrome (SARS) coronavirus PUMC02 (organism)
C1532902|T005|SY|415420003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus PUMC02|Severe acute respiratory syndrome coronavirus PUMC02
C1532902|T005|FN|415420003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus PUMC02 (organism)|Severe acute respiratory syndrome coronavirus PUMC02 (organism)
C1532903|T005|PT|415421004|SNOMEDCT_US|SARS coronavirus PUMC03|SARS coronavirus PUMC03
C1532903|T005|OF|415421004|SNOMEDCT_US|SARS coronavirus PUMC03 (organism)|SARS coronavirus PUMC03 (organism)
C1532903|T005|SY|415421004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus PUMC03|Severe acute respiratory syndrome (SARS) coronavirus PUMC03
C1532903|T005|OF|415421004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus PUMC03 (organism)|Severe acute respiratory syndrome (SARS) coronavirus PUMC03 (organism)
C1532903|T005|SY|415421004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus PUMC03|Severe acute respiratory syndrome coronavirus PUMC03
C1532903|T005|FN|415421004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus PUMC03 (organism)|Severe acute respiratory syndrome coronavirus PUMC03 (organism)
C1532904|T005|PT|415422006|SNOMEDCT_US|SARS coronavirus sf098|SARS coronavirus sf098
C1532904|T005|OF|415422006|SNOMEDCT_US|SARS coronavirus sf098 (organism)|SARS coronavirus sf098 (organism)
C1532904|T005|SY|415422006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus sf098|Severe acute respiratory syndrome (SARS) coronavirus sf098
C1532904|T005|OF|415422006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus sf098 (organism)|Severe acute respiratory syndrome (SARS) coronavirus sf098 (organism)
C1532904|T005|SY|415422006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus sf098|Severe acute respiratory syndrome coronavirus sf098
C1532904|T005|FN|415422006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus sf098 (organism)|Severe acute respiratory syndrome coronavirus sf098 (organism)
C1532905|T005|PT|415423001|SNOMEDCT_US|SARS coronavirus sf099|SARS coronavirus sf099
C1532905|T005|OF|415423001|SNOMEDCT_US|SARS coronavirus sf099 (organism)|SARS coronavirus sf099 (organism)
C1532905|T005|SY|415423001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus sf099|Severe acute respiratory syndrome (SARS) coronavirus sf099
C1532905|T005|OF|415423001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus sf099 (organism)|Severe acute respiratory syndrome (SARS) coronavirus sf099 (organism)
C1532905|T005|SY|415423001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus sf099|Severe acute respiratory syndrome coronavirus sf099
C1532905|T005|FN|415423001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus sf099 (organism)|Severe acute respiratory syndrome coronavirus sf099 (organism)
C1532906|T005|SY|415424007|SNOMEDCT_US|SARS coronavirus Shanghai LY|SARS coronavirus Shanghai LY
C1532906|T005|OF|415424007|SNOMEDCT_US|SARS coronavirus Shanghai LY (organism)|SARS coronavirus Shanghai LY (organism)
C1532906|T005|IS|415424007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Shanghai LY|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Shanghai LY
C1532906|T005|OF|415424007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Shanghai LY (organism)|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Shanghai LY (organism)
C1532906|T005|PT|415424007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Shanghai LY|Severe acute respiratory syndrome (SARS) coronavirus Shanghai LY
C1532906|T005|OF|415424007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Shanghai LY (organism)|Severe acute respiratory syndrome (SARS) coronavirus Shanghai LY (organism)
C1532906|T005|SY|415424007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Shanghai LY|Severe acute respiratory syndrome coronavirus Shanghai LY
C1532906|T005|FN|415424007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Shanghai LY (organism)|Severe acute respiratory syndrome coronavirus Shanghai LY (organism)
C1532907|T005|SY|415425008|SNOMEDCT_US|SARS coronavirus ShanghaiQXC1|SARS coronavirus ShanghaiQXC1
C1532907|T005|OF|415425008|SNOMEDCT_US|SARS coronavirus ShanghaiQXC1 (organism)|SARS coronavirus ShanghaiQXC1 (organism)
C1532907|T005|IS|415425008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus coronavirus ShanghaiQXC1|Severe acute respiratory syndrome (SARS) coronavirus coronavirus ShanghaiQXC1
C1532907|T005|OF|415425008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus coronavirus ShanghaiQXC1 (organism)|Severe acute respiratory syndrome (SARS) coronavirus coronavirus ShanghaiQXC1 (organism)
C1532907|T005|PT|415425008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus ShanghaiQXC1|Severe acute respiratory syndrome (SARS) coronavirus ShanghaiQXC1
C1532907|T005|OF|415425008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus ShanghaiQXC1 (organism)|Severe acute respiratory syndrome (SARS) coronavirus ShanghaiQXC1 (organism)
C1532907|T005|SY|415425008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus ShanghaiQXC1|Severe acute respiratory syndrome coronavirus ShanghaiQXC1
C1532907|T005|FN|415425008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus ShanghaiQXC1 (organism)|Severe acute respiratory syndrome coronavirus ShanghaiQXC1 (organism)
C1532908|T005|SY|415426009|SNOMEDCT_US|SARS coronavirus ShanghaiQXC2|SARS coronavirus ShanghaiQXC2
C1532908|T005|OF|415426009|SNOMEDCT_US|SARS coronavirus ShanghaiQXC2 (organism)|SARS coronavirus ShanghaiQXC2 (organism)
C1532908|T005|IS|415426009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus coronavirus ShanghaiQXC2|Severe acute respiratory syndrome (SARS) coronavirus coronavirus ShanghaiQXC2
C1532908|T005|OF|415426009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus coronavirus ShanghaiQXC2 (organism)|Severe acute respiratory syndrome (SARS) coronavirus coronavirus ShanghaiQXC2 (organism)
C1532908|T005|PT|415426009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus ShanghaiQXC2|Severe acute respiratory syndrome (SARS) coronavirus ShanghaiQXC2
C1532908|T005|OF|415426009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus ShanghaiQXC2 (organism)|Severe acute respiratory syndrome (SARS) coronavirus ShanghaiQXC2 (organism)
C1532908|T005|SY|415426009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus ShanghaiQXC2|Severe acute respiratory syndrome coronavirus ShanghaiQXC2
C1532908|T005|FN|415426009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus ShanghaiQXC2 (organism)|Severe acute respiratory syndrome coronavirus ShanghaiQXC2 (organism)
C1532909|T005|PT|415427000|SNOMEDCT_US|SARS coronavirus Sin 3765V|SARS coronavirus Sin 3765V
C1532909|T005|OF|415427000|SNOMEDCT_US|SARS coronavirus Sin 3765V (organism)|SARS coronavirus Sin 3765V (organism)
C1532909|T005|SY|415427000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin 3765V|Severe acute respiratory syndrome (SARS) coronavirus Sin 3765V
C1532909|T005|OF|415427000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin 3765V (organism)|Severe acute respiratory syndrome (SARS) coronavirus Sin 3765V (organism)
C1532909|T005|SY|415427000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin 3765V|Severe acute respiratory syndrome coronavirus Sin 3765V
C1532909|T005|FN|415427000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin 3765V (organism)|Severe acute respiratory syndrome coronavirus Sin 3765V (organism)
C1532910|T005|SY|415428005|SNOMEDCT_US|SARS coronavirus Sin0409|SARS coronavirus Sin0409
C1532910|T005|OF|415428005|SNOMEDCT_US|SARS coronavirus Sin0409 (organism)|SARS coronavirus Sin0409 (organism)
C1532910|T005|IS|415428005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin0409|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin0409
C1532910|T005|OF|415428005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin0409 (organism)|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin0409 (organism)
C1532910|T005|PT|415428005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin0409|Severe acute respiratory syndrome (SARS) coronavirus Sin0409
C1532910|T005|OF|415428005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin0409 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Sin0409 (organism)
C1532910|T005|SY|415428005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin0409|Severe acute respiratory syndrome coronavirus Sin0409
C1532910|T005|FN|415428005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin0409 (organism)|Severe acute respiratory syndrome coronavirus Sin0409 (organism)
C1532911|T005|PT|415429002|SNOMEDCT_US|SARS coronavirus Sin1-11|SARS coronavirus Sin1-11
C1532911|T005|OF|415429002|SNOMEDCT_US|SARS coronavirus Sin1-11 (organism)|SARS coronavirus Sin1-11 (organism)
C1532911|T005|SY|415429002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin1-11|Severe acute respiratory syndrome (SARS) coronavirus Sin1-11
C1532911|T005|OF|415429002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin1-11 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Sin1-11 (organism)
C1532911|T005|SY|415429002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin1-11|Severe acute respiratory syndrome coronavirus Sin1-11
C1532911|T005|FN|415429002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin1-11 (organism)|Severe acute respiratory syndrome coronavirus Sin1-11 (organism)
C1532912|T005|PT|415430007|SNOMEDCT_US|SARS coronavirus Sin2500|SARS coronavirus Sin2500
C1532912|T005|OF|415430007|SNOMEDCT_US|SARS coronavirus Sin2500 (organism)|SARS coronavirus Sin2500 (organism)
C1532912|T005|IS|415430007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin2500|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin2500
C1532912|T005|OF|415430007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin2500 (organism)|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin2500 (organism)
C1532912|T005|SY|415430007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin2500|Severe acute respiratory syndrome (SARS) coronavirus Sin2500
C1532912|T005|OF|415430007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin2500 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Sin2500 (organism)
C1532912|T005|SY|415430007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin2500|Severe acute respiratory syndrome coronavirus Sin2500
C1532912|T005|FN|415430007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin2500 (organism)|Severe acute respiratory syndrome coronavirus Sin2500 (organism)
C1532913|T005|SY|415431006|SNOMEDCT_US|SARS coronavirus Sin2677|SARS coronavirus Sin2677
C1532913|T005|OF|415431006|SNOMEDCT_US|SARS coronavirus Sin2677 (organism)|SARS coronavirus Sin2677 (organism)
C1532913|T005|IS|415431006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin2677|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin2677
C1532913|T005|OF|415431006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin2677 (organism)|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin2677 (organism)
C1532913|T005|PT|415431006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin2677|Severe acute respiratory syndrome (SARS) coronavirus Sin2677
C1532913|T005|OF|415431006|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin2677 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Sin2677 (organism)
C1532913|T005|SY|415431006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin2677|Severe acute respiratory syndrome coronavirus Sin2677
C1532913|T005|FN|415431006|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin2677 (organism)|Severe acute respiratory syndrome coronavirus Sin2677 (organism)
C1532914|T005|SY|415432004|SNOMEDCT_US|SARS coronavirus Sin2679|SARS coronavirus Sin2679
C1532914|T005|OF|415432004|SNOMEDCT_US|SARS coronavirus Sin2679 (organism)|SARS coronavirus Sin2679 (organism)
C1532914|T005|IS|415432004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin2679|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin2679
C1532914|T005|OF|415432004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin2679 (organism)|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin2679 (organism)
C1532914|T005|PT|415432004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin2679|Severe acute respiratory syndrome (SARS) coronavirus Sin2679
C1532914|T005|OF|415432004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin2679 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Sin2679 (organism)
C1532914|T005|SY|415432004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin2679|Severe acute respiratory syndrome coronavirus Sin2679
C1532914|T005|FN|415432004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin2679 (organism)|Severe acute respiratory syndrome coronavirus Sin2679 (organism)
C1532915|T005|SY|415433009|SNOMEDCT_US|SARS coronavirus Sin2748|SARS coronavirus Sin2748
C1532915|T005|OF|415433009|SNOMEDCT_US|SARS coronavirus Sin2748 (organism)|SARS coronavirus Sin2748 (organism)
C1532915|T005|IS|415433009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin2748|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin2748
C1532915|T005|OF|415433009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin2748 (organism)|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin2748 (organism)
C1532915|T005|PT|415433009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin2748|Severe acute respiratory syndrome (SARS) coronavirus Sin2748
C1532915|T005|OF|415433009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin2748 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Sin2748 (organism)
C1532915|T005|SY|415433009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin2748|Severe acute respiratory syndrome coronavirus Sin2748
C1532915|T005|FN|415433009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin2748 (organism)|Severe acute respiratory syndrome coronavirus Sin2748 (organism)
C1532916|T005|SY|415434003|SNOMEDCT_US|SARS coronavirus Sin2774|SARS coronavirus Sin2774
C1532916|T005|OF|415434003|SNOMEDCT_US|SARS coronavirus Sin2774 (organism)|SARS coronavirus Sin2774 (organism)
C1532916|T005|IS|415434003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin2774|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin2774
C1532916|T005|OF|415434003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin2774 (organism)|Severe acute respiratory syndrome (SARS) coronavirus coronavirus Sin2774 (organism)
C1532916|T005|PT|415434003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin2774|Severe acute respiratory syndrome (SARS) coronavirus Sin2774
C1532916|T005|OF|415434003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin2774 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Sin2774 (organism)
C1532916|T005|SY|415434003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin2774|Severe acute respiratory syndrome coronavirus Sin2774
C1532916|T005|FN|415434003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin2774 (organism)|Severe acute respiratory syndrome coronavirus Sin2774 (organism)
C1532917|T005|PT|415435002|SNOMEDCT_US|SARS coronavirus Sin3-11|SARS coronavirus Sin3-11
C1532917|T005|OF|415435002|SNOMEDCT_US|SARS coronavirus Sin3-11 (organism)|SARS coronavirus Sin3-11 (organism)
C1532917|T005|SY|415435002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin3-11|Severe acute respiratory syndrome (SARS) coronavirus Sin3-11
C1532917|T005|OF|415435002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin3-11 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Sin3-11 (organism)
C1532917|T005|SY|415435002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin3-11|Severe acute respiratory syndrome coronavirus Sin3-11
C1532917|T005|FN|415435002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin3-11 (organism)|Severe acute respiratory syndrome coronavirus Sin3-11 (organism)
C1532918|T005|PT|415436001|SNOMEDCT_US|SARS coronavirus Sin3408|SARS coronavirus Sin3408
C1532918|T005|OF|415436001|SNOMEDCT_US|SARS coronavirus Sin3408 (organism)|SARS coronavirus Sin3408 (organism)
C1532918|T005|SY|415436001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin3408|Severe acute respiratory syndrome (SARS) coronavirus Sin3408
C1532918|T005|OF|415436001|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin3408 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Sin3408 (organism)
C1532918|T005|SY|415436001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin3408|Severe acute respiratory syndrome coronavirus Sin3408
C1532918|T005|FN|415436001|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin3408 (organism)|Severe acute respiratory syndrome coronavirus Sin3408 (organism)
C1532919|T005|PT|415437005|SNOMEDCT_US|SARS coronavirus Sin3725V|SARS coronavirus Sin3725V
C1532919|T005|OF|415437005|SNOMEDCT_US|SARS coronavirus Sin3725V (organism)|SARS coronavirus Sin3725V (organism)
C1532919|T005|SY|415437005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin3725V|Severe acute respiratory syndrome (SARS) coronavirus Sin3725V
C1532919|T005|OF|415437005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin3725V (organism)|Severe acute respiratory syndrome (SARS) coronavirus Sin3725V (organism)
C1532919|T005|SY|415437005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin3725V|Severe acute respiratory syndrome coronavirus Sin3725V
C1532919|T005|FN|415437005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin3725V (organism)|Severe acute respiratory syndrome coronavirus Sin3725V (organism)
C1532920|T005|PT|415438000|SNOMEDCT_US|SARS coronavirus Sin842|SARS coronavirus Sin842
C1532920|T005|OF|415438000|SNOMEDCT_US|SARS coronavirus Sin842 (organism)|SARS coronavirus Sin842 (organism)
C1532920|T005|SY|415438000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin842|Severe acute respiratory syndrome (SARS) coronavirus Sin842
C1532920|T005|OF|415438000|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin842 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Sin842 (organism)
C1532920|T005|SY|415438000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin842|Severe acute respiratory syndrome coronavirus Sin842
C1532920|T005|FN|415438000|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin842 (organism)|Severe acute respiratory syndrome coronavirus Sin842 (organism)
C1532921|T005|PT|415439008|SNOMEDCT_US|SARS coronavirus Sin845|SARS coronavirus Sin845
C1532921|T005|OF|415439008|SNOMEDCT_US|SARS coronavirus Sin845 (organism)|SARS coronavirus Sin845 (organism)
C1532921|T005|SY|415439008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin845|Severe acute respiratory syndrome (SARS) coronavirus Sin845
C1532921|T005|OF|415439008|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin845 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Sin845 (organism)
C1532921|T005|SY|415439008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin845|Severe acute respiratory syndrome coronavirus Sin845
C1532921|T005|FN|415439008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin845 (organism)|Severe acute respiratory syndrome coronavirus Sin845 (organism)
C1532922|T005|PT|415440005|SNOMEDCT_US|SARS coronavirus Sin846|SARS coronavirus Sin846
C1532922|T005|OF|415440005|SNOMEDCT_US|SARS coronavirus Sin846 (organism)|SARS coronavirus Sin846 (organism)
C1532922|T005|SY|415440005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin846|Severe acute respiratory syndrome (SARS) coronavirus Sin846
C1532922|T005|OF|415440005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin846 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Sin846 (organism)
C1532922|T005|SY|415440005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin846|Severe acute respiratory syndrome coronavirus Sin846
C1532922|T005|FN|415440005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin846 (organism)|Severe acute respiratory syndrome coronavirus Sin846 (organism)
C1532923|T005|PT|415441009|SNOMEDCT_US|SARS coronavirus Sin847|SARS coronavirus Sin847
C1532923|T005|OF|415441009|SNOMEDCT_US|SARS coronavirus Sin847 (organism)|SARS coronavirus Sin847 (organism)
C1532923|T005|SY|415441009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin847|Severe acute respiratory syndrome (SARS) coronavirus Sin847
C1532923|T005|OF|415441009|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin847 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Sin847 (organism)
C1532923|T005|SY|415441009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin847|Severe acute respiratory syndrome coronavirus Sin847
C1532923|T005|FN|415441009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin847 (organism)|Severe acute respiratory syndrome coronavirus Sin847 (organism)
C1532924|T005|PT|415442002|SNOMEDCT_US|SARS coronavirus Sin848|SARS coronavirus Sin848
C1532924|T005|OF|415442002|SNOMEDCT_US|SARS coronavirus Sin848 (organism)|SARS coronavirus Sin848 (organism)
C1532924|T005|SY|415442002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin848|Severe acute respiratory syndrome (SARS) coronavirus Sin848
C1532924|T005|OF|415442002|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin848 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Sin848 (organism)
C1532924|T005|SY|415442002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin848|Severe acute respiratory syndrome coronavirus Sin848
C1532924|T005|FN|415442002|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin848 (organism)|Severe acute respiratory syndrome coronavirus Sin848 (organism)
C1532925|T005|PT|415443007|SNOMEDCT_US|SARS coronavirus Sin849|SARS coronavirus Sin849
C1532925|T005|OF|415443007|SNOMEDCT_US|SARS coronavirus Sin849 (organism)|SARS coronavirus Sin849 (organism)
C1532925|T005|SY|415443007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin849|Severe acute respiratory syndrome (SARS) coronavirus Sin849
C1532925|T005|OF|415443007|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Sin849 (organism)|Severe acute respiratory syndrome (SARS) coronavirus Sin849 (organism)
C1532925|T005|SY|415443007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin849|Severe acute respiratory syndrome coronavirus Sin849
C1532925|T005|FN|415443007|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Sin849 (organism)|Severe acute respiratory syndrome coronavirus Sin849 (organism)
C1533184|T005|LPN|LP31724-5|LNC|SARS coronavirus Urbani|SARS coronavirus Urbani
C1533184|T005|PT|415495004|SNOMEDCT_US|SARS coronavirus Urbani|SARS coronavirus Urbani
C1533184|T005|PN|NOCODE|MTH|SARS coronavirus Urbani|SARS coronavirus Urbani
C1533184|T005|OF|415495004|SNOMEDCT_US|SARS coronavirus Urbani (organism)|SARS coronavirus Urbani (organism)
C1533184|T005|SY|415495004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Urbani|Severe acute respiratory syndrome (SARS) coronavirus Urbani
C1533184|T005|OF|415495004|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus Urbani (organism)|Severe acute respiratory syndrome (SARS) coronavirus Urbani (organism)
C1533184|T005|SY|415495004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Urbani|Severe acute respiratory syndrome coronavirus Urbani
C1533184|T005|FN|415495004|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Urbani (organism)|Severe acute respiratory syndrome coronavirus Urbani (organism)
C1544947|T201|DN|41000-1|LNC|HCoV RNA NAA+probe Nom (Unsp spec)|HCoV RNA NAA+probe Nom (Unsp spec)
C1544947|T201|OSN|41000-1|LNC|HCoV RNA XXX NAA+probe|HCoV RNA XXX NAA+probe
C1544947|T201|MTH_LN|41000-1|LNC|Human coronavirus ribonucleic acid:Presence or Identity:Point in time:To be specified in another part of the message:Nominal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus ribonucleic acid:Presence or Identity:Point in time:To be specified in another part of the message:Nominal:DNA Nucleic Acid Probe.amp.tar
C1544947|T201|LC|41000-1|LNC|Human coronavirus RNA [Identifier] in Unspecified specimen by NAA with probe detection|Human coronavirus RNA [Identifier] in Unspecified specimen by NAA with probe detection
C1544947|T201|LN|41000-1|LNC|Human coronavirus RNA:Prid:Pt:XXX:Nom:Probe.amp.tar|Human coronavirus RNA:Prid:Pt:XXX:Nom:Probe.amp.tar
C1544948|T201|DN|41001-9|LNC|HCoV RNA NAA+probe Ql (Unsp spec)|HCoV RNA NAA+probe Ql (Unsp spec)
C1544948|T201|OSN|41001-9|LNC|HCoV RNA XXX Ql NAA+probe|HCoV RNA XXX Ql NAA+probe
C1544948|T201|MTH_LN|41001-9|LNC|Human coronavirus ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar
C1544948|T201|LC|41001-9|LNC|Human coronavirus RNA [Presence] in Unspecified specimen by NAA with probe detection|Human coronavirus RNA [Presence] in Unspecified specimen by NAA with probe detection
C1544948|T201|LN|41001-9|LNC|Human coronavirus RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar|Human coronavirus RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar
C1544949|T201|DN|41002-7|LNC|HCoV 229E IgG IA Ql (S)|HCoV 229E IgG IA Ql (S)
C1544949|T201|OSN|41002-7|LNC|HCoV 229E IgG Ser Ql IA|HCoV 229E IgG Ser Ql IA
C1544949|T201|LN|41002-7|LNC|Human coronavirus 229E Ab.IgG:PrThr:Pt:Ser:Ord:IA|Human coronavirus 229E Ab.IgG:PrThr:Pt:Ser:Ord:IA
C1544949|T201|MTH_LN|41002-7|LNC|Human coronavirus 229E Antibody.immunoglobulin G:Presence or Threshold:Point in time:Serum:Ordinal:Enzyme Immunoassay|Human coronavirus 229E Antibody.immunoglobulin G:Presence or Threshold:Point in time:Serum:Ordinal:Enzyme Immunoassay
C1544949|T201|LC|41002-7|LNC|Human coronavirus 229E IgG Ab [Presence] in Serum by Immunoassay|Human coronavirus 229E IgG Ab [Presence] in Serum by Immunoassay
C1544950|T201|DN|41003-5|LNC|HCoV 229E RNA NAA+probe Ql (Unsp spec)|HCoV 229E RNA NAA+probe Ql (Unsp spec)
C1544950|T201|OSN|41003-5|LNC|HCoV 229E RNA XXX Ql NAA+probe|HCoV 229E RNA XXX Ql NAA+probe
C1544950|T201|MTH_LN|41003-5|LNC|Human coronavirus 229E ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus 229E ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar
C1544950|T201|LC|41003-5|LNC|Human coronavirus 229E RNA [Presence] in Unspecified specimen by NAA with probe detection|Human coronavirus 229E RNA [Presence] in Unspecified specimen by NAA with probe detection
C1544950|T201|LN|41003-5|LNC|Human coronavirus 229E RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar|Human coronavirus 229E RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar
C1544951|T201|DN|41004-3|LNC|HCoV 229E Ag IF Ql (Unsp spec)|HCoV 229E Ag IF Ql (Unsp spec)
C1544951|T201|OSN|41004-3|LNC|HCoV 229E Ag XXX Ql IF|HCoV 229E Ag XXX Ql IF
C1544951|T201|LC|41004-3|LNC|Human coronavirus 229E Ag [Presence] in Unspecified specimen by Immunofluorescence|Human coronavirus 229E Ag [Presence] in Unspecified specimen by Immunofluorescence
C1544951|T201|LN|41004-3|LNC|Human coronavirus 229E Ag:PrThr:Pt:XXX:Ord:IF|Human coronavirus 229E Ag:PrThr:Pt:XXX:Ord:IF
C1544951|T201|MTH_LN|41004-3|LNC|Human coronavirus 229E Antigen:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:Immune Fluorescence|Human coronavirus 229E Antigen:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:Immune Fluorescence
C1544952|T201|DN|41005-0|LNC|HCoV NL63 RNA NAA+probe Ql (Unsp spec)|HCoV NL63 RNA NAA+probe Ql (Unsp spec)
C1544952|T201|OSN|41005-0|LNC|HCoV NL63 RNA XXX Ql NAA+probe|HCoV NL63 RNA XXX Ql NAA+probe
C1544952|T201|MTH_LN|41005-0|LNC|Human coronavirus NL63 ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus NL63 ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar
C1544952|T201|LC|41005-0|LNC|Human coronavirus NL63 RNA [Presence] in Unspecified specimen by NAA with probe detection|Human coronavirus NL63 RNA [Presence] in Unspecified specimen by NAA with probe detection
C1544952|T201|LN|41005-0|LNC|Human coronavirus NL63 RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar|Human coronavirus NL63 RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar
C1544953|T201|DN|41006-8|LNC|HCoV NL63 IgG IA Ql (S)|HCoV NL63 IgG IA Ql (S)
C1544953|T201|OSN|41006-8|LNC|HCoV NL63 IgG Ser Ql IA|HCoV NL63 IgG Ser Ql IA
C1544953|T201|LN|41006-8|LNC|Human coronavirus NL63 Ab.IgG:PrThr:Pt:Ser:Ord:IA|Human coronavirus NL63 Ab.IgG:PrThr:Pt:Ser:Ord:IA
C1544953|T201|MTH_LN|41006-8|LNC|Human coronavirus NL63 Antibody.immunoglobulin G:Presence or Threshold:Point in time:Serum:Ordinal:Enzyme Immunoassay|Human coronavirus NL63 Antibody.immunoglobulin G:Presence or Threshold:Point in time:Serum:Ordinal:Enzyme Immunoassay
C1544953|T201|LC|41006-8|LNC|Human coronavirus NL63 IgG Ab [Presence] in Serum by Immunoassay|Human coronavirus NL63 IgG Ab [Presence] in Serum by Immunoassay
C1544954|T201|DN|41007-6|LNC|HCoV OC43 Ag IF Ql (Unsp spec)|HCoV OC43 Ag IF Ql (Unsp spec)
C1544954|T201|OSN|41007-6|LNC|HCoV OC43 Ag XXX Ql IF|HCoV OC43 Ag XXX Ql IF
C1544954|T201|LC|41007-6|LNC|Human coronavirus OC43 Ag [Presence] in Unspecified specimen by Immunofluorescence|Human coronavirus OC43 Ag [Presence] in Unspecified specimen by Immunofluorescence
C1544954|T201|LN|41007-6|LNC|Human coronavirus OC43 Ag:PrThr:Pt:XXX:Ord:IF|Human coronavirus OC43 Ag:PrThr:Pt:XXX:Ord:IF
C1544954|T201|MTH_LN|41007-6|LNC|Human coronavirus OC43 Antigen:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:Immune Fluorescence|Human coronavirus OC43 Antigen:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:Immune Fluorescence
C1544955|T201|DN|41008-4|LNC|HCoV OC43 IgG IA Ql (S)|HCoV OC43 IgG IA Ql (S)
C1544955|T201|OSN|41008-4|LNC|HCoV OC43 IgG Ser Ql IA|HCoV OC43 IgG Ser Ql IA
C1544955|T201|LN|41008-4|LNC|Human coronavirus OC43 Ab.IgG:PrThr:Pt:Ser:Ord:IA|Human coronavirus OC43 Ab.IgG:PrThr:Pt:Ser:Ord:IA
C1544955|T201|MTH_LN|41008-4|LNC|Human coronavirus OC43 Antibody.immunoglobulin G:Presence or Threshold:Point in time:Serum:Ordinal:Enzyme Immunoassay|Human coronavirus OC43 Antibody.immunoglobulin G:Presence or Threshold:Point in time:Serum:Ordinal:Enzyme Immunoassay
C1544955|T201|LC|41008-4|LNC|Human coronavirus OC43 IgG Ab [Presence] in Serum by Immunoassay|Human coronavirus OC43 IgG Ab [Presence] in Serum by Immunoassay
C1544956|T201|DN|41009-2|LNC|HCoV OC43 RNA NAA+probe Ql (Unsp spec)|HCoV OC43 RNA NAA+probe Ql (Unsp spec)
C1544956|T201|OSN|41009-2|LNC|HCoV OC43 RNA XXX Ql NAA+probe|HCoV OC43 RNA XXX Ql NAA+probe
C1544956|T201|MTH_LN|41009-2|LNC|Human coronavirus OC43 ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus OC43 ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar
C1544956|T201|LC|41009-2|LNC|Human coronavirus OC43 RNA [Presence] in Unspecified specimen by NAA with probe detection|Human coronavirus OC43 RNA [Presence] in Unspecified specimen by NAA with probe detection
C1544956|T201|LN|41009-2|LNC|Human coronavirus OC43 RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar|Human coronavirus OC43 RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar
C1544960|T201|DN|41013-4|LNC|HCoV 229E IgG Ql (S)|HCoV 229E IgG Ql (S)
C1544960|T201|OSN|41013-4|LNC|HCoV 229E IgG Ser Ql|HCoV 229E IgG Ser Ql
C1544960|T201|LN|41013-4|LNC|Human coronavirus 229E Ab.IgG:PrThr:Pt:Ser:Ord|Human coronavirus 229E Ab.IgG:PrThr:Pt:Ser:Ord
C1544960|T201|MTH_LN|41013-4|LNC|Human coronavirus 229E Antibody.immunoglobulin G:Presence or Threshold:Point in time:Serum:Ordinal|Human coronavirus 229E Antibody.immunoglobulin G:Presence or Threshold:Point in time:Serum:Ordinal
C1544960|T201|LC|41013-4|LNC|Human coronavirus 229E IgG Ab [Presence] in Serum|Human coronavirus 229E IgG Ab [Presence] in Serum
C1544961|T201|DN|41014-2|LNC|HCoV NL63 IgG Ql (S)|HCoV NL63 IgG Ql (S)
C1544961|T201|OSN|41014-2|LNC|HCoV NL63 IgG Ser Ql|HCoV NL63 IgG Ser Ql
C1544961|T201|LN|41014-2|LNC|Human coronavirus NL63 Ab.IgG:PrThr:Pt:Ser:Ord|Human coronavirus NL63 Ab.IgG:PrThr:Pt:Ser:Ord
C1544961|T201|MTH_LN|41014-2|LNC|Human coronavirus NL63 Antibody.immunoglobulin G:Presence or Threshold:Point in time:Serum:Ordinal|Human coronavirus NL63 Antibody.immunoglobulin G:Presence or Threshold:Point in time:Serum:Ordinal
C1544961|T201|LC|41014-2|LNC|Human coronavirus NL63 IgG Ab [Presence] in Serum|Human coronavirus NL63 IgG Ab [Presence] in Serum
C1544962|T201|DN|41015-9|LNC|HCoV OC43 IgG Ql (S)|HCoV OC43 IgG Ql (S)
C1544962|T201|OSN|41015-9|LNC|HCoV OC43 IgG Ser Ql|HCoV OC43 IgG Ser Ql
C1544962|T201|LN|41015-9|LNC|Human coronavirus OC43 Ab.IgG:PrThr:Pt:Ser:Ord|Human coronavirus OC43 Ab.IgG:PrThr:Pt:Ser:Ord
C1544962|T201|MTH_LN|41015-9|LNC|Human coronavirus OC43 Antibody.immunoglobulin G:Presence or Threshold:Point in time:Serum:Ordinal|Human coronavirus OC43 Antibody.immunoglobulin G:Presence or Threshold:Point in time:Serum:Ordinal
C1544962|T201|LC|41015-9|LNC|Human coronavirus OC43 IgG Ab [Presence] in Serum|Human coronavirus OC43 IgG Ab [Presence] in Serum
C1545336|T116|SY|720062006|SNOMEDCT_US|Anti-Human coronavirus 229E IgG|Anti-Human coronavirus 229E IgG
C1545336|T129|SY|720062006|SNOMEDCT_US|Anti-Human coronavirus 229E IgG|Anti-Human coronavirus 229E IgG
C1545336|T116|LPN|LP38551-5|LNC|Human coronavirus 229E Ab.IgG|Human coronavirus 229E Ab.IgG
C1545336|T129|LPN|LP38551-5|LNC|Human coronavirus 229E Ab.IgG|Human coronavirus 229E Ab.IgG
C1545336|T116|CN|MTHU018542|LNC|Human coronavirus 229E Ab.IgG|Human coronavirus 229E Ab.IgG
C1545336|T129|CN|MTHU018542|LNC|Human coronavirus 229E Ab.IgG|Human coronavirus 229E Ab.IgG
C1545336|T116|MTH_CN|MTHU018542|LNC|Human coronavirus 229E Antibody.immunoglobulin G|Human coronavirus 229E Antibody.immunoglobulin G
C1545336|T129|MTH_CN|MTHU018542|LNC|Human coronavirus 229E Antibody.immunoglobulin G|Human coronavirus 229E Antibody.immunoglobulin G
C1545336|T116|PT|720062006|SNOMEDCT_US|Human coronavirus 229E IgG|Human coronavirus 229E IgG
C1545336|T129|PT|720062006|SNOMEDCT_US|Human coronavirus 229E IgG|Human coronavirus 229E IgG
C1545336|T116|SY|720062006|SNOMEDCT_US|Immunoglobulin G antibody to Human coronavirus 229E|Immunoglobulin G antibody to Human coronavirus 229E
C1545336|T129|SY|720062006|SNOMEDCT_US|Immunoglobulin G antibody to Human coronavirus 229E|Immunoglobulin G antibody to Human coronavirus 229E
C1545336|T116|FN|720062006|SNOMEDCT_US|Immunoglobulin G antibody to Human coronavirus 229E (substance)|Immunoglobulin G antibody to Human coronavirus 229E (substance)
C1545336|T129|FN|720062006|SNOMEDCT_US|Immunoglobulin G antibody to Human coronavirus 229E (substance)|Immunoglobulin G antibody to Human coronavirus 229E (substance)
C1545337|T114|MTH_CN|MTHU018544|LNC|Human coronavirus 229E ribonucleic acid|Human coronavirus 229E ribonucleic acid
C1545337|T114|LPN|LP38554-9|LNC|Human coronavirus 229E RNA|Human coronavirus 229E RNA
C1545337|T114|CN|MTHU018544|LNC|Human coronavirus 229E RNA|Human coronavirus 229E RNA
C1545337|T114|PT|707892006|SNOMEDCT_US|Human coronavirus 229E RNA|Human coronavirus 229E RNA
C1545337|T114|SY|707892006|SNOMEDCT_US|Ribonucleic acid of Human coronavirus 229E|Ribonucleic acid of Human coronavirus 229E
C1545337|T114|FN|707892006|SNOMEDCT_US|Ribonucleic acid of Human coronavirus 229E (substance)|Ribonucleic acid of Human coronavirus 229E (substance)
C1545338|T116|SY|720063001|SNOMEDCT_US|Anti-Human coronavirus NL63 IgG|Anti-Human coronavirus NL63 IgG
C1545338|T129|SY|720063001|SNOMEDCT_US|Anti-Human coronavirus NL63 IgG|Anti-Human coronavirus NL63 IgG
C1545338|T116|LPN|LP38555-6|LNC|Human coronavirus NL63 Ab.IgG|Human coronavirus NL63 Ab.IgG
C1545338|T129|LPN|LP38555-6|LNC|Human coronavirus NL63 Ab.IgG|Human coronavirus NL63 Ab.IgG
C1545338|T116|CN|MTHU018550|LNC|Human coronavirus NL63 Ab.IgG|Human coronavirus NL63 Ab.IgG
C1545338|T129|CN|MTHU018550|LNC|Human coronavirus NL63 Ab.IgG|Human coronavirus NL63 Ab.IgG
C1545338|T116|MTH_CN|MTHU018550|LNC|Human coronavirus NL63 Antibody.immunoglobulin G|Human coronavirus NL63 Antibody.immunoglobulin G
C1545338|T129|MTH_CN|MTHU018550|LNC|Human coronavirus NL63 Antibody.immunoglobulin G|Human coronavirus NL63 Antibody.immunoglobulin G
C1545338|T116|PT|720063001|SNOMEDCT_US|Human coronavirus NL63 IgG|Human coronavirus NL63 IgG
C1545338|T129|PT|720063001|SNOMEDCT_US|Human coronavirus NL63 IgG|Human coronavirus NL63 IgG
C1545338|T116|SY|720063001|SNOMEDCT_US|Immunoglobulin G antibody to Human coronavirus NL63|Immunoglobulin G antibody to Human coronavirus NL63
C1545338|T129|SY|720063001|SNOMEDCT_US|Immunoglobulin G antibody to Human coronavirus NL63|Immunoglobulin G antibody to Human coronavirus NL63
C1545338|T116|FN|720063001|SNOMEDCT_US|Immunoglobulin G antibody to Human coronavirus NL63 (substance)|Immunoglobulin G antibody to Human coronavirus NL63 (substance)
C1545338|T129|FN|720063001|SNOMEDCT_US|Immunoglobulin G antibody to Human coronavirus NL63 (substance)|Immunoglobulin G antibody to Human coronavirus NL63 (substance)
C1545339|T114|MTH_CN|MTHU018548|LNC|Human coronavirus NL63 ribonucleic acid|Human coronavirus NL63 ribonucleic acid
C1545339|T114|LPN|LP38557-2|LNC|Human coronavirus NL63 RNA|Human coronavirus NL63 RNA
C1545339|T114|CN|MTHU018548|LNC|Human coronavirus NL63 RNA|Human coronavirus NL63 RNA
C1545339|T114|PT|707894007|SNOMEDCT_US|Human coronavirus NL63 RNA|Human coronavirus NL63 RNA
C1545339|T114|SY|707894007|SNOMEDCT_US|Ribonucleic acid of Human coronavirus NL63|Ribonucleic acid of Human coronavirus NL63
C1545339|T114|FN|707894007|SNOMEDCT_US|Ribonucleic acid of Human coronavirus NL63 (substance)|Ribonucleic acid of Human coronavirus NL63 (substance)
C1545340|T116|SY|720064007|SNOMEDCT_US|Anti-Human coronavirus OC43 IgG|Anti-Human coronavirus OC43 IgG
C1545340|T129|SY|720064007|SNOMEDCT_US|Anti-Human coronavirus OC43 IgG|Anti-Human coronavirus OC43 IgG
C1545340|T116|LPN|LP38558-0|LNC|Human coronavirus OC43 Ab.IgG|Human coronavirus OC43 Ab.IgG
C1545340|T129|LPN|LP38558-0|LNC|Human coronavirus OC43 Ab.IgG|Human coronavirus OC43 Ab.IgG
C1545340|T116|CN|MTHU018554|LNC|Human coronavirus OC43 Ab.IgG|Human coronavirus OC43 Ab.IgG
C1545340|T129|CN|MTHU018554|LNC|Human coronavirus OC43 Ab.IgG|Human coronavirus OC43 Ab.IgG
C1545340|T116|MTH_CN|MTHU018554|LNC|Human coronavirus OC43 Antibody.immunoglobulin G|Human coronavirus OC43 Antibody.immunoglobulin G
C1545340|T129|MTH_CN|MTHU018554|LNC|Human coronavirus OC43 Antibody.immunoglobulin G|Human coronavirus OC43 Antibody.immunoglobulin G
C1545340|T116|PT|720064007|SNOMEDCT_US|Human coronavirus OC43 IgG|Human coronavirus OC43 IgG
C1545340|T129|PT|720064007|SNOMEDCT_US|Human coronavirus OC43 IgG|Human coronavirus OC43 IgG
C1545340|T116|SY|720064007|SNOMEDCT_US|Immunoglobulin G antibody to Human coronavirus OC43|Immunoglobulin G antibody to Human coronavirus OC43
C1545340|T129|SY|720064007|SNOMEDCT_US|Immunoglobulin G antibody to Human coronavirus OC43|Immunoglobulin G antibody to Human coronavirus OC43
C1545340|T116|FN|720064007|SNOMEDCT_US|Immunoglobulin G antibody to Human coronavirus OC43 (substance)|Immunoglobulin G antibody to Human coronavirus OC43 (substance)
C1545340|T129|FN|720064007|SNOMEDCT_US|Immunoglobulin G antibody to Human coronavirus OC43 (substance)|Immunoglobulin G antibody to Human coronavirus OC43 (substance)
C1545341|T116|SY|709346006|SNOMEDCT_US|Antigen of Human coronavirus OC43|Antigen of Human coronavirus OC43
C1545341|T129|SY|709346006|SNOMEDCT_US|Antigen of Human coronavirus OC43|Antigen of Human coronavirus OC43
C1545341|T116|FN|709346006|SNOMEDCT_US|Antigen of Human coronavirus OC43 (substance)|Antigen of Human coronavirus OC43 (substance)
C1545341|T129|FN|709346006|SNOMEDCT_US|Antigen of Human coronavirus OC43 (substance)|Antigen of Human coronavirus OC43 (substance)
C1545341|T116|LPN|LP38560-6|LNC|Human coronavirus OC43 Ag|Human coronavirus OC43 Ag
C1545341|T129|LPN|LP38560-6|LNC|Human coronavirus OC43 Ag|Human coronavirus OC43 Ag
C1545341|T116|CN|MTHU018552|LNC|Human coronavirus OC43 Ag|Human coronavirus OC43 Ag
C1545341|T129|CN|MTHU018552|LNC|Human coronavirus OC43 Ag|Human coronavirus OC43 Ag
C1545341|T116|PT|709346006|SNOMEDCT_US|Human coronavirus OC43 Ag|Human coronavirus OC43 Ag
C1545341|T129|PT|709346006|SNOMEDCT_US|Human coronavirus OC43 Ag|Human coronavirus OC43 Ag
C1545341|T116|SY|709346006|SNOMEDCT_US|Human coronavirus OC43 antigen|Human coronavirus OC43 antigen
C1545341|T129|SY|709346006|SNOMEDCT_US|Human coronavirus OC43 antigen|Human coronavirus OC43 antigen
C1545341|T116|MTH_CN|MTHU018552|LNC|Human coronavirus OC43 Antigen|Human coronavirus OC43 Antigen
C1545341|T129|MTH_CN|MTHU018552|LNC|Human coronavirus OC43 Antigen|Human coronavirus OC43 Antigen
C1545342|T114|MTH_CN|MTHU018556|LNC|Human coronavirus OC43 ribonucleic acid|Human coronavirus OC43 ribonucleic acid
C1545342|T114|LPN|LP38561-4|LNC|Human coronavirus OC43 RNA|Human coronavirus OC43 RNA
C1545342|T114|CN|MTHU018556|LNC|Human coronavirus OC43 RNA|Human coronavirus OC43 RNA
C1545342|T114|PT|707895008|SNOMEDCT_US|Human coronavirus OC43 RNA|Human coronavirus OC43 RNA
C1545342|T114|SY|707895008|SNOMEDCT_US|Ribonucleic acid of Human coronavirus OC43|Ribonucleic acid of Human coronavirus OC43
C1545342|T114|FN|707895008|SNOMEDCT_US|Ribonucleic acid of Human coronavirus OC43 (substance)|Ribonucleic acid of Human coronavirus OC43 (substance)
C1545343|T114|MTH_CN|MTHU062870|LNC|Human Coronavirus ribonucleic acid|Human Coronavirus ribonucleic acid
C1545343|T114|MTH_CN|MTHU018540|LNC|Human coronavirus ribonucleic acid|Human coronavirus ribonucleic acid
C1545343|T114|LPN|LP38550-7|LNC|Human coronavirus RNA|Human coronavirus RNA
C1545343|T114|CN|MTHU018540|LNC|Human coronavirus RNA|Human coronavirus RNA
C1545343|T114|PT|720112004|SNOMEDCT_US|Human coronavirus RNA|Human coronavirus RNA
C1545343|T114|CN|MTHU062870|LNC|Human Coronavirus RNA|Human Coronavirus RNA
C1545343|T114|SY|720112004|SNOMEDCT_US|Ribonucleic acid of Human coronavirus|Ribonucleic acid of Human coronavirus
C1545343|T114|FN|720112004|SNOMEDCT_US|Ribonucleic acid of Human coronavirus (substance)|Ribonucleic acid of Human coronavirus (substance)
C1546317|T116|SY|709344009|SNOMEDCT_US|Antigen of Human coronavirus 229E|Antigen of Human coronavirus 229E
C1546317|T129|SY|709344009|SNOMEDCT_US|Antigen of Human coronavirus 229E|Antigen of Human coronavirus 229E
C1546317|T116|FN|709344009|SNOMEDCT_US|Antigen of Human coronavirus 229E (substance)|Antigen of Human coronavirus 229E (substance)
C1546317|T129|FN|709344009|SNOMEDCT_US|Antigen of Human coronavirus 229E (substance)|Antigen of Human coronavirus 229E (substance)
C1546317|T116|LPN|LP38553-1|LNC|Human coronavirus 229E Ag|Human coronavirus 229E Ag
C1546317|T129|LPN|LP38553-1|LNC|Human coronavirus 229E Ag|Human coronavirus 229E Ag
C1546317|T116|CN|MTHU018546|LNC|Human coronavirus 229E Ag|Human coronavirus 229E Ag
C1546317|T129|CN|MTHU018546|LNC|Human coronavirus 229E Ag|Human coronavirus 229E Ag
C1546317|T116|PT|709344009|SNOMEDCT_US|Human coronavirus 229E Ag|Human coronavirus 229E Ag
C1546317|T129|PT|709344009|SNOMEDCT_US|Human coronavirus 229E Ag|Human coronavirus 229E Ag
C1546317|T116|SY|709344009|SNOMEDCT_US|Human coronavirus 229E antigen|Human coronavirus 229E antigen
C1546317|T129|SY|709344009|SNOMEDCT_US|Human coronavirus 229E antigen|Human coronavirus 229E antigen
C1546317|T116|PN|NOCODE|MTH|Human coronavirus 229E antigen|Human coronavirus 229E antigen
C1546317|T129|PN|NOCODE|MTH|Human coronavirus 229E antigen|Human coronavirus 229E antigen
C1546317|T116|MTH_CN|MTHU018546|LNC|Human coronavirus 229E Antigen|Human coronavirus 229E Antigen
C1546317|T129|MTH_CN|MTHU018546|LNC|Human coronavirus 229E Antigen|Human coronavirus 229E Antigen
C1567331|T116|NM|C498660|MSH|protein C, SARS virus|protein C, SARS virus
C1567331|T129|NM|C498660|MSH|protein C, SARS virus|protein C, SARS virus
C1567331|T116|CE|C498660|MSH|protein C, severe acute respiratory syndrome virus|protein C, severe acute respiratory syndrome virus
C1567331|T129|CE|C498660|MSH|protein C, severe acute respiratory syndrome virus|protein C, severe acute respiratory syndrome virus
C1570531|T116|NM|C501689|MSH|E protein, SARS coronavirus|E protein, SARS coronavirus
C1570531|T123|NM|C501689|MSH|E protein, SARS coronavirus|E protein, SARS coronavirus
C1570531|T116|CE|C501689|MSH|protein E, SARS coronavirus|protein E, SARS coronavirus
C1570531|T123|CE|C501689|MSH|protein E, SARS coronavirus|protein E, SARS coronavirus
C1570531|T116|CE|C501689|MSH|protein E, SCoVE|protein E, SCoVE
C1570531|T123|CE|C501689|MSH|protein E, SCoVE|protein E, SCoVE
C1615569|T116|NM|C504965|MSH|Nps13 protein, SARS-CoV|Nps13 protein, SARS-CoV
C1615569|T126|NM|C504965|MSH|Nps13 protein, SARS-CoV|Nps13 protein, SARS-CoV
C1615569|T116|CE|C504965|MSH|SARS-VoV nsp13 protein, SARS-associated coronavirus|SARS-VoV nsp13 protein, SARS-associated coronavirus
C1615569|T126|CE|C504965|MSH|SARS-VoV nsp13 protein, SARS-associated coronavirus|SARS-VoV nsp13 protein, SARS-associated coronavirus
C1621889|T116|PCE|C067997|MSH|M protein, Human coronavirus OC43|M protein, Human coronavirus OC43
C1621889|T123|PCE|C067997|MSH|M protein, Human coronavirus OC43|M protein, Human coronavirus OC43
C1621889|T116|CE|C067997|MSH|membrane protein, Human coronavirus OC43|membrane protein, Human coronavirus OC43
C1621889|T123|CE|C067997|MSH|membrane protein, Human coronavirus OC43|membrane protein, Human coronavirus OC43
C1623644|T116|SY|709345005|SNOMEDCT_US|Antigen of Human coronavirus|Antigen of Human coronavirus
C1623644|T129|SY|709345005|SNOMEDCT_US|Antigen of Human coronavirus|Antigen of Human coronavirus
C1623644|T116|FN|709345005|SNOMEDCT_US|Antigen of Human coronavirus (substance)|Antigen of Human coronavirus (substance)
C1623644|T129|FN|709345005|SNOMEDCT_US|Antigen of Human coronavirus (substance)|Antigen of Human coronavirus (substance)
C1623644|T116|LPN|LP38548-1|LNC|Human coronavirus Ag|Human coronavirus Ag
C1623644|T129|LPN|LP38548-1|LNC|Human coronavirus Ag|Human coronavirus Ag
C1623644|T116|CN|MTHU018678|LNC|Human coronavirus Ag|Human coronavirus Ag
C1623644|T129|CN|MTHU018678|LNC|Human coronavirus Ag|Human coronavirus Ag
C1623644|T116|PT|709345005|SNOMEDCT_US|Human coronavirus Ag|Human coronavirus Ag
C1623644|T129|PT|709345005|SNOMEDCT_US|Human coronavirus Ag|Human coronavirus Ag
C1623644|T116|SY|709345005|SNOMEDCT_US|Human coronavirus antigen|Human coronavirus antigen
C1623644|T129|SY|709345005|SNOMEDCT_US|Human coronavirus antigen|Human coronavirus antigen
C1623644|T116|MTH_CN|MTHU018678|LNC|Human coronavirus Antigen|Human coronavirus Antigen
C1623644|T129|MTH_CN|MTHU018678|LNC|Human coronavirus Antigen|Human coronavirus Antigen
C1625777|T034|LPN|LP38549-9|LNC|Human coronavirus identified|Human coronavirus identified
C1625777|T034|CN|MTHU018680|LNC|Human coronavirus identified|Human coronavirus identified
C1627946|T116|SY|720294006|SNOMEDCT_US|Anti-SARS coronavirus IgM|Anti-SARS coronavirus IgM
C1627946|T129|SY|720294006|SNOMEDCT_US|Anti-SARS coronavirus IgM|Anti-SARS coronavirus IgM
C1627946|T116|SY|720294006|SNOMEDCT_US|Immunoglobulin M antibody to SARS coronavirus|Immunoglobulin M antibody to SARS coronavirus
C1627946|T129|SY|720294006|SNOMEDCT_US|Immunoglobulin M antibody to SARS coronavirus|Immunoglobulin M antibody to SARS coronavirus
C1627946|T116|SY|720294006|SNOMEDCT_US|Immunoglobulin M antibody to severe acute respiratory syndrome-related coronavirus|Immunoglobulin M antibody to severe acute respiratory syndrome-related coronavirus
C1627946|T129|SY|720294006|SNOMEDCT_US|Immunoglobulin M antibody to severe acute respiratory syndrome-related coronavirus|Immunoglobulin M antibody to severe acute respiratory syndrome-related coronavirus
C1627946|T116|FN|720294006|SNOMEDCT_US|Immunoglobulin M antibody to severe acute respiratory syndrome-related coronavirus (substance)|Immunoglobulin M antibody to severe acute respiratory syndrome-related coronavirus (substance)
C1627946|T129|FN|720294006|SNOMEDCT_US|Immunoglobulin M antibody to severe acute respiratory syndrome-related coronavirus (substance)|Immunoglobulin M antibody to severe acute respiratory syndrome-related coronavirus (substance)
C1627946|T116|LPN|LP39709-8|LNC|SARS coronavirus Ab.IgM|SARS coronavirus Ab.IgM
C1627946|T129|LPN|LP39709-8|LNC|SARS coronavirus Ab.IgM|SARS coronavirus Ab.IgM
C1627946|T116|CN|MTHU018887|LNC|SARS coronavirus Ab.IgM|SARS coronavirus Ab.IgM
C1627946|T129|CN|MTHU018887|LNC|SARS coronavirus Ab.IgM|SARS coronavirus Ab.IgM
C1627946|T116|MTH_CN|MTHU018887|LNC|SARS coronavirus Antibody.immunoglobulin M|SARS coronavirus Antibody.immunoglobulin M
C1627946|T129|MTH_CN|MTHU018887|LNC|SARS coronavirus Antibody.immunoglobulin M|SARS coronavirus Antibody.immunoglobulin M
C1627946|T116|PT|720294006|SNOMEDCT_US|SARS coronavirus IgM|SARS coronavirus IgM
C1627946|T129|PT|720294006|SNOMEDCT_US|SARS coronavirus IgM|SARS coronavirus IgM
C1628478|T116|SY|720293000|SNOMEDCT_US|Anti-SARS coronavirus IgG|Anti-SARS coronavirus IgG
C1628478|T129|SY|720293000|SNOMEDCT_US|Anti-SARS coronavirus IgG|Anti-SARS coronavirus IgG
C1628478|T116|SY|720293000|SNOMEDCT_US|Immunoglobulin G antibody to SARS coronavirus|Immunoglobulin G antibody to SARS coronavirus
C1628478|T129|SY|720293000|SNOMEDCT_US|Immunoglobulin G antibody to SARS coronavirus|Immunoglobulin G antibody to SARS coronavirus
C1628478|T116|SY|720293000|SNOMEDCT_US|Immunoglobulin G antibody to severe acute respiratory syndrome-related coronavirus|Immunoglobulin G antibody to severe acute respiratory syndrome-related coronavirus
C1628478|T129|SY|720293000|SNOMEDCT_US|Immunoglobulin G antibody to severe acute respiratory syndrome-related coronavirus|Immunoglobulin G antibody to severe acute respiratory syndrome-related coronavirus
C1628478|T116|FN|720293000|SNOMEDCT_US|Immunoglobulin G antibody to severe acute respiratory syndrome-related coronavirus (substance)|Immunoglobulin G antibody to severe acute respiratory syndrome-related coronavirus (substance)
C1628478|T129|FN|720293000|SNOMEDCT_US|Immunoglobulin G antibody to severe acute respiratory syndrome-related coronavirus (substance)|Immunoglobulin G antibody to severe acute respiratory syndrome-related coronavirus (substance)
C1628478|T116|LPN|LP39707-2|LNC|SARS coronavirus Ab.IgG|SARS coronavirus Ab.IgG
C1628478|T129|LPN|LP39707-2|LNC|SARS coronavirus Ab.IgG|SARS coronavirus Ab.IgG
C1628478|T116|CN|MTHU018687|LNC|SARS coronavirus Ab.IgG|SARS coronavirus Ab.IgG
C1628478|T129|CN|MTHU018687|LNC|SARS coronavirus Ab.IgG|SARS coronavirus Ab.IgG
C1628478|T116|MTH_CN|MTHU018687|LNC|SARS coronavirus Antibody.immunoglobulin G|SARS coronavirus Antibody.immunoglobulin G
C1628478|T129|MTH_CN|MTHU018687|LNC|SARS coronavirus Antibody.immunoglobulin G|SARS coronavirus Antibody.immunoglobulin G
C1628478|T116|PT|720293000|SNOMEDCT_US|SARS coronavirus IgG|SARS coronavirus IgG
C1628478|T129|PT|720293000|SNOMEDCT_US|SARS coronavirus IgG|SARS coronavirus IgG
C1628999|T114|SY|707784009|SNOMEDCT_US|Ribonucleic acid of Severe acute respiratory syndrome coronavirus|Ribonucleic acid of Severe acute respiratory syndrome coronavirus
C1628999|T114|FN|707784009|SNOMEDCT_US|Ribonucleic acid of Severe acute respiratory syndrome coronavirus (substance)|Ribonucleic acid of Severe acute respiratory syndrome coronavirus (substance)
C1628999|T114|SY|707784009|SNOMEDCT_US|SARS (severe acute respiratory syndrome) coronavirus RNA|SARS (severe acute respiratory syndrome) coronavirus RNA
C1628999|T114|MTH_CN|MTHU018684|LNC|SARS coronavirus ribonucleic acid|SARS coronavirus ribonucleic acid
C1628999|T114|LPN|LP39711-4|LNC|SARS coronavirus RNA|SARS coronavirus RNA
C1628999|T114|OP|707784009|SNOMEDCT_US|SARS coronavirus RNA|SARS coronavirus RNA
C1628999|T114|CN|MTHU018684|LNC|SARS coronavirus RNA|SARS coronavirus RNA
C1628999|T114|PT|707784009|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus RNA|Severe acute respiratory syndrome coronavirus RNA
C1631820|T201|LN|42957-1|LNC|SARS coronavirus Ab.IgG:PrThr:Pt:Ser:Ord|SARS coronavirus Ab.IgG:PrThr:Pt:Ser:Ord
C1631820|T201|MTH_LN|42957-1|LNC|SARS coronavirus Antibody.immunoglobulin G:Presence or Threshold:Point in time:Serum:Ordinal|SARS coronavirus Antibody.immunoglobulin G:Presence or Threshold:Point in time:Serum:Ordinal
C1631820|T201|LC|42957-1|LNC|SARS coronavirus IgG Ab [Presence] in Serum|SARS coronavirus IgG Ab [Presence] in Serum
C1631820|T201|DN|42957-1|LNC|SARS coronavirus IgG Ql (S)|SARS coronavirus IgG Ql (S)
C1631820|T201|OSN|42957-1|LNC|SARS-CoV IgG Ser Ql|SARS-CoV IgG Ser Ql
C1632362|T201|LN|42956-3|LNC|SARS coronavirus Ab.IgM:PrThr:Pt:Ser:Ord|SARS coronavirus Ab.IgM:PrThr:Pt:Ser:Ord
C1632362|T201|MTH_LN|42956-3|LNC|SARS coronavirus Antibody.immunoglobulin M:Presence or Threshold:Point in time:Serum:Ordinal|SARS coronavirus Antibody.immunoglobulin M:Presence or Threshold:Point in time:Serum:Ordinal
C1632362|T201|LC|42956-3|LNC|SARS coronavirus IgM Ab [Presence] in Serum|SARS coronavirus IgM Ab [Presence] in Serum
C1632362|T201|DN|42956-3|LNC|SARS coronavirus IgM Ql (S)|SARS coronavirus IgM Ql (S)
C1632362|T201|OSN|42956-3|LNC|SARS-CoV IgM Ser Ql|SARS-CoV IgM Ser Ql
C1641503|T201|DN|41453-2|LNC|HCoV Ag IF Ql (Unsp spec)|HCoV Ag IF Ql (Unsp spec)
C1641503|T201|OSN|41453-2|LNC|HCoV Ag XXX Ql IF|HCoV Ag XXX Ql IF
C1641503|T201|LC|41453-2|LNC|Human coronavirus Ag [Presence] in Unspecified specimen by Immunofluorescence|Human coronavirus Ag [Presence] in Unspecified specimen by Immunofluorescence
C1641503|T201|LN|41453-2|LNC|Human coronavirus Ag:PrThr:Pt:XXX:Ord:IF|Human coronavirus Ag:PrThr:Pt:XXX:Ord:IF
C1641503|T201|MTH_LN|41453-2|LNC|Human coronavirus Antigen:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:Immune Fluorescence|Human coronavirus Antigen:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:Immune Fluorescence
C1642052|T201|MTH_LN|41458-1|LNC|SARS coronavirus ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar|SARS coronavirus ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar
C1642052|T201|LC|41458-1|LNC|SARS coronavirus RNA [Presence] in Unspecified specimen by NAA with probe detection|SARS coronavirus RNA [Presence] in Unspecified specimen by NAA with probe detection
C1642052|T201|DN|41458-1|LNC|SARS coronavirus RNA NAA+probe Ql (Unsp spec)|SARS coronavirus RNA NAA+probe Ql (Unsp spec)
C1642052|T201|LN|41458-1|LNC|SARS coronavirus RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar|SARS coronavirus RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar
C1642052|T201|OSN|41458-1|LNC|SARS-CoV RNA XXX Ql NAA+probe|SARS-CoV RNA XXX Ql NAA+probe
C1642546|T201|DN|41454-0|LNC|HCoV identified Nom (Unsp spec)|HCoV identified Nom (Unsp spec)
C1642546|T201|OSN|41454-0|LNC|HCoV XXX|HCoV XXX
C1642546|T201|LC|41454-0|LNC|Human coronavirus identified in Unspecified specimen|Human coronavirus identified in Unspecified specimen
C1642546|T201|MTH_LN|41454-0|LNC|Human coronavirus identified:Presence or Identity:Point in time:To be specified in another part of the message:Nominal|Human coronavirus identified:Presence or Identity:Point in time:To be specified in another part of the message:Nominal
C1642546|T201|LN|41454-0|LNC|Human coronavirus identified:Prid:Pt:XXX:Nom|Human coronavirus identified:Prid:Pt:XXX:Nom
C1642839|T005|LA|LA19210-6|LNC|HK1|HK1
C1642839|T005|OAP|417819004|SNOMEDCT_US|Human coronavirus HK1|Human coronavirus HK1
C1642839|T005|PN|NOCODE|MTH|Human coronavirus HK1|Human coronavirus HK1
C1642839|T005|OAF|417819004|SNOMEDCT_US|Human coronavirus HK1 (organism)|Human coronavirus HK1 (organism)
C1643178|T201|LC|41459-9|LNC|SARS coronavirus [Presence] in Unspecified specimen|SARS coronavirus [Presence] in Unspecified specimen
C1643178|T201|DN|41459-9|LNC|SARS coronavirus Ql (Unsp spec)|SARS coronavirus Ql (Unsp spec)
C1643178|T201|MTH_LN|41459-9|LNC|SARS coronavirus:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal|SARS coronavirus:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal
C1643178|T201|LN|41459-9|LNC|SARS coronavirus:PrThr:Pt:XXX:Ord|SARS coronavirus:PrThr:Pt:XXX:Ord
C1643178|T201|OSN|41459-9|LNC|SARS-CoV XXX Ql|SARS-CoV XXX Ql
C1643179|T201|LN|41460-7|LNC|SARS coronavirus Ab.IgG:PrThr:Pt:Ser:Ord:IA|SARS coronavirus Ab.IgG:PrThr:Pt:Ser:Ord:IA
C1643179|T201|MTH_LN|41460-7|LNC|SARS coronavirus Antibody.immunoglobulin G:Presence or Threshold:Point in time:Serum:Ordinal:Enzyme Immunoassay|SARS coronavirus Antibody.immunoglobulin G:Presence or Threshold:Point in time:Serum:Ordinal:Enzyme Immunoassay
C1643179|T201|LC|41460-7|LNC|SARS coronavirus IgG Ab [Presence] in Serum by Immunoassay|SARS coronavirus IgG Ab [Presence] in Serum by Immunoassay
C1643179|T201|DN|41460-7|LNC|SARS coronavirus IgG IA Ql (S)|SARS coronavirus IgG IA Ql (S)
C1643179|T201|OSN|41460-7|LNC|SARS-CoV IgG Ser Ql IA|SARS-CoV IgG Ser Ql IA
C1654324|T201|LN|41991-1|LNC|SARS coronavirus Ab.IgM:PrThr:Pt:Ser:Ord:IA|SARS coronavirus Ab.IgM:PrThr:Pt:Ser:Ord:IA
C1654324|T201|MTH_LN|41991-1|LNC|SARS coronavirus Antibody.immunoglobulin M:Presence or Threshold:Point in time:Serum:Ordinal:Enzyme Immunoassay|SARS coronavirus Antibody.immunoglobulin M:Presence or Threshold:Point in time:Serum:Ordinal:Enzyme Immunoassay
C1654324|T201|LC|41991-1|LNC|SARS coronavirus IgM Ab [Presence] in Serum by Immunoassay|SARS coronavirus IgM Ab [Presence] in Serum by Immunoassay
C1654324|T201|DN|41991-1|LNC|SARS coronavirus IgM IA Ql (S)|SARS coronavirus IgM IA Ql (S)
C1654324|T201|OSN|41991-1|LNC|SARS-CoV IgM Ser Ql IA|SARS-CoV IgM Ser Ql IA
C1676985|T005|ET|D000073640|MSH|HCoV-HKU1|HCoV-HKU1
C1676985|T005|LPN|LP111518-9|LNC|Human coronavirus HKU1|Human coronavirus HKU1
C1676985|T005|PEP|D000073640|MSH|Human coronavirus HKU1|Human coronavirus HKU1
C1676985|T005|PT|697942007|SNOMEDCT_US|Human coronavirus HKU1|Human coronavirus HKU1
C1676985|T005|FN|697942007|SNOMEDCT_US|Human coronavirus HKU1 (organism)|Human coronavirus HKU1 (organism)
C1689295|T116|CE|C507223|MSH|ORF-6 protein, SARS coronovirus|ORF-6 protein, SARS coronovirus
C1689295|T123|CE|C507223|MSH|ORF-6 protein, SARS coronovirus|ORF-6 protein, SARS coronovirus
C1689295|T116|NM|C507223|MSH|protein 6, SARS virus|protein 6, SARS virus
C1689295|T123|NM|C507223|MSH|protein 6, SARS virus|protein 6, SARS virus
C1689295|T116|CE|C507223|MSH|SARS-CoV ORF6 protein|SARS-CoV ORF6 protein
C1689295|T123|CE|C507223|MSH|SARS-CoV ORF6 protein|SARS-CoV ORF6 protein
C1689295|T116|CE|C507223|MSH|X3 protein, SARS-CoV|X3 protein, SARS-CoV
C1689295|T123|CE|C507223|MSH|X3 protein, SARS-CoV|X3 protein, SARS-CoV
C1718836|T116|LPN|LP38552-3|LNC|Human coronavirus 229E Ab|Human coronavirus 229E Ab
C1718836|T129|LPN|LP38552-3|LNC|Human coronavirus 229E Ab|Human coronavirus 229E Ab
C1718837|T116|LPN|LP38556-4|LNC|Human coronavirus NL63 Ab|Human coronavirus NL63 Ab
C1718837|T129|LPN|LP38556-4|LNC|Human coronavirus NL63 Ab|Human coronavirus NL63 Ab
C1718953|T116|SY|709904008|SNOMEDCT_US|Anti-Severe acute respiratory syndrome coronavirus antibody|Anti-Severe acute respiratory syndrome coronavirus antibody
C1718953|T129|SY|709904008|SNOMEDCT_US|Anti-Severe acute respiratory syndrome coronavirus antibody|Anti-Severe acute respiratory syndrome coronavirus antibody
C1718953|T116|SY|709904008|SNOMEDCT_US|Antibody to Severe acute respiratory syndrome coronavirus|Antibody to Severe acute respiratory syndrome coronavirus
C1718953|T129|SY|709904008|SNOMEDCT_US|Antibody to Severe acute respiratory syndrome coronavirus|Antibody to Severe acute respiratory syndrome coronavirus
C1718953|T116|FN|709904008|SNOMEDCT_US|Antibody to Severe acute respiratory syndrome coronavirus (substance)|Antibody to Severe acute respiratory syndrome coronavirus (substance)
C1718953|T129|FN|709904008|SNOMEDCT_US|Antibody to Severe acute respiratory syndrome coronavirus (substance)|Antibody to Severe acute respiratory syndrome coronavirus (substance)
C1718953|T116|LPN|LP39708-0|LNC|SARS coronavirus Ab|SARS coronavirus Ab
C1718953|T129|LPN|LP39708-0|LNC|SARS coronavirus Ab|SARS coronavirus Ab
C1718953|T116|CN|MTHU036263|LNC|SARS coronavirus Ab|SARS coronavirus Ab
C1718953|T129|CN|MTHU036263|LNC|SARS coronavirus Ab|SARS coronavirus Ab
C1718953|T116|SY|709904008|SNOMEDCT_US|SARS coronavirus Ab|SARS coronavirus Ab
C1718953|T129|SY|709904008|SNOMEDCT_US|SARS coronavirus Ab|SARS coronavirus Ab
C1718953|T116|MTH_CN|MTHU036263|LNC|SARS coronavirus Antibody|SARS coronavirus Antibody
C1718953|T129|MTH_CN|MTHU036263|LNC|SARS coronavirus Antibody|SARS coronavirus Antibody
C1718953|T116|PT|709904008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Ab|Severe acute respiratory syndrome coronavirus Ab
C1718953|T129|PT|709904008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Ab|Severe acute respiratory syndrome coronavirus Ab
C1718953|T116|SY|709904008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus antibody|Severe acute respiratory syndrome coronavirus antibody
C1718953|T129|SY|709904008|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus antibody|Severe acute respiratory syndrome coronavirus antibody
C1719193|T116|LPN|LP38559-8|LNC|Human coronavirus OC43 Ab|Human coronavirus OC43 Ab
C1719193|T129|LPN|LP38559-8|LNC|Human coronavirus OC43 Ab|Human coronavirus OC43 Ab
C1722447|T116|NM|C510959|MSH|nonstructural protein 3, SARS coronovirus|nonstructural protein 3, SARS coronovirus
C1722447|T126|NM|C510959|MSH|nonstructural protein 3, SARS coronovirus|nonstructural protein 3, SARS coronovirus
C1722447|T116|CE|C510959|MSH|Nsp3 protein, SARS-CoV|Nsp3 protein, SARS-CoV
C1722447|T126|CE|C510959|MSH|Nsp3 protein, SARS-CoV|Nsp3 protein, SARS-CoV
C1722448|T116|NM|C510960|MSH|nonstructural protein 15, SARS coronovirus|nonstructural protein 15, SARS coronovirus
C1722448|T126|NM|C510960|MSH|nonstructural protein 15, SARS coronovirus|nonstructural protein 15, SARS coronovirus
C1722448|T116|CE|C510960|MSH|Nsp15 protein, SARS-CoV|Nsp15 protein, SARS-CoV
C1722448|T126|CE|C510960|MSH|Nsp15 protein, SARS-CoV|Nsp15 protein, SARS-CoV
C1737633|T130|ET|31-988|UMD|Reagents, Molecular Assay, Infection, Virus, Severe Acute Respiratory Syndrome Coronavirus, RNA|Reagents, Molecular Assay, Infection, Virus, Severe Acute Respiratory Syndrome Coronavirus, RNA
C1740657|T130|ET|32-608|UMD|Reagents, Serology, Virus, Severe Acute Respiratory Syndrome Coronavirus, IgG Antibody|Reagents, Serology, Virus, Severe Acute Respiratory Syndrome Coronavirus, IgG Antibody
C1852539|T033|PN|NOCODE|MTH|CORONAVIRUS 229E SUSCEPTIBILITY|CORONAVIRUS 229E SUSCEPTIBILITY
C1852539|T033|PT|HP:0005396|HPO|Susceptibility to coronavirus 229e|Susceptibility to coronavirus 229e
C1870542|T116|NM|C515313|MSH|ORF3A protein, SARS coronavirus|ORF3A protein, SARS coronavirus
C1870542|T123|NM|C515313|MSH|ORF3A protein, SARS coronavirus|ORF3A protein, SARS coronavirus
C1870542|T116|CE|C515313|MSH|ORF3A protein, SARS-CoV|ORF3A protein, SARS-CoV
C1870542|T123|CE|C515313|MSH|ORF3A protein, SARS-CoV|ORF3A protein, SARS-CoV
C1871553|T116|CE|C515314|MSH|accessory protein 7b, SARS coronavirus|accessory protein 7b, SARS coronavirus
C1871553|T123|CE|C515314|MSH|accessory protein 7b, SARS coronavirus|accessory protein 7b, SARS coronavirus
C1871553|T116|NM|C515314|MSH|ORF7b protein, SARS coronavirus|ORF7b protein, SARS coronavirus
C1871553|T123|NM|C515314|MSH|ORF7b protein, SARS coronavirus|ORF7b protein, SARS coronavirus
C1958909|T116|NM|C521592|MSH|Nsp1 protein, SARS coronavirus|Nsp1 protein, SARS coronavirus
C1958909|T126|NM|C521592|MSH|Nsp1 protein, SARS coronavirus|Nsp1 protein, SARS coronavirus
C1958909|T116|CE|C521592|MSH|Nsp1 protein, SARS-CoV|Nsp1 protein, SARS-CoV
C1958909|T126|CE|C521592|MSH|Nsp1 protein, SARS-CoV|Nsp1 protein, SARS-CoV
C2003364|T116|NM|C525596|MSH|nsp14 protein, SARS coronavirus|nsp14 protein, SARS coronavirus
C2022391|T034|PT|19504|MEDCIN|nasopharyngeal culture coronavirus|nasopharyngeal culture coronavirus
C2022391|T034|FN|19504|MEDCIN|nasopharyngeal culture coronavirus (lab test)|nasopharyngeal culture coronavirus (lab test)
C2207719|T059|SY|223662|MEDCIN|serum PCR for SARS|serum PCR for SARS
C2207719|T059|SY|223662|MEDCIN|serum polymerase chain reactions for SARS (available july, 2|serum polymerase chain reactions for SARS (available july, 2
C2207719|T059|PT|223662|MEDCIN|serum SARS coronavirus detection by polymerase chain reaction test|serum SARS coronavirus detection by polymerase chain reaction test
C2207719|T059|FN|223662|MEDCIN|serum SARS coronavirus detection by polymerase chain reaction test (lab test)|serum SARS coronavirus detection by polymerase chain reaction test (lab test)
C2229919|T047|SY|272883|MEDCIN|SARS pneumonia|SARS pneumonia
C2229919|T047|PT|272883|MEDCIN|severe acute respiratory syndrome (SARS) pneumonia|severe acute respiratory syndrome (SARS) pneumonia
C2229919|T047|FN|272883|MEDCIN|severe acute respiratory syndrome (SARS) pneumonia (diagnosis)|severe acute respiratory syndrome (SARS) pneumonia (diagnosis)
C2321692|T033|PT|321197|MEDCIN|left tonsil culture for coronavirus|left tonsil culture for coronavirus
C2321692|T033|FN|321197|MEDCIN|left tonsil culture for coronavirus (lab test)|left tonsil culture for coronavirus (lab test)
C2322051|T033|PT|321156|MEDCIN|right tonsil culture for coronavirus|right tonsil culture for coronavirus
C2322051|T033|FN|321156|MEDCIN|right tonsil culture for coronavirus (lab test)|right tonsil culture for coronavirus (lab test)
C2604739|T116|PCE|C479931|MSH|Nsp5, SARS coronavirus|Nsp5, SARS coronavirus
C2604739|T126|PCE|C479931|MSH|Nsp5, SARS coronavirus|Nsp5, SARS coronavirus
C2718208|T201|OLC|23375-9|LNC|Deprecated Porcine respiratory coronavirus Ab [Presence] in Serum|Deprecated Porcine respiratory coronavirus Ab [Presence] in Serum
C2718208|T201|PN|NOCODE|MTH|Deprecated Porcine respiratory coronavirus Ab [Presence] in Serum|Deprecated Porcine respiratory coronavirus Ab [Presence] in Serum
C2718208|T201|OOSN|23375-9|LNC|Deprecated PRCoV Ab Ser Ql|Deprecated PRCoV Ab Ser Ql
C2718208|T201|DN|23375-9|LNC|Porcine respiratory coronavirus Ab Ql (S)|Porcine respiratory coronavirus Ab Ql (S)
C2718208|T201|LO|23375-9|LNC|Porcine respiratory coronavirus Ab:ACnc:Pt:Ser:Ord|Porcine respiratory coronavirus Ab:ACnc:Pt:Ser:Ord
C2718208|T201|MTH_LO|23375-9|LNC|Porcine respiratory coronavirus Antibody:Arbitrary Concentration:Point in time:Serum:Ordinal|Porcine respiratory coronavirus Antibody:Arbitrary Concentration:Point in time:Serum:Ordinal
C2733460|T051|PT|444482005|SNOMEDCT_US|Exposure to severe acute respiratory syndrome coronavirus|Exposure to severe acute respiratory syndrome coronavirus
C2733460|T051|OP|444482005|SNOMEDCT_US|Exposure to Severe acute respiratory syndrome coronavirus|Exposure to Severe acute respiratory syndrome coronavirus
C2733460|T051|FN|444482005|SNOMEDCT_US|Exposure to severe acute respiratory syndrome coronavirus (event)|Exposure to severe acute respiratory syndrome coronavirus (event)
C2733460|T051|OF|444482005|SNOMEDCT_US|Exposure to Severe acute respiratory syndrome coronavirus (event)|Exposure to Severe acute respiratory syndrome coronavirus (event)
C2748216|T034|PT|10070255|MDR|Coronavirus test positive|Coronavirus test positive
C2748216|T034|LLT|10070255|MDR|Coronavirus test positive|Coronavirus test positive
C2748226|T034|LLT|10070268|MDR|Severe acute respiratory syndrome virus test positive|Severe acute respiratory syndrome virus test positive
C2806447|T005|PT|C119319|NCI|Alphacoronavirus|Alphacoronavirus
C2806447|T005|MH|D000073638|MSH|Alphacoronavirus|Alphacoronavirus
C2806447|T005|PT|C119319|NCI_CDISC|ALPHACORONAVIRUS|ALPHACORONAVIRUS
C2806447|T005|PM|D000073638|MSH|Alphacoronaviruses|Alphacoronaviruses
C2806447|T005|SY|C119319|NCI_CDISC|Coronavirus Group 1|Coronavirus Group 1
C2806448|T005|SY|697941000|SNOMEDCT_US|ACoV-1|ACoV-1
C2806448|T005|MH|D000073639|MSH|Alphacoronavirus 1|Alphacoronavirus 1
C2806448|T005|PT|697941000|SNOMEDCT_US|Alphacoronavirus 1|Alphacoronavirus 1
C2806448|T005|FN|697941000|SNOMEDCT_US|Alphacoronavirus 1 (organism)|Alphacoronavirus 1 (organism)
C2806449|T005|SY|709681004|SNOMEDCT_US|Coronavirus HKU2|Coronavirus HKU2
C2806449|T005|PEP|D000073638|MSH|Rhinolophus bat coronavirus HKU2|Rhinolophus bat coronavirus HKU2
C2806449|T005|PT|709681004|SNOMEDCT_US|Rhinolophus bat coronavirus HKU2|Rhinolophus bat coronavirus HKU2
C2806449|T005|FN|709681004|SNOMEDCT_US|Rhinolophus bat coronavirus HKU2 (organism)|Rhinolophus bat coronavirus HKU2 (organism)
C2806450|T005|PEP|D000073638|MSH|Scotophilus bat coronavirus 512|Scotophilus bat coronavirus 512
C2806451|T005|PEP|D000073638|MSH|Miniopterus bat coronavirus 1|Miniopterus bat coronavirus 1
C2806452|T005|PEP|D000073638|MSH|Miniopterus bat coronavirus HKU8|Miniopterus bat coronavirus HKU8
C2806453|T005|SY|C113207|NCI|Beta-CoV|Beta-CoV
C2806453|T005|PT|C113207|NCI|Betacoronavirus|Betacoronavirus
C2806453|T005|MH|D000073640|MSH|Betacoronavirus|Betacoronavirus
C2806453|T005|PT|C113207|NCI_CDISC|BETACORONAVIRUS|BETACORONAVIRUS
C2806453|T005|PM|D000073640|MSH|Betacoronaviruses|Betacoronaviruses
C2806453|T005|SY|C113207|NCI_CDISC|Coronavirus Group 2|Coronavirus Group 2
C2806454|T005|SY|697940004|SNOMEDCT_US|BCoV-1|BCoV-1
C2806454|T005|MH|D000073641|MSH|Betacoronavirus 1|Betacoronavirus 1
C2806454|T005|PT|697940004|SNOMEDCT_US|Betacoronavirus 1|Betacoronavirus 1
C2806454|T005|FN|697940004|SNOMEDCT_US|Betacoronavirus 1 (organism)|Betacoronavirus 1 (organism)
C2806456|T005|PEP|D000073640|MSH|Rousettus bat coronavirus HKU9|Rousettus bat coronavirus HKU9
C2806457|T005|PEP|D000073640|MSH|Tylonycteris bat coronavirus HKU4|Tylonycteris bat coronavirus HKU4
C2806458|T005|PEP|D000073640|MSH|Pipistrellus bat coronavirus HKU5|Pipistrellus bat coronavirus HKU5
C2806460|T005|SY|C122313|NCI_CDISC|Coronavirus group 3|Coronavirus group 3
C2806460|T005|PT|C122313|NCI|Gammacoronavirus|Gammacoronavirus
C2806460|T005|MH|D000073642|MSH|Gammacoronavirus|Gammacoronavirus
C2806460|T005|PN|NOCODE|MTH|Gammacoronavirus|Gammacoronavirus
C2806460|T005|PT|C122313|NCI_CDISC|GAMMACORONAVIRUS|GAMMACORONAVIRUS
C2806460|T005|PM|D000073642|MSH|Gammacoronaviruses|Gammacoronaviruses
C2806461|T005|PEP|D000073642|MSH|Avian coronavirus|Avian coronavirus
C2806461|T005|PT|697939001|SNOMEDCT_US|Avian coronavirus|Avian coronavirus
C2806461|T005|FN|697939001|SNOMEDCT_US|Avian coronavirus (organism)|Avian coronavirus (organism)
C2806461|T005|PM|D000073642|MSH|Avian coronaviruses|Avian coronaviruses
C2833819|T047|SY|330009|MEDCIN|coronavirus sars-associated as cause of disease classified elsewhere|coronavirus sars-associated as cause of disease classified elsewhere
C2833819|T047|PT|330009|MEDCIN|SARS-associated coronavirus as cause of disease classified elsewhere|SARS-associated coronavirus as cause of disease classified elsewhere
C2833819|T047|FN|330009|MEDCIN|SARS-associated coronavirus as cause of disease classified elsewhere (diagnosis)|SARS-associated coronavirus as cause of disease classified elsewhere (diagnosis)
C2833819|T047|PT|B97.21|ICD10CM|SARS-associated coronavirus as the cause of diseases classified elsewhere|SARS-associated coronavirus as the cause of diseases classified elsewhere
C2833819|T047|AB|B97.21|ICD10CM|SARS-associated coronavirus causing diseases classd elswhr|SARS-associated coronavirus causing diseases classd elswhr
C2833820|T047|AB|B97.29|ICD10CM|Oth coronavirus as the cause of diseases classd elswhr|Oth coronavirus as the cause of diseases classd elswhr
C2833820|T047|PT|B97.29|ICD10CM|Other coronavirus as the cause of diseases classified elsewhere|Other coronavirus as the cause of diseases classified elsewhere
C2939460|T005|PT|415462005|SNOMEDCT_US|SARS coronavirus TW|SARS coronavirus TW
C2939460|T005|OF|415462005|SNOMEDCT_US|SARS coronavirus TW (organism)|SARS coronavirus TW (organism)
C2939460|T005|SY|415462005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW|Severe acute respiratory syndrome (SARS) coronavirus TW
C2939460|T005|OF|415462005|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus TW (organism)|Severe acute respiratory syndrome (SARS) coronavirus TW (organism)
C2939460|T005|SY|415462005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW|Severe acute respiratory syndrome coronavirus TW
C2939460|T005|FN|415462005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus TW (organism)|Severe acute respiratory syndrome coronavirus TW (organism)
C2970108|T201|DN|60265-6|LNC|HCoV RNA NAA+probe Ql|HCoV RNA NAA+probe Ql
C2970108|T201|OSN|60265-6|LNC|HCoV RNA SerPl Ql NAA+probe|HCoV RNA SerPl Ql NAA+probe
C2970108|T201|MTH_LN|60265-6|LNC|Human coronavirus ribonucleic acid:Presence or Threshold:Point in time:Serum/Plasma:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus ribonucleic acid:Presence or Threshold:Point in time:Serum/Plasma:Ordinal:DNA Nucleic Acid Probe.amp.tar
C2970108|T201|LC|60265-6|LNC|Human coronavirus RNA [Presence] in Serum or Plasma by NAA with probe detection|Human coronavirus RNA [Presence] in Serum or Plasma by NAA with probe detection
C2970108|T201|LN|60265-6|LNC|Human coronavirus RNA:PrThr:Pt:Ser/Plas:Ord:Probe.amp.tar|Human coronavirus RNA:PrThr:Pt:Ser/Plas:Ord:Probe.amp.tar
C2970118|T201|MTH_LN|60275-5|LNC|SARS coronavirus ribonucleic acid:Presence or Threshold:Point in time:Isolate:Ordinal:DNA Nucleic Acid Probe.amp.tar|SARS coronavirus ribonucleic acid:Presence or Threshold:Point in time:Isolate:Ordinal:DNA Nucleic Acid Probe.amp.tar
C2970118|T201|LC|60275-5|LNC|SARS coronavirus RNA [Presence] in Isolate by NAA with probe detection|SARS coronavirus RNA [Presence] in Isolate by NAA with probe detection
C2970118|T201|DN|60275-5|LNC|SARS coronavirus RNA NAA+probe Ql (Isol)|SARS coronavirus RNA NAA+probe Ql (Isol)
C2970118|T201|LN|60275-5|LNC|SARS coronavirus RNA:PrThr:Pt:Isolate:Ord:Probe.amp.tar|SARS coronavirus RNA:PrThr:Pt:Isolate:Ord:Probe.amp.tar
C2970118|T201|OSN|60275-5|LNC|SARS-CoV RNA Islt Ql NAA+probe|SARS-CoV RNA Islt Ql NAA+probe
C2970236|T201|DN|60426-4|LNC|SARS coronavirus Ab (S) [Titer]|SARS coronavirus Ab (S) [Titer]
C2970236|T201|LC|60426-4|LNC|SARS coronavirus Ab [Titer] in Serum|SARS coronavirus Ab [Titer] in Serum
C2970236|T201|LN|60426-4|LNC|SARS coronavirus Ab:Titr:Pt:Ser:Qn|SARS coronavirus Ab:Titr:Pt:Ser:Qn
C2970236|T201|MTH_LN|60426-4|LNC|SARS coronavirus Antibody:Dilution Factor (Titer):Point in time:Serum:Quantitative|SARS coronavirus Antibody:Dilution Factor (Titer):Point in time:Serum:Quantitative
C2970236|T201|OSN|60426-4|LNC|SARS-CoV Ab Titr Ser|SARS-CoV Ab Titr Ser
C2970316|T201|MTH_LN|60534-5|LNC|SARS coronavirus ribonucleic acid:Presence or Threshold:Point in time:Serum/Plasma:Ordinal:DNA Nucleic Acid Probe.amp.tar|SARS coronavirus ribonucleic acid:Presence or Threshold:Point in time:Serum/Plasma:Ordinal:DNA Nucleic Acid Probe.amp.tar
C2970316|T201|LC|60534-5|LNC|SARS coronavirus RNA [Presence] in Serum or Plasma by NAA with probe detection|SARS coronavirus RNA [Presence] in Serum or Plasma by NAA with probe detection
C2970316|T201|DN|60534-5|LNC|SARS coronavirus RNA NAA+probe Ql|SARS coronavirus RNA NAA+probe Ql
C2970316|T201|LN|60534-5|LNC|SARS coronavirus RNA:PrThr:Pt:Ser/Plas:Ord:Probe.amp.tar|SARS coronavirus RNA:PrThr:Pt:Ser/Plas:Ord:Probe.amp.tar
C2970316|T201|OSN|60534-5|LNC|SARS-CoV RNA SerPl Ql NAA+probe|SARS-CoV RNA SerPl Ql NAA+probe
C3169505|T201|DN|62423-9|LNC|HCoV HKU1 RNA NAA+probe Ql (Unsp spec)|HCoV HKU1 RNA NAA+probe Ql (Unsp spec)
C3169505|T201|OSN|62423-9|LNC|HCoV HKU1 RNA XXX Ql NAA+probe|HCoV HKU1 RNA XXX Ql NAA+probe
C3169505|T201|MTH_LN|62423-9|LNC|Human coronavirus HKU1 ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus HKU1 ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar
C3169505|T201|LC|62423-9|LNC|Human coronavirus HKU1 RNA [Presence] in Unspecified specimen by NAA with probe detection|Human coronavirus HKU1 RNA [Presence] in Unspecified specimen by NAA with probe detection
C3169505|T201|LN|62423-9|LNC|Human coronavirus HKU1 RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar|Human coronavirus HKU1 RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar
C3169506|T114|MTH_CN|MTHU037034|LNC|Human coronavirus HKU1 ribonucleic acid|Human coronavirus HKU1 ribonucleic acid
C3169506|T114|LPN|LP111517-1|LNC|Human coronavirus HKU1 RNA|Human coronavirus HKU1 RNA
C3169506|T114|CN|MTHU037034|LNC|Human coronavirus HKU1 RNA|Human coronavirus HKU1 RNA
C3169506|T114|PT|707893001|SNOMEDCT_US|Human coronavirus HKU1 RNA|Human coronavirus HKU1 RNA
C3169506|T114|SY|707893001|SNOMEDCT_US|Ribonucleic acid of Human coronavirus HKU1|Ribonucleic acid of Human coronavirus HKU1
C3169506|T114|FN|707893001|SNOMEDCT_US|Ribonucleic acid of Human coronavirus HKU1 (substance)|Ribonucleic acid of Human coronavirus HKU1 (substance)
C3172513|T201|OSN|63430-3|LNC|HCoV pnl XXX NAA+probe|HCoV pnl XXX NAA+probe
C3172513|T201|DN|63430-3|LNC|HCoV RNA panel NAA+probe (Unsp spec)|HCoV RNA panel NAA+probe (Unsp spec)
C3172513|T201|MTH_LN|63430-3|LNC|Human coronavirus ribonucleic acid panel:-:Point in time:To be specified in another part of the message:-:DNA Nucleic Acid Probe.amp.tar|Human coronavirus ribonucleic acid panel:-:Point in time:To be specified in another part of the message:-:DNA Nucleic Acid Probe.amp.tar
C3172513|T201|LC|63430-3|LNC|Human coronavirus RNA panel - Unspecified specimen by NAA with probe detection|Human coronavirus RNA panel - Unspecified specimen by NAA with probe detection
C3172513|T201|LN|63430-3|LNC|Human coronavirus RNA panel:-:Pt:XXX:-:Probe.amp.tar|Human coronavirus RNA panel:-:Pt:XXX:-:Probe.amp.tar
C3172514|T059|MTH_CN|MTHU037695|LNC|Human coronavirus ribonucleic acid panel|Human coronavirus ribonucleic acid panel
C3172514|T059|LPN|LP113746-4|LNC|Human coronavirus RNA panel|Human coronavirus RNA panel
C3172514|T059|CN|MTHU037695|LNC|Human coronavirus RNA panel|Human coronavirus RNA panel
C3441987|T005|SY|C122279|NCI_CDISC|Coronavirus Group 3|Coronavirus Group 3
C3441987|T005|PT|C122279|NCI|Deltacoronavirus|Deltacoronavirus
C3441987|T005|PEP|D017934|MSH|Deltacoronavirus|Deltacoronavirus
C3441987|T005|PN|NOCODE|MTH|Deltacoronavirus|Deltacoronavirus
C3441987|T005|PT|C122279|NCI_CDISC|DELTACORONAVIRUS|DELTACORONAVIRUS
C3441987|T005|PM|D017934|MSH|Deltacoronaviruses|Deltacoronaviruses
C3463158|T005|PEP|D017934|MSH|Bulbul coronavirus HKU11|Bulbul coronavirus HKU11
C3598902|T005|PEP|D000073638|MSH|Bat coronavirus HKU10|Bat coronavirus HKU10
C3598902|T005|PM|D000073638|MSH|HKU10, Bat coronavirus|HKU10, Bat coronavirus
C3627024|T005|PEP|D017934|MSH|Munia coronavirus HKU13|Munia coronavirus HKU13
C3627025|T005|PEP|D017934|MSH|Thrush coronavirus HKU12|Thrush coronavirus HKU12
C3658241|T116|ET|D064370|MSH|E2 Spike Glycoprotein, Coronavirus|E2 Spike Glycoprotein, Coronavirus
C3658241|T123|ET|D064370|MSH|E2 Spike Glycoprotein, Coronavirus|E2 Spike Glycoprotein, Coronavirus
C3658241|T116|PEP|D064370|MSH|Spike Protein S2, Coronavirus|Spike Protein S2, Coronavirus
C3658241|T123|PEP|D064370|MSH|Spike Protein S2, Coronavirus|Spike Protein S2, Coronavirus
C3658242|T116|PEP|D064370|MSH|Spike Glycoprotein S1, Coronavirus|Spike Glycoprotein S1, Coronavirus
C3658242|T123|PEP|D064370|MSH|Spike Glycoprotein S1, Coronavirus|Spike Glycoprotein S1, Coronavirus
C3658242|T116|ET|D064370|MSH|Spike Gp S1, Cor|Spike Gp S1, Cor
C3658242|T123|ET|D064370|MSH|Spike Gp S1, Cor|Spike Gp S1, Cor
C3658243|T116|PM|D064370|MSH|Coronavirus Spike Glycoprotein|Coronavirus Spike Glycoprotein
C3658243|T123|PM|D064370|MSH|Coronavirus Spike Glycoprotein|Coronavirus Spike Glycoprotein
C3658243|T116|PM|D064370|MSH|Coronavirus Spike Protein|Coronavirus Spike Protein
C3658243|T123|PM|D064370|MSH|Coronavirus Spike Protein|Coronavirus Spike Protein
C3658243|T116|ET|D064370|MSH|Glycoprotein S, Coronavirus|Glycoprotein S, Coronavirus
C3658243|T123|ET|D064370|MSH|Glycoprotein S, Coronavirus|Glycoprotein S, Coronavirus
C3658243|T116|MH|D064370|MSH|Spike Glycoprotein, Coronavirus|Spike Glycoprotein, Coronavirus
C3658243|T123|MH|D064370|MSH|Spike Glycoprotein, Coronavirus|Spike Glycoprotein, Coronavirus
C3658243|T116|ET|D064370|MSH|Spike Glycoproteins, Coronavirus|Spike Glycoproteins, Coronavirus
C3658243|T123|ET|D064370|MSH|Spike Glycoproteins, Coronavirus|Spike Glycoproteins, Coronavirus
C3658243|T116|ET|D064370|MSH|Spike Protein, Coronavirus|Spike Protein, Coronavirus
C3658243|T123|ET|D064370|MSH|Spike Protein, Coronavirus|Spike Protein, Coronavirus
C3686947|T005|PEP|D000073641|MSH|Equine coronavirus|Equine coronavirus
C3686947|T005|PM|D000073641|MSH|Equine coronaviruses|Equine coronaviruses
C3690073|T074|PT|22-441|UMD|IVD Test Reagent/Kits, Serology, Virus, Severe Acute Respiratory Syndrome Coronavirus, IgG Antibody|IVD Test Reagent/Kits, Serology, Virus, Severe Acute Respiratory Syndrome Coronavirus, IgG Antibody
C3690175|T074|PT|22-339|UMD|IVD Test Reagent/Kits, Molecular Assay, Infection, Virus, Severe Acute Respiratory Syndrome Coronavirus, RNA|IVD Test Reagent/Kits, Molecular Assay, Infection, Virus, Severe Acute Respiratory Syndrome Coronavirus, RNA
C3697412|T005|PT|697938009|SNOMEDCT_US|Genus Gammacoronavirus|Genus Gammacoronavirus
C3697412|T005|FN|697938009|SNOMEDCT_US|Genus Gammacoronavirus (organism)|Genus Gammacoronavirus (organism)
C3697502|T005|PT|697937004|SNOMEDCT_US|Genus Deltacoronavirus|Genus Deltacoronavirus
C3697502|T005|FN|697937004|SNOMEDCT_US|Genus Deltacoronavirus (organism)|Genus Deltacoronavirus (organism)
C3697872|T005|PT|697936008|SNOMEDCT_US|Genus Betacoronavirus|Genus Betacoronavirus
C3697872|T005|FN|697936008|SNOMEDCT_US|Genus Betacoronavirus (organism)|Genus Betacoronavirus (organism)
C3698297|T005|PT|697935007|SNOMEDCT_US|Genus Alphacoronavirus|Genus Alphacoronavirus
C3698297|T005|FN|697935007|SNOMEDCT_US|Genus Alphacoronavirus (organism)|Genus Alphacoronavirus (organism)
C3698360|T005|SY|697932005|SNOMEDCT_US|MERS coronavirus|MERS coronavirus
C3698360|T005|ET|D065207|MSH|MERS Virus|MERS Virus
C3698360|T005|PM|D065207|MSH|MERS Viruses|MERS Viruses
C3698360|T005|LA|LA26151-3|LNC|MERS- CoV|MERS- CoV
C3698360|T005|ET|D065207|MSH|MERS-CoV|MERS-CoV
C3698360|T005|PT|697932005|SNOMEDCT_US|MERS-CoV|MERS-CoV
C3698360|T005|MH|D065207|MSH|Middle East Respiratory Syndrome Coronavirus|Middle East Respiratory Syndrome Coronavirus
C3698360|T005|SY|697932005|SNOMEDCT_US|Middle East Respiratory Syndrome Coronavirus|Middle East Respiratory Syndrome Coronavirus
C3698360|T005|LPN|LP173753-7|LNC|Middle East respiratory syndrome coronavirus|Middle East respiratory syndrome coronavirus
C3698360|T005|SY|697932005|SNOMEDCT_US|Middle East respiratory syndrome coronavirus|Middle East respiratory syndrome coronavirus
C3698360|T005|FN|697932005|SNOMEDCT_US|Middle East respiratory syndrome coronavirus (organism)|Middle East respiratory syndrome coronavirus (organism)
C3698360|T005|PM|D065207|MSH|Middle East respiratory syndrome related coronavirus|Middle East respiratory syndrome related coronavirus
C3698360|T005|ET|D065207|MSH|Middle East respiratory syndrome-related coronavirus|Middle East respiratory syndrome-related coronavirus
C3698360|T005|PM|D065207|MSH|Virus, MERS|Virus, MERS
C3698360|T005|PM|D065207|MSH|Viruses, MERS|Viruses, MERS
C3699854|T201|DN|74408-6|LNC|MERS-CoV RNA panel (Unsp spec)|MERS-CoV RNA panel (Unsp spec)
C3699854|T201|OSN|74408-6|LNC|MERS-CoV RNA Pnl XXX|MERS-CoV RNA Pnl XXX
C3699854|T201|LC|74408-6|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA panel - Unspecified specimen|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA panel - Unspecified specimen
C3699854|T201|MTH_LN|74408-6|LNC|Middle east respiratory syndrome coronavirus ribonucleic acid panel:-:Point in time:To be specified in another part of the message:-|Middle east respiratory syndrome coronavirus ribonucleic acid panel:-:Point in time:To be specified in another part of the message:-
C3699854|T201|LN|74408-6|LNC|Middle east respiratory syndrome coronavirus RNA panel:-:Pt:XXX:-|Middle east respiratory syndrome coronavirus RNA panel:-:Pt:XXX:-
C3699855|T059|MTH_CN|MTHU047597|LNC|Middle east respiratory syndrome coronavirus ribonucleic acid panel|Middle east respiratory syndrome coronavirus ribonucleic acid panel
C3699855|T059|CN|MTHU047597|LNC|Middle east respiratory syndrome coronavirus RNA panel|Middle east respiratory syndrome coronavirus RNA panel
C3699855|T059|LPN|LP175722-0|LNC|Middle East respiratory syndrome coronavirus RNA panel|Middle East respiratory syndrome coronavirus RNA panel
C3699926|T201|DN|74472-2|LNC|MERS-CoV N3 gene RNA NAA+probe Ql (Unsp spec)|MERS-CoV N3 gene RNA NAA+probe Ql (Unsp spec)
C3699926|T201|OSN|74472-2|LNC|MERS-CoV N3 RNA XXX Ql NAA+probe|MERS-CoV N3 RNA XXX Ql NAA+probe
C3699926|T201|LC|74472-2|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) N3 gene RNA [Presence] in Unspecified specimen by NAA with probe detection|Middle East respiratory syndrome coronavirus (MERS-CoV) N3 gene RNA [Presence] in Unspecified specimen by NAA with probe detection
C3699926|T201|MTH_LN|74472-2|LNC|Middle east respiratory syndrome coronavirus N3 gene ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar|Middle east respiratory syndrome coronavirus N3 gene ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar
C3699926|T201|LN|74472-2|LNC|Middle east respiratory syndrome coronavirus N3 gene RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar|Middle east respiratory syndrome coronavirus N3 gene RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar
C3699927|T114|MTH_CN|MTHU047620|LNC|Middle east respiratory syndrome coronavirus N3 gene ribonucleic acid|Middle east respiratory syndrome coronavirus N3 gene ribonucleic acid
C3699927|T123|MTH_CN|MTHU047620|LNC|Middle east respiratory syndrome coronavirus N3 gene ribonucleic acid|Middle east respiratory syndrome coronavirus N3 gene ribonucleic acid
C3699927|T114|CN|MTHU047620|LNC|Middle east respiratory syndrome coronavirus N3 gene RNA|Middle east respiratory syndrome coronavirus N3 gene RNA
C3699927|T123|CN|MTHU047620|LNC|Middle east respiratory syndrome coronavirus N3 gene RNA|Middle east respiratory syndrome coronavirus N3 gene RNA
C3699927|T114|LPN|LP175710-5|LNC|Middle East respiratory syndrome coronavirus N3 gene RNA|Middle East respiratory syndrome coronavirus N3 gene RNA
C3699927|T123|LPN|LP175710-5|LNC|Middle East respiratory syndrome coronavirus N3 gene RNA|Middle East respiratory syndrome coronavirus N3 gene RNA
C3699928|T201|DN|74473-0|LNC|MERS-CoV N2 gene RNA NAA+probe Ql (Unsp spec)|MERS-CoV N2 gene RNA NAA+probe Ql (Unsp spec)
C3699928|T201|OSN|74473-0|LNC|MERS-CoV N2 RNA XXX Ql NAA+probe|MERS-CoV N2 RNA XXX Ql NAA+probe
C3699928|T201|LC|74473-0|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) N2 gene RNA [Presence] in Unspecified specimen by NAA with probe detection|Middle East respiratory syndrome coronavirus (MERS-CoV) N2 gene RNA [Presence] in Unspecified specimen by NAA with probe detection
C3699928|T201|MTH_LN|74473-0|LNC|Middle east respiratory syndrome coronavirus N2 gene ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar|Middle east respiratory syndrome coronavirus N2 gene ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar
C3699928|T201|LN|74473-0|LNC|Middle east respiratory syndrome coronavirus N2 gene RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar|Middle east respiratory syndrome coronavirus N2 gene RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar
C3699929|T114|MTH_CN|MTHU047621|LNC|Middle east respiratory syndrome coronavirus N2 gene ribonucleic acid|Middle east respiratory syndrome coronavirus N2 gene ribonucleic acid
C3699929|T123|MTH_CN|MTHU047621|LNC|Middle east respiratory syndrome coronavirus N2 gene ribonucleic acid|Middle east respiratory syndrome coronavirus N2 gene ribonucleic acid
C3699929|T114|CN|MTHU047621|LNC|Middle east respiratory syndrome coronavirus N2 gene RNA|Middle east respiratory syndrome coronavirus N2 gene RNA
C3699929|T123|CN|MTHU047621|LNC|Middle east respiratory syndrome coronavirus N2 gene RNA|Middle east respiratory syndrome coronavirus N2 gene RNA
C3699929|T114|LPN|LP175711-3|LNC|Middle East respiratory syndrome coronavirus N2 gene RNA|Middle East respiratory syndrome coronavirus N2 gene RNA
C3699929|T123|LPN|LP175711-3|LNC|Middle East respiratory syndrome coronavirus N2 gene RNA|Middle East respiratory syndrome coronavirus N2 gene RNA
C3699930|T201|DN|74474-8|LNC|MERS-CoV upE gene RNA NAA+probe Ql (Unsp spec)|MERS-CoV upE gene RNA NAA+probe Ql (Unsp spec)
C3699930|T201|OSN|74474-8|LNC|MERS-CoV upE RNA XXX Ql NAA+probe|MERS-CoV upE RNA XXX Ql NAA+probe
C3699930|T201|LC|74474-8|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) upE gene RNA [Presence] in Unspecified specimen by NAA with probe detection|Middle East respiratory syndrome coronavirus (MERS-CoV) upE gene RNA [Presence] in Unspecified specimen by NAA with probe detection
C3699930|T201|MTH_LN|74474-8|LNC|Middle east respiratory syndrome coronavirus upE gene ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar|Middle east respiratory syndrome coronavirus upE gene ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar
C3699930|T201|LN|74474-8|LNC|Middle east respiratory syndrome coronavirus upE gene RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar|Middle east respiratory syndrome coronavirus upE gene RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar
C3699931|T114|MTH_CN|MTHU047622|LNC|Middle east respiratory syndrome coronavirus upE gene ribonucleic acid|Middle east respiratory syndrome coronavirus upE gene ribonucleic acid
C3699931|T123|MTH_CN|MTHU047622|LNC|Middle east respiratory syndrome coronavirus upE gene ribonucleic acid|Middle east respiratory syndrome coronavirus upE gene ribonucleic acid
C3699931|T114|CN|MTHU047622|LNC|Middle east respiratory syndrome coronavirus upE gene RNA|Middle east respiratory syndrome coronavirus upE gene RNA
C3699931|T123|CN|MTHU047622|LNC|Middle east respiratory syndrome coronavirus upE gene RNA|Middle east respiratory syndrome coronavirus upE gene RNA
C3699931|T114|LPN|LP175712-1|LNC|Middle East respiratory syndrome coronavirus upE gene RNA|Middle East respiratory syndrome coronavirus upE gene RNA
C3699931|T123|LPN|LP175712-1|LNC|Middle East respiratory syndrome coronavirus upE gene RNA|Middle East respiratory syndrome coronavirus upE gene RNA
C3699932|T201|DN|74475-5|LNC|MERS-CoV RNA NAA+probe Ql (Unsp spec) [Interp]|MERS-CoV RNA NAA+probe Ql (Unsp spec) [Interp]
C3699932|T201|OSN|74475-5|LNC|MERS-CoV RNA XXX NAA+probe-Imp|MERS-CoV RNA XXX NAA+probe-Imp
C3699932|T201|LC|74475-5|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Interpretation] in Unspecified specimen Qualitative by NAA with probe detection|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Interpretation] in Unspecified specimen Qualitative by NAA with probe detection
C3699932|T201|MTH_LN|74475-5|LNC|Middle east respiratory syndrome coronavirus ribonucleic acid:Impression/interpretation of study:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar|Middle east respiratory syndrome coronavirus ribonucleic acid:Impression/interpretation of study:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar
C3699932|T201|LN|74475-5|LNC|Middle east respiratory syndrome coronavirus RNA:Imp:Pt:XXX:Ord:Probe.amp.tar|Middle east respiratory syndrome coronavirus RNA:Imp:Pt:XXX:Ord:Probe.amp.tar
C3699933|T114|MTH_CN|MTHU047623|LNC|Middle east respiratory syndrome coronavirus ribonucleic acid|Middle east respiratory syndrome coronavirus ribonucleic acid
C3699933|T123|MTH_CN|MTHU047623|LNC|Middle east respiratory syndrome coronavirus ribonucleic acid|Middle east respiratory syndrome coronavirus ribonucleic acid
C3699933|T114|MTH_CN|MTHU056753|LNC|Middle East respiratory syndrome coronavirus ribonucleic acid|Middle East respiratory syndrome coronavirus ribonucleic acid
C3699933|T123|MTH_CN|MTHU056753|LNC|Middle East respiratory syndrome coronavirus ribonucleic acid|Middle East respiratory syndrome coronavirus ribonucleic acid
C3699933|T114|CN|MTHU047623|LNC|Middle east respiratory syndrome coronavirus RNA|Middle east respiratory syndrome coronavirus RNA
C3699933|T123|CN|MTHU047623|LNC|Middle east respiratory syndrome coronavirus RNA|Middle east respiratory syndrome coronavirus RNA
C3699933|T114|LPN|LP173752-9|LNC|Middle East respiratory syndrome coronavirus RNA|Middle East respiratory syndrome coronavirus RNA
C3699933|T123|LPN|LP173752-9|LNC|Middle East respiratory syndrome coronavirus RNA|Middle East respiratory syndrome coronavirus RNA
C3699933|T114|CN|MTHU056753|LNC|Middle East respiratory syndrome coronavirus RNA|Middle East respiratory syndrome coronavirus RNA
C3699933|T123|CN|MTHU056753|LNC|Middle East respiratory syndrome coronavirus RNA|Middle East respiratory syndrome coronavirus RNA
C3700012|T028|LPN|LP175714-7|LNC|Middle East respiratory syndrome coronavirus N2 gene|Middle East respiratory syndrome coronavirus N2 gene
C3700013|T028|LPN|LP175715-4|LNC|Middle East respiratory syndrome coronavirus N3 gene|Middle East respiratory syndrome coronavirus N3 gene
C3700014|T028|LPN|LP175713-9|LNC|Middle East respiratory syndrome coronavirus upE gene|Middle East respiratory syndrome coronavirus upE gene
C3711684|T116|CE|C578557|MSH|S protein, SARS-CoV|S protein, SARS-CoV
C3711684|T123|CE|C578557|MSH|S protein, SARS-CoV|S protein, SARS-CoV
C3711684|T116|NM|C578557|MSH|S protein, severe acute respiratory syndrome coronavirus|S protein, severe acute respiratory syndrome coronavirus
C3711684|T123|NM|C578557|MSH|S protein, severe acute respiratory syndrome coronavirus|S protein, severe acute respiratory syndrome coronavirus
C3711684|T116|CE|C578557|MSH|SARS S protein, SARS-CoV|SARS S protein, SARS-CoV
C3711684|T123|CE|C578557|MSH|SARS S protein, SARS-CoV|SARS S protein, SARS-CoV
C3713754|T116|NM|C578555|MSH|S protein, canine coronavirus (CCV)|S protein, canine coronavirus (CCV)
C3713754|T123|NM|C578555|MSH|S protein, canine coronavirus (CCV)|S protein, canine coronavirus (CCV)
C3713755|T116|NM|C578559|MSH|spike glycoprotein, human coronavirus (HCV)|spike glycoprotein, human coronavirus (HCV)
C3713755|T123|NM|C578559|MSH|spike glycoprotein, human coronavirus (HCV)|spike glycoprotein, human coronavirus (HCV)
C3713756|T116|NM|C578558|MSH|spike glycoprotein, bovine coronavirus (BCV)|spike glycoprotein, bovine coronavirus (BCV)
C3713756|T123|NM|C578558|MSH|spike glycoprotein, bovine coronavirus (BCV)|spike glycoprotein, bovine coronavirus (BCV)
C3838696|T033|PT|700217006|SNOMEDCT_US|Suspected coronavirus infection|Suspected coronavirus infection
C3838696|T033|FN|700217006|SNOMEDCT_US|Suspected coronavirus infection (situation)|Suspected coronavirus infection (situation)
C3839253|T033|PT|702547000|SNOMEDCT_US|Exposure to coronavirus infection|Exposure to coronavirus infection
C3839253|T033|FN|702547000|SNOMEDCT_US|Exposure to coronavirus infection (event)|Exposure to coronavirus infection (event)
C3872915|T114|SY|707785005|SNOMEDCT_US|Ribonucleic acid of Severe acute respiratory syndrome coronavirus Urbani|Ribonucleic acid of Severe acute respiratory syndrome coronavirus Urbani
C3872915|T114|FN|707785005|SNOMEDCT_US|Ribonucleic acid of Severe acute respiratory syndrome coronavirus Urbani (substance)|Ribonucleic acid of Severe acute respiratory syndrome coronavirus Urbani (substance)
C3872915|T114|SY|707785005|SNOMEDCT_US|SARS (severe acute respiratory syndrome) coronavirus Urbani RNA|SARS (severe acute respiratory syndrome) coronavirus Urbani RNA
C3872915|T114|OP|707785005|SNOMEDCT_US|SARS Urbani RNA|SARS Urbani RNA
C3872915|T114|PT|707785005|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus Urbani RNA|Severe acute respiratory syndrome coronavirus Urbani RNA
C3873497|T047|PT|707224005|SNOMEDCT_US|Severe acute respiratory infection|Severe acute respiratory infection
C3873497|T047|FN|707224005|SNOMEDCT_US|Severe acute respiratory infection (disorder)|Severe acute respiratory infection (disorder)
C3873497|T047|SY|707224005|SNOMEDCT_US|Severe acute respiratory infection (SARI)|Severe acute respiratory infection (SARI)
C3884565|T116|CE|C000593134|MSH|open reading frame-9b, SARS coronavirus|open reading frame-9b, SARS coronavirus
C3884565|T123|CE|C000593134|MSH|open reading frame-9b, SARS coronavirus|open reading frame-9b, SARS coronavirus
C3884565|T116|NM|C000593134|MSH|ORF-9b protein, SARS coronavirus|ORF-9b protein, SARS coronavirus
C3884565|T123|NM|C000593134|MSH|ORF-9b protein, SARS coronavirus|ORF-9b protein, SARS coronavirus
C4034672|T116|LPN|LP189868-5|LNC|Human coronavirus 229E+OC43|Human coronavirus 229E+OC43
C4034672|T129|LPN|LP189868-5|LNC|Human coronavirus 229E+OC43|Human coronavirus 229E+OC43
C4035026|T114|MTH_CN|MTHU055965|LNC|Porcine deltacoronavirus ribonucleic acid|Porcine deltacoronavirus ribonucleic acid
C4035026|T123|MTH_CN|MTHU055965|LNC|Porcine deltacoronavirus ribonucleic acid|Porcine deltacoronavirus ribonucleic acid
C4035026|T114|LPN|LP188527-8|LNC|Porcine deltacoronavirus RNA|Porcine deltacoronavirus RNA
C4035026|T123|LPN|LP188527-8|LNC|Porcine deltacoronavirus RNA|Porcine deltacoronavirus RNA
C4035026|T114|CN|MTHU055965|LNC|Porcine deltacoronavirus RNA|Porcine deltacoronavirus RNA
C4035026|T123|CN|MTHU055965|LNC|Porcine deltacoronavirus RNA|Porcine deltacoronavirus RNA
C4037273|T201|DN|77008-1|LNC|HCoV 229E+OC43 RNA NAA+probe Ql (Nph)|HCoV 229E+OC43 RNA NAA+probe Ql (Nph)
C4037273|T201|OSN|77008-1|LNC|HCoV 229E+OC43 RNA Nph Ql NAA+probe|HCoV 229E+OC43 RNA Nph Ql NAA+probe
C4037273|T201|MTH_LN|77008-1|LNC|Human coronavirus 229E+OC43 ribonucleic acid:Presence or Threshold:Point in time:Naspopharynx:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus 229E+OC43 ribonucleic acid:Presence or Threshold:Point in time:Naspopharynx:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4037273|T201|LC|77008-1|LNC|Human coronavirus 229E+OC43 RNA [Presence] in Nasopharynx by NAA with probe detection|Human coronavirus 229E+OC43 RNA [Presence] in Nasopharynx by NAA with probe detection
C4037273|T201|LN|77008-1|LNC|Human coronavirus 229E+OC43 RNA:PrThr:Pt:Nph:Ord:Probe.amp.tar|Human coronavirus 229E+OC43 RNA:PrThr:Pt:Nph:Ord:Probe.amp.tar
C4037838|T201|OSN|76340-9|LNC|PDCoV RNA Ct XXX Qn NAA+probe|PDCoV RNA Ct XXX Qn NAA+probe
C4037838|T201|MTH_LN|76340-9|LNC|Porcine deltacoronavirus ribonucleic acid:Threshold Number:Point in time:To be specified in another part of the message:Quantitative:DNA Nucleic Acid Probe.amp.tar|Porcine deltacoronavirus ribonucleic acid:Threshold Number:Point in time:To be specified in another part of the message:Quantitative:DNA Nucleic Acid Probe.amp.tar
C4037838|T201|LC|76340-9|LNC|Porcine deltacoronavirus RNA [Cycle Threshold #] in Unspecified specimen by NAA with probe detection|Porcine deltacoronavirus RNA [Cycle Threshold #] in Unspecified specimen by NAA with probe detection
C4037838|T201|DN|76340-9|LNC|Porcine deltacoronavirus RNA NAA+probe (Unsp spec) [ThreshNum]|Porcine deltacoronavirus RNA NAA+probe (Unsp spec) [ThreshNum]
C4037838|T201|LN|76340-9|LNC|Porcine deltacoronavirus RNA:ThreshNum:Pt:XXX:Qn:Probe.amp.tar|Porcine deltacoronavirus RNA:ThreshNum:Pt:XXX:Qn:Probe.amp.tar
C4037839|T201|OSN|76339-1|LNC|PDCoV RNA XXX Ql NAA+probe|PDCoV RNA XXX Ql NAA+probe
C4037839|T201|MTH_LN|76339-1|LNC|Porcine deltacoronavirus ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar|Porcine deltacoronavirus ribonucleic acid:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4037839|T201|LC|76339-1|LNC|Porcine deltacoronavirus RNA [Presence] in Unspecified specimen by NAA with probe detection|Porcine deltacoronavirus RNA [Presence] in Unspecified specimen by NAA with probe detection
C4037839|T201|DN|76339-1|LNC|Porcine deltacoronavirus RNA NAA+probe Ql (Unsp spec)|Porcine deltacoronavirus RNA NAA+probe Ql (Unsp spec)
C4037839|T201|LN|76339-1|LNC|Porcine deltacoronavirus RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar|Porcine deltacoronavirus RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar
C4038448|T005|LPN|LP188420-6|LNC|Porcine deltacoronavirus|Porcine deltacoronavirus
C4038448|T005|CN|MTHU056613|LNC|Porcine deltacoronavirus|Porcine deltacoronavirus
C4042621|T116|CE|C000595202|MSH|Nsp3 protein, MERS-CoV|Nsp3 protein, MERS-CoV
C4042621|T116|NM|C000595202|MSH|Nsp3 protein, Middle East respiratory syndrome coronavirus|Nsp3 protein, Middle East respiratory syndrome coronavirus
C4075701|T047|PT|713084008|SNOMEDCT_US|Pneumonia caused by Human coronavirus|Pneumonia caused by Human coronavirus
C4075701|T047|FN|713084008|SNOMEDCT_US|Pneumonia caused by Human coronavirus (disorder)|Pneumonia caused by Human coronavirus (disorder)
C4263799|T114|MTH_CN|MTHU052570|LNC|Human coronavirus 229E+OC43 ribonucleic acid|Human coronavirus 229E+OC43 ribonucleic acid
C4263799|T123|MTH_CN|MTHU052570|LNC|Human coronavirus 229E+OC43 ribonucleic acid|Human coronavirus 229E+OC43 ribonucleic acid
C4263799|T114|LPN|LP189803-2|LNC|Human coronavirus 229E+OC43 RNA|Human coronavirus 229E+OC43 RNA
C4263799|T123|LPN|LP189803-2|LNC|Human coronavirus 229E+OC43 RNA|Human coronavirus 229E+OC43 RNA
C4263799|T114|CN|MTHU052570|LNC|Human coronavirus 229E+OC43 RNA|Human coronavirus 229E+OC43 RNA
C4263799|T123|CN|MTHU052570|LNC|Human coronavirus 229E+OC43 RNA|Human coronavirus 229E+OC43 RNA
C4264757|T201|DN|82162-9|LNC|HCoV NL63 RNA NAA+non-probe Ql (Nph)|HCoV NL63 RNA NAA+non-probe Ql (Nph)
C4264757|T201|OSN|82162-9|LNC|HCoV NL63 RNA Nph Ql NAA+non-probe|HCoV NL63 RNA Nph Ql NAA+non-probe
C4264757|T201|MTH_LN|82162-9|LNC|Human coronavirus NL63 ribonucleic acid:Presence or Threshold:Point in time:Naspopharynx:Ordinal:Non-probe.amp.tar|Human coronavirus NL63 ribonucleic acid:Presence or Threshold:Point in time:Naspopharynx:Ordinal:Non-probe.amp.tar
C4264757|T201|LC|82162-9|LNC|Human coronavirus NL63 RNA [Presence] in Nasopharynx by NAA with non-probe detection|Human coronavirus NL63 RNA [Presence] in Nasopharynx by NAA with non-probe detection
C4264757|T201|LN|82162-9|LNC|Human coronavirus NL63 RNA:PrThr:Pt:Nph:Ord:Non-probe.amp.tar|Human coronavirus NL63 RNA:PrThr:Pt:Nph:Ord:Non-probe.amp.tar
C4264758|T201|DN|82161-1|LNC|HCoV HKU1 RNA NAA+non-probe Ql (Nph)|HCoV HKU1 RNA NAA+non-probe Ql (Nph)
C4264758|T201|OSN|82161-1|LNC|HCoV HKU1 RNA Nph Ql NAA+non-probe|HCoV HKU1 RNA Nph Ql NAA+non-probe
C4264758|T201|MTH_LN|82161-1|LNC|Human coronavirus HKU1 ribonucleic acid:Presence or Threshold:Point in time:Naspopharynx:Ordinal:Non-probe.amp.tar|Human coronavirus HKU1 ribonucleic acid:Presence or Threshold:Point in time:Naspopharynx:Ordinal:Non-probe.amp.tar
C4264758|T201|LC|82161-1|LNC|Human coronavirus HKU1 RNA [Presence] in Nasopharynx by NAA with non-probe detection|Human coronavirus HKU1 RNA [Presence] in Nasopharynx by NAA with non-probe detection
C4264758|T201|LN|82161-1|LNC|Human coronavirus HKU1 RNA:PrThr:Pt:Nph:Ord:Non-probe.amp.tar|Human coronavirus HKU1 RNA:PrThr:Pt:Nph:Ord:Non-probe.amp.tar
C4265422|T201|DN|82164-5|LNC|HCoV OC43 RNA NAA+non-probe Ql (Nph)|HCoV OC43 RNA NAA+non-probe Ql (Nph)
C4265422|T201|OSN|82164-5|LNC|HCoV OC43 RNA Nph Ql NAA+non-probe|HCoV OC43 RNA Nph Ql NAA+non-probe
C4265422|T201|MTH_LN|82164-5|LNC|Human coronavirus OC43 ribonucleic acid:Presence or Threshold:Point in time:Naspopharynx:Ordinal:Non-probe.amp.tar|Human coronavirus OC43 ribonucleic acid:Presence or Threshold:Point in time:Naspopharynx:Ordinal:Non-probe.amp.tar
C4265422|T201|LC|82164-5|LNC|Human coronavirus OC43 RNA [Presence] in Nasopharynx by NAA with non-probe detection|Human coronavirus OC43 RNA [Presence] in Nasopharynx by NAA with non-probe detection
C4265422|T201|LN|82164-5|LNC|Human coronavirus OC43 RNA:PrThr:Pt:Nph:Ord:Non-probe.amp.tar|Human coronavirus OC43 RNA:PrThr:Pt:Nph:Ord:Non-probe.amp.tar
C4265423|T201|DN|82163-7|LNC|HCoV 229E RNA NAA+non-probe Ql (Nph)|HCoV 229E RNA NAA+non-probe Ql (Nph)
C4265423|T201|OSN|82163-7|LNC|HCoV 229E RNA Nph Ql NAA+non-probe|HCoV 229E RNA Nph Ql NAA+non-probe
C4265423|T201|MTH_LN|82163-7|LNC|Human coronavirus 229E ribonucleic acid:Presence or Threshold:Point in time:Naspopharynx:Ordinal:Non-probe.amp.tar|Human coronavirus 229E ribonucleic acid:Presence or Threshold:Point in time:Naspopharynx:Ordinal:Non-probe.amp.tar
C4265423|T201|LC|82163-7|LNC|Human coronavirus 229E RNA [Presence] in Nasopharynx by NAA with non-probe detection|Human coronavirus 229E RNA [Presence] in Nasopharynx by NAA with non-probe detection
C4265423|T201|LN|82163-7|LNC|Human coronavirus 229E RNA:PrThr:Pt:Nph:Ord:Non-probe.amp.tar|Human coronavirus 229E RNA:PrThr:Pt:Nph:Ord:Non-probe.amp.tar
C4274956|T047|PT|715882005|SNOMEDCT_US|Severe acute respiratory syndrome of upper respiratory tract|Severe acute respiratory syndrome of upper respiratory tract
C4274956|T047|FN|715882005|SNOMEDCT_US|Severe acute respiratory syndrome of upper respiratory tract (disorder)|Severe acute respiratory syndrome of upper respiratory tract (disorder)
C4302012|T033|PT|12601000132105|SNOMEDCT_US|Probable SARS (severe acute respiratory syndrome)|Probable SARS (severe acute respiratory syndrome)
C4302012|T033|SY|12601000132105|SNOMEDCT_US|Probable severe acute respiratory syndrome|Probable severe acute respiratory syndrome
C4302012|T033|FN|12601000132105|SNOMEDCT_US|Probable severe acute respiratory syndrome (situation)|Probable severe acute respiratory syndrome (situation)
C4302019|T033|PT|12611000132107|SNOMEDCT_US|SARS (severe acute respiratory syndrome) confirmed|SARS (severe acute respiratory syndrome) confirmed
C4302019|T033|SY|12611000132107|SNOMEDCT_US|Severe acute respiratory syndrome confirmed|Severe acute respiratory syndrome confirmed
C4302019|T033|FN|12611000132107|SNOMEDCT_US|Severe acute respiratory syndrome confirmed (situation)|Severe acute respiratory syndrome confirmed (situation)
C4302020|T033|PT|12591000132100|SNOMEDCT_US|Suspected SARS (severe acute respiratory syndrome)|Suspected SARS (severe acute respiratory syndrome)
C4302020|T033|SY|12591000132100|SNOMEDCT_US|Suspected severe acute respiratory syndrome|Suspected severe acute respiratory syndrome
C4302020|T033|FN|12591000132100|SNOMEDCT_US|Suspected severe acute respiratory syndrome (situation)|Suspected severe acute respiratory syndrome (situation)
C4303065|T005|PT|721884000|SNOMEDCT_US|Bat coronavirus HKU3|Bat coronavirus HKU3
C4303065|T005|FN|721884000|SNOMEDCT_US|Bat coronavirus HKU3 (organism)|Bat coronavirus HKU3 (organism)
C4434726|T005|PEP|D000073638|MSH|Mink coronavirus 1|Mink coronavirus 1
C4434727|T005|PEP|D000073638|MSH|Bat coronavirus CDPHE15|Bat coronavirus CDPHE15
C4434727|T005|PM|D000073638|MSH|Bat coronavirus CDPHE15s|Bat coronavirus CDPHE15s
C4434727|T005|PM|D000073638|MSH|CDPHE15, Bat coronavirus|CDPHE15, Bat coronavirus
C4461651|T005|PEP|D017934|MSH|Coronavirus HKU15|Coronavirus HKU15
C4483677|T201|OSN|86204-5|LNC|PDCoV XXX Ql Cult|PDCoV XXX Ql Cult
C4483677|T201|LC|86204-5|LNC|Porcine deltacoronavirus [Presence] in Unspecified specimen by Organism specific culture|Porcine deltacoronavirus [Presence] in Unspecified specimen by Organism specific culture
C4483677|T201|DN|86204-5|LNC|Porcine deltacoronavirus Org specific cx Ql (Unsp spec)|Porcine deltacoronavirus Org specific cx Ql (Unsp spec)
C4483677|T201|MTH_LN|86204-5|LNC|Porcine deltacoronavirus:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:Organism specific culture|Porcine deltacoronavirus:Presence or Threshold:Point in time:To be specified in another part of the message:Ordinal:Organism specific culture
C4483677|T201|LN|86204-5|LNC|Porcine deltacoronavirus:PrThr:Pt:XXX:Ord:Organism specific culture|Porcine deltacoronavirus:PrThr:Pt:XXX:Ord:Organism specific culture
C4483989|T201|OSN|86578-2|LNC|MERS-CoV RNA Bld Ql NAA+probe|MERS-CoV RNA Bld Ql NAA+probe
C4483989|T201|DN|86578-2|LNC|MERS-CoV RNA NAA+probe Ql (Bld)|MERS-CoV RNA NAA+probe Ql (Bld)
C4483989|T201|LC|86578-2|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Blood by NAA with probe detection|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Blood by NAA with probe detection
C4483989|T201|MTH_LN|86578-2|LNC|Middle East respiratory syndrome coronavirus ribonucleic acid:Presence or Threshold:Point in time:Whole blood:Ordinal:DNA Nucleic Acid Probe.amp.tar|Middle East respiratory syndrome coronavirus ribonucleic acid:Presence or Threshold:Point in time:Whole blood:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4483989|T201|LN|86578-2|LNC|Middle East respiratory syndrome coronavirus RNA:PrThr:Pt:Bld:Ord:Probe.amp.tar|Middle East respiratory syndrome coronavirus RNA:PrThr:Pt:Bld:Ord:Probe.amp.tar
C4483990|T201|DN|86579-0|LNC|MERS-CoV RNA NAA+probe Ql (U)|MERS-CoV RNA NAA+probe Ql (U)
C4483990|T201|OSN|86579-0|LNC|MERS-CoV RNA Ur Ql NAA+probe|MERS-CoV RNA Ur Ql NAA+probe
C4483990|T201|LC|86579-0|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Urine by NAA with probe detection|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Urine by NAA with probe detection
C4483990|T201|MTH_LN|86579-0|LNC|Middle East respiratory syndrome coronavirus ribonucleic acid:Presence or Threshold:Point in time:Urine:Ordinal:DNA Nucleic Acid Probe.amp.tar|Middle East respiratory syndrome coronavirus ribonucleic acid:Presence or Threshold:Point in time:Urine:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4483990|T201|LN|86579-0|LNC|Middle East respiratory syndrome coronavirus RNA:PrThr:Pt:Urine:Ord:Probe.amp.tar|Middle East respiratory syndrome coronavirus RNA:PrThr:Pt:Urine:Ord:Probe.amp.tar
C4484060|T201|MTH_LN|86703-6|LNC|Porcine respiratory coronavirus ribonucleic acid:Threshold Number:Point in time:To be specified in another part of the message:Quantitative:DNA Nucleic Acid Probe.amp.tar|Porcine respiratory coronavirus ribonucleic acid:Threshold Number:Point in time:To be specified in another part of the message:Quantitative:DNA Nucleic Acid Probe.amp.tar
C4484060|T201|LC|86703-6|LNC|Porcine respiratory coronavirus RNA [Cycle Threshold #] in Unspecified specimen by NAA with probe detection|Porcine respiratory coronavirus RNA [Cycle Threshold #] in Unspecified specimen by NAA with probe detection
C4484060|T201|DN|86703-6|LNC|Porcine respiratory coronavirus RNA NAA+probe (Unsp spec) [ThreshNum]|Porcine respiratory coronavirus RNA NAA+probe (Unsp spec) [ThreshNum]
C4484060|T201|LN|86703-6|LNC|Porcine respiratory coronavirus RNA:ThreshNum:Pt:XXX:Qn:Probe.amp.tar|Porcine respiratory coronavirus RNA:ThreshNum:Pt:XXX:Qn:Probe.amp.tar
C4484060|T201|OSN|86703-6|LNC|PRCoV RNA Ct XXX Qn NAA+probe|PRCoV RNA Ct XXX Qn NAA+probe
C4484064|T201|OSN|86711-9|LNC|PDCoV Ag Tiss Ql ImStn|PDCoV Ag Tiss Ql ImStn
C4484064|T201|LC|86711-9|LNC|Porcine deltacoronavirus Ag [Presence] in Tissue by Immune stain|Porcine deltacoronavirus Ag [Presence] in Tissue by Immune stain
C4484064|T201|DN|86711-9|LNC|Porcine deltacoronavirus Ag Immune stain Ql (Tiss)|Porcine deltacoronavirus Ag Immune stain Ql (Tiss)
C4484064|T201|LN|86711-9|LNC|Porcine deltacoronavirus Ag:PrThr:Pt:Tiss:Ord:Immune stain|Porcine deltacoronavirus Ag:PrThr:Pt:Tiss:Ord:Immune stain
C4484064|T201|MTH_LN|86711-9|LNC|Porcine deltacoronavirus Antigen:Presence or Threshold:Point in time:Tissue, unspecified:Ordinal:Immune stain|Porcine deltacoronavirus Antigen:Presence or Threshold:Point in time:Tissue, unspecified:Ordinal:Immune stain
C4484065|T116|LPN|LP248607-6|LNC|Porcine deltacoronavirus Ag|Porcine deltacoronavirus Ag
C4484065|T129|LPN|LP248607-6|LNC|Porcine deltacoronavirus Ag|Porcine deltacoronavirus Ag
C4484065|T116|CN|MTHU056806|LNC|Porcine deltacoronavirus Ag|Porcine deltacoronavirus Ag
C4484065|T129|CN|MTHU056806|LNC|Porcine deltacoronavirus Ag|Porcine deltacoronavirus Ag
C4484065|T116|MTH_CN|MTHU056806|LNC|Porcine deltacoronavirus Antigen|Porcine deltacoronavirus Antigen
C4484065|T129|MTH_CN|MTHU056806|LNC|Porcine deltacoronavirus Antigen|Porcine deltacoronavirus Antigen
C4531941|T201|DN|86927-1|LNC|Porcine respiratory coronavirus Ab/Negative control IA (S) [Relative ratio]|Porcine respiratory coronavirus Ab/Negative control IA (S) [Relative ratio]
C4531941|T201|LC|86927-1|LNC|Porcine respiratory coronavirus Ab/Negative control in Serum by Immunoassay|Porcine respiratory coronavirus Ab/Negative control in Serum by Immunoassay
C4531941|T201|LN|86927-1|LNC|Porcine respiratory coronavirus Ab/Negative control:RelRto:Pt:Ser:Qn:IA|Porcine respiratory coronavirus Ab/Negative control:RelRto:Pt:Ser:Qn:IA
C4531941|T201|MTH_LN|86927-1|LNC|Porcine respiratory coronavirus Antibody/Negative control:Relative Ratio:Point in time:Serum:Quantitative:Enzyme Immunoassay|Porcine respiratory coronavirus Antibody/Negative control:Relative Ratio:Point in time:Serum:Quantitative:Enzyme Immunoassay
C4531941|T201|OSN|86927-1|LNC|PRCoV Ab Ser IA|PRCoV Ab Ser IA
C4531942|T081|LPN|LP286872-9|LNC|Porcine respiratory coronavirus Ab/Negative control|Porcine respiratory coronavirus Ab/Negative control
C4531942|T081|CN|MTHU057282|LNC|Porcine respiratory coronavirus Ab/Negative control|Porcine respiratory coronavirus Ab/Negative control
C4531942|T081|MTH_CN|MTHU057282|LNC|Porcine respiratory coronavirus Antibody/Negative control|Porcine respiratory coronavirus Antibody/Negative control
C4533027|T201|DN|88196-1|LNC|MERS-CoV RNA NAA+probe Ql (Stl)|MERS-CoV RNA NAA+probe Ql (Stl)
C4533027|T201|OSN|88196-1|LNC|MERS-CoV RNA Stl Ql NAA+probe|MERS-CoV RNA Stl Ql NAA+probe
C4533027|T201|LC|88196-1|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Stool by NAA with probe detection|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Stool by NAA with probe detection
C4533027|T201|MTH_LN|88196-1|LNC|Middle East respiratory syndrome coronavirus ribonucleic acid:Presence or Threshold:Point in time:Stool = Fecal:Ordinal:DNA Nucleic Acid Probe.amp.tar|Middle East respiratory syndrome coronavirus ribonucleic acid:Presence or Threshold:Point in time:Stool = Fecal:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4533027|T201|LN|88196-1|LNC|Middle East respiratory syndrome coronavirus RNA:PrThr:Pt:Stool:Ord:Probe.amp.tar|Middle East respiratory syndrome coronavirus RNA:PrThr:Pt:Stool:Ord:Probe.amp.tar
C4533028|T201|DN|88197-9|LNC|MERS-CoV RNA NAA+probe Ql (Nph)|MERS-CoV RNA NAA+probe Ql (Nph)
C4533028|T201|OSN|88197-9|LNC|MERS-CoV RNA Nph Ql NAA+probe|MERS-CoV RNA Nph Ql NAA+probe
C4533028|T201|LC|88197-9|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Nasopharynx by NAA with probe detection|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Nasopharynx by NAA with probe detection
C4533028|T201|MTH_LN|88197-9|LNC|Middle East respiratory syndrome coronavirus ribonucleic acid:Presence or Threshold:Point in time:Naspopharynx:Ordinal:DNA Nucleic Acid Probe.amp.tar|Middle East respiratory syndrome coronavirus ribonucleic acid:Presence or Threshold:Point in time:Naspopharynx:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4533028|T201|LN|88197-9|LNC|Middle East respiratory syndrome coronavirus RNA:PrThr:Pt:Nph:Ord:Probe.amp.tar|Middle East respiratory syndrome coronavirus RNA:PrThr:Pt:Nph:Ord:Probe.amp.tar
C4533029|T201|OSN|88198-7|LNC|MERS-CoV RNA Corn/Cnjt Ql NAA+probe|MERS-CoV RNA Corn/Cnjt Ql NAA+probe
C4533029|T201|DN|88198-7|LNC|MERS-CoV RNA NAA+probe Ql (Corn/Cnjt)|MERS-CoV RNA NAA+probe Ql (Corn/Cnjt)
C4533029|T201|LC|88198-7|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Cornea or Conjunctiva by NAA with probe detection|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Cornea or Conjunctiva by NAA with probe detection
C4533029|T201|MTH_LN|88198-7|LNC|Middle East respiratory syndrome coronavirus ribonucleic acid:Presence or Threshold:Point in time:Cornea/Conjunctiva:Ordinal:DNA Nucleic Acid Probe.amp.tar|Middle East respiratory syndrome coronavirus ribonucleic acid:Presence or Threshold:Point in time:Cornea/Conjunctiva:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4533029|T201|LN|88198-7|LNC|Middle East respiratory syndrome coronavirus RNA:PrThr:Pt:Cornea/Conjunctiva:Ord:Probe.amp.tar|Middle East respiratory syndrome coronavirus RNA:PrThr:Pt:Cornea/Conjunctiva:Ord:Probe.amp.tar
C4533599|T201|OSN|88199-5|LNC|MERS-CoV RNA Aspirate Ql NAA+probe|MERS-CoV RNA Aspirate Ql NAA+probe
C4533599|T201|DN|88199-5|LNC|MERS-CoV RNA NAA+probe Ql (Asp)|MERS-CoV RNA NAA+probe Ql (Asp)
C4533599|T201|LC|88199-5|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Aspirate by NAA with probe detection|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Aspirate by NAA with probe detection
C4533599|T201|MTH_LN|88199-5|LNC|Middle East respiratory syndrome coronavirus ribonucleic acid:Presence or Threshold:Point in time:Aspirate:Ordinal:DNA Nucleic Acid Probe.amp.tar|Middle East respiratory syndrome coronavirus ribonucleic acid:Presence or Threshold:Point in time:Aspirate:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4533599|T201|LN|88199-5|LNC|Middle East respiratory syndrome coronavirus RNA:PrThr:Pt:Asp:Ord:Probe.amp.tar|Middle East respiratory syndrome coronavirus RNA:PrThr:Pt:Asp:Ord:Probe.amp.tar
C4536544|T047|PT|366307|MEDCIN|human coronavirus pneumonia|human coronavirus pneumonia
C4536544|T047|FN|366307|MEDCIN|human coronavirus pneumonia (diagnosis)|human coronavirus pneumonia (diagnosis)
C4536544|T047|SY|366307|MEDCIN|viral pneumonia human coronavirus|viral pneumonia human coronavirus
C4609501|T005|CE|C000627033|MSH|SADS-CoV|SADS-CoV
C4609501|T005|NM|C000627033|MSH|Swine acute diarrhea syndrome coronavirus|Swine acute diarrhea syndrome coronavirus
C4695210|T201|DN|88604-4|LNC|HCoV HKU1 RNA NAA+probe Ql (Upper resp)|HCoV HKU1 RNA NAA+probe Ql (Upper resp)
C4695210|T201|OSN|88604-4|LNC|HCoV HKU1 RNA Up resp Ql NAA+probe|HCoV HKU1 RNA Up resp Ql NAA+probe
C4695210|T201|MTH_LN|88604-4|LNC|Human coronavirus HKU1 ribonucleic acid:Presence or Threshold:Point in time:Respiratory.upper:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus HKU1 ribonucleic acid:Presence or Threshold:Point in time:Respiratory.upper:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4695210|T201|LC|88604-4|LNC|Human coronavirus HKU1 RNA [Presence] in Upper respiratory specimen by NAA with probe detection|Human coronavirus HKU1 RNA [Presence] in Upper respiratory specimen by NAA with probe detection
C4695210|T201|LN|88604-4|LNC|Human coronavirus HKU1 RNA:PrThr:Pt:Respiratory.upper:Ord:Probe.amp.tar|Human coronavirus HKU1 RNA:PrThr:Pt:Respiratory.upper:Ord:Probe.amp.tar
C4695211|T201|OSN|88605-1|LNC|HCoV OC43 RNA Lower Resp Ql NAA+probe|HCoV OC43 RNA Lower Resp Ql NAA+probe
C4695211|T201|DN|88605-1|LNC|HCoV OC43 RNA NAA+probe Ql (Lower resp)|HCoV OC43 RNA NAA+probe Ql (Lower resp)
C4695211|T201|MTH_LN|88605-1|LNC|Human coronavirus OC43 ribonucleic acid:Presence or Threshold:Point in time:Respiratory.lower:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus OC43 ribonucleic acid:Presence or Threshold:Point in time:Respiratory.lower:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4695211|T201|LC|88605-1|LNC|Human coronavirus OC43 RNA [Presence] in Lower respiratory specimen by NAA with probe detection|Human coronavirus OC43 RNA [Presence] in Lower respiratory specimen by NAA with probe detection
C4695211|T201|LN|88605-1|LNC|Human coronavirus OC43 RNA:PrThr:Pt:Respiratory.lower:Ord:Probe.amp.tar|Human coronavirus OC43 RNA:PrThr:Pt:Respiratory.lower:Ord:Probe.amp.tar
C4695213|T201|OSN|88607-7|LNC|HCoV 229E RNA Aspirate Ql NAA+probe|HCoV 229E RNA Aspirate Ql NAA+probe
C4695213|T201|DN|88607-7|LNC|HCoV 229E RNA NAA+probe Ql (Asp)|HCoV 229E RNA NAA+probe Ql (Asp)
C4695213|T201|MTH_LN|88607-7|LNC|Human coronavirus 229E ribonucleic acid:Presence or Threshold:Point in time:Aspirate:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus 229E ribonucleic acid:Presence or Threshold:Point in time:Aspirate:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4695213|T201|LC|88607-7|LNC|Human coronavirus 229E RNA [Presence] in Aspirate by NAA with probe detection|Human coronavirus 229E RNA [Presence] in Aspirate by NAA with probe detection
C4695213|T201|LN|88607-7|LNC|Human coronavirus 229E RNA:PrThr:Pt:Asp:Ord:Probe.amp.tar|Human coronavirus 229E RNA:PrThr:Pt:Asp:Ord:Probe.amp.tar
C4695214|T201|OSN|88608-5|LNC|HCoV 229E RNA Lower Resp Ql NAA+probe|HCoV 229E RNA Lower Resp Ql NAA+probe
C4695214|T201|DN|88608-5|LNC|HCoV 229E RNA NAA+probe Ql (Lower resp)|HCoV 229E RNA NAA+probe Ql (Lower resp)
C4695214|T201|MTH_LN|88608-5|LNC|Human coronavirus 229E ribonucleic acid:Presence or Threshold:Point in time:Respiratory.lower:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus 229E ribonucleic acid:Presence or Threshold:Point in time:Respiratory.lower:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4695214|T201|LC|88608-5|LNC|Human coronavirus 229E RNA [Presence] in Lower respiratory specimen by NAA with probe detection|Human coronavirus 229E RNA [Presence] in Lower respiratory specimen by NAA with probe detection
C4695214|T201|LN|88608-5|LNC|Human coronavirus 229E RNA:PrThr:Pt:Respiratory.lower:Ord:Probe.amp.tar|Human coronavirus 229E RNA:PrThr:Pt:Respiratory.lower:Ord:Probe.amp.tar
C4695736|T201|OSN|88594-7|LNC|HCoV HKU1 RNA Lower Resp Ql NAA+probe|HCoV HKU1 RNA Lower Resp Ql NAA+probe
C4695736|T201|DN|88594-7|LNC|HCoV HKU1 RNA NAA+probe Ql (Lower resp)|HCoV HKU1 RNA NAA+probe Ql (Lower resp)
C4695736|T201|MTH_LN|88594-7|LNC|Human coronavirus HKU1 ribonucleic acid:Presence or Threshold:Point in time:Respiratory.lower:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus HKU1 ribonucleic acid:Presence or Threshold:Point in time:Respiratory.lower:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4695736|T201|LC|88594-7|LNC|Human coronavirus HKU1 RNA [Presence] in Lower respiratory specimen by NAA with probe detection|Human coronavirus HKU1 RNA [Presence] in Lower respiratory specimen by NAA with probe detection
C4695736|T201|LN|88594-7|LNC|Human coronavirus HKU1 RNA:PrThr:Pt:Respiratory.lower:Ord:Probe.amp.tar|Human coronavirus HKU1 RNA:PrThr:Pt:Respiratory.lower:Ord:Probe.amp.tar
C4695746|T201|OSN|88609-3|LNC|HCoV 229E RNA Corn/Cnjt Ql NAA+probe|HCoV 229E RNA Corn/Cnjt Ql NAA+probe
C4695746|T201|DN|88609-3|LNC|HCoV 229E RNA NAA+probe Ql (Corn/Cnjt)|HCoV 229E RNA NAA+probe Ql (Corn/Cnjt)
C4695746|T201|MTH_LN|88609-3|LNC|Human coronavirus 229E ribonucleic acid:Presence or Threshold:Point in time:Cornea/Conjunctiva:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus 229E ribonucleic acid:Presence or Threshold:Point in time:Cornea/Conjunctiva:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4695746|T201|LC|88609-3|LNC|Human coronavirus 229E RNA [Presence] in Cornea or Conjunctiva by NAA with probe detection|Human coronavirus 229E RNA [Presence] in Cornea or Conjunctiva by NAA with probe detection
C4695746|T201|LN|88609-3|LNC|Human coronavirus 229E RNA:PrThr:Pt:Cornea/Conjunctiva:Ord:Probe.amp.tar|Human coronavirus 229E RNA:PrThr:Pt:Cornea/Conjunctiva:Ord:Probe.amp.tar
C4695747|T201|DN|88610-1|LNC|HCoV 229E RNA NAA+probe Ql (Upper resp)|HCoV 229E RNA NAA+probe Ql (Upper resp)
C4695747|T201|OSN|88610-1|LNC|HCoV 229E RNA Up resp Ql NAA+probe|HCoV 229E RNA Up resp Ql NAA+probe
C4695747|T201|MTH_LN|88610-1|LNC|Human coronavirus 229E ribonucleic acid:Presence or Threshold:Point in time:Respiratory.upper:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus 229E ribonucleic acid:Presence or Threshold:Point in time:Respiratory.upper:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4695747|T201|LC|88610-1|LNC|Human coronavirus 229E RNA [Presence] in Upper respiratory specimen by NAA with probe detection|Human coronavirus 229E RNA [Presence] in Upper respiratory specimen by NAA with probe detection
C4695747|T201|LN|88610-1|LNC|Human coronavirus 229E RNA:PrThr:Pt:Respiratory.upper:Ord:Probe.amp.tar|Human coronavirus 229E RNA:PrThr:Pt:Respiratory.upper:Ord:Probe.amp.tar
C4695748|T201|OSN|88611-9|LNC|HCoV HKU1 RNA Aspirate Ql NAA+probe|HCoV HKU1 RNA Aspirate Ql NAA+probe
C4695748|T201|DN|88611-9|LNC|HCoV HKU1 RNA NAA+probe Ql (Asp)|HCoV HKU1 RNA NAA+probe Ql (Asp)
C4695748|T201|MTH_LN|88611-9|LNC|Human coronavirus HKU1 ribonucleic acid:Presence or Threshold:Point in time:Aspirate:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus HKU1 ribonucleic acid:Presence or Threshold:Point in time:Aspirate:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4695748|T201|LC|88611-9|LNC|Human coronavirus HKU1 RNA [Presence] in Aspirate by NAA with probe detection|Human coronavirus HKU1 RNA [Presence] in Aspirate by NAA with probe detection
C4695748|T201|LN|88611-9|LNC|Human coronavirus HKU1 RNA:PrThr:Pt:Asp:Ord:Probe.amp.tar|Human coronavirus HKU1 RNA:PrThr:Pt:Asp:Ord:Probe.amp.tar
C4695749|T201|OSN|88612-7|LNC|HCoV HKU1 RNA Corn/Cnjt Ql NAA+probe|HCoV HKU1 RNA Corn/Cnjt Ql NAA+probe
C4695749|T201|DN|88612-7|LNC|HCoV HKU1 RNA NAA+probe Ql (Corn/Cnjt)|HCoV HKU1 RNA NAA+probe Ql (Corn/Cnjt)
C4695749|T201|MTH_LN|88612-7|LNC|Human coronavirus HKU1 ribonucleic acid:Presence or Threshold:Point in time:Cornea/Conjunctiva:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus HKU1 ribonucleic acid:Presence or Threshold:Point in time:Cornea/Conjunctiva:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4695749|T201|LC|88612-7|LNC|Human coronavirus HKU1 RNA [Presence] in Cornea or Conjunctiva by NAA with probe detection|Human coronavirus HKU1 RNA [Presence] in Cornea or Conjunctiva by NAA with probe detection
C4695749|T201|LN|88612-7|LNC|Human coronavirus HKU1 RNA:PrThr:Pt:Cornea/Conjunctiva:Ord:Probe.amp.tar|Human coronavirus HKU1 RNA:PrThr:Pt:Cornea/Conjunctiva:Ord:Probe.amp.tar
C4695751|T201|OSN|88614-3|LNC|HCoV RNA Aspirate Ql NAA+probe|HCoV RNA Aspirate Ql NAA+probe
C4695751|T201|DN|88614-3|LNC|HCoV RNA NAA+probe Ql (Asp)|HCoV RNA NAA+probe Ql (Asp)
C4695751|T201|MTH_LN|88614-3|LNC|Human coronavirus ribonucleic acid:Presence or Threshold:Point in time:Aspirate:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus ribonucleic acid:Presence or Threshold:Point in time:Aspirate:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4695751|T201|LC|88614-3|LNC|Human coronavirus RNA [Presence] in Aspirate by NAA with probe detection|Human coronavirus RNA [Presence] in Aspirate by NAA with probe detection
C4695751|T201|LN|88614-3|LNC|Human coronavirus RNA:PrThr:Pt:Asp:Ord:Probe.amp.tar|Human coronavirus RNA:PrThr:Pt:Asp:Ord:Probe.amp.tar
C4695752|T201|OSN|88615-0|LNC|HCoV NL63 RNA Aspirate Ql NAA+probe|HCoV NL63 RNA Aspirate Ql NAA+probe
C4695752|T201|DN|88615-0|LNC|HCoV NL63 RNA NAA+probe Ql (Asp)|HCoV NL63 RNA NAA+probe Ql (Asp)
C4695752|T201|MTH_LN|88615-0|LNC|Human coronavirus NL63 ribonucleic acid:Presence or Threshold:Point in time:Aspirate:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus NL63 ribonucleic acid:Presence or Threshold:Point in time:Aspirate:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4695752|T201|LC|88615-0|LNC|Human coronavirus NL63 RNA [Presence] in Aspirate by NAA with probe detection|Human coronavirus NL63 RNA [Presence] in Aspirate by NAA with probe detection
C4695752|T201|LN|88615-0|LNC|Human coronavirus NL63 RNA:PrThr:Pt:Asp:Ord:Probe.amp.tar|Human coronavirus NL63 RNA:PrThr:Pt:Asp:Ord:Probe.amp.tar
C4695753|T201|OSN|88616-8|LNC|HCoV NL63 RNA Lower Resp Ql NAA+probe|HCoV NL63 RNA Lower Resp Ql NAA+probe
C4695753|T201|DN|88616-8|LNC|HCoV NL63 RNA NAA+probe Ql (Lower resp)|HCoV NL63 RNA NAA+probe Ql (Lower resp)
C4695753|T201|MTH_LN|88616-8|LNC|Human coronavirus NL63 ribonucleic acid:Presence or Threshold:Point in time:Respiratory.lower:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus NL63 ribonucleic acid:Presence or Threshold:Point in time:Respiratory.lower:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4695753|T201|LC|88616-8|LNC|Human coronavirus NL63 RNA [Presence] in Lower respiratory specimen by NAA with probe detection|Human coronavirus NL63 RNA [Presence] in Lower respiratory specimen by NAA with probe detection
C4695753|T201|LN|88616-8|LNC|Human coronavirus NL63 RNA:PrThr:Pt:Respiratory.lower:Ord:Probe.amp.tar|Human coronavirus NL63 RNA:PrThr:Pt:Respiratory.lower:Ord:Probe.amp.tar
C4695754|T201|OSN|88617-6|LNC|HCoV NL63 RNA Corn/Cnjt Ql NAA+probe|HCoV NL63 RNA Corn/Cnjt Ql NAA+probe
C4695754|T201|DN|88617-6|LNC|HCoV NL63 RNA NAA+probe Ql (Corn/Cnjt)|HCoV NL63 RNA NAA+probe Ql (Corn/Cnjt)
C4695754|T201|MTH_LN|88617-6|LNC|Human coronavirus NL63 ribonucleic acid:Presence or Threshold:Point in time:Cornea/Conjunctiva:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus NL63 ribonucleic acid:Presence or Threshold:Point in time:Cornea/Conjunctiva:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4695754|T201|LC|88617-6|LNC|Human coronavirus NL63 RNA [Presence] in Cornea or Conjunctiva by NAA with probe detection|Human coronavirus NL63 RNA [Presence] in Cornea or Conjunctiva by NAA with probe detection
C4695754|T201|LN|88617-6|LNC|Human coronavirus NL63 RNA:PrThr:Pt:Cornea/Conjunctiva:Ord:Probe.amp.tar|Human coronavirus NL63 RNA:PrThr:Pt:Cornea/Conjunctiva:Ord:Probe.amp.tar
C4695755|T201|DN|88618-4|LNC|HCoV NL63 RNA NAA+probe Ql (Upper resp)|HCoV NL63 RNA NAA+probe Ql (Upper resp)
C4695755|T201|OSN|88618-4|LNC|HCoV NL63 RNA Up resp Ql NAA+probe|HCoV NL63 RNA Up resp Ql NAA+probe
C4695755|T201|MTH_LN|88618-4|LNC|Human coronavirus NL63 ribonucleic acid:Presence or Threshold:Point in time:Respiratory.upper:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus NL63 ribonucleic acid:Presence or Threshold:Point in time:Respiratory.upper:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4695755|T201|LC|88618-4|LNC|Human coronavirus NL63 RNA [Presence] in Upper respiratory specimen by NAA with probe detection|Human coronavirus NL63 RNA [Presence] in Upper respiratory specimen by NAA with probe detection
C4695755|T201|LN|88618-4|LNC|Human coronavirus NL63 RNA:PrThr:Pt:Respiratory.upper:Ord:Probe.amp.tar|Human coronavirus NL63 RNA:PrThr:Pt:Respiratory.upper:Ord:Probe.amp.tar
C4695756|T201|OSN|88619-2|LNC|HCoV OC43 RNA Aspirate Ql NAA+probe|HCoV OC43 RNA Aspirate Ql NAA+probe
C4695756|T201|DN|88619-2|LNC|HCoV OC43 RNA NAA+probe Ql (Asp)|HCoV OC43 RNA NAA+probe Ql (Asp)
C4695756|T201|MTH_LN|88619-2|LNC|Human coronavirus OC43 ribonucleic acid:Presence or Threshold:Point in time:Aspirate:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus OC43 ribonucleic acid:Presence or Threshold:Point in time:Aspirate:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4695756|T201|LC|88619-2|LNC|Human coronavirus OC43 RNA [Presence] in Aspirate by NAA with probe detection|Human coronavirus OC43 RNA [Presence] in Aspirate by NAA with probe detection
C4695756|T201|LN|88619-2|LNC|Human coronavirus OC43 RNA:PrThr:Pt:Asp:Ord:Probe.amp.tar|Human coronavirus OC43 RNA:PrThr:Pt:Asp:Ord:Probe.amp.tar
C4695757|T201|OSN|88620-0|LNC|HCoV RNA Lower Resp Ql NAA+probe|HCoV RNA Lower Resp Ql NAA+probe
C4695757|T201|DN|88620-0|LNC|HCoV RNA NAA+probe Ql (Lower resp)|HCoV RNA NAA+probe Ql (Lower resp)
C4695757|T201|MTH_LN|88620-0|LNC|Human coronavirus ribonucleic acid:Presence or Threshold:Point in time:Respiratory.lower:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus ribonucleic acid:Presence or Threshold:Point in time:Respiratory.lower:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4695757|T201|LC|88620-0|LNC|Human coronavirus RNA [Presence] in Lower respiratory specimen by NAA with probe detection|Human coronavirus RNA [Presence] in Lower respiratory specimen by NAA with probe detection
C4695757|T201|LN|88620-0|LNC|Human coronavirus RNA:PrThr:Pt:Respiratory.lower:Ord:Probe.amp.tar|Human coronavirus RNA:PrThr:Pt:Respiratory.lower:Ord:Probe.amp.tar
C4695758|T201|OSN|88621-8|LNC|HCoV OC43 RNA Corn/Cnjt Ql NAA+probe|HCoV OC43 RNA Corn/Cnjt Ql NAA+probe
C4695758|T201|DN|88621-8|LNC|HCoV OC43 RNA NAA+probe Ql (Corn/Cnjt)|HCoV OC43 RNA NAA+probe Ql (Corn/Cnjt)
C4695758|T201|MTH_LN|88621-8|LNC|Human coronavirus OC43 ribonucleic acid:Presence or Threshold:Point in time:Cornea/Conjunctiva:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus OC43 ribonucleic acid:Presence or Threshold:Point in time:Cornea/Conjunctiva:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4695758|T201|LC|88621-8|LNC|Human coronavirus OC43 RNA [Presence] in Cornea or Conjunctiva by NAA with probe detection|Human coronavirus OC43 RNA [Presence] in Cornea or Conjunctiva by NAA with probe detection
C4695758|T201|LN|88621-8|LNC|Human coronavirus OC43 RNA:PrThr:Pt:Cornea/Conjunctiva:Ord:Probe.amp.tar|Human coronavirus OC43 RNA:PrThr:Pt:Cornea/Conjunctiva:Ord:Probe.amp.tar
C4695763|T201|DN|88626-7|LNC|HCoV OC43 RNA NAA+probe Ql (Upper resp)|HCoV OC43 RNA NAA+probe Ql (Upper resp)
C4695763|T201|OSN|88626-7|LNC|HCoV OC43 RNA Up resp Ql NAA+probe|HCoV OC43 RNA Up resp Ql NAA+probe
C4695763|T201|MTH_LN|88626-7|LNC|Human coronavirus OC43 ribonucleic acid:Presence or Threshold:Point in time:Respiratory.upper:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus OC43 ribonucleic acid:Presence or Threshold:Point in time:Respiratory.upper:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4695763|T201|LC|88626-7|LNC|Human coronavirus OC43 RNA [Presence] in Upper respiratory specimen by NAA with probe detection|Human coronavirus OC43 RNA [Presence] in Upper respiratory specimen by NAA with probe detection
C4695763|T201|LN|88626-7|LNC|Human coronavirus OC43 RNA:PrThr:Pt:Respiratory.upper:Ord:Probe.amp.tar|Human coronavirus OC43 RNA:PrThr:Pt:Respiratory.upper:Ord:Probe.amp.tar
C4695764|T201|DN|88627-5|LNC|HCoV RNA NAA+probe Ql (Upper resp)|HCoV RNA NAA+probe Ql (Upper resp)
C4695764|T201|OSN|88627-5|LNC|HCoV RNA Up resp Ql NAA+probe|HCoV RNA Up resp Ql NAA+probe
C4695764|T201|MTH_LN|88627-5|LNC|Human coronavirus ribonucleic acid:Presence or Threshold:Point in time:Respiratory.upper:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus ribonucleic acid:Presence or Threshold:Point in time:Respiratory.upper:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4695764|T201|LC|88627-5|LNC|Human coronavirus RNA [Presence] in Upper respiratory specimen by NAA with probe detection|Human coronavirus RNA [Presence] in Upper respiratory specimen by NAA with probe detection
C4695764|T201|LN|88627-5|LNC|Human coronavirus RNA:PrThr:Pt:Respiratory.upper:Ord:Probe.amp.tar|Human coronavirus RNA:PrThr:Pt:Respiratory.upper:Ord:Probe.amp.tar
C4695765|T201|OSN|88628-3|LNC|HCoV RNA Corn/Cnjt Ql NAA+probe|HCoV RNA Corn/Cnjt Ql NAA+probe
C4695765|T201|DN|88628-3|LNC|HCoV RNA NAA+probe Ql (Corn/Cnjt)|HCoV RNA NAA+probe Ql (Corn/Cnjt)
C4695765|T201|MTH_LN|88628-3|LNC|Human coronavirus ribonucleic acid:Presence or Threshold:Point in time:Cornea/Conjunctiva:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus ribonucleic acid:Presence or Threshold:Point in time:Cornea/Conjunctiva:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4695765|T201|LC|88628-3|LNC|Human coronavirus RNA [Presence] in Cornea or Conjunctiva by NAA with probe detection|Human coronavirus RNA [Presence] in Cornea or Conjunctiva by NAA with probe detection
C4695765|T201|LN|88628-3|LNC|Human coronavirus RNA:PrThr:Pt:Cornea/Conjunctiva:Ord:Probe.amp.tar|Human coronavirus RNA:PrThr:Pt:Cornea/Conjunctiva:Ord:Probe.amp.tar
C4695840|T201|OSN|88719-0|LNC|HCoV 229E+HKU1+NL63+OC43 Nph Ql NAA+Pr|HCoV 229E+HKU1+NL63+OC43 Nph Ql NAA+Pr
C4695840|T201|DN|88719-0|LNC|HCoV 229E+HKU1+NL63+OC43 RNA NAA+probe Ql (Nph)|HCoV 229E+HKU1+NL63+OC43 RNA NAA+probe Ql (Nph)
C4695840|T201|MTH_LN|88719-0|LNC|Human coronavirus 229E+HKU1+NL63+OC43 ribonucleic acid:Presence or Threshold:Point in time:Naspopharynx:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus 229E+HKU1+NL63+OC43 ribonucleic acid:Presence or Threshold:Point in time:Naspopharynx:Ordinal:DNA Nucleic Acid Probe.amp.tar
C4695840|T201|LC|88719-0|LNC|Human coronavirus 229E+HKU1+NL63+OC43 RNA [Presence] in Nasopharynx by NAA with probe detection|Human coronavirus 229E+HKU1+NL63+OC43 RNA [Presence] in Nasopharynx by NAA with probe detection
C4695840|T201|LN|88719-0|LNC|Human coronavirus 229E+HKU1+NL63+OC43 RNA:PrThr:Pt:Nph:Ord:Probe.amp.tar|Human coronavirus 229E+HKU1+NL63+OC43 RNA:PrThr:Pt:Nph:Ord:Probe.amp.tar
C4695841|T114|MTH_CN|MTHU058503|LNC|Human coronavirus 229E+HKU1+NL63+OC43 ribonucleic acid|Human coronavirus 229E+HKU1+NL63+OC43 ribonucleic acid
C4695841|T114|LPN|LP263694-4|LNC|Human coronavirus 229E+HKU1+NL63+OC43 RNA|Human coronavirus 229E+HKU1+NL63+OC43 RNA
C4695841|T114|CN|MTHU058503|LNC|Human coronavirus 229E+HKU1+NL63+OC43 RNA|Human coronavirus 229E+HKU1+NL63+OC43 RNA
C4696149|T201|DN|88889-1|LNC|MERS-CoV RNA NAA+non-probe Ql (Nph)|MERS-CoV RNA NAA+non-probe Ql (Nph)
C4696149|T201|OSN|88889-1|LNC|MERS-CoV RNA Nph Ql NAA+non-probe|MERS-CoV RNA Nph Ql NAA+non-probe
C4696149|T201|LC|88889-1|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Nasopharynx by NAA with non-probe detection|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Nasopharynx by NAA with non-probe detection
C4696149|T201|MTH_LN|88889-1|LNC|Middle east respiratory syndrome coronavirus ribonucleic acid:Presence or Threshold:Point in time:Naspopharynx:Ordinal:Non-probe.amp.tar|Middle east respiratory syndrome coronavirus ribonucleic acid:Presence or Threshold:Point in time:Naspopharynx:Ordinal:Non-probe.amp.tar
C4696149|T201|LN|88889-1|LNC|Middle east respiratory syndrome coronavirus RNA:PrThr:Pt:Nph:Ord:Non-probe.amp.tar|Middle east respiratory syndrome coronavirus RNA:PrThr:Pt:Nph:Ord:Non-probe.amp.tar
C4696152|T201|OSN|88891-7|LNC|HCoV 229E+HKU1+NL63+OC43 Np Ql NAA+nonpr|HCoV 229E+HKU1+NL63+OC43 Np Ql NAA+nonpr
C4696152|T201|DN|88891-7|LNC|HCoV 229E+HKU1+NL63+OC43 RNA NAA+non-probe Ql (Nph)|HCoV 229E+HKU1+NL63+OC43 RNA NAA+non-probe Ql (Nph)
C4696152|T201|MTH_LN|88891-7|LNC|Human coronavirus 229E+HKU1+NL63+OC43 ribonucleic acid:Presence or Threshold:Point in time:Naspopharynx:Ordinal:Non-probe.amp.tar|Human coronavirus 229E+HKU1+NL63+OC43 ribonucleic acid:Presence or Threshold:Point in time:Naspopharynx:Ordinal:Non-probe.amp.tar
C4696152|T201|LC|88891-7|LNC|Human coronavirus 229E+HKU1+NL63+OC43 RNA [Presence] in Nasopharynx by NAA with non-probe detection|Human coronavirus 229E+HKU1+NL63+OC43 RNA [Presence] in Nasopharynx by NAA with non-probe detection
C4696152|T201|LN|88891-7|LNC|Human coronavirus 229E+HKU1+NL63+OC43 RNA:PrThr:Pt:Nph:Ord:Non-probe.amp.tar|Human coronavirus 229E+HKU1+NL63+OC43 RNA:PrThr:Pt:Nph:Ord:Non-probe.amp.tar
C4697044|T005|LPN|LP263700-9|LNC|Human coronavirus 229E+HKU1+NL63+OC43|Human coronavirus 229E+HKU1+NL63+OC43
C4699345|T005|LA|LA26148-9|LNC|Coronavirus OC43|Coronavirus OC43
C4699346|T005|LA|LA26150-5|LNC|Coronavirus HKU1|Coronavirus HKU1
C4739655|T201|OSN|90329-4|LNC|PDCoV IgG/Pos cntrl XXX IA|PDCoV IgG/Pos cntrl XXX IA
C4739655|T201|LN|90329-4|LNC|Porcine deltacoronavirus Ab.IgG/Positive control:RelRto:Pt:XXX:Qn:IA|Porcine deltacoronavirus Ab.IgG/Positive control:RelRto:Pt:XXX:Qn:IA
C4739655|T201|MTH_LN|90329-4|LNC|Porcine deltacoronavirus Antibody.immunoglobulin G/Positive control:Relative Ratio:Point in time:To be specified in another part of the message:Quantitative:Enzyme Immunoassay|Porcine deltacoronavirus Antibody.immunoglobulin G/Positive control:Relative Ratio:Point in time:To be specified in another part of the message:Quantitative:Enzyme Immunoassay
C4739655|T201|LC|90329-4|LNC|Porcine deltacoronavirus IgG Ab/Positive control in Unspecified specimen by Immunoassay|Porcine deltacoronavirus IgG Ab/Positive control in Unspecified specimen by Immunoassay
C4739655|T201|DN|90329-4|LNC|Porcine deltacoronavirus IgG/Positive control IA (Unsp spec) [Relative ratio]|Porcine deltacoronavirus IgG/Positive control IA (Unsp spec) [Relative ratio]
C4739656|T081|LPN|LP286860-4|LNC|Porcine deltacoronavirus Ab.IgG/Positive control|Porcine deltacoronavirus Ab.IgG/Positive control
C4739656|T081|CN|MTHU060187|LNC|Porcine deltacoronavirus Ab.IgG/Positive control|Porcine deltacoronavirus Ab.IgG/Positive control
C4739656|T081|MTH_CN|MTHU060187|LNC|Porcine deltacoronavirus Antibody.immunoglobulin G/Positive control|Porcine deltacoronavirus Antibody.immunoglobulin G/Positive control
C4740230|T116|LPN|LP267191-7|LNC|Porcine deltacoronavirus Ab|Porcine deltacoronavirus Ab
C4740230|T129|LPN|LP267191-7|LNC|Porcine deltacoronavirus Ab|Porcine deltacoronavirus Ab
C4740760|T116|LPN|LP267190-9|LNC|Porcine deltacoronavirus Ab.IgG|Porcine deltacoronavirus Ab.IgG
C4740760|T129|LPN|LP267190-9|LNC|Porcine deltacoronavirus Ab.IgG|Porcine deltacoronavirus Ab.IgG
C5142245|T114|MTH_CN|MTHU062283|LNC|Human coronavirus 229E+NL63 ribonucleic acid|Human coronavirus 229E+NL63 ribonucleic acid
C5142245|T114|LPN|LP341566-0|LNC|Human coronavirus 229E+NL63 RNA|Human coronavirus 229E+NL63 RNA
C5142245|T114|CN|MTHU062283|LNC|Human coronavirus 229E+NL63 RNA|Human coronavirus 229E+NL63 RNA
C5142246|T114|MTH_CN|MTHU062284|LNC|Human coronavirus HKU1+OC43 ribonucleic acid|Human coronavirus HKU1+OC43 ribonucleic acid
C5142246|T114|LPN|LP341563-7|LNC|Human coronavirus HKU1+OC43 RNA|Human coronavirus HKU1+OC43 RNA
C5142246|T114|CN|MTHU062284|LNC|Human coronavirus HKU1+OC43 RNA|Human coronavirus HKU1+OC43 RNA
C5142650|T059|MTH_CN|MTHU062830|LNC|Human coronavirus 229E+HKU1+NL63+OC43 & Parainfluenza virus 1+2+3+4 ribonucleic acid panel|Human coronavirus 229E+HKU1+NL63+OC43 & Parainfluenza virus 1+2+3+4 ribonucleic acid panel
C5142650|T059|LPN|LP344992-5|LNC|Human coronavirus 229E+HKU1+NL63+OC43 & Parainfluenza virus 1+2+3+4 RNA panel|Human coronavirus 229E+HKU1+NL63+OC43 & Parainfluenza virus 1+2+3+4 RNA panel
C5142650|T059|CN|MTHU062830|LNC|Human coronavirus 229E+HKU1+NL63+OC43 & Parainfluenza virus 1+2+3+4 RNA panel|Human coronavirus 229E+HKU1+NL63+OC43 & Parainfluenza virus 1+2+3+4 RNA panel
C5143877|T201|DN|91807-8|LNC|MERS-CoV RNA NAA+probe Ql (Upper resp)|MERS-CoV RNA NAA+probe Ql (Upper resp)
C5143877|T201|OSN|91807-8|LNC|MERS-CoV RNA Up resp Ql NAA+probe|MERS-CoV RNA Up resp Ql NAA+probe
C5143877|T201|LC|91807-8|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Upper respiratory specimen by NAA with probe detection|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Upper respiratory specimen by NAA with probe detection
C5143877|T201|MTH_LN|91807-8|LNC|Middle east respiratory syndrome coronavirus ribonucleic acid:Presence or Threshold:Point in time:Respiratory.upper:Ordinal:DNA Nucleic Acid Probe.amp.tar|Middle east respiratory syndrome coronavirus ribonucleic acid:Presence or Threshold:Point in time:Respiratory.upper:Ordinal:DNA Nucleic Acid Probe.amp.tar
C5143877|T201|LN|91807-8|LNC|Middle east respiratory syndrome coronavirus RNA:PrThr:Pt:Respiratory.upper:Ord:Probe.amp.tar|Middle east respiratory syndrome coronavirus RNA:PrThr:Pt:Respiratory.upper:Ord:Probe.amp.tar
C5143900|T201|OSN|91830-0|LNC|MERS-CoV RNA Lower Resp Ql NAA+probe|MERS-CoV RNA Lower Resp Ql NAA+probe
C5143900|T201|DN|91830-0|LNC|MERS-CoV RNA NAA+probe Ql (Lower resp)|MERS-CoV RNA NAA+probe Ql (Lower resp)
C5143900|T201|LC|91830-0|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Lower respiratory specimen by NAA with probe detection|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Lower respiratory specimen by NAA with probe detection
C5143900|T201|MTH_LN|91830-0|LNC|Middle east respiratory syndrome coronavirus ribonucleic acid:Presence or Threshold:Point in time:Respiratory.lower:Ordinal:DNA Nucleic Acid Probe.amp.tar|Middle east respiratory syndrome coronavirus ribonucleic acid:Presence or Threshold:Point in time:Respiratory.lower:Ordinal:DNA Nucleic Acid Probe.amp.tar
C5143900|T201|LN|91830-0|LNC|Middle east respiratory syndrome coronavirus RNA:PrThr:Pt:Respiratory.lower:Ord:Probe.amp.tar|Middle east respiratory syndrome coronavirus RNA:PrThr:Pt:Respiratory.lower:Ord:Probe.amp.tar
C5144175|T201|DN|92146-0|LNC|HCoV 229E+NL63 RNA NAA+probe Ql (Resp)|HCoV 229E+NL63 RNA NAA+probe Ql (Resp)
C5144175|T201|OSN|92146-0|LNC|HCoV 229E+NL63 RNA Resp Ql NAA+probe|HCoV 229E+NL63 RNA Resp Ql NAA+probe
C5144175|T201|MTH_LN|92146-0|LNC|Human coronavirus 229E+NL63 ribonucleic acid:Presence or Threshold:Point in time:Respiratory:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus 229E+NL63 ribonucleic acid:Presence or Threshold:Point in time:Respiratory:Ordinal:DNA Nucleic Acid Probe.amp.tar
C5144175|T201|LC|92146-0|LNC|Human coronavirus 229E+NL63 RNA [Presence] in Respiratory specimen by NAA with probe detection|Human coronavirus 229E+NL63 RNA [Presence] in Respiratory specimen by NAA with probe detection
C5144175|T201|LN|92146-0|LNC|Human coronavirus 229E+NL63 RNA:PrThr:Pt:Respiratory:Ord:Probe.amp.tar|Human coronavirus 229E+NL63 RNA:PrThr:Pt:Respiratory:Ord:Probe.amp.tar
C5144176|T201|DN|92147-8|LNC|HCoV HKU1+OC43 RNA NAA+probe Ql (Resp)|HCoV HKU1+OC43 RNA NAA+probe Ql (Resp)
C5144176|T201|OSN|92147-8|LNC|HCoV HKU1+OC43 RNA Resp Ql NAA+probe|HCoV HKU1+OC43 RNA Resp Ql NAA+probe
C5144176|T201|MTH_LN|92147-8|LNC|Human coronavirus HKU1+OC43 ribonucleic acid:Presence or Threshold:Point in time:Respiratory:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus HKU1+OC43 ribonucleic acid:Presence or Threshold:Point in time:Respiratory:Ordinal:DNA Nucleic Acid Probe.amp.tar
C5144176|T201|LC|92147-8|LNC|Human coronavirus HKU1+OC43 RNA [Presence] in Respiratory specimen by NAA with probe detection|Human coronavirus HKU1+OC43 RNA [Presence] in Respiratory specimen by NAA with probe detection
C5144176|T201|LN|92147-8|LNC|Human coronavirus HKU1+OC43 RNA:PrThr:Pt:Respiratory:Ord:Probe.amp.tar|Human coronavirus HKU1+OC43 RNA:PrThr:Pt:Respiratory:Ord:Probe.amp.tar
C5144760|T201|OSN|92876-2|LNC|4 HCoVs + HPIV1-4 RNA Pnl LowResp NAA+Pr|4 HCoVs + HPIV1-4 RNA Pnl LowResp NAA+Pr
C5144760|T201|DN|92876-2|LNC|HCoV 229E+HKU1+NL63+OC43 and Parainfluenza virus 1+2+3+4 RNA panel NAA+probe (Lower resp)|HCoV 229E+HKU1+NL63+OC43 and Parainfluenza virus 1+2+3+4 RNA panel NAA+probe (Lower resp)
C5144760|T201|MTH_LN|92876-2|LNC|Human coronavirus 229E+HKU1+NL63+OC43 & Parainfluenza virus 1+2+3+4 ribonucleic acid panel:-:Point in time:Respiratory.lower:-:DNA Nucleic Acid Probe.amp.tar|Human coronavirus 229E+HKU1+NL63+OC43 & Parainfluenza virus 1+2+3+4 ribonucleic acid panel:-:Point in time:Respiratory.lower:-:DNA Nucleic Acid Probe.amp.tar
C5144760|T201|LN|92876-2|LNC|Human coronavirus 229E+HKU1+NL63+OC43 & Parainfluenza virus 1+2+3+4 RNA panel:-:Pt:Respiratory.lower:-:Probe.amp.tar|Human coronavirus 229E+HKU1+NL63+OC43 & Parainfluenza virus 1+2+3+4 RNA panel:-:Pt:Respiratory.lower:-:Probe.amp.tar
C5144760|T201|LC|92876-2|LNC|Human coronavirus 229E+HKU1+NL63+OC43 and Parainfluenza virus 1+2+3+4 RNA panel - Lower respiratory specimen by NAA with probe detection|Human coronavirus 229E+HKU1+NL63+OC43 and Parainfluenza virus 1+2+3+4 RNA panel - Lower respiratory specimen by NAA with probe detection
C5144761|T201|OSN|92877-0|LNC|4 HCoVs + HPIV1-4 RNA Pnl Up resp NAA+pr|4 HCoVs + HPIV1-4 RNA Pnl Up resp NAA+pr
C5144761|T201|DN|92877-0|LNC|HCoV 229E+HKU1+NL63+OC43 and Parainfluenza virus 1+2+3+4 RNA panel NAA+probe (Upper resp)|HCoV 229E+HKU1+NL63+OC43 and Parainfluenza virus 1+2+3+4 RNA panel NAA+probe (Upper resp)
C5144761|T201|MTH_LN|92877-0|LNC|Human coronavirus 229E+HKU1+NL63+OC43 & Parainfluenza virus 1+2+3+4 ribonucleic acid panel:-:Point in time:Respiratory.upper:-:DNA Nucleic Acid Probe.amp.tar|Human coronavirus 229E+HKU1+NL63+OC43 & Parainfluenza virus 1+2+3+4 ribonucleic acid panel:-:Point in time:Respiratory.upper:-:DNA Nucleic Acid Probe.amp.tar
C5144761|T201|LN|92877-0|LNC|Human coronavirus 229E+HKU1+NL63+OC43 & Parainfluenza virus 1+2+3+4 RNA panel:-:Pt:Respiratory.upper:-:Probe.amp.tar|Human coronavirus 229E+HKU1+NL63+OC43 & Parainfluenza virus 1+2+3+4 RNA panel:-:Pt:Respiratory.upper:-:Probe.amp.tar
C5144761|T201|LC|92877-0|LNC|Human coronavirus 229E+HKU1+NL63+OC43 and Parainfluenza virus 1+2+3+4 RNA panel - Upper respiratory specimen by NAA with probe detection|Human coronavirus 229E+HKU1+NL63+OC43 and Parainfluenza virus 1+2+3+4 RNA panel - Upper respiratory specimen by NAA with probe detection
C5144762|T201|OSN|92878-8|LNC|4 HCoVs RNA Lower resp Ql NAA+probe|4 HCoVs RNA Lower resp Ql NAA+probe
C5144762|T201|DN|92878-8|LNC|HCoV 229E+HKU1+NL63+OC43 RNA NAA+probe Ql (Lower resp)|HCoV 229E+HKU1+NL63+OC43 RNA NAA+probe Ql (Lower resp)
C5144762|T201|MTH_LN|92878-8|LNC|Human coronavirus 229E+HKU1+NL63+OC43 ribonucleic acid:Presence or Threshold:Point in time:Respiratory.lower:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus 229E+HKU1+NL63+OC43 ribonucleic acid:Presence or Threshold:Point in time:Respiratory.lower:Ordinal:DNA Nucleic Acid Probe.amp.tar
C5144762|T201|LC|92878-8|LNC|Human coronavirus 229E+HKU1+NL63+OC43 RNA [Presence] in Lower respiratory specimen by NAA with probe detection|Human coronavirus 229E+HKU1+NL63+OC43 RNA [Presence] in Lower respiratory specimen by NAA with probe detection
C5144762|T201|LN|92878-8|LNC|Human coronavirus 229E+HKU1+NL63+OC43 RNA:PrThr:Pt:Respiratory.lower:Ord:Probe.amp.tar|Human coronavirus 229E+HKU1+NL63+OC43 RNA:PrThr:Pt:Respiratory.lower:Ord:Probe.amp.tar
C5144763|T201|OSN|92879-6|LNC|4 HCoVs RNA Up resp Ql NAA+probe|4 HCoVs RNA Up resp Ql NAA+probe
C5144763|T201|DN|92879-6|LNC|HCoV 229E+HKU1+NL63+OC43 RNA NAA+probe Ql (Upper resp)|HCoV 229E+HKU1+NL63+OC43 RNA NAA+probe Ql (Upper resp)
C5144763|T201|MTH_LN|92879-6|LNC|Human coronavirus 229E+HKU1+NL63+OC43 ribonucleic acid:Presence or Threshold:Point in time:Respiratory.upper:Ordinal:DNA Nucleic Acid Probe.amp.tar|Human coronavirus 229E+HKU1+NL63+OC43 ribonucleic acid:Presence or Threshold:Point in time:Respiratory.upper:Ordinal:DNA Nucleic Acid Probe.amp.tar
C5144763|T201|LC|92879-6|LNC|Human coronavirus 229E+HKU1+NL63+OC43 RNA [Presence] in Upper respiratory specimen by NAA with probe detection|Human coronavirus 229E+HKU1+NL63+OC43 RNA [Presence] in Upper respiratory specimen by NAA with probe detection
C5144763|T201|LN|92879-6|LNC|Human coronavirus 229E+HKU1+NL63+OC43 RNA:PrThr:Pt:Respiratory.upper:Ord:Probe.amp.tar|Human coronavirus 229E+HKU1+NL63+OC43 RNA:PrThr:Pt:Respiratory.upper:Ord:Probe.amp.tar
C5144842|T201|OSN|92967-9|LNC|MERS-CoV RNA Lower Resp Ql NAA+non-probe|MERS-CoV RNA Lower Resp Ql NAA+non-probe
C5144842|T201|DN|92967-9|LNC|MERS-CoV RNA NAA+non-probe Ql (Lower resp)|MERS-CoV RNA NAA+non-probe Ql (Lower resp)
C5144842|T201|LC|92967-9|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Lower respiratory specimen by NAA with non-probe detection|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Lower respiratory specimen by NAA with non-probe detection
C5144842|T201|MTH_LN|92967-9|LNC|Middle East respiratory syndrome coronavirus ribonucleic acid:Presence or Threshold:Point in time:Respiratory.lower:Ordinal:Non-probe.amp.tar|Middle East respiratory syndrome coronavirus ribonucleic acid:Presence or Threshold:Point in time:Respiratory.lower:Ordinal:Non-probe.amp.tar
C5144842|T201|LN|92967-9|LNC|Middle East respiratory syndrome coronavirus RNA:PrThr:Pt:Respiratory.lower:Ord:Non-probe.amp.tar|Middle East respiratory syndrome coronavirus RNA:PrThr:Pt:Respiratory.lower:Ord:Non-probe.amp.tar
C5144854|T201|OSN|92979-4|LNC|HCoV RNA Lower Resp Ql NAA+non-probe|HCoV RNA Lower Resp Ql NAA+non-probe
C5144854|T201|DN|92979-4|LNC|HCoV RNA NAA+non-probe Ql (Lower resp)|HCoV RNA NAA+non-probe Ql (Lower resp)
C5144854|T201|MTH_LN|92979-4|LNC|Human Coronavirus ribonucleic acid:Presence or Threshold:Point in time:Respiratory.lower:Ordinal:Non-probe.amp.tar|Human Coronavirus ribonucleic acid:Presence or Threshold:Point in time:Respiratory.lower:Ordinal:Non-probe.amp.tar
C5144854|T201|LC|92979-4|LNC|Human coronavirus RNA [Presence] in Lower respiratory specimen by NAA with non-probe detection|Human coronavirus RNA [Presence] in Lower respiratory specimen by NAA with non-probe detection
C5144854|T201|LN|92979-4|LNC|Human Coronavirus RNA:PrThr:Pt:Respiratory.lower:Ord:Non-probe.amp.tar|Human Coronavirus RNA:PrThr:Pt:Respiratory.lower:Ord:Non-probe.amp.tar
C5147436|T005|LPN|LP341565-2|LNC|Human coronavirus 229E+NL63|Human coronavirus 229E+NL63
C5147437|T005|LPN|LP341564-5|LNC|Human coronavirus HKU1+OC43|Human coronavirus HKU1+OC43
C5155811|T129|LPN|LP379206-8|LNC|Bovine coronavirus Ag &#x7C; Tissue and Smears &#x7C; Microbiology|Bovine coronavirus Ag &#x7C; Tissue and Smears &#x7C; Microbiology
C5156670|T116|LPN|LP379254-8|LNC|Canine coronavirus Ab &#x7C; Serum &#x7C; Microbiology|Canine coronavirus Ab &#x7C; Serum &#x7C; Microbiology
C5156670|T129|LPN|LP379254-8|LNC|Canine coronavirus Ab &#x7C; Serum &#x7C; Microbiology|Canine coronavirus Ab &#x7C; Serum &#x7C; Microbiology
C5156671|T116|LPN|LP379255-5|LNC|Canine coronavirus Ag &#x7C; Tissue and Smears &#x7C; Microbiology|Canine coronavirus Ag &#x7C; Tissue and Smears &#x7C; Microbiology
C5156671|T129|LPN|LP379255-5|LNC|Canine coronavirus Ag &#x7C; Tissue and Smears &#x7C; Microbiology|Canine coronavirus Ag &#x7C; Tissue and Smears &#x7C; Microbiology
C5160916|T116|LPN|LP377158-3|LNC|Coronavirus Ab &#x7C; Serum &#x7C; Microbiology|Coronavirus Ab &#x7C; Serum &#x7C; Microbiology
C5160916|T129|LPN|LP377158-3|LNC|Coronavirus Ab &#x7C; Serum &#x7C; Microbiology|Coronavirus Ab &#x7C; Serum &#x7C; Microbiology
C5164382|T116|LPN|LP379356-1|LNC|Feline coronavirus Ab &#x7C; Serum &#x7C; Microbiology|Feline coronavirus Ab &#x7C; Serum &#x7C; Microbiology
C5164382|T129|LPN|LP379356-1|LNC|Feline coronavirus Ab &#x7C; Serum &#x7C; Microbiology|Feline coronavirus Ab &#x7C; Serum &#x7C; Microbiology
C5168314|T116|LPN|LP377160-9|LNC|Human coronavirus 229E Ag &#x7C; XXX &#x7C; Microbiology|Human coronavirus 229E Ag &#x7C; XXX &#x7C; Microbiology
C5168314|T129|LPN|LP377160-9|LNC|Human coronavirus 229E Ag &#x7C; XXX &#x7C; Microbiology|Human coronavirus 229E Ag &#x7C; XXX &#x7C; Microbiology
C5168315|T114|LPN|LP377197-1|LNC|Human coronavirus 229E and OC43 RNA &#x7C; Nasopharynx &#x7C; Microbiology|Human coronavirus 229E and OC43 RNA &#x7C; Nasopharynx &#x7C; Microbiology
C5168315|T123|LPN|LP377197-1|LNC|Human coronavirus 229E and OC43 RNA &#x7C; Nasopharynx &#x7C; Microbiology|Human coronavirus 229E and OC43 RNA &#x7C; Nasopharynx &#x7C; Microbiology
C5168316|T116|LPN|LP377159-1|LNC|Human coronavirus 229E IgG &#x7C; Serum &#x7C; Microbiology|Human coronavirus 229E IgG &#x7C; Serum &#x7C; Microbiology
C5168316|T129|LPN|LP377159-1|LNC|Human coronavirus 229E IgG &#x7C; Serum &#x7C; Microbiology|Human coronavirus 229E IgG &#x7C; Serum &#x7C; Microbiology
C5168317|T114|LPN|LP377161-7|LNC|Human coronavirus 229E RNA &#x7C; Aspirate &#x7C; Microbiology|Human coronavirus 229E RNA &#x7C; Aspirate &#x7C; Microbiology
C5168318|T114|LPN|LP377162-5|LNC|Human coronavirus 229E RNA &#x7C; Cornea or Conjunctiva &#x7C; Microbiology|Human coronavirus 229E RNA &#x7C; Cornea or Conjunctiva &#x7C; Microbiology
C5168319|T114|LPN|LP377164-1|LNC|Human coronavirus 229E RNA &#x7C; Lower respiratory specimen &#x7C; Microbiology|Human coronavirus 229E RNA &#x7C; Lower respiratory specimen &#x7C; Microbiology
C5168320|T114|LPN|LP377163-3|LNC|Human coronavirus 229E RNA &#x7C; Nasopharynx &#x7C; Microbiology|Human coronavirus 229E RNA &#x7C; Nasopharynx &#x7C; Microbiology
C5168321|T114|LPN|LP377165-8|LNC|Human coronavirus 229E RNA &#x7C; Upper respiratory specimen &#x7C; Microbiology|Human coronavirus 229E RNA &#x7C; Upper respiratory specimen &#x7C; Microbiology
C5168322|T114|LPN|LP377166-6|LNC|Human coronavirus 229E RNA &#x7C; XXX &#x7C; Microbiology|Human coronavirus 229E RNA &#x7C; XXX &#x7C; Microbiology
C5168323|T114|LPN|LP377199-7|LNC|Human coronavirus 229E+HKU1+NL63+OC43 RNA &#x7C; Lower respiratory specimen &#x7C; Microbiology|Human coronavirus 229E+HKU1+NL63+OC43 RNA &#x7C; Lower respiratory specimen &#x7C; Microbiology
C5168324|T114|LPN|LP377198-9|LNC|Human coronavirus 229E+HKU1+NL63+OC43 RNA &#x7C; Nasopharynx &#x7C; Microbiology|Human coronavirus 229E+HKU1+NL63+OC43 RNA &#x7C; Nasopharynx &#x7C; Microbiology
C5168325|T114|LPN|LP377200-3|LNC|Human coronavirus 229E+HKU1+NL63+OC43 RNA &#x7C; Upper respiratory specimen &#x7C; Microbiology|Human coronavirus 229E+HKU1+NL63+OC43 RNA &#x7C; Upper respiratory specimen &#x7C; Microbiology
C5168326|T114|LPN|LP377196-3|LNC|Human coronavirus 229E+NL63 RNA &#x7C; Respiratory specimen &#x7C; Microbiology|Human coronavirus 229E+NL63 RNA &#x7C; Respiratory specimen &#x7C; Microbiology
C5168327|T116|LPN|LP377167-4|LNC|Human coronavirus Ag &#x7C; XXX &#x7C; Microbiology|Human coronavirus Ag &#x7C; XXX &#x7C; Microbiology
C5168327|T129|LPN|LP377167-4|LNC|Human coronavirus Ag &#x7C; XXX &#x7C; Microbiology|Human coronavirus Ag &#x7C; XXX &#x7C; Microbiology
C5168328|T114|LPN|LP377169-0|LNC|Human coronavirus HKU1 RNA &#x7C; Aspirate &#x7C; Microbiology|Human coronavirus HKU1 RNA &#x7C; Aspirate &#x7C; Microbiology
C5168329|T114|LPN|LP377170-8|LNC|Human coronavirus HKU1 RNA &#x7C; Cornea or Conjunctiva &#x7C; Microbiology|Human coronavirus HKU1 RNA &#x7C; Cornea or Conjunctiva &#x7C; Microbiology
C5168330|T114|LPN|LP377172-4|LNC|Human coronavirus HKU1 RNA &#x7C; Lower respiratory specimen &#x7C; Microbiology|Human coronavirus HKU1 RNA &#x7C; Lower respiratory specimen &#x7C; Microbiology
C5168331|T114|LPN|LP377171-6|LNC|Human coronavirus HKU1 RNA &#x7C; Nasopharynx &#x7C; Microbiology|Human coronavirus HKU1 RNA &#x7C; Nasopharynx &#x7C; Microbiology
C5168332|T114|LPN|LP377173-2|LNC|Human coronavirus HKU1 RNA &#x7C; Upper respiratory specimen &#x7C; Microbiology|Human coronavirus HKU1 RNA &#x7C; Upper respiratory specimen &#x7C; Microbiology
C5168333|T114|LPN|LP377174-0|LNC|Human coronavirus HKU1 RNA &#x7C; XXX &#x7C; Microbiology|Human coronavirus HKU1 RNA &#x7C; XXX &#x7C; Microbiology
C5168334|T114|LPN|LP377201-1|LNC|Human coronavirus HKU1+OC43 RNA &#x7C; Respiratory specimen &#x7C; Microbiology|Human coronavirus HKU1+OC43 RNA &#x7C; Respiratory specimen &#x7C; Microbiology
C5168335|T034|LPN|LP377168-2|LNC|Human coronavirus identified &#x7C; XXX &#x7C; Microbiology|Human coronavirus identified &#x7C; XXX &#x7C; Microbiology
C5168336|T116|LPN|LP377175-7|LNC|Human coronavirus NL63 IgG &#x7C; Serum &#x7C; Microbiology|Human coronavirus NL63 IgG &#x7C; Serum &#x7C; Microbiology
C5168336|T129|LPN|LP377175-7|LNC|Human coronavirus NL63 IgG &#x7C; Serum &#x7C; Microbiology|Human coronavirus NL63 IgG &#x7C; Serum &#x7C; Microbiology
C5168337|T114|LPN|LP377176-5|LNC|Human coronavirus NL63 RNA &#x7C; Aspirate &#x7C; Microbiology|Human coronavirus NL63 RNA &#x7C; Aspirate &#x7C; Microbiology
C5168338|T114|LPN|LP377177-3|LNC|Human coronavirus NL63 RNA &#x7C; Cornea or Conjunctiva &#x7C; Microbiology|Human coronavirus NL63 RNA &#x7C; Cornea or Conjunctiva &#x7C; Microbiology
C5168339|T114|LPN|LP377179-9|LNC|Human coronavirus NL63 RNA &#x7C; Lower respiratory specimen &#x7C; Microbiology|Human coronavirus NL63 RNA &#x7C; Lower respiratory specimen &#x7C; Microbiology
C5168340|T114|LPN|LP377178-1|LNC|Human coronavirus NL63 RNA &#x7C; Nasopharynx &#x7C; Microbiology|Human coronavirus NL63 RNA &#x7C; Nasopharynx &#x7C; Microbiology
C5168341|T114|LPN|LP377180-7|LNC|Human coronavirus NL63 RNA &#x7C; Upper respiratory specimen &#x7C; Microbiology|Human coronavirus NL63 RNA &#x7C; Upper respiratory specimen &#x7C; Microbiology
C5168342|T114|LPN|LP377181-5|LNC|Human coronavirus NL63 RNA &#x7C; XXX &#x7C; Microbiology|Human coronavirus NL63 RNA &#x7C; XXX &#x7C; Microbiology
C5168343|T116|LPN|LP377183-1|LNC|Human coronavirus OC43 Ag &#x7C; XXX &#x7C; Microbiology|Human coronavirus OC43 Ag &#x7C; XXX &#x7C; Microbiology
C5168343|T129|LPN|LP377183-1|LNC|Human coronavirus OC43 Ag &#x7C; XXX &#x7C; Microbiology|Human coronavirus OC43 Ag &#x7C; XXX &#x7C; Microbiology
C5168344|T116|LPN|LP377182-3|LNC|Human coronavirus OC43 IgG &#x7C; Serum &#x7C; Microbiology|Human coronavirus OC43 IgG &#x7C; Serum &#x7C; Microbiology
C5168344|T129|LPN|LP377182-3|LNC|Human coronavirus OC43 IgG &#x7C; Serum &#x7C; Microbiology|Human coronavirus OC43 IgG &#x7C; Serum &#x7C; Microbiology
C5168345|T114|LPN|LP377184-9|LNC|Human coronavirus OC43 RNA &#x7C; Aspirate &#x7C; Microbiology|Human coronavirus OC43 RNA &#x7C; Aspirate &#x7C; Microbiology
C5168346|T114|LPN|LP377185-6|LNC|Human coronavirus OC43 RNA &#x7C; Cornea or Conjunctiva &#x7C; Microbiology|Human coronavirus OC43 RNA &#x7C; Cornea or Conjunctiva &#x7C; Microbiology
C5168347|T114|LPN|LP377187-2|LNC|Human coronavirus OC43 RNA &#x7C; Lower respiratory specimen &#x7C; Microbiology|Human coronavirus OC43 RNA &#x7C; Lower respiratory specimen &#x7C; Microbiology
C5168348|T114|LPN|LP377186-4|LNC|Human coronavirus OC43 RNA &#x7C; Nasopharynx &#x7C; Microbiology|Human coronavirus OC43 RNA &#x7C; Nasopharynx &#x7C; Microbiology
C5168349|T114|LPN|LP377188-0|LNC|Human coronavirus OC43 RNA &#x7C; Upper respiratory specimen &#x7C; Microbiology|Human coronavirus OC43 RNA &#x7C; Upper respiratory specimen &#x7C; Microbiology
C5168350|T114|LPN|LP377189-8|LNC|Human coronavirus OC43 RNA &#x7C; XXX &#x7C; Microbiology|Human coronavirus OC43 RNA &#x7C; XXX &#x7C; Microbiology
C5168351|T114|LPN|LP377190-6|LNC|Human coronavirus RNA &#x7C; Aspirate &#x7C; Microbiology|Human coronavirus RNA &#x7C; Aspirate &#x7C; Microbiology
C5168351|T123|LPN|LP377190-6|LNC|Human coronavirus RNA &#x7C; Aspirate &#x7C; Microbiology|Human coronavirus RNA &#x7C; Aspirate &#x7C; Microbiology
C5168352|T114|LPN|LP377191-4|LNC|Human coronavirus RNA &#x7C; Cornea or Conjunctiva &#x7C; Microbiology|Human coronavirus RNA &#x7C; Cornea or Conjunctiva &#x7C; Microbiology
C5168352|T123|LPN|LP377191-4|LNC|Human coronavirus RNA &#x7C; Cornea or Conjunctiva &#x7C; Microbiology|Human coronavirus RNA &#x7C; Cornea or Conjunctiva &#x7C; Microbiology
C5168353|T114|LPN|LP377192-2|LNC|Human coronavirus RNA &#x7C; Lower respiratory specimen &#x7C; Microbiology|Human coronavirus RNA &#x7C; Lower respiratory specimen &#x7C; Microbiology
C5168353|T123|LPN|LP377192-2|LNC|Human coronavirus RNA &#x7C; Lower respiratory specimen &#x7C; Microbiology|Human coronavirus RNA &#x7C; Lower respiratory specimen &#x7C; Microbiology
C5168354|T114|LPN|LP377194-8|LNC|Human coronavirus RNA &#x7C; Serum or Plasma &#x7C; Microbiology|Human coronavirus RNA &#x7C; Serum or Plasma &#x7C; Microbiology
C5168354|T123|LPN|LP377194-8|LNC|Human coronavirus RNA &#x7C; Serum or Plasma &#x7C; Microbiology|Human coronavirus RNA &#x7C; Serum or Plasma &#x7C; Microbiology
C5168355|T114|LPN|LP377193-0|LNC|Human coronavirus RNA &#x7C; Upper respiratory specimen &#x7C; Microbiology|Human coronavirus RNA &#x7C; Upper respiratory specimen &#x7C; Microbiology
C5168355|T123|LPN|LP377193-0|LNC|Human coronavirus RNA &#x7C; Upper respiratory specimen &#x7C; Microbiology|Human coronavirus RNA &#x7C; Upper respiratory specimen &#x7C; Microbiology
C5168356|T114|LPN|LP377195-5|LNC|Human coronavirus RNA &#x7C; XXX &#x7C; Microbiology|Human coronavirus RNA &#x7C; XXX &#x7C; Microbiology
C5168356|T123|LPN|LP377195-5|LNC|Human coronavirus RNA &#x7C; XXX &#x7C; Microbiology|Human coronavirus RNA &#x7C; XXX &#x7C; Microbiology
C5168357|T059|LPN|LP380015-0|LNC|Human coronavirus RNA panel &#x7C; XXX &#x7C; Microbiology Panels|Human coronavirus RNA panel &#x7C; XXX &#x7C; Microbiology Panels
C5173236|T114|LPN|LP377211-0|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) N2 gene RNA &#x7C; XXX &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) N2 gene RNA &#x7C; XXX &#x7C; Microbiology
C5173236|T123|LPN|LP377211-0|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) N2 gene RNA &#x7C; XXX &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) N2 gene RNA &#x7C; XXX &#x7C; Microbiology
C5173237|T114|LPN|LP377212-8|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) N3 gene RNA &#x7C; XXX &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) N3 gene RNA &#x7C; XXX &#x7C; Microbiology
C5173237|T123|LPN|LP377212-8|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) N3 gene RNA &#x7C; XXX &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) N3 gene RNA &#x7C; XXX &#x7C; Microbiology
C5173238|T114|LPN|LP377202-9|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Aspirate &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Aspirate &#x7C; Microbiology
C5173238|T123|LPN|LP377202-9|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Aspirate &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Aspirate &#x7C; Microbiology
C5173239|T114|LPN|LP377203-7|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Blood &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Blood &#x7C; Microbiology
C5173239|T123|LPN|LP377203-7|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Blood &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Blood &#x7C; Microbiology
C5173240|T114|LPN|LP377204-5|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Cornea or Conjunctiva &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Cornea or Conjunctiva &#x7C; Microbiology
C5173240|T123|LPN|LP377204-5|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Cornea or Conjunctiva &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Cornea or Conjunctiva &#x7C; Microbiology
C5173241|T114|LPN|LP377206-0|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Lower respiratory specimen &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Lower respiratory specimen &#x7C; Microbiology
C5173241|T123|LPN|LP377206-0|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Lower respiratory specimen &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Lower respiratory specimen &#x7C; Microbiology
C5173242|T114|LPN|LP377205-2|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Nasopharynx &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Nasopharynx &#x7C; Microbiology
C5173242|T123|LPN|LP377205-2|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Nasopharynx &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Nasopharynx &#x7C; Microbiology
C5173243|T114|LPN|LP377208-6|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Stool &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Stool &#x7C; Microbiology
C5173243|T123|LPN|LP377208-6|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Stool &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Stool &#x7C; Microbiology
C5173244|T114|LPN|LP377207-8|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Upper respiratory specimen &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Upper respiratory specimen &#x7C; Microbiology
C5173244|T123|LPN|LP377207-8|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Upper respiratory specimen &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Upper respiratory specimen &#x7C; Microbiology
C5173245|T114|LPN|LP377209-4|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Urine &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Urine &#x7C; Microbiology
C5173245|T123|LPN|LP377209-4|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Urine &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; Urine &#x7C; Microbiology
C5173246|T114|LPN|LP377210-2|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; XXX &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; XXX &#x7C; Microbiology
C5173246|T123|LPN|LP377210-2|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; XXX &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA &#x7C; XXX &#x7C; Microbiology
C5173247|T059|LPN|LP380060-6|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA panel &#x7C; XXX &#x7C; Microbiology Panels|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA panel &#x7C; XXX &#x7C; Microbiology Panels
C5173248|T114|LPN|LP377213-6|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) upE gene RNA &#x7C; XXX &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) upE gene RNA &#x7C; XXX &#x7C; Microbiology
C5173248|T123|LPN|LP377213-6|LNC|Middle East respiratory syndrome coronavirus (MERS-CoV) upE gene RNA &#x7C; XXX &#x7C; Microbiology|Middle East respiratory syndrome coronavirus (MERS-CoV) upE gene RNA &#x7C; XXX &#x7C; Microbiology
C5177858|T005|LPN|LP379476-7|LNC|Porcine deltacoronavirus &#x7C; XXX &#x7C; Microbiology|Porcine deltacoronavirus &#x7C; XXX &#x7C; Microbiology
C5177859|T081|LPN|LP379478-3|LNC|Porcine deltacoronavirus Ab.IgG/Positive control &#x7C; XXX &#x7C; Microbiology|Porcine deltacoronavirus Ab.IgG/Positive control &#x7C; XXX &#x7C; Microbiology
C5177860|T116|LPN|LP379479-1|LNC|Porcine deltacoronavirus Ag &#x7C; Tissue and Smears &#x7C; Microbiology|Porcine deltacoronavirus Ag &#x7C; Tissue and Smears &#x7C; Microbiology
C5177860|T129|LPN|LP379479-1|LNC|Porcine deltacoronavirus Ag &#x7C; Tissue and Smears &#x7C; Microbiology|Porcine deltacoronavirus Ag &#x7C; Tissue and Smears &#x7C; Microbiology
C5177861|T114|LPN|LP379477-5|LNC|Porcine deltacoronavirus RNA &#x7C; XXX &#x7C; Microbiology|Porcine deltacoronavirus RNA &#x7C; XXX &#x7C; Microbiology
C5177861|T123|LPN|LP379477-5|LNC|Porcine deltacoronavirus RNA &#x7C; XXX &#x7C; Microbiology|Porcine deltacoronavirus RNA &#x7C; XXX &#x7C; Microbiology
C5177897|T116|LPN|LP379537-6|LNC|Porcine respiratory coronavirus Ab &#x7C; Serum &#x7C; Microbiology|Porcine respiratory coronavirus Ab &#x7C; Serum &#x7C; Microbiology
C5177897|T129|LPN|LP379537-6|LNC|Porcine respiratory coronavirus Ab &#x7C; Serum &#x7C; Microbiology|Porcine respiratory coronavirus Ab &#x7C; Serum &#x7C; Microbiology
C5177898|T081|LPN|LP379541-8|LNC|Porcine respiratory coronavirus Ab/Negative control &#x7C; Serum &#x7C; Microbiology|Porcine respiratory coronavirus Ab/Negative control &#x7C; Serum &#x7C; Microbiology
C5177899|T116|LPN|LP379538-4|LNC|Porcine respiratory coronavirus Ag &#x7C; Small intestine Tissue &#x7C; Microbiology|Porcine respiratory coronavirus Ag &#x7C; Small intestine Tissue &#x7C; Microbiology
C5177899|T129|LPN|LP379538-4|LNC|Porcine respiratory coronavirus Ag &#x7C; Small intestine Tissue &#x7C; Microbiology|Porcine respiratory coronavirus Ag &#x7C; Small intestine Tissue &#x7C; Microbiology
C5177900|T116|LPN|LP379539-2|LNC|Porcine respiratory coronavirus Ag &#x7C; XXX &#x7C; Microbiology|Porcine respiratory coronavirus Ag &#x7C; XXX &#x7C; Microbiology
C5177900|T129|LPN|LP379539-2|LNC|Porcine respiratory coronavirus Ag &#x7C; XXX &#x7C; Microbiology|Porcine respiratory coronavirus Ag &#x7C; XXX &#x7C; Microbiology
C5177901|T114|LPN|LP379540-0|LNC|Porcine respiratory coronavirus RNA &#x7C; XXX &#x7C; Microbiology|Porcine respiratory coronavirus RNA &#x7C; XXX &#x7C; Microbiology
C5180353|T005|LPN|LP377214-4|LNC|SARS coronavirus &#x7C; XXX &#x7C; Microbiology|SARS coronavirus &#x7C; XXX &#x7C; Microbiology
C5180354|T116|LPN|LP377215-1|LNC|SARS coronavirus Ab &#x7C; Serum &#x7C; Microbiology|SARS coronavirus Ab &#x7C; Serum &#x7C; Microbiology
C5180354|T129|LPN|LP377215-1|LNC|SARS coronavirus Ab &#x7C; Serum &#x7C; Microbiology|SARS coronavirus Ab &#x7C; Serum &#x7C; Microbiology
C5180355|T116|LPN|LP377216-9|LNC|SARS Coronavirus IgG &#x7C; Serum &#x7C; Microbiology|SARS Coronavirus IgG &#x7C; Serum &#x7C; Microbiology
C5180355|T129|LPN|LP377216-9|LNC|SARS Coronavirus IgG &#x7C; Serum &#x7C; Microbiology|SARS Coronavirus IgG &#x7C; Serum &#x7C; Microbiology
C5180356|T116|LPN|LP377217-7|LNC|SARS Coronavirus IgM &#x7C; Serum &#x7C; Microbiology|SARS Coronavirus IgM &#x7C; Serum &#x7C; Microbiology
C5180356|T129|LPN|LP377217-7|LNC|SARS Coronavirus IgM &#x7C; Serum &#x7C; Microbiology|SARS Coronavirus IgM &#x7C; Serum &#x7C; Microbiology
C5180357|T114|LPN|LP377218-5|LNC|SARS coronavirus RNA &#x7C; Isolate &#x7C; Microbiology|SARS coronavirus RNA &#x7C; Isolate &#x7C; Microbiology
C5180358|T114|LPN|LP377219-3|LNC|SARS coronavirus RNA &#x7C; Serum or Plasma &#x7C; Microbiology|SARS coronavirus RNA &#x7C; Serum or Plasma &#x7C; Microbiology
C5180359|T114|LPN|LP377220-1|LNC|SARS coronavirus RNA &#x7C; XXX &#x7C; Microbiology|SARS coronavirus RNA &#x7C; XXX &#x7C; Microbiology
C5180360|T116|LPN|LP377221-9|LNC|SARS coronavirus Urbani Ab &#x7C; Serum &#x7C; Microbiology|SARS coronavirus Urbani Ab &#x7C; Serum &#x7C; Microbiology
C5180360|T129|LPN|LP377221-9|LNC|SARS coronavirus Urbani Ab &#x7C; Serum &#x7C; Microbiology|SARS coronavirus Urbani Ab &#x7C; Serum &#x7C; Microbiology
C5180361|T114|LPN|LP377222-7|LNC|SARS coronavirus Urbani RNA &#x7C; Nose &#x7C; Microbiology|SARS coronavirus Urbani RNA &#x7C; Nose &#x7C; Microbiology
C5180361|T123|LPN|LP377222-7|LNC|SARS coronavirus Urbani RNA &#x7C; Nose &#x7C; Microbiology|SARS coronavirus Urbani RNA &#x7C; Nose &#x7C; Microbiology
C5180362|T114|LPN|LP377223-5|LNC|SARS coronavirus Urbani RNA &#x7C; Serum or Plasma &#x7C; Microbiology|SARS coronavirus Urbani RNA &#x7C; Serum or Plasma &#x7C; Microbiology
C5180362|T123|LPN|LP377223-5|LNC|SARS coronavirus Urbani RNA &#x7C; Serum or Plasma &#x7C; Microbiology|SARS coronavirus Urbani RNA &#x7C; Serum or Plasma &#x7C; Microbiology
C5180363|T114|LPN|LP377224-3|LNC|SARS coronavirus Urbani RNA &#x7C; Sputum &#x7C; Microbiology|SARS coronavirus Urbani RNA &#x7C; Sputum &#x7C; Microbiology
C5180363|T123|LPN|LP377224-3|LNC|SARS coronavirus Urbani RNA &#x7C; Sputum &#x7C; Microbiology|SARS coronavirus Urbani RNA &#x7C; Sputum &#x7C; Microbiology
C5180364|T114|LPN|LP377225-0|LNC|SARS coronavirus Urbani RNA &#x7C; Stool &#x7C; Microbiology|SARS coronavirus Urbani RNA &#x7C; Stool &#x7C; Microbiology
C5180364|T123|LPN|LP377225-0|LNC|SARS coronavirus Urbani RNA &#x7C; Stool &#x7C; Microbiology|SARS coronavirus Urbani RNA &#x7C; Stool &#x7C; Microbiology
C5180365|T114|LPN|LP377226-8|LNC|SARS coronavirus Urbani RNA &#x7C; XXX &#x7C; Microbiology|SARS coronavirus Urbani RNA &#x7C; XXX &#x7C; Microbiology
C5180365|T123|LPN|LP377226-8|LNC|SARS coronavirus Urbani RNA &#x7C; XXX &#x7C; Microbiology|SARS coronavirus Urbani RNA &#x7C; XXX &#x7C; Microbiology
C5184304|T005|LPN|LP379594-7|LNC|Turkey enteritis coronavirus &#x7C; Serum &#x7C; Microbiology|Turkey enteritis coronavirus &#x7C; Serum &#x7C; Microbiology
C5203670|T047|PN|NOCODE|MTH|COVID-19|COVID-19
C5203670|T047|SY|840539006|SNOMEDCT_US|Disease caused by 2019 novel coronavirus|Disease caused by 2019 novel coronavirus
C5203670|T047|FN|840539006|SNOMEDCT_US|Disease caused by 2019 novel coronavirus (disorder)|Disease caused by 2019 novel coronavirus (disorder)
C5203670|T047|PT|840539006|SNOMEDCT_US|Disease caused by 2019-nCoV|Disease caused by 2019-nCoV
C5203670|T047|SY|840539006|SNOMEDCT_US|Disease caused by Wuhan coronavirus|Disease caused by Wuhan coronavirus
C5203671|T033|PN|NOCODE|MTH|Suspected COVID-19|Suspected COVID-19
C5203671|T033|SY|840544004|SNOMEDCT_US|Suspected disease caused by 2019 novel coronavirus|Suspected disease caused by 2019 novel coronavirus
C5203671|T033|FN|840544004|SNOMEDCT_US|Suspected disease caused by 2019 novel coronavirus (situation)|Suspected disease caused by 2019 novel coronavirus (situation)
C5203671|T033|PT|840544004|SNOMEDCT_US|Suspected disease caused by 2019-nCoV|Suspected disease caused by 2019-nCoV
C5203671|T033|SY|840544004|SNOMEDCT_US|Suspected disease caused by Wuhan coronavirus|Suspected disease caused by Wuhan coronavirus
C5203672|T061|SY|840534001|SNOMEDCT_US|2019 novel coronavirus vaccination|2019 novel coronavirus vaccination
C5203672|T061|FN|840534001|SNOMEDCT_US|2019 novel coronavirus vaccination (procedure)|2019 novel coronavirus vaccination (procedure)
C5203672|T061|PT|840534001|SNOMEDCT_US|2019-nCoV vaccination|2019-nCoV vaccination
C5203672|T061|PN|NOCODE|MTH|SARS-CoV-2 vaccination|SARS-CoV-2 vaccination
C5203672|T061|SY|840534001|SNOMEDCT_US|Wuhan coronavirus vaccination|Wuhan coronavirus vaccination
C5203673|T116|SY|840536004|SNOMEDCT_US|Antigen of 2019 novel coronavirus|Antigen of 2019 novel coronavirus
C5203673|T129|SY|840536004|SNOMEDCT_US|Antigen of 2019 novel coronavirus|Antigen of 2019 novel coronavirus
C5203673|T116|FN|840536004|SNOMEDCT_US|Antigen of 2019 novel coronavirus (substance)|Antigen of 2019 novel coronavirus (substance)
C5203673|T129|FN|840536004|SNOMEDCT_US|Antigen of 2019 novel coronavirus (substance)|Antigen of 2019 novel coronavirus (substance)
C5203673|T116|PT|840536004|SNOMEDCT_US|Antigen of 2019-nCoV|Antigen of 2019-nCoV
C5203673|T129|PT|840536004|SNOMEDCT_US|Antigen of 2019-nCoV|Antigen of 2019-nCoV
C5203673|T116|PN|NOCODE|MTH|Antigen of SARS-CoV-2|Antigen of SARS-CoV-2
C5203673|T129|PN|NOCODE|MTH|Antigen of SARS-CoV-2|Antigen of SARS-CoV-2
C5203673|T116|SY|840536004|SNOMEDCT_US|Antigen of Wuhan coronavirus|Antigen of Wuhan coronavirus
C5203673|T129|SY|840536004|SNOMEDCT_US|Antigen of Wuhan coronavirus|Antigen of Wuhan coronavirus
C5203674|T116|SY|840535000|SNOMEDCT_US|Antibody to 2019 novel coronavirus|Antibody to 2019 novel coronavirus
C5203674|T129|SY|840535000|SNOMEDCT_US|Antibody to 2019 novel coronavirus|Antibody to 2019 novel coronavirus
C5203674|T116|FN|840535000|SNOMEDCT_US|Antibody to 2019 novel coronavirus (substance)|Antibody to 2019 novel coronavirus (substance)
C5203674|T129|FN|840535000|SNOMEDCT_US|Antibody to 2019 novel coronavirus (substance)|Antibody to 2019 novel coronavirus (substance)
C5203674|T116|PT|840535000|SNOMEDCT_US|Antibody to 2019-nCoV|Antibody to 2019-nCoV
C5203674|T129|PT|840535000|SNOMEDCT_US|Antibody to 2019-nCoV|Antibody to 2019-nCoV
C5203674|T116|PN|NOCODE|MTH|Antibody to SARS-CoV-2|Antibody to SARS-CoV-2
C5203674|T129|PN|NOCODE|MTH|Antibody to SARS-CoV-2|Antibody to SARS-CoV-2
C5203674|T116|SY|840535000|SNOMEDCT_US|Antibody to Wuhan coronavirus|Antibody to Wuhan coronavirus
C5203674|T129|SY|840535000|SNOMEDCT_US|Antibody to Wuhan coronavirus|Antibody to Wuhan coronavirus
C5203675|T033|PT|840546002|SNOMEDCT_US|Exposure to 2019 novel coronavirus|Exposure to 2019 novel coronavirus
C5203675|T033|FN|840546002|SNOMEDCT_US|Exposure to 2019 novel coronavirus (event)|Exposure to 2019 novel coronavirus (event)
C5203675|T033|SY|840546002|SNOMEDCT_US|Exposure to 2019-nCoV|Exposure to 2019-nCoV
C5203675|T033|PN|NOCODE|MTH|Exposure to SARS-CoV-2|Exposure to SARS-CoV-2
C5203675|T033|SY|840546002|SNOMEDCT_US|Exposure to Wuhan coronavirus|Exposure to Wuhan coronavirus
C5203676|T005|SY|840533007|SNOMEDCT_US|2019 novel coronavirus|2019 novel coronavirus
C5203676|T005|FN|840533007|SNOMEDCT_US|2019 novel coronavirus (organism)|2019 novel coronavirus (organism)
C5203676|T005|PT|840533007|SNOMEDCT_US|2019-nCoV|2019-nCoV
C5203676|T005|PN|NOCODE|MTH|SARS-CoV-2|SARS-CoV-2
C5203676|T005|SY|840533007|SNOMEDCT_US|Wuhan coronavirus|Wuhan coronavirus
C5213519|T059|LPN|LP417136-1|LNC|Human coronavirus 229E+HKU1+NL63+OC43 and Parainfluenza virus 1+2+3+4 RNA panel &#x7C; Lower respiratory specimen &#x7C; Microbiology Panels|Human coronavirus 229E+HKU1+NL63+OC43 and Parainfluenza virus 1+2+3+4 RNA panel &#x7C; Lower respiratory specimen &#x7C; Microbiology Panels
C5213520|T059|LPN|LP417137-9|LNC|Human coronavirus 229E+HKU1+NL63+OC43 and Parainfluenza virus 1+2+3+4 RNA panel &#x7C; Upper respiratory specimen &#x7C; Microbiology Panels|Human coronavirus 229E+HKU1+NL63+OC43 and Parainfluenza virus 1+2+3+4 RNA panel &#x7C; Upper respiratory specimen &#x7C; Microbiology Panels
C5218549|T114|LG|LG34137-6|LNC|Human coronavirus 229E RNA&#x7C;PrThr&#x7C;Sys:ANYResp|Human coronavirus 229E RNA&#x7C;PrThr&#x7C;Sys:ANYResp
C5218550|T114|LG|LG50873-5|LNC|Human coronavirus 229E+HKU1+NL63+OC43 RNA&#x7C;PrThr&#x7C;Sys:ANYResp|Human coronavirus 229E+HKU1+NL63+OC43 RNA&#x7C;PrThr&#x7C;Sys:ANYResp
C5218551|T114|LG|LG34135-0|LNC|Human coronavirus HKU1 RNA&#x7C;PrThr&#x7C;Sys:ANYResp|Human coronavirus HKU1 RNA&#x7C;PrThr&#x7C;Sys:ANYResp
C5218552|T114|LG|LG34136-8|LNC|Human coronavirus NL63 RNA&#x7C;PrThr&#x7C;Sys:ANYResp|Human coronavirus NL63 RNA&#x7C;PrThr&#x7C;Sys:ANYResp
C5218553|T114|LG|LG34138-4|LNC|Human coronavirus OC43 RNA&#x7C;PrThr&#x7C;Sys:ANYResp|Human coronavirus OC43 RNA&#x7C;PrThr&#x7C;Sys:ANYResp
C5218554|T114|LG|LG41760-6|LNC|Human coronavirus RNA&#x7C;PrThr&#x7C;Sys:ANYResp|Human coronavirus RNA&#x7C;PrThr&#x7C;Sys:ANYResp
C5218582|T114|LG|LG50060-9|LNC|Middle East respiratory syndrome coronavirus RNA&#x7C;PrThr&#x7C;Sys:ANYResp|Middle East respiratory syndrome coronavirus RNA&#x7C;PrThr&#x7C;Sys:ANYResp
C5218582|T123|LG|LG50060-9|LNC|Middle East respiratory syndrome coronavirus RNA&#x7C;PrThr&#x7C;Sys:ANYResp|Middle East respiratory syndrome coronavirus RNA&#x7C;PrThr&#x7C;Sys:ANYResp
C5218621|T114|LG|LG34001-4|LNC|SARS coronavirus Urbani RNA&#x7C;PrThr&#x7C;Sys:ANYResp|SARS coronavirus Urbani RNA&#x7C;PrThr&#x7C;Sys:ANYResp
C5225060|T059|PT|393049|MEDCIN|NAA with probe detection for human coronavirus 229E + OC43 RNA|NAA with probe detection for human coronavirus 229E + OC43 RNA
C5225060|T059|FN|393049|MEDCIN|NAA with probe detection for human coronavirus 229E + OC43 RNA (lab test)|NAA with probe detection for human coronavirus 229E + OC43 RNA (lab test)
C5225060|T059|SY|393049|MEDCIN|NAA with probe detection human coronavirus RNA 229E + OC43 RNA|NAA with probe detection human coronavirus RNA 229E + OC43 RNA
C5225061|T059|PT|393050|MEDCIN|NAA with probe detection for human coronavirus 229E + OC43 RNA in nasopharynx|NAA with probe detection for human coronavirus 229E + OC43 RNA in nasopharynx
C5225061|T059|FN|393050|MEDCIN|NAA with probe detection for human coronavirus 229E + OC43 RNA in nasopharynx (lab test)|NAA with probe detection for human coronavirus 229E + OC43 RNA in nasopharynx (lab test)
C5225061|T059|SY|393050|MEDCIN|NAA with probe detection human coronavirus 229E + OC43 RNA in nasopharynx|NAA with probe detection human coronavirus 229E + OC43 RNA in nasopharynx
C5225062|T059|PT|393048|MEDCIN|NAA with probe detection for human coronavirus RNA|NAA with probe detection for human coronavirus RNA
C5225062|T059|FN|393048|MEDCIN|NAA with probe detection for human coronavirus RNA (lab test)|NAA with probe detection for human coronavirus RNA (lab test)
C5225062|T059|SY|393048|MEDCIN|NAA with probe detection human coronavirus RNA|NAA with probe detection human coronavirus RNA
C5234677|T201|LC|94531-1|LNC_SPECIAL_USE|SARS Coronavirus 2 RNA panel - Respiratory specimen by NAA with probe detection|SARS Coronavirus 2 RNA panel - Respiratory specimen by NAA with probe detection
C5234677|T201|LN|94531-1|LNC_SPECIAL_USE|SARS coronavirus 2 RNA panel:-:Pt:Respiratory:-:Probe.amp.tar|SARS coronavirus 2 RNA panel:-:Pt:Respiratory:-:Probe.amp.tar
C5234677|T201|OSN|94531-1|LNC_SPECIAL_USE|SARS-CoV-2 RNA Pnl Resp NAA+probe|SARS-CoV-2 RNA Pnl Resp NAA+probe
C5234678|T201|LC|94532-9|LNC_SPECIAL_USE|SARS coronavirus+SARS-like coronavirus+SARS coronavirus 2+MERS coronavirus RNA [Presence] in Respiratory specimen by NAA with probe detection|SARS coronavirus+SARS-like coronavirus+SARS coronavirus 2+MERS coronavirus RNA [Presence] in Respiratory specimen by NAA with probe detection
C5234678|T201|LN|94532-9|LNC_SPECIAL_USE|SARS coronavirus+SARS-like coronavirus+SARS coronavirus 2+MERS coronavirus RNA:PrThr:Pt:Respiratory:Ord:Probe.amp.tar|SARS coronavirus+SARS-like coronavirus+SARS coronavirus 2+MERS coronavirus RNA:PrThr:Pt:Respiratory:Ord:Probe.amp.tar
C5234678|T201|OSN|94532-9|LNC_SPECIAL_USE|SARS+SARS-Lk+SARS-CoV-2+MERS Ql NAA-prb|SARS+SARS-Lk+SARS-CoV-2+MERS Ql NAA-prb
C5234679|T201|LC|94534-5|LNC_SPECIAL_USE|SARS coronavirus 2 RdRp gene [Presence] in Respiratory specimen by NAA with probe detection|SARS coronavirus 2 RdRp gene [Presence] in Respiratory specimen by NAA with probe detection
C5234679|T201|LN|94534-5|LNC_SPECIAL_USE|SARS coronavirus 2 RdRp gene:PrThr:Pt:Respiratory:Ord:Probe.amp.tar|SARS coronavirus 2 RdRp gene:PrThr:Pt:Respiratory:Ord:Probe.amp.tar
C5234679|T201|OSN|94534-5|LNC_SPECIAL_USE|SARS-CoV-2 RdRp gene Resp Ql NAA+probe|SARS-CoV-2 RdRp gene Resp Ql NAA+probe
C5234680|T201|LC|94533-7|LNC_SPECIAL_USE|SARS coronavirus 2 N gene [Presence] in Respiratory specimen by NAA with probe detection|SARS coronavirus 2 N gene [Presence] in Respiratory specimen by NAA with probe detection
C5234680|T201|LN|94533-7|LNC_SPECIAL_USE|SARS coronavirus 2 N gene:PrThr:Pt:Respiratory:Ord:Probe.amp.tar|SARS coronavirus 2 N gene:PrThr:Pt:Respiratory:Ord:Probe.amp.tar
C5234680|T201|OSN|94533-7|LNC_SPECIAL_USE|SARS-CoV-2 N gene Resp Ql NAA+probe|SARS-CoV-2 N gene Resp Ql NAA+probe
C5234682|T201|LC|94500-6|LNC_SPECIAL_USE|SARS coronavirus 2 RNA [Presence] in Respiratory specimen by NAA with probe detection|SARS coronavirus 2 RNA [Presence] in Respiratory specimen by NAA with probe detection
C5234682|T201|LN|94500-6|LNC_SPECIAL_USE|SARS coronavirus 2 RNA:PrThr:Pt:Respiratory:Ord:Probe.amp.tar|SARS coronavirus 2 RNA:PrThr:Pt:Respiratory:Ord:Probe.amp.tar
C5234682|T201|OSN|94500-6|LNC_SPECIAL_USE|SARS-CoV-2 RNA Resp Ql NAA+probe|SARS-CoV-2 RNA Resp Ql NAA+probe
C5234683|T201|OSN|94501-4|LNC_SPECIAL_USE|MERS-CoV RNA Resp Ql NAA+probe|MERS-CoV RNA Resp Ql NAA+probe
C5234683|T201|LC|94501-4|LNC_SPECIAL_USE|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Respiratory specimen by NAA with probe detection|Middle East respiratory syndrome coronavirus (MERS-CoV) RNA [Presence] in Respiratory specimen by NAA with probe detection
C5234683|T201|LN|94501-4|LNC_SPECIAL_USE|Middle east respiratory syndrome coronavirus RNA:PrThr:Pt:Respiratory:Ord:Probe.amp.tar|Middle east respiratory syndrome coronavirus RNA:PrThr:Pt:Respiratory:Ord:Probe.amp.tar
C5234684|T201|LC|94502-2|LNC_SPECIAL_USE|SARS coronavirus+SARS-like coronavirus+SARS coronavirus 2 RNA [Presence] in Respiratory specimen by NAA with probe detection|SARS coronavirus+SARS-like coronavirus+SARS coronavirus 2 RNA [Presence] in Respiratory specimen by NAA with probe detection
C5234684|T201|LN|94502-2|LNC_SPECIAL_USE|SARS coronavirus+SARS-like coronavirus+SARS coronavirus 2 RNA:PrThr:Pt:Respiratory:Ord:Probe.amp.tar|SARS coronavirus+SARS-like coronavirus+SARS coronavirus 2 RNA:PrThr:Pt:Respiratory:Ord:Probe.amp.tar
C5234684|T201|OSN|94502-2|LNC_SPECIAL_USE|SARS+SARS-Lk+SARS-CoV-2 RNA Resp Ql NAA|SARS+SARS-Lk+SARS-CoV-2 RNA Resp Ql NAA
C5234685|T201|LN|94503-0|LNC_SPECIAL_USE|SARS coronavirus 2 Ab.IgG & IgM panel:-:Pt:Ser/Plas:Ord:IA|SARS coronavirus 2 Ab.IgG & IgM panel:-:Pt:Ser/Plas:Ord:IA
C5234685|T201|LC|94503-0|LNC_SPECIAL_USE|SARS coronavirus 2 IgG and IgM panel - Serum or Plasma Qualitative by Immunoassay|SARS coronavirus 2 IgG and IgM panel - Serum or Plasma Qualitative by Immunoassay
C5234685|T201|OSN|94503-0|LNC_SPECIAL_USE|SARS-CoV-2 IgG+IgM Pnl SerPl IA|SARS-CoV-2 IgG+IgM Pnl SerPl IA
C5234686|T201|LN|94505-5|LNC_SPECIAL_USE|SARS coronavirus 2 Ab.IgG:ACnc:Pt:Ser/Plas:Qn:IA|SARS coronavirus 2 Ab.IgG:ACnc:Pt:Ser/Plas:Qn:IA
C5234686|T201|LC|94505-5|LNC_SPECIAL_USE|SARS coronavirus 2 IgG Ab [Units/volume] in Serum or Plasma by Immunoassay|SARS coronavirus 2 IgG Ab [Units/volume] in Serum or Plasma by Immunoassay
C5234686|T201|OSN|94505-5|LNC_SPECIAL_USE|SARS-CoV-2 IgG SerPl IA-aCnc|SARS-CoV-2 IgG SerPl IA-aCnc
C5234687|T201|LN|94506-3|LNC_SPECIAL_USE|SARS coronavirus 2 Ab.IgM:ACnc:Pt:Ser/Plas:Qn:IA|SARS coronavirus 2 Ab.IgM:ACnc:Pt:Ser/Plas:Qn:IA
C5234687|T201|LC|94506-3|LNC_SPECIAL_USE|SARS coronavirus 2 IgM Ab [Units/volume] in Serum or Plasma by Immunoassay|SARS coronavirus 2 IgM Ab [Units/volume] in Serum or Plasma by Immunoassay
C5234687|T201|OSN|94506-3|LNC_SPECIAL_USE|SARS-CoV-2 IgM SerPl IA-aCnc|SARS-CoV-2 IgM SerPl IA-aCnc
C5234688|T201|LN|94504-8|LNC_SPECIAL_USE|SARS coronavirus 2 Ab.IgG & IgM panel:-:Pt:Ser/Plas:Qn:IA|SARS coronavirus 2 Ab.IgG & IgM panel:-:Pt:Ser/Plas:Qn:IA
C5234688|T201|LC|94504-8|LNC_SPECIAL_USE|SARS coronavirus 2 IgG and IgM panel - Serum or Plasma by Immunoassay|SARS coronavirus 2 IgG and IgM panel - Serum or Plasma by Immunoassay
C5234688|T201|OSN|94504-8|LNC_SPECIAL_USE|SARS-CoV-2 IgG+IgM Pnl SerPl IA-aCnc|SARS-CoV-2 IgG+IgM Pnl SerPl IA-aCnc
C5234689|T201|LN|94508-9|LNC_SPECIAL_USE|SARS coronavirus 2 Ab.IgM:PrThr:Pt:Ser/Plas:Ord:IA|SARS coronavirus 2 Ab.IgM:PrThr:Pt:Ser/Plas:Ord:IA
C5234689|T201|LC|94508-9|LNC_SPECIAL_USE|SARS coronavirus 2 IgM Ab [Presence] in Serum or Plasma by Immunoassay|SARS coronavirus 2 IgM Ab [Presence] in Serum or Plasma by Immunoassay
C5234689|T201|OSN|94508-9|LNC_SPECIAL_USE|SARS-CoV-2 IgM SerPl Ql IA|SARS-CoV-2 IgM SerPl Ql IA
C5234690|T201|LC|94509-7|LNC_SPECIAL_USE|SARS coronavirus 2 E gene [Cycle Threshold #] in Unspecified specimen by NAA with probe detection|SARS coronavirus 2 E gene [Cycle Threshold #] in Unspecified specimen by NAA with probe detection
C5234690|T201|LN|94509-7|LNC_SPECIAL_USE|SARS coronavirus 2 E gene:ThreshNum:Pt:XXX:Qn:Probe.amp.tar|SARS coronavirus 2 E gene:ThreshNum:Pt:XXX:Qn:Probe.amp.tar
C5234690|T201|OSN|94509-7|LNC_SPECIAL_USE|SARS-CoV-2 E gene Ct XXX Qn NAA+probe|SARS-CoV-2 E gene Ct XXX Qn NAA+probe
C5234691|T201|LN|94507-1|LNC_SPECIAL_USE|SARS coronavirus 2 Ab.IgG:PrThr:Pt:Ser/Plas:Ord:IA|SARS coronavirus 2 Ab.IgG:PrThr:Pt:Ser/Plas:Ord:IA
C5234691|T201|LC|94507-1|LNC_SPECIAL_USE|SARS coronavirus 2 IgG Ab [Presence] in Serum or Plasma by Immunoassay|SARS coronavirus 2 IgG Ab [Presence] in Serum or Plasma by Immunoassay
C5234691|T201|OSN|94507-1|LNC_SPECIAL_USE|SARS-CoV-2 IgG SerPl Ql IA|SARS-CoV-2 IgG SerPl Ql IA
C5234692|T201|LC|94510-5|LNC_SPECIAL_USE|SARS coronavirus 2 N gene [Cycle Threshold #] in Unspecified specimen by NAA with probe detection|SARS coronavirus 2 N gene [Cycle Threshold #] in Unspecified specimen by NAA with probe detection
C5234692|T201|LN|94510-5|LNC_SPECIAL_USE|SARS coronavirus 2 N gene:ThreshNum:Pt:XXX:Qn:Probe.amp.tar|SARS coronavirus 2 N gene:ThreshNum:Pt:XXX:Qn:Probe.amp.tar
C5234692|T201|OSN|94510-5|LNC_SPECIAL_USE|SARS-CoV-2 N gene Ct XXX Qn NAA+probe|SARS-CoV-2 N gene Ct XXX Qn NAA+probe
C5234693|T201|LC|94511-3|LNC_SPECIAL_USE|SARS coronavirus 2 ORF1ab region [Cycle Threshold #] in Unspecified specimen by NAA with probe detection|SARS coronavirus 2 ORF1ab region [Cycle Threshold #] in Unspecified specimen by NAA with probe detection
C5234693|T201|LN|94511-3|LNC_SPECIAL_USE|SARS coronavirus 2 ORF1ab region:ThreshNum:Pt:XXX:Qn:Probe.amp.tar|SARS coronavirus 2 ORF1ab region:ThreshNum:Pt:XXX:Qn:Probe.amp.tar
C5234693|T201|OSN|94511-3|LNC_SPECIAL_USE|SARS-CoV-2 ORF1ab Ct XXX Qn NAA+probe|SARS-CoV-2 ORF1ab Ct XXX Qn NAA+probe
C5234694|T201|LC|94306-8|LNC_SPECIAL_USE|SARS Coronavirus 2 RNA panel - Unspecified specimen by NAA with probe detection|SARS Coronavirus 2 RNA panel - Unspecified specimen by NAA with probe detection
C5234694|T201|LN|94306-8|LNC_SPECIAL_USE|SARS coronavirus 2 RNA panel:-:Pt:XXX:-:Probe.amp.tar|SARS coronavirus 2 RNA panel:-:Pt:XXX:-:Probe.amp.tar
C5234694|T201|OSN|94306-8|LNC_SPECIAL_USE|SARS-CoV-2 RNA Pnl XXX NAA+probe|SARS-CoV-2 RNA Pnl XXX NAA+probe
C5234695|T201|LC|94307-6|LNC_SPECIAL_USE|SARS coronavirus 2 N gene [Presence] in Unspecified specimen by Nucleic acid amplification using primer-probe set N1|SARS coronavirus 2 N gene [Presence] in Unspecified specimen by Nucleic acid amplification using primer-probe set N1
C5234695|T201|LN|94307-6|LNC_SPECIAL_USE|SARS coronavirus 2 N gene:PrThr:Pt:XXX:Ord:Probe.amp.tar.primer-probe set N1|SARS coronavirus 2 N gene:PrThr:Pt:XXX:Ord:Probe.amp.tar.primer-probe set N1
C5234695|T201|OSN|94307-6|LNC_SPECIAL_USE|SARS-CoV-2 N gene XXX Ql NAA N1|SARS-CoV-2 N gene XXX Ql NAA N1
C5234696|T201|LC|94308-4|LNC_SPECIAL_USE|SARS coronavirus 2 N gene [Presence] in Unspecified specimen by Nucleic acid amplification using primer-probe set N2|SARS coronavirus 2 N gene [Presence] in Unspecified specimen by Nucleic acid amplification using primer-probe set N2
C5234696|T201|LN|94308-4|LNC_SPECIAL_USE|SARS coronavirus 2 N gene:PrThr:Pt:XXX:Ord:Probe.amp.tar.primer-probe set N2|SARS coronavirus 2 N gene:PrThr:Pt:XXX:Ord:Probe.amp.tar.primer-probe set N2
C5234696|T201|OSN|94308-4|LNC_SPECIAL_USE|SARS-CoV-2 N gene XXX Ql NAA N2|SARS-CoV-2 N gene XXX Ql NAA N2
C5234697|T201|LC|94309-2|LNC_SPECIAL_USE|SARS coronavirus 2 RNA [Presence] in Unspecified specimen by NAA with probe detection|SARS coronavirus 2 RNA [Presence] in Unspecified specimen by NAA with probe detection
C5234697|T201|LN|94309-2|LNC_SPECIAL_USE|SARS coronavirus 2 RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar|SARS coronavirus 2 RNA:PrThr:Pt:XXX:Ord:Probe.amp.tar
C5234697|T201|OSN|94309-2|LNC_SPECIAL_USE|SARS-CoV-2 RNA XXX Ql NAA+probe|SARS-CoV-2 RNA XXX Ql NAA+probe
C5234698|T201|LC|94312-6|LNC_SPECIAL_USE|SARS coronavirus 2 N gene [Cycle Threshold #] in Unspecified specimen by Nucleic acid amplification using primer-probe set N2|SARS coronavirus 2 N gene [Cycle Threshold #] in Unspecified specimen by Nucleic acid amplification using primer-probe set N2
C5234698|T201|LN|94312-6|LNC_SPECIAL_USE|SARS coronavirus 2 N gene:ThreshNum:Pt:XXX:Qn:Probe.amp.tar.primer-probe set N2|SARS coronavirus 2 N gene:ThreshNum:Pt:XXX:Qn:Probe.amp.tar.primer-probe set N2
C5234698|T201|OSN|94312-6|LNC_SPECIAL_USE|SARS-CoV-2 N gene Ct XXX Qn NAA N2|SARS-CoV-2 N gene Ct XXX Qn NAA N2
C5234699|T201|LC|94310-0|LNC_SPECIAL_USE|SARS-like Coronavirus N gene [Presence] in Unspecified specimen by NAA with probe detection|SARS-like Coronavirus N gene [Presence] in Unspecified specimen by NAA with probe detection
C5234699|T201|LN|94310-0|LNC_SPECIAL_USE|SARS-like Coronavirus N gene:PrThr:Pt:XXX:Ord:Probe.amp.tar|SARS-like Coronavirus N gene:PrThr:Pt:XXX:Ord:Probe.amp.tar
C5234699|T201|OSN|94310-0|LNC_SPECIAL_USE|SARS-like CoV N XXX Ql NAA+probe|SARS-like CoV N XXX Ql NAA+probe
C5234700|T201|LC|94311-8|LNC_SPECIAL_USE|SARS coronavirus 2 N gene [Cycle Threshold #] in Unspecified specimen by Nucleic acid amplification using primer-probe set N1|SARS coronavirus 2 N gene [Cycle Threshold #] in Unspecified specimen by Nucleic acid amplification using primer-probe set N1
C5234700|T201|LN|94311-8|LNC_SPECIAL_USE|SARS coronavirus 2 N gene:ThreshNum:Pt:XXX:Qn:Probe.amp.tar.primer-probe set N1|SARS coronavirus 2 N gene:ThreshNum:Pt:XXX:Qn:Probe.amp.tar.primer-probe set N1
C5234700|T201|OSN|94311-8|LNC_SPECIAL_USE|SARS-CoV-2 N gene Ct XXX Qn NAA N1|SARS-CoV-2 N gene Ct XXX Qn NAA N1
C5234701|T201|LC|94313-4|LNC_SPECIAL_USE|SARS-like Coronavirus N gene [Cycle Threshold #] in Unspecified specimen by NAA with probe detection|SARS-like Coronavirus N gene [Cycle Threshold #] in Unspecified specimen by NAA with probe detection
C5234701|T201|LN|94313-4|LNC_SPECIAL_USE|SARS-like Coronavirus N gene:ThreshNum:Pt:XXX:Qn:Probe.amp.tar|SARS-like Coronavirus N gene:ThreshNum:Pt:XXX:Qn:Probe.amp.tar
C5234701|T201|OSN|94313-4|LNC_SPECIAL_USE|SARS-like CoV N Ct XXX Qn NAA+probe|SARS-like CoV N Ct XXX Qn NAA+probe
C5234702|T201|LC|94314-2|LNC_SPECIAL_USE|SARS coronavirus 2 RdRp gene [Presence] in Unspecified specimen by NAA with probe detection|SARS coronavirus 2 RdRp gene [Presence] in Unspecified specimen by NAA with probe detection
C5234702|T201|LN|94314-2|LNC_SPECIAL_USE|SARS coronavirus 2 RdRp gene:PrThr:Pt:XXX:Ord:Probe.amp.tar|SARS coronavirus 2 RdRp gene:PrThr:Pt:XXX:Ord:Probe.amp.tar
C5234702|T201|OSN|94314-2|LNC_SPECIAL_USE|SARS-CoV-2 RdRp gene XXX Ql NAA+probe|SARS-CoV-2 RdRp gene XXX Ql NAA+probe
C5234703|T201|LC|94315-9|LNC_SPECIAL_USE|SARS coronavirus 2 E gene [Presence] in Unspecified specimen by NAA with probe detection|SARS coronavirus 2 E gene [Presence] in Unspecified specimen by NAA with probe detection
C5234703|T201|LN|94315-9|LNC_SPECIAL_USE|SARS coronavirus 2 E gene:PrThr:Pt:XXX:Ord:Probe.amp.tar|SARS coronavirus 2 E gene:PrThr:Pt:XXX:Ord:Probe.amp.tar
C5234703|T201|OSN|94315-9|LNC_SPECIAL_USE|SARS-CoV-2 E gene XXX Ql NAA+probe|SARS-CoV-2 E gene XXX Ql NAA+probe
C5234704|T201|LC|94316-7|LNC_SPECIAL_USE|SARS coronavirus 2 N gene [Presence] in Unspecified specimen by NAA with probe detection|SARS coronavirus 2 N gene [Presence] in Unspecified specimen by NAA with probe detection
C5234704|T201|LN|94316-7|LNC_SPECIAL_USE|SARS coronavirus 2 N gene:PrThr:Pt:XXX:Ord:Probe.amp.tar|SARS coronavirus 2 N gene:PrThr:Pt:XXX:Ord:Probe.amp.tar
C5234704|T201|OSN|94316-7|LNC_SPECIAL_USE|SARS-CoV-2 N gene XXX Ql NAA+probe|SARS-CoV-2 N gene XXX Ql NAA+probe
C0949880|T005|ET|D028941|MSH|HCoV229E|HCoV-229E
C1312200|T116|CE|C477905|MSH|PLP2, coronavirus|PLP-2, coronavirus
C1312200|T126|CE|C477905|MSH|PLP2, coronavirus|PLP-2, coronavirus
C1532880|T005|PT|415398003|SNOMEDCT_US|SARS coronavirus HPZ2003|SARS coronavirus HPZ-2003
C1532880|T005|OF|415398003|SNOMEDCT_US|SARS coronavirus HPZ2003 (organism)|SARS coronavirus HPZ-2003 (organism)
C1532880|T005|SY|415398003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HPZ2003|Severe acute respiratory syndrome (SARS) coronavirus HPZ-2003
C1532880|T005|OF|415398003|SNOMEDCT_US|Severe acute respiratory syndrome (SARS) coronavirus HPZ2003 (organism)|Severe acute respiratory syndrome (SARS) coronavirus HPZ-2003 (organism)
C1532880|T005|SY|415398003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HPZ2003|Severe acute respiratory syndrome coronavirus HPZ-2003
C1532880|T005|FN|415398003|SNOMEDCT_US|Severe acute respiratory syndrome coronavirus HPZ2003 (organism)|Severe acute respiratory syndrome coronavirus HPZ-2003 (organism)
C5203672|T061|PN|NOCODE|MTH|SARS-CoV2 vaccination|SARS-CoV-2 vaccination
C5203673|T116|PN|NOCODE|MTH|Antigen of SARS-CoV2|Antigen of SARS-CoV-2
C5203673|T129|PN|NOCODE|MTH|Antigen of SARS-CoV2|Antigen of SARS-CoV-2
C5203674|T116|PN|NOCODE|MTH|Antibody to SARS-CoV2|Antibody to SARS-CoV-2
C5203674|T129|PN|NOCODE|MTH|Antibody to SARS-CoV2|Antibody to SARS-CoV-2
C5203675|T033|PN|NOCODE|MTH|Exposure to SARS-CoV2|Exposure to SARS-CoV-2
C5203676|T005|PN|NOCODE|MTH|SARS-CoV2|SARS-CoV-2
C5234677|T201|OSN|94531-1|LNC_SPECIAL_USE|SARS-CoV2 RNA Pnl Resp NAA+probe|SARS-CoV-2 RNA Pnl Resp NAA+probe
C5234678|T201|OSN|94532-9|LNC_SPECIAL_USE|SARS+SARS-Lk+SARS-CoV2+MERS Ql NAA-prb|SARS+SARS-Lk+SARS-CoV-2+MERS Ql NAA-prb
C5234679|T201|OSN|94534-5|LNC_SPECIAL_USE|SARS-CoV2 RdRp gene Resp Ql NAA+probe|SARS-CoV-2 RdRp gene Resp Ql NAA+probe
C5234680|T201|OSN|94533-7|LNC_SPECIAL_USE|SARS-CoV2 N gene Resp Ql NAA+probe|SARS-CoV-2 N gene Resp Ql NAA+probe
C5234682|T201|OSN|94500-6|LNC_SPECIAL_USE|SARS-CoV2 RNA Resp Ql NAA+probe|SARS-CoV-2 RNA Resp Ql NAA+probe
C5234684|T201|OSN|94502-2|LNC_SPECIAL_USE|SARS+SARS-Lk+SARS-CoV2 RNA Resp Ql NAA|SARS+SARS-Lk+SARS-CoV-2 RNA Resp Ql NAA
C5234685|T201|OSN|94503-0|LNC_SPECIAL_USE|SARS-CoV2 IgG+IgM Pnl SerPl IA|SARS-CoV-2 IgG+IgM Pnl SerPl IA
C5234686|T201|OSN|94505-5|LNC_SPECIAL_USE|SARS-CoV2 IgG SerPl IA-aCnc|SARS-CoV-2 IgG SerPl IA-aCnc
C5234687|T201|OSN|94506-3|LNC_SPECIAL_USE|SARS-CoV2 IgM SerPl IA-aCnc|SARS-CoV-2 IgM SerPl IA-aCnc
C5234688|T201|OSN|94504-8|LNC_SPECIAL_USE|SARS-CoV2 IgG+IgM Pnl SerPl IA-aCnc|SARS-CoV-2 IgG+IgM Pnl SerPl IA-aCnc
C5234689|T201|OSN|94508-9|LNC_SPECIAL_USE|SARS-CoV2 IgM SerPl Ql IA|SARS-CoV-2 IgM SerPl Ql IA
C5234690|T201|OSN|94509-7|LNC_SPECIAL_USE|SARS-CoV2 E gene Ct XXX Qn NAA+probe|SARS-CoV-2 E gene Ct XXX Qn NAA+probe
C5234691|T201|OSN|94507-1|LNC_SPECIAL_USE|SARS-CoV2 IgG SerPl Ql IA|SARS-CoV-2 IgG SerPl Ql IA
C5234692|T201|OSN|94510-5|LNC_SPECIAL_USE|SARS-CoV2 N gene Ct XXX Qn NAA+probe|SARS-CoV-2 N gene Ct XXX Qn NAA+probe
C5234693|T201|OSN|94511-3|LNC_SPECIAL_USE|SARS-CoV2 ORF1ab Ct XXX Qn NAA+probe|SARS-CoV-2 ORF1ab Ct XXX Qn NAA+probe
C5234694|T201|OSN|94306-8|LNC_SPECIAL_USE|SARS-CoV2 RNA Pnl XXX NAA+probe|SARS-CoV-2 RNA Pnl XXX NAA+probe
C5234695|T201|OSN|94307-6|LNC_SPECIAL_USE|SARS-CoV2 N gene XXX Ql NAA N1|SARS-CoV-2 N gene XXX Ql NAA N1
C5234696|T201|OSN|94308-4|LNC_SPECIAL_USE|SARS-CoV2 N gene XXX Ql NAA N2|SARS-CoV-2 N gene XXX Ql NAA N2
C5234697|T201|OSN|94309-2|LNC_SPECIAL_USE|SARS-CoV2 RNA XXX Ql NAA+probe|SARS-CoV-2 RNA XXX Ql NAA+probe
C5234698|T201|OSN|94312-6|LNC_SPECIAL_USE|SARS-CoV2 N gene Ct XXX Qn NAA N2|SARS-CoV-2 N gene Ct XXX Qn NAA N2
C5234700|T201|OSN|94311-8|LNC_SPECIAL_USE|SARS-CoV2 N gene Ct XXX Qn NAA N1|SARS-CoV-2 N gene Ct XXX Qn NAA N1
C5234702|T201|OSN|94314-2|LNC_SPECIAL_USE|SARS-CoV2 RdRp gene XXX Ql NAA+probe|SARS-CoV-2 RdRp gene XXX Ql NAA+probe
C5234703|T201|OSN|94315-9|LNC_SPECIAL_USE|SARS-CoV2 E gene XXX Ql NAA+probe|SARS-CoV-2 E gene XXX Ql NAA+probe
C5234704|T201|OSN|94316-7|LNC_SPECIAL_USE|SARS-CoV2 N gene XXX Ql NAA+probe|SARS-CoV-2 N gene XXX Ql NAA+probe
C5203670|T047|PN|NOCODE|MTH|COVID19|COVID-19
C5203671|T033|PN|NOCODE|MTH|Suspected COVID19|Suspected COVID-19
