C0002210|T034||LNC|ALPHA-FETOPROTEINS
C0201539|T034||LNC|ALPHA ONE FETOPROTEIN MEASUREMENT
C0002210|T034||LNC|ALPHA FETOPROTEIN
C0002210|T034||LNC|ALPHA FETOPROTEINS
C0002210|T034||LNC|ALPHA-FETOPROTEINS
C0002210|T034||LNC|ALPHA FOETOPROTEIN
C0002210|T034||LNC|ALPHA-FETOPROTEIN
C0002210|T034||LNC|ALPHA-FETOPROTEINS [CHEMICAL/INGREDIENT]
C0002210|T034||LNC|ALPHA-1-FETOPROTEIN
C0002210|T034||LNC|AFP
C0002210|T034||LNC|ALPHA FETAL PROTEIN
C0002210|T034||LNC|AFP - ALPHA-FETOPROTEIN
C0002210|T034||LNC|ALPHA FETOPROTEIN 
C0002210|T034||LNC|ALPHA-FETOGLOBULIN
C1981150|T034|LP43503-9|LNC|ALPHA-1-FETOPROTEIN AMNIOTIC FLUID|ALPHA-1-FETOPROTEIN &#X7C; AMNIOTIC FLUID
C2600377|T034|LP89453-2|LNC|ALPHA-1-FETOPROTEIN BLOOD CORD|ALPHA-1-FETOPROTEIN &#X7C; BLOOD CORD
C1981155|T034|LP64841-7|LNC|ALPHA-1-FETOPROTEIN PERITONEAL FLUID|ALPHA-1-FETOPROTEIN &#X7C; PERITONEAL FLUID
C1981152|T034|LP41454-7|LNC|ALPHA-1-FETOPROTEIN BODY FLUID|ALPHA-1-FETOPROTEIN &#X7C; BODY FLUID
C1981151|T034|LP45776-9|LNC|ALPHA-1-FETOPROTEIN BLD-SER-PLAS|ALPHA-1-FETOPROTEIN &#X7C; BLD-SER-PLAS
C2600378|T034|LP71676-8|LNC|ALPHA-1-FETOPROTEIN TUMOR MARKER BLD-SER-PLAS|ALPHA-1-FETOPROTEIN.TUMOR MARKER &#X7C; BLD-SER-PLAS
C1981156|T034|LP46116-7|LNC|ALPHA-1-FETOPROTEIN &#X7C; PLEURAL FLUID|ALPHA-1-FETOPROTEIN &#X7C; PLEURAL FLUID
C1307640|T034||LNC|AFP PROTEIN, HUMAN
C1307640|T034||LNC|ALPHA-FETOPROTEIN, HUMAN
# C1307640|T034||LNC| CAN'T FIND ANYTHING THAT CONFIRMS OR DENYS THAT ALPHA GLYCOPROTEIN FETOSPECIFIC IS AFP, LEAVING ON FOR NOW, BUT MAY CONSIDER EXCLUDING (THE CHANCES YOU SEE THIS EXACT MATCH IN A MEDICAL RECORD IS VERY LOW)
C1307640|T034||LNC|ALPHA-GLYCOPROTEIN, FETOSPECIFIC, HUMAN
C1307640|T034||LNC|AF GLYCOPROTEIN, HUMAN
C0201539|T034||LNC|AFP
C0201539|T034||LNC|ALPHA 1 FOETOPROTEIN
C0201539|T034||LNC|AFP ALPHAFOETOPROTEIN
C0201539|T034||LNC|ALPHA-FETOPROTEIN MEASUREMENT
C0201539|T034||LNC|ALPHA-1-FOETOPROTEIN MEASUREMENT
C0201539|T034||LNC|ALPHA FOETOPROTEIN MEASUREMENT
C0201539|T034||LNC|ALPHA ONE FETOPROTEIN MEASUREMENT
C0201539|T034||LNC|TEST;ALPHA FETOPROTEIN
C0201539|T034||LNC|ALPHA-FETOPROTEIN NOS
C0201539|T034||LNC|ALPHA-FETOPROTEIN NOS 
C0201539|T034||LNC|ALPHA-FETOPROTEIN (AFP)
C0201539|T034||LNC|ALPHA FETOPROTEIN
C0201539|T034||LNC|ALPHA-1-FETOPROTEIN MEASUREMENT
C0201539|T034||LNC|ALPHAFETOPROTEIN
C0201539|T034||LNC|ALPHA 1 FETOPROTEIN
C0201539|T034||LNC|ALPHAFOETOPROTEIN
C0201539|T034||LNC|AFP MEASUREMENT
C0201539|T034||LNC|ALPHA FETOPROTEIN MEASUREMENT
C0201539|T034||LNC|ALPHA-1-FETOPROTEIN MEASUREMENT 
C0201539|T034||LNC|ALPHA FETOPROTEIN TEST
C2711551|T034||LNC|MEASUREMENT OF ALPHA FETOPROTEIN AS MARKER FOR MALIGNANT NEOPLASM 
C2711551|T034||LNC|MEASUREMENT OF ALPHA FETOPROTEIN AS MARKER FOR MALIGNANT NEOPLASM
C2368140|T034||LNC|BODY FLUID ALPHA-FETOPROTEIN
C2368140|T034||LNC|BODY FLUID AFP
C2368140|T034||LNC|BODY FLUID ALPHA-FETOPROTEIN MEASUREMENT
C2368140|T034||LNC|BODY FLUID ALPHA-FETOPROTEIN MEASUREMENT 
C0546833|T034||LNC|ALPHA-FETOPROTEIN (AFP); SERUM
C0546833|T034||LNC|SERUM ALPHA-FETOPROTEIN MEASUREMENT 
C0546833|T034||LNC|SERUM AFP
C0546833|T034||LNC|SERUM ALPHA-FETOPROTEIN
C0546833|T034||LNC|SERUM ALPHA-FETOPROTEIN MEASUREMENT
C0546833|T034||LNC|SERUM ALPHA-FETOPROTEIN (AFP) MEASUREMENT
C0546833|T034||LNC|ALPHA-FETOPROTEIN SERUM
C0546833|T034||LNC|ALPHA-FETOPROTEIN (AFP) LEVEL, SERUM
C0546833|T034||LNC|MEASUREMENT OF ALPHA-FETOPROTEIN (AFP) IN SERUM
C0546833|T034||LNC|ALPHA-FETOPROTEIN (AFP) LEVEL, SERUM"
C0419584|T034||LNC|ALPHA-FETOPROTEIN BLOOD TEST
C0419584|T034||LNC|ALPHA-FETOPROTEIN BLOOD TEST 
C1271788|T034||LNC|FLUID SAMPLE AFP LEVEL 
C1271788|T034||LNC|FLUID SAMPLE ALPHA FETOPROTEIN LEVEL
C1271788|T034||LNC|FLUID SAMPLE ALPHA FETOPROTEIN LEVEL 
C1271788|T034||LNC|FLUID SAMPLE AFP LEVEL
