// CUI|STR|TTY|CODE|SAB|TUI|PREF
C0004096|ASTHMA|BN|195979001|SNOMEDCT_US|T047|ASTHMA UNSPECIFIED (DISORDER)