C0201916|T034||LNC|BILI
C0201916|T034||LNC|BILIRUBIN
C0201916|T034||LNC|BILIRUBIN, DIRECT MEASUREMENT
C0201916|T034||LNC|DIRECT BILI
C0236556|T034||LNC|DIRECT BILIRUBIN
C0236556|T034||LNC|DIRECT REACTING BILIRUBIN
C1883011|T034||LNC|SERUM DIRECT BILIRUBIN MEASUREMENT
C0428439|T034||LNC|CONJUGATED BILIRUBIN LEVEL 
C1278035|T034||LNC|PLASMA CONJUGATED BILIRUBIN LEVEL 
C1278035|T034||LNC|PLASMA CONJUGATED BILIRUBIN MEASUREMENT
C1278038|T034||LNC|SERUM CONJUGATED BILIRUBIN LEVEL 
C1278038|T034||LNC|SERUM DIRECT (CONJUGATED) BILIRUBIN TEST
C1278038|T034||LNC|SERUM CONJUGATED BILIRUBIN MEASUREMENT
