C0555903|T034||LNC|TOTAL PROTEIN MEASUREMENT
C1261360|T034||LNC|TOTAL PROTEIN RESULT
C0036836|T034||LNC|SERUM TOTAL PROTEIN MEASUREMENT
C0580563|T034||LNC|SERUM TOTAL PROTEIN NORMAL
C0580564|T034||LNC|SERUM TOTAL PROTEIN ABNORMAL
C0555903|T034||LNC|TOTAL PROTEIN MEASUREMENT
C0555903|T034||LNC|PROTEIN TOTAL
C0555903|T034||LNC|MEASUREMENT OF TOTAL PROTEIN
C0555903|T034||LNC|PROTEIN
C0555903|T034||LNC|PROT
C0555903|T034||LNC|TOTAL PROTEIN
C0555903|T034||LNC|TP - TOTAL PROTEIN
C0555903|T034||LNC|TPR - TOTAL PROTEIN
C0555903|T034||LNC|TOTAL PROTEIN MEASUREMENT 
C2097239|T034||LNC|SERUM TOTAL PROTEIN BY REFRACTOMETRY 
C2097239|T034||LNC|SERUM TOTAL PROTEIN BY REFRACTOMETRY
C2097239|T034||LNC|TOTAL SERUM PROTEIN LEVEL BY REFRACTOMETRY
C0036836|T034||LNC|SERUM TOTAL PROTEIN MEASUREMENT
C0036836|T034||LNC|TOTAL SERUM PROTEIN LEVEL
C0036836|T034||LNC|SERUM TOTAL PROTEIN MEASUREMENT 
C0036836|T034||LNC|SERUM TOTAL PROTEIN
C0036836|T034||LNC|SERUM PROTEIN TOTAL MEASUREMENT
C0036836|T034||LNC|TOTAL SERUM PROTEIN MEASUREMENT
C0036836|T034||LNC|MEASUREMENT OF TOTAL PROTEIN IN SERUM
C0036836|T034||LNC|SERUM TOTAL PROTEIN (& LEVEL) 
C0036836|T034||LNC|SERUM TOTAL PROTEIN (& LEVEL)
C0036836|T034||LNC|SERUM TOTAL PROTEIN TEST
C0036836|T034||LNC|SERUM TOTAL PROTEIN LEVEL
C0036836|T034||LNC|SERUM TOTAL PROTEIN MEASUREMENT 
C0855756|T034||LNC|PROTEIN TOTAL ABNORMAL
C0855756|T034||LNC|PROTEIN TOTAL ABNORMAL NOS
C0855757|T034||LNC|PROTEIN TOTAL NORMAL
C0855757|T034||LNC|TOTAL PROTEIN NORMAL
C0859351|T034||LNC|SERUM TOTAL PROTEIN INCREASED
C0855758|T034||LNC|PROTEIN TOTAL INCREASED
C0855758|T034||LNC|TOTAL PROTEIN HIGH
C0855758|T034||LNC|PROTEIN TOTAL HIGH
C0860703|T034||LNC|SERUM TOTAL PROTEIN DECREASED
C0860901|T034||LNC|PROTEIN TOTAL DECREASED
C0860901|T034||LNC|DECREASED TOTAL PROTEIN
C0860901|T034||LNC|TOTAL PROTEIN LOW
