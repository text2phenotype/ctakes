C0489786|T034|6071|MEDCIN|HEIGHT|HEIGHT (PHYSICAL FINDING)
C0005890|T034||MEDCIN|BODY HEIGHT
C0424645|T034|297814|MEDCIN|STANDING HEIGHT|STANDING HEIGHT (PHYSICAL FINDING)
C0487985|T034||MEDCIN|BODY HEIGHT:LENGTH:POINT IN TIME:^PATIENT:QUANTITATIVE
C0424639|T034||MEDCIN|HEIGHT / GROWTH MEASURE
C2030323|T034|209270|MEDCIN|HEIGHT ___ PERCENTILE FOR AGE|HEIGHT PERCENTILE FOR AGE (PHYSICAL FINDING)
C2030323|T034|209270|MEDCIN|HEIGHT PERCENTILE FOR AGE|HEIGHT PERCENTILE FOR AGE (PHYSICAL FINDING)
C2030323|T034|209270|MEDCIN|HEIGHT PERCENTILE FOR AGE (PHYSICAL FINDING)|HEIGHT PERCENTILE FOR AGE (PHYSICAL FINDING)
C0424639|T034||MEDCIN|HEIGHT / GROWTH MEASURE
C0424639|T034||MEDCIN|HEIGHT AND GROWTH
C0424639|T034||MEDCIN|LENGTH AND GROWTH
C0424639|T034||MEDCIN|OBSERVATION OF HEIGHT AND GROWTH
C0424639|T034||MEDCIN|HEIGHT / GROWTH MEASURE (OBSERVABLE ENTITY)
C3836210|T034|297815|MEDCIN|RECUMBENT HEIGHT ___|RECUMBENT HEIGHT (PHYSICAL FINDING)
C3836210|T034|297815|MEDCIN|RECUMBENT HEIGHT|RECUMBENT HEIGHT (PHYSICAL FINDING)
C3836210|T034|297815|MEDCIN|RECUMBENT HEIGHT (PHYSICAL FINDING)|RECUMBENT HEIGHT (PHYSICAL FINDING)
C3836390|T034|297816|MEDCIN|PRE-OPERATIVE HEIGHT (PHYSICAL FINDING)|PRE-OPERATIVE HEIGHT (PHYSICAL FINDING)
C3836390|T034|297816|MEDCIN|PRE-OPERATIVE HEIGHT|PRE-OPERATIVE HEIGHT (PHYSICAL FINDING)
C3835668|T034|283414|MEDCIN|STATED HEIGHT|STATED HEIGHT (SYMPTOM)
C3835668|T034|283414|MEDCIN|STATED HEIGHT |STATED HEIGHT (SYMPTOM)
C0424645|T034|297814|MEDCIN|STANDING HEIGHT|STANDING HEIGHT (PHYSICAL FINDING)
C0424645|T034|297814|MEDCIN|STANDING HEIGHT ___|STANDING HEIGHT (PHYSICAL FINDING)
C0424645|T034|297814|MEDCIN|STANDING HEIGHT (PHYSICAL FINDING)|STANDING HEIGHT (PHYSICAL FINDING)
C0424645|T034|297814|MEDCIN|STANDING HEIGHT (OBSERVABLE ENTITY)|STANDING HEIGHT (PHYSICAL FINDING)
C0424646|T034|298056|MEDCIN|SITTING HEIGHT ___|SITTING HEIGHT ___ (PHYSICAL FINDING)
C0424646|T034|298056|MEDCIN|SITTING HEIGHT ___ (PHYSICAL FINDING)|SITTING HEIGHT ___ (PHYSICAL FINDING)
C0424646|T034|298056|MEDCIN|SITTING HEIGHT|SITTING HEIGHT ___ (PHYSICAL FINDING)
C0424646|T034|298056|MEDCIN|SITTING HEIGHT (OBSERVABLE ENTITY)|SITTING HEIGHT ___ (PHYSICAL FINDING)
C1842215|T034||MEDCIN|ADULT MALE HEIGHT 142-169 CM
C1850172|T034||MEDCIN|ADULT HEIGHT 92-108 CM
C1854762|T034||MEDCIN|ADULT HEIGHT 110-140 CM
C1854812|T034||MEDCIN|ADULT HEIGHT 82 TO 115 CM
C1854812|T034||MEDCIN|ADULT HEIGHT 82-115 CM
C1834972|T034||MEDCIN|ADULT HEIGHT 130-160CM
C1865835|T034||MEDCIN|ADULT FEMALE HEIGHT 152-167CM
C1840336|T034||MEDCIN|FINAL HEIGHT, 125 TO 160 CM
C1866721|T034||MEDCIN|FINAL ADULT HEIGHT, 84-128CM
C1851987|T034||MEDCIN|ADULT HEIGHT 135CM TO NORMAL
C1834951|T034||MEDCIN|FINAL ADULT HEIGHT 106-145CM
C1867125|T034||MEDCIN|AVERAGE ADULT FEMALE HEIGHT 147 CM
C1849528|T034||MEDCIN|AVERAGE ADULT FEMALE HEIGHT 135 (4'5")
C1864359|T034||MEDCIN|FINAL ADULT HEIGHT 38-49 INCHES
C1865834|T034||MEDCIN|ADULT MALE HEIGHT 167-173CM
C1839692|T034||MEDCIN|ADULT HEIGHT 120-150CM
C1857182|T034||MEDCIN|ADULT HEIGHT 98-127 CM
C1855747|T034||MEDCIN|ADULT MALE HEIGHT 136-157 CM
C1839249|T034||MEDCIN|FINAL ADULT HEIGHT 131-156 CM
C1849935|T034||MEDCIN|ADULT MALE HEIGHT 141-155CM
C1842216|T034||MEDCIN|ADULT FEMALE HEIGHT 130-157 CM
C0221097|T034||MEDCIN|TOTAL BODY LENGTH
C0221097|T034||MEDCIN|BODY LENGTH
C0221097|T034||MEDCIN|BODLNGTH
C0221097|T034||MEDCIN|LENGTH OF BODY
C0221097|T034||MEDCIN|LENGTH OF BODY (OBSERVABLE ENTITY)
C0005890|T034||MEDCIN|BODY HEIGHT
C0005890|T034||MEDCIN|BODY HEIGHTS
C0005890|T034||MEDCIN|HEIGHT, BODY
C0005890|T034||MEDCIN|HEIGHTS, BODY
C0005890|T034||MEDCIN|STATURE
C0005890|T034||MEDCIN|BODY HEIGHT MEASURE (OBSERVABLE ENTITY)
C0005890|T034||MEDCIN|BODY HEIGHT MEASURE
C0005890|T034||MEDCIN|BODY HEIGHT, NOS
C0005890|T034||MEDCIN|BODY LENGTH
C0005890|T034||MEDCIN|BODY LENGTH, NOS
C0005890|T034||MEDCIN|HEIGHT (BODY)
C0424648|T034||MEDCIN|HEIGHT FROM DEMISPAN
C0424648|T034||MEDCIN|HEIGHT FROM DEMISPAN (OBSERVABLE ENTITY)
C1827986|T034||MEDCIN|METHOD FOR MEASURING HEIGHT
C1827986|T034||MEDCIN|METHOD FOR MEASURING HEIGHT (OBSERVABLE ENTITY)
C0487985|T034||MEDCIN|BODY HEIGHT:LENGTH:POINT IN TIME:^PATIENT:QUANTITATIVE
C0487985|T034||MEDCIN|BODY HEIGHT
C0487985|T034||MEDCIN|BODY HEIGHT:LEN:PT:^PATIENT:QN
C0424649|T034||MEDCIN|HEIGHT CENTILE
C0424649|T034||MEDCIN|LENGTH CENTILE
C0424649|T034||MEDCIN|HEIGHT CENTILE (OBSERVABLE ENTITY)
C0419485|T034||MEDCIN|CHILD HEIGHT CENTILES
C0419485|T034||MEDCIN|HEIGHT CENTILES - CHILD
C0419485|T034||MEDCIN|CHILD HEIGHT CENTILES NOS
C0419485|T034||MEDCIN|CHILD HEIGHT CENTILES NOS 
C0419485|T034||MEDCIN|CHILD HEIGHT CENTILES NOS (OBSERVABLE ENTITY)
C0419485|T034||MEDCIN|CHILD HEIGHT CENTILE (OBSERVABLE ENTITY)
C0419485|T034||MEDCIN|CHILD HEIGHT CENTILE
C1156245|T034||MEDCIN|GROWTH PATTERN (OBSERVABLE ENTITY)
C1156245|T034||MEDCIN|GROWTH PATTERN
C0424638|T034||MEDCIN|HEIGHT AND WEIGHT
C0424638|T034||MEDCIN|HEIGHT AND WEIGHT (OBSERVABLE ENTITY)
C0424638|T034||MEDCIN|HEIGHT & WEIGHT
