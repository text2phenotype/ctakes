C0021682|T058||CSP|HEALTH INSURANCE
C0018717|T058|1385-6531|CSP|MEDICARE|MEDICARE
C0018717|T058|1385-6531|CSP|MEDICARE COVERAGE|MEDICARE
C3530230|T058||CSP|PRIVATE HEALTH INSURANCE
C3530230|T058||CSP|PRIVATE HEALTH INSURANCE--OTHER COMMERCIAL INDEMNITY
C4069202|T058||CSP|PRIVATE INSURANCE (INCLUDES "NO-FAULT", BCBS, UNITED HEALTH, ETC)
C2347682|T058||CSP|PRIVATE HEALTH INSURANCE
C1955981|T058||CSP|BLUE CROSS BLUE SHIELD
C1955981|T058||CSP|BLUE CROSS BLUE SHIELD INSURANCE
C1955981|T058||CSP|BLUE CROSS BLUE SHIELD INSURANCE PLANS
C0005864|T058||CSP|BLUE CROSS
C0021681|T058|1385-6500|CSP|INSURANCE, DENTAL|DENTAL HEALTH INSURANCE
C0021681|T058|1385-6500|CSP|DENTAL HEALTH INSURANCE|DENTAL HEALTH INSURANCE
C0021681|T058|1385-6500|CSP|INSURANCE DENT|DENTAL HEALTH INSURANCE
C0021681|T058|1385-6500|CSP|DENT INSURANCE|DENTAL HEALTH INSURANCE
C0021681|T058|1385-6500|CSP|DENTAL INSURANCE|DENTAL HEALTH INSURANCE
C0596896|T058||CSP|MEDICARE/MEDICAID
C0018717|T058|1385-6531|CSP|MEDICARE|MEDICARE
C0018717|T058|1385-6531|CSP|HEALTH INSURANCE AGED DISABLED|MEDICARE
C0018717|T058|1385-6531|CSP|HEALTH INSURANCE AGED DISABLED TITLE 18|MEDICARE
C0018717|T058|1385-6531|CSP|HEALTH INSURANCE AGED TITLE 18|MEDICARE
C0018717|T058|1385-6531|CSP|MEDICARE PROGRAM|MEDICARE
C0018717|T058|1385-6531|CSP|MEDICARE COVERAGE |MEDICARE
C0018717|T058|1385-6531|CSP|MEDICARE COVERAGE|MEDICARE
C0018717|T058|1385-6531|CSP|HEALTH INSURANCE FOR AGED, DISABLED, TITLE 18|MEDICARE
C0018717|T058|1385-6531|CSP|HEALTH INSURANCE FOR AGED, TITLE 18|MEDICARE
C0018717|T058|1385-6531|CSP|HEALTH INSURANCE FOR AGED AND DISABLED, TITLE 18|MEDICARE
C0018720|T058|1385-3793|CSP|HEALTH MAINTENANCE ORGANIZATIONS|HMO
C0018720|T058|1385-3793|CSP|HMO|HMO
C0018720|T058|1385-3793|CSP|ORGANIZATION, HEALTH MAINTENANCE|HMO
C0018720|T058|1385-3793|CSP|HEALTH MAINTENANCE ORGANIZATION|HMO
C0018720|T058|1385-3793|CSP|GROUP HEALTH ORGAN PREPAID|HMO
C0018720|T058|1385-3793|CSP|ORGAN HEALTH MAINTENANCE|HMO
C0018720|T058|1385-3793|CSP|HEALTH MAINTENANCE ORGAN|HMO
C0018720|T058|1385-3793|CSP|PREPAID GROUP HEALTH ORGAN|HMO
C0018720|T058|1385-3793|CSP|ORGANIZATIONS, HEALTH MAINTENANCE|HMO
C0018720|T058|1385-3793|CSP|PREPAID GROUP HEALTH ORGANIZATIONS|HMO
C0018720|T058|1385-3793|CSP|GROUP HEALTH ORGANIZATIONS, PREPAID|HMO
C0018720|T058|1385-3793|CSP|PREPAID HEALTHCARE ORGANIZATION|HMO
C0018720|T058|1385-3793|CSP|HEALTH MAINTENANCE ORGANISATION|HMO
C0018720|T058|1385-3793|CSP|HEALTH MAINTENANCE ORGANIZATION |HMO
C0018720|T058|1385-3793|CSP|PREPAID HEALTHCARE ORGANISATION|HMO
C0021684|T058||CSP|HEALTH INSURANCE REIMBURSEMENTS
C0021684|T058||CSP|INSURANCE REIMBURSEMENT, HEALTH
C0021684|T058||CSP|INSURANCE REIMBURSEMENTS, HEALTH
C0021684|T058||CSP|INSURANCE, HEALTH, REIMBURSEMENT
C0021684|T058||CSP|PAYMENT, THIRD-PARTY
C0021684|T058||CSP|PAYMENTS, THIRD-PARTY
C0021684|T058||CSP|REIMBURSEMENTS, HEALTH INSURANCE
C0021684|T058||CSP|THIRD PARTY PAYMENTS
C0021684|T058||CSP|THIRD-PARTY PAYMENT
C0021684|T058||CSP|HEALTH INSURANCE REIMBURSEMENT
C0021684|T058||CSP|THIRD-PARTY PAYMENTS
C0021684|T058||CSP|REIMBURSEMENT, HEALTH INSURANCE
C0021684|T058||CSP|THIRD PARTY PAYMENT
C0021694|T058||CSP|INSURANCE, PSYCHIATRIC
C0021694|T058||CSP|INSURANCES, PSYCHIATRIC
C0021694|T058||CSP|PSYCHIATRIC INSURANCE
C0021694|T058||CSP|PSYCHIATRIC INSURANCES
C0021694|T058||CSP|MENTAL HEALTH INSURANCE
C0025071|T058|1385-6531|CSP|MEDICAID|MEDICAID
C0025071|T058|1385-6531|CSP|MEDICAID PROGRAM|MEDICAID
C0025071|T058|1385-6531|CSP|MEDICAID COVERAGE |MEDICAID
C0025071|T058|1385-6531|CSP|MEDICAID COVERAGE|MEDICAID
C0042613|T058||CSP|CLAIM, VETERANS DISABILITY
C0042613|T058||CSP|CLAIMS, VETERANS DISABILITY
C0042613|T058||CSP|DISABILITY CLAIM, VETERANS
C0042613|T058||CSP|DISABILITY CLAIMS, VETERANS
C0042613|T058||CSP|VETERANS DISABILITY CLAIM
C0042613|T058||CSP|VETERANS DISABILITY CLAIMS
C0043233|T058||CSP|COMPENSATION, WORKMAN'S
C0043233|T058||CSP|COMPENSATION, WORKMEN'S
C0043233|T058||CSP|COMPENSATIONS, WORKMAN'S
C0043233|T058||CSP|COMPENSATIONS, WORKMEN'S
C0043233|T058||CSP|WORKMAN COMPENSATION
C0043233|T058||CSP|WORKMAN'S COMPENSATIONS
C0043233|T058||CSP|WORKMANS COMPENSATION
C0043233|T058||CSP|WORKMEN COMPENSATION
C0043233|T058||CSP|WORKMEN'S COMPENSATIONS
C0043233|T058||CSP|WORKMENS COMPENSATION
C0043233|T058||CSP|WORKERS' COMPENSATION
C0043233|T058||CSP|COMPENSATION, WORKER'S
C0043233|T058||CSP|COMPENSATION, WORKERS'
C0043233|T058||CSP|COMPENSATIONS, WORKER'S
C0043233|T058||CSP|COMPENSATIONS, WORKERS'
C0043233|T058||CSP|WORKER COMPENSATION
C0043233|T058||CSP|WORKER'S COMPENSATIONS
C0043233|T058||CSP|WORKERS COMPENSATION
C0043233|T058||CSP|WORKERS' COMPENSATIONS
C0043233|T058||CSP|WORKMEN'S COMPENSATION
C0043233|T058||CSP|WORKERS COMPENSATION PLAN
C0043233|T058||CSP|WORKER'S COMPENSATION
C0043233|T058||CSP|WORKMAN'S COMPENSATION
C0242816|T058||CSP|FEE FOR SERVICE PLANS
C0242816|T058||CSP|FEE FOR SERVICES
C0242816|T058||CSP|FEE-FOR-SERVICE PLAN
C0242816|T058||CSP|FEE-FOR-SERVICE PLANS
C0242816|T058||CSP|FEES FOR SERVICES
C0242816|T058||CSP|PLAN, FEE-FOR-SERVICE
C0242816|T058||CSP|PLANS, FEE-FOR-SERVICE
C0242816|T058||CSP|SERVICE, FEE FOR
C0242816|T058||CSP|SERVICE, FEES FOR
C0242816|T058||CSP|SERVICES, FEE FOR
C0242816|T058||CSP|SERVICES, FEES FOR
C0242816|T058||CSP|FEE SERV
C0242816|T058||CSP|FEE FOR SERVICE PAYMENT METHOD
C0242816|T058||CSP|FEE-FOR-SERVICE
C0242816|T058||CSP|FEE FOR SERVICE
C0242816|T058||CSP|FFS
C0242816|T058||CSP|FEES FOR SERVICE
C0242816|T058||CSP|FEE FOR SERVICE PAYMENT PLAN
C0681104|T058||CSP|EMPLOYEE HEALTH INSURANCE
C0086599|T058||CSP|MED ASSISTANCE TITLE 19
C0086599|T058||CSP|MEDICAL ASSISTANCE, TITLE 19
C0021680|T058||CSP|ACCIDENT INSURANCES
C0021680|T058||CSP|INSURANCE, ACCIDENT
C0021680|T058||CSP|INSURANCES, ACCIDENT
C0021680|T058||CSP|ACCIDENT INSURANCE
C0021685|T058||CSP|INSURANCE, HOSPITALIZATION
C0021685|T058||CSP|HOSPITALIZATION INSURANCE
C0024679|T058||CSP|MANAGED CARE PROGRAM
C0024679|T058||CSP|MANAGED CARE PROGRAMS
C0024679|T058||CSP|PROGRAM, MANAGED CARE
C0024679|T058||CSP|PROGRAMS, MANAGED CARE
C0024679|T058||CSP|MANAGED HEALTH CARE INSURANCE PLANS
C0085563|T058||CSP|HEALTH PLAN, PREPAID
C0085563|T058||CSP|PLAN, PREPAID HEALTH
C0085563|T058||CSP|PLANS, PREPAID HEALTH
C0085563|T058||CSP|PREPAID HEALTH PLAN
C0085563|T058||CSP|PREPAID HEALTH PLANS
C0085563|T058||CSP|HEALTH PLANS, PREPAID
C0282485|T058||CSP|MANAGED COMPETITION
C0282485|T058||CSP|COMPETITION, MANAGED
C0600593|T058|5004-0021|CSP|PUBLIC LAW 104 191|HEALTH INSURANCE PORTABILITY AND ACCOUNTABILITY ACT
C0600593|T058|5004-0021|CSP|PL 104 191|HEALTH INSURANCE PORTABILITY AND ACCOUNTABILITY ACT
C0600593|T058|5004-0021|CSP|KASSEBAUM KENNEDY ACT|HEALTH INSURANCE PORTABILITY AND ACCOUNTABILITY ACT
C0600593|T058|5004-0021|CSP|PL 104-191|HEALTH INSURANCE PORTABILITY AND ACCOUNTABILITY ACT
C0600593|T058|5004-0021|CSP|HIPAA|HEALTH INSURANCE PORTABILITY AND ACCOUNTABILITY ACT
C0600593|T058|5004-0021|CSP|PUBLIC LAW 104-191|HEALTH INSURANCE PORTABILITY AND ACCOUNTABILITY ACT
C0600593|T058|5004-0021|CSP|UNITED STATES HEALTH INSURANCE PORTABILITY AND ACCOUNTABILITY ACT|HEALTH INSURANCE PORTABILITY AND ACCOUNTABILITY ACT
C0600593|T058|5004-0021|CSP|HEALTH INSURANCE PORTABILITY AND ACCOUNTABILITY ACT|HEALTH INSURANCE PORTABILITY AND ACCOUNTABILITY ACT
C0600593|T058|5004-0021|CSP|PL104 191|HEALTH INSURANCE PORTABILITY AND ACCOUNTABILITY ACT
C0600593|T058|5004-0021|CSP|KENNEDY KASSEBAUM ACT|HEALTH INSURANCE PORTABILITY AND ACCOUNTABILITY ACT
C0600593|T058|5004-0021|CSP|PL104-191|HEALTH INSURANCE PORTABILITY AND ACCOUNTABILITY ACT
C0021682|T058||CSP|INSURANCE, HEALTH
C0021682|T058||CSP|HEALTH INSURANCE
C0018688|T058||CSP|HEALTH BENEFIT PLANS, EMPLOYEE
C0018688|T058||CSP|EMPLOYEE HEALTH BENEFIT PLANS
C0021688|T058||CSP|INSURANCE, LONG TERM CARE
C0021688|T058||CSP|INSURANCE, LONG-TERM CARE
C0021688|T058||CSP|LONG TERM CARE INSURANCE
C0021688|T058||CSP|LONG-TERM CARE INSURANCE
C0021690|T058||CSP|INSURANCE, NURSING SERVICES
C0021690|T058||CSP|INSURANCES, NURSING SERVICES
C0021690|T058||CSP|NURSING SERVICES INSURANCES
C0021690|T058||CSP|SERVICES INSURANCE, NURSING
C0021690|T058||CSP|SERVICES INSURANCES, NURSING
C0021690|T058||CSP|INSURANCE NURS SERV
C0021690|T058||CSP|NURS SERV INSURANCE
C0021690|T058||CSP|NURSING SERVICES INSURANCE
C0021691|T058||CSP|INSURANCE, PHARMACEUTICAL SERVICES
C0021691|T058||CSP|PHARM SERV INSURANCE
C0021691|T058||CSP|INSURANCE PHARM SERV
C0021691|T058||CSP|PHARMACEUTICAL SERVICES INSURANCE
C0021691|T058||CSP|INSURANCE, PHARMACY SERVICES
C0021691|T058||CSP|PHARMACY SERVICES INSURANCE
C0021691|T058||CSP|INSURANCE, PHARMACEUTIC SERVICES
C0021691|T058||CSP|PHARMACEUTIC SERVICES INSURANCE
C0085558|T058||CSP|INSURANCE, MEDIGAP
C0085558|T058||CSP|MEDIGAP POLICIES
C0085558|T058||CSP|POLICIES, MEDIGAP
C0085558|T058||CSP|POLICY, MEDIGAP
C0085558|T058||CSP|MEDIGAP INSURANCE
C0085558|T058||CSP|MEDIGAP POLICY
C0600588|T058||CSP|SAVINGS ACCOUNTS MED
C0600588|T058||CSP|ACCOUNTS MED SAVINGS
C0600588|T058||CSP|MED SAVINGS ACCOUNTS
C0600588|T058||CSP|ACCOUNT, MEDICAL SAVINGS
C0600588|T058||CSP|MEDICAL SAVINGS ACCOUNT
C0600588|T058||CSP|MEDICAL SAVINGS ACCOUNTS
C0600588|T058||CSP|SAVINGS ACCOUNT, MEDICAL
C0600588|T058||CSP|ACCOUNTS, MEDICAL SAVINGS
C0600588|T058||CSP|SAVINGS ACCOUNTS, MEDICAL
C0021689|T058||CSP|INSURANCE, MAJOR MEDICAL
C0021689|T058||CSP|INSURANCE MAJOR MED
C0021689|T058||CSP|MAJOR MED INSURANCE
C0021689|T058||CSP|MED INSURANCE MAJOR
C0021689|T058||CSP|MEDICAL INSURANCE, MAJOR
C0021689|T058||CSP|MAJOR MEDICAL INSURANCE
C0021693|T058||CSP|INSURANCE, PHYSICIAN SERVICES
C0021693|T058||CSP|INSURANCES, PHYSICIAN SERVICES
C0021693|T058||CSP|PHYSICIAN SERVICES INSURANCE
C0021693|T058||CSP|PHYSICIAN SERVICES INSURANCES
C0021693|T058||CSP|SERVICES INSURANCES, PHYSICIAN
C0021693|T058||CSP|INSURANCE PHYSICIAN SERVICE
C0021693|T058||CSP|INSURANCE PHYSICIAN SERVICES
C0021693|T058||CSP|PHYSICIAN SERVICE, INSURANCE
C0021693|T058||CSP|SERVICE, INSURANCE PHYSICIAN
C0021693|T058||CSP|SERVICES, INSURANCE PHYSICIAN
C0021693|T058||CSP|INSURANCE PHYSICIAN SERV
C0021693|T058||CSP|SERV INSURANCE PHYSICIAN
C0021693|T058||CSP|PHYSICIAN SERV INSURANCE
C0021693|T058||CSP|SERVICES INSURANCE, PHYSICIAN
C0021693|T058||CSP|PHYSICIAN SERVICES, INSURANCE
C0021695|T058||CSP|INSURANCE, SURGICAL
C0021695|T058||CSP|INSURANCES, SURGICAL
C0021695|T058||CSP|SURGICAL INSURANCES
C0021695|T058||CSP|INSURANCE SURG
C0021695|T058||CSP|SURG INSURANCE
C0021695|T058||CSP|SURGICAL INSURANCE
C0027454|T058||CSP|NATIONAL HEALTH INSURANCE, UNITED STATES
C0027454|T058||CSP|NATL HEALTH INSUR US
C0027454|T058||CSP|NATIONAL HEALTH INSURANCE--UNITED STATES
C0027454|T058||CSP|UNITED STATES NATIONAL HEALTH INSURANCE
C0027454|T058||CSP|FEDERAL HEALTH INSURANCE PLANS, UNITED STATES
C0282487|T058||CSP|SINGLE PAYER SYSTEM
C0282487|T058||CSP|SINGLE-PAYER SYSTEM
C0282487|T058||CSP|SINGLE-PAYER SYSTEMS
C0282487|T058||CSP|SYSTEM, SINGLE-PAYER
C0282487|T058||CSP|SYSTEMS, SINGLE-PAYER
C0018256|T058||CSP|HEALTH INSURANCE, GROUP
C0018256|T058||CSP|INSURANCE, GROUP HEALTH
C0018256|T058||CSP|GROUP HEALTH INSURANCE
C0018718|T058||CSP|INSURANCE, VOLUNTARY HEALTH
C0018718|T058||CSP|VOLUNTARY HEALTH INSURANCE
C0018718|T058||CSP|HEALTH INSURANCE, VOLUNTARY
C2936611|T058||CSP|PL111 148
C2936611|T058||CSP|111-148, PL
C2936611|T058||CSP|PUBLIC LAW 111 148
C2936611|T058||CSP|PATIENT PROTECTION AND AFFORDABLE CARE ACT
C2936611|T058||CSP|PL 111 148
C2936611|T058||CSP|CARE ACT, AFFORDABLE (ACA)
C2936611|T058||CSP|ACTS, AFFORDABLE CARE (ACA)
C2936611|T058||CSP|CARE ACT, AFFORDABLE
C2936611|T058||CSP|ACTS, AFFORDABLE CARE
C2936611|T058||CSP|ACT, AFFORDABLE CARE
C2936611|T058||CSP|AFFORDABLE CARE ACTS
C2936611|T058||CSP|CARE ACTS, AFFORDABLE
C2936611|T058||CSP|AFFORDABLE CARE ACT
C2936611|T058||CSP|PL 111-148
C2936611|T058||CSP|OBAMACARE
C2936611|T058||CSP|PUBLIC LAW 111-148
C2936611|T058||CSP|AFFORDABLE CARE ACT (ACA)
C2936611|T058||CSP|HEALTH CARE REFORM ACT
C2936611|T058||CSP|PL111-148
C2936638|T058||CSP|FOR PROFIT INSURANCE PLANS
C2936638|T058||CSP|INSURANCE PLANS, FOR-PROFIT
C2936638|T058||CSP|INSURANCE PLAN, FOR-PROFIT
C2936638|T058||CSP|FOR-PROFIT INSURANCE PLAN
C2936638|T058||CSP|PLANS, FOR-PROFIT INSURANCE
C2936638|T058||CSP|FOR-PROFIT INSURANCE PLANS
C2936639|T058||CSP|PLANS, NOT-FOR-PROFIT INSURANCE
C2936639|T058||CSP|NOT-FOR-PROFIT INSURANCE PLAN
C2936639|T058||CSP|NOT-FOR-PROFIT INSURANCE PLANS
C2936639|T058||CSP|INSURANCE PLAN, NOT-FOR-PROFIT
C2936639|T058||CSP|INSURANCE PLANS, NOT-FOR-PROFIT
C2936639|T058||CSP|PLAN, NOT-FOR-PROFIT INSURANCE
C2936639|T058||CSP|NOT FOR PROFIT INSURANCE PLANS
C2347682|T058||CSP|PRIVATE HEALTH INSURANCE
C2347682|T058||CSP|HEALTH INSURANCE
C3494321|T058||CSP|PURCHASINGS, VALUE-BASED
C3494321|T058||CSP|VALUE-BASED PURCHASING
C3494321|T058||CSP|VALUE BASED PURCHASING
C3494321|T058||CSP|VALUE-BASED PURCHASINGS
C3494321|T058||CSP|PURCHASING, VALUE-BASED
C4042889|T058||CSP|CHILDREN'S HEALTH INSURANCE PROGRAM
C0079817|T058||CSP|MEDICARE PART A
C0079817|T058||CSP|PART A, MEDICARE
C0079817|T058||CSP|MEDICARE HOSP INSURANCE PROGRAM
C0079817|T058||CSP|MEDICARE A
C0079817|T058||CSP|HOSP INSURANCE PROGRAM MEDICARE
C0079817|T058||CSP|HOSPITAL INSURANCE PROGRAM, MEDICARE
C0079817|T058||CSP|MEDICARE HOSPITAL INSURANCE PROGRAM
C0079818|T058||CSP|MEDICARE PART B
C0079818|T058||CSP|PART B, MEDICARE
C0079818|T058||CSP|PROGRAM, SMI
C0079818|T058||CSP|PROGRAMS, SMI
C0079818|T058||CSP|SMI PROGRAMS
C0079818|T058||CSP|MEDICARE SUPPLEMENTARY MED INSURANCE PROGRAM
C0079818|T058||CSP|MEDICARE B
C0079818|T058||CSP|SUPPLEMENTARY MED INSURANCE PROGRAM MEDICARE
C0079818|T058||CSP|SUPPLEMENTARY MEDICAL INSURANCE PROGRAM, MEDICARE
C0079818|T058||CSP|SMI PROGRAM
C0079818|T058||CSP|MEDICARE SUPPLEMENTARY MEDICAL INSURANCE PROGRAM
C0025114|T058||CSP|ASSIGNMENT, MEDICARE
C0025114|T058||CSP|ASSIGNMENTS, MEDICARE
C0025114|T058||CSP|MEDICARE ASSIGNMENT
C0025114|T058||CSP|MEDICARE ASSIGNMENTS
C0600580|T058||CSP|MEDICARE C
C0600580|T058||CSP|MEDICARE PART C
C0600580|T058||CSP|PART C, MEDICARE
C0600580|T058||CSP|CHOICE, MEDICARE PLUS
C0600580|T058||CSP|PLUS CHOICE, MEDICARE
C0600580|T058||CSP|PROGRAMS, MEDICARE+CHOICE (US)
C0600580|T058||CSP|MEDICARE+CHOICE PROGRAMS (US)
C0600580|T058||CSP|PROGRAM, MEDICARE+CHOICE (US)
C0600580|T058||CSP|MEDICARE+CHOICE PROGRAM (US)
C0600580|T058||CSP|MEDICARE PLUS CHOICE PROGRAM (US)
C0600580|T058||CSP|MEDICARE CHOICE
C0600580|T058||CSP|MEDICARE PLUS CHOICE
C1955953|T058||CSP|MEDICARE PART D
C1955953|T058||CSP|PART D, MEDICARE
C3530305|T058||CSP|MEDICARE (MANAGED CARE)
C3530300|T058||CSP|MEDICARE (NON-MANAGED CARE)
C3530295|T058||CSP|MEDICARE OTHER
C3530238|T058||CSP|MANAGED CARE (PRIVATE)
C3530234|T058||CSP|PRIVATE HEALTH INSURANCE - INDEMNITY
C3530229|T058||CSP|MANAGED CARE (PRIVATE) OR PRIVATE HEALTH INSURANCE (INDEMNITY), NOT OTHERWISE SPECIFIED
C3530228|T058||CSP|ORGANIZED DELIVERY SYSTEM
C3530227|T058||CSP|SMALL EMPLOYER PURCHASING GROUP
C3530226|T058||CSP|OTHER PRIVATE INSURANCE
C1955981|T058||CSP|BLUE CROSS BLUE SHIELD INSURANCE PLANS
C1955981|T058||CSP|BLUE CROSS/BLUE SHIELD
C0005864|T058||CSP|BLUE CROSS
C0005864|T058||CSP|BLUE CROSSES
C0005864|T058||CSP|CROSS, BLUE
C0005864|T058||CSP|CROSSES, BLUE
C0005865|T058||CSP|SHIELDS, BLUE
C0005865|T058||CSP|SHIELD, BLUE
C0005865|T058||CSP|BLUE SHIELD
C0005865|T058||CSP|BLUE SHIELDS
C3530225|T058||CSP|BC MANAGED CARE
C3530220|T058||CSP|BC INDEMNITY
C3530219|T058||CSP|BC (INDEMNITY OR MANAGED CARE) - OUT OF STATE
C3530218|T058||CSP|BC (INDEMNITY OR MANAGED CARE) - UNSPECIFIED
C3530217|T058||CSP|BC (INDEMNITY OR MANAGED CARE) - OTHER
