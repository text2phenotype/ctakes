C0809969|T047|33|CCS_10|CANCER OF KIDNEY AND RENAL PELVIS|CANCER OF KIDNEY AND RENAL PELVIS
C0809971|T047|35|CCS_10|CANCER OF BRAIN AND NERVOUS SYSTEM|CANCER OF BRAIN AND NERVOUS SYSTEM
C0809972|T047|41|CCS_10|CANCER; OTHER AND UNSPECIFIED PRIMARY|CANCER; OTHER AND UNSPECIFIED PRIMARY
C0810239|T047|2.7|CCS_10|CANCER OF OVARY AND OTHER FEMALE GENITAL ORGANS|CANCER OF OVARY AND OTHER FEMALE GENITAL ORGANS
C0810243|T047|2.11|CCS_10|CANCER; OTHER PRIMARY|CANCER; OTHER PRIMARY
C1140680|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY
C4048328|T047||CCS_10|CERVICAL CANCER
C4048331|T047|2.3|CCS_10|CANCER OF BRONCHUS; LUNG|CANCER OF BRONCHUS; LUNG
C0005684|T047||CCS_10|MALIGNANT NEOPLASM OF URINARY BLADDER
C0006142|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST
C0007102|T047||CCS_10|MALIGNANT TUMOR OF COLON
C0007114|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN
C0007115|T047||CCS_10|MALIGNANT NEOPLASM OF THYROID
C0153448|T047|16|CCS_10|MALIGNANT NEOPLASM OF LIVER AND INTRAHEPATIC BILE DUCTS|CANCER OF LIVER AND INTRAHEPATIC BILE DUCT
C0153567|T047||CCS_10|UTERINE CANCER
C0153594|T047||CCS_10|MALIGNANT NEOPLASM OF TESTIS
C0153606|T047|2.8|CCS_10|MALIGNANT TUMOR OF MALE GENITAL ORGAN|CANCER OF MALE GENITAL ORGANS
C0278996|T047||CCS_10|CANCER OF HEAD AND NECK
C0346647|T047||CCS_10|MALIGNANT NEOPLASM OF PANCREAS
C0346890|T047|34|CCS_10|MALIGNANT NEOPLASM OF OTHER AND UNSPECIFIED URINARY ORGANS|CANCER OF OTHER URINARY ORGANS
C0348371|T047||CCS_10|MALIGNANT NEOPLASM OF URINARY ORGAN, UNSPECIFIED
C0348393|T047|2.10|CCS_10|MALIGNANT TUMOR OF LYMPHOID HEMOPOIETIC AND RELATED TISSUE|CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0376358|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE
C0392920|T047||CCS_10|CHEMOTHERAPY REGIMEN
C0497581|T047|31|CCS_10|OTHER MALE GENITAL MALIGNANT NEOPLASM|CANCER OF OTHER MALE GENITAL ORGANS
C0546837|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS
C0699791|T047||CCS_10|STOMACH CARCINOMA
C0740458|T047||CCS_10|CANCER OF UTERUS AND CERVIX
C0809960|T047|15|CCS_10|CANCER OF RECTUM AND ANUS|CANCER OF RECTUM AND ANUS
C0809962|T047|18|CCS_10|CANCER OF OTHER GI ORGANS; PERITONEUM|CANCER OF OTHER GI ORGANS; PERITONEUM
C0809964|T047|20|CCS_10|CANCER; OTHER RESPIRATORY AND INTRATHORACIC|CANCER; OTHER RESPIRATORY AND INTRATHORACIC
C0809965|T047|21|CCS_10|CANCER OF BONE AND CONNECTIVE TISSUE|CANCER OF BONE AND CONNECTIVE TISSUE
C0809967|T047|28|CCS_10|CANCER OF OTHER FEMALE GENITAL ORGANS|CANCER OF OTHER FEMALE GENITAL ORGANS
C0809969|T047|33|CCS_10|CANCER OF KIDNEY AND RENAL PELVIS|CANCER OF KIDNEY AND RENAL PELVIS
C0809971|T047|35|CCS_10|CANCER OF BRAIN AND NERVOUS SYSTEM|CANCER OF BRAIN AND NERVOUS SYSTEM
C0809972|T047|41|CCS_10|CANCER; OTHER AND UNSPECIFIED PRIMARY|CANCER; OTHER AND UNSPECIFIED PRIMARY
C1140680|T047||CCS_10|CANCER, OVARIAN
C1140680|T047||CCS_10|CANCERS, OVARIAN
C1140680|T047||CCS_10|OVARIAN CANCERS
C1140680|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY
C1140680|T047||CCS_10|OVARIAN CANCER
C1140680|T047||CCS_10|CANCER OF OVARY
C1140680|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY 
C1140680|T047||CCS_10|OVARIAN CANCER 
C1140680|T047||CCS_10|CA OVARY
C1140680|T047||CCS_10|CANCERS, OVARY
C1140680|T047||CCS_10|OVARY CANCERS
C1140680|T047||CCS_10|MALIGNANT TUMOR OF OVARY
C1140680|T047||CCS_10|MALIGN NEOPL OVARY
C1140680|T047||CCS_10|CANCER, OVARY
C1140680|T047||CCS_10|MALIGNANT TUMOUR OF OVARY
C1140680|T047||CCS_10|MALIGNANT TUMOUR OF OVARY 
C1140680|T047||CCS_10|OVARIES--CANCER
C1140680|T047||CCS_10|OVARIAN CANCER, NOS
C1140680|T047||CCS_10|-- OVARIAN CANCER
C1140680|T047||CCS_10|OVARIAN CA
C1140680|T047||CCS_10|OVARIAN CANCER NOS
C1140680|T047||CCS_10|CANCER OF THE OVARY
C1140680|T047||CCS_10|OVARY CANCER
C1140680|T047||CCS_10|CA - CANCER OF OVARY
C1140680|T047||CCS_10|MALIGNANT TUMOR OF OVARY 
C1140680|T047||CCS_10|MALIGNANT NEOPLASM OF THE OVARY
C1140680|T047||CCS_10|MALIGNANT OVARIAN NEOPLASM
C1140680|T047||CCS_10|MALIGNANT OVARIAN TUMOR
C1140680|T047||CCS_10|MALIGNANT TUMOR OF THE OVARY
C0809967|T047|28|CCS_10|CANCER OF OTHER FEMALE GENITAL ORGANS|CANCER OF OTHER FEMALE GENITAL ORGANS
C0809965|T047|21|CCS_10|CANCER OF BONE AND CONNECTIVE TISSUE|CANCER OF BONE AND CONNECTIVE TISSUE
C0278996|T047||CCS_10|MALIGNANT TUMOR OF HEAD AND NECK 
C0278996|T047||CCS_10|MALIGNANT TUMOR OF HEAD AND/OR NECK 
C0278996|T047||CCS_10|HEAD AND NECK CANCER
C0278996|T047||CCS_10|MALIGNANT TUMOUR OF HEAD AND/OR NECK
C0278996|T047||CCS_10|MALIGNANT TUMOR OF HEAD AND/OR NECK
C0278996|T047||CCS_10|CANCER OF HEAD AND NECK
C0278996|T047||CCS_10|MALIGNANT NEOPLASM OF HEAD AND/OR NECK 
C0278996|T047||CCS_10|MALIGNANT NEOPLASM OF HEAD AND/OR NECK
C0278996|T047||CCS_10|HEAD AND NECK CANCER, NOS
C0278996|T047||CCS_10|CANCER OF THE HEAD AND NECK
C0278996|T047||CCS_10|MALIGNANT TUMOR OF HEAD AND NECK
C0278996|T047||CCS_10|MALIGNANT TUMOUR OF HEAD AND NECK
C0278996|T047||CCS_10|MALIGNANT HEAD AND NECK NEOPLASM
C0278996|T047||CCS_10|MALIGNANT HEAD AND NECK TUMOR
C0278996|T047||CCS_10|MALIGNANT NEOPLASM OF HEAD AND NECK
C0278996|T047||CCS_10|MALIGNANT NEOPLASM OF THE HEAD AND NECK
C0278996|T047||CCS_10|MALIGNANT TUMOR OF THE HEAD AND NECK
C0007115|T047||CCS_10|MALIGNANT NEOPLASM OF THYROID GLAND
C0007115|T047||CCS_10|MALIGNANT THYROID GLAND NEOPLASM
C0007115|T047||CCS_10|MALIGNANT THYROID NEOPLASM
C0007115|T047||CCS_10|THYROID CANCER
C0007115|T047||CCS_10|MALIGNANT NEOPLASM OF THYROID GLAND 
C0007115|T047||CCS_10|THYROID NEOPLASMS MALIGNANT
C0007115|T047||CCS_10|MALIGNANT TUMOR OF THYROID GLAND
C0007115|T047||CCS_10|MALIGN NEOPL THYROID
C0007115|T047||CCS_10|CANCER OF THYROID
C0007115|T047||CCS_10|MALIGNANT TUMOUR OF THYROID GLAND
C0007115|T047||CCS_10|MALIGNANT TUMOUR OF THYROID GLAND 
C0007115|T047||CCS_10|-- THYROID CANCER
C0007115|T047||CCS_10|THYROID NEOPLASM MALIGNANT
C0007115|T047||CCS_10|THYROID GLAND CANCER
C0007115|T047||CCS_10|THYROID CA
C0007115|T047||CCS_10|MALIGNANT TUMOR OF THYROID GLAND 
C0007115|T047||CCS_10|MALIGNANT NEOPLASM OF THYROID
C0007115|T047||CCS_10|MALIGNANT NEOPLASM OF THE THYROID GLAND
C0007115|T047||CCS_10|MALIGNANT NEOPLASM OF THE THYROID
C0007115|T047||CCS_10|MALIGNANT THYROID GLAND TUMOR
C0007115|T047||CCS_10|MALIGNANT THYROID TUMOR
C0007115|T047||CCS_10|MALIGNANT TUMOR OF THYROID
C0007115|T047||CCS_10|MALIGNANT TUMOR OF THE THYROID GLAND
C0007115|T047||CCS_10|MALIGNANT TUMOR OF THE THYROID
C0007115|T047||CCS_10|NEOPLASM MALIG;THYROID GLAND
C0007115|T047||CCS_10|MALIGNANT NEOSPLASM OF THE THYROID GLAND
C0809964|T047|20|CCS_10|CANCER; OTHER RESPIRATORY AND INTRATHORACIC|CANCER; OTHER RESPIRATORY AND INTRATHORACIC
C0948216|T047||CCS_10|ADENOCARCINOMA OF OVARY 
C0948216|T047||CCS_10|ADENOCARCINOMA OF OVARY
C0948216|T047||CCS_10|OVARIAN ADENOCARCINOMA
C0948216|T047||CCS_10|ADENOCARCINOMA OF THE OVARY
C0334495|T047||CCS_10|MALIGNANT BRENNER TUMOR OF OVARY 
C0334495|T047||CCS_10|MALIGNANT BRENNER TUMOR OF OVARY
C0334495|T047||CCS_10|MALIGNANT BRENNER TUMOR
C0334495|T047||CCS_10|BRENNER TUMOR, MALIGNANT
C0334495|T047||CCS_10|MALIGNANT BRENNER TUMOUR
C0334495|T047||CCS_10|BRENNER TUMOUR, MALIGNANT
C0334495|T047||CCS_10|BRENNER TUMOR, MALIGNANT (MORPHOLOGIC ABNORMALITY)
C0334495|T047||CCS_10|BRENNER; TUMOR, MALIGNANT
C0334495|T047||CCS_10|TUMOR; BRENNER, MALIGNANT
C0334495|T047||CCS_10|MALIGNANT BRENNER TUMOR OF THE OVARY
C0334495|T047||CCS_10|MALIGNANT OVARIAN BRENNER TUMOR
C1297991|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM ENDOMETRIUM
C1297991|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM ENDOMETRIUM 
C1297991|T047||CCS_10|OVARIAN NEOPLASM LEFT BY DIRECT EXTENSION FROM ENDOMETRIUM
C1297991|T047||CCS_10|MALIGNANT TUMOR INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM ENDOMETRIUM 
C1297991|T047||CCS_10|MALIGNANT TUMOR INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM ENDOMETRIUM
C1297991|T047||CCS_10|MALIGNANT TUMOUR INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM ENDOMETRIUM
C1297992|T047||CCS_10|MALIGNANT TUMOR INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM FALLOPIAN TUBE 
C1297992|T047||CCS_10|MALIGNANT TUMOR INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM FALLOPIAN TUBE
C1297992|T047||CCS_10|MALIGNANT TUMOUR INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM FALLOPIAN TUBE
C1297993|T047||CCS_10|MALIGNANT TUMOR INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM RIGHT OVARY 
C1297993|T047||CCS_10|MALIGNANT TUMOR INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM RIGHT OVARY
C1297993|T047||CCS_10|MALIGNANT TUMOUR INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM RIGHT OVARY
C1297994|T047||CCS_10|MALIGNANT TUMOR INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM UTERINE CERVIX 
C1297994|T047||CCS_10|MALIGNANT TUMOR INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM UTERINE CERVIX
C1297994|T047||CCS_10|MALIGNANT TUMOUR INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM UTERINE CERVIX
C1297995|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM UTERUS
C1297995|T047||CCS_10|OVARIAN NEOPLASM LEFT BY DIRECT EXTENSION FROM UTERUS
C1297995|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM UTERUS 
C1297995|T047||CCS_10|MALIGNANT TUMOR INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM UTERUS 
C1297995|T047||CCS_10|MALIGNANT TUMOR INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM UTERUS
C1297995|T047||CCS_10|MALIGNANT TUMOUR INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM UTERUS
C1297998|T047||CCS_10|MALIGNANT TUMOR INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM ENDOMETRIUM 
C1297998|T047||CCS_10|MALIGNANT TUMOR INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM ENDOMETRIUM
C1297998|T047||CCS_10|MALIGNANT TUMOUR INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM ENDOMETRIUM
C1297999|T047||CCS_10|OVARIAN NEOPLASM RIGHT BY DIRECT EXTENSION FROM FALLOPIAN TUBE
C1297999|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM FALLOPIAN TUBE 
C1297999|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM FALLOPIAN TUBE
C1297999|T047||CCS_10|MALIGNANT TUMOR INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM FALLOPIAN TUBE 
C1297999|T047||CCS_10|MALIGNANT TUMOR INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM FALLOPIAN TUBE
C1297999|T047||CCS_10|MALIGNANT TUMOUR INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM FALLOPIAN TUBE
C1298000|T047||CCS_10|MALIGNANT TUMOR INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM LEFT OVARY 
C1298000|T047||CCS_10|MALIGNANT TUMOR INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM LEFT OVARY
C1298000|T047||CCS_10|MALIGNANT TUMOUR INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM LEFT OVARY
C1298001|T047||CCS_10|OVARIAN NEOPLASM RIGHT BY DIRECT EXTENSION FROM UTERINE CERVIX
C1298001|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM UTERINE CERVIX 
C1298001|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM UTERINE CERVIX
C1298001|T047||CCS_10|MALIGNANT TUMOR INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM UTERINE CERVIX 
C1298001|T047||CCS_10|MALIGNANT TUMOR INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM UTERINE CERVIX
C1298001|T047||CCS_10|MALIGNANT TUMOUR INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM UTERINE CERVIX
C1298026|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM VAGINA 
C1298026|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM VAGINA
C1298026|T047||CCS_10|OVARIAN NEOPLASM LEFT BY DIRECT EXTENSION FROM VAGINA
C1298026|T047||CCS_10|MALIGNANT TUMOR INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM VAGINA 
C1298026|T047||CCS_10|MALIGNANT TUMOR INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM VAGINA
C1298026|T047||CCS_10|MALIGNANT TUMOUR INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM VAGINA
C1298033|T047||CCS_10|MALIGNANT TUMOR INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM UTERUS 
C1298033|T047||CCS_10|MALIGNANT TUMOR INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM UTERUS
C1298033|T047||CCS_10|MALIGNANT TUMOUR INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM UTERUS
C1298034|T047||CCS_10|MALIGNANT TUMOR INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM VAGINA 
C1298034|T047||CCS_10|MALIGNANT TUMOR INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM VAGINA
C1298034|T047||CCS_10|MALIGNANT TUMOUR INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM VAGINA
C0346182|T047||CCS_10|MALIGNANT TERATOMA OF OVARY 
C0346182|T047||CCS_10|MALIGNANT TERATOMA OF OVARY
C0346182|T047||CCS_10|IMMATURE TERATOMA OF OVARY
C0346182|T047||CCS_10|IMMATURE TERATOMA OF OVARY 
C0346182|T047||CCS_10|OVARIAN NEOPLASM MALIGNANT IMMATURE TERATOMA
C0346182|T047||CCS_10|IMMATURE TERATOMA OF OVARY 
C0346182|T047||CCS_10|OVARIAN GERM CELL IMMATURE TERATOMA
C0346182|T047||CCS_10|IMMATURE TERATOMA, OVARIAN GERM CELL
C0346182|T047||CCS_10|TERATOMA, IMMATURE, OVARIAN GERM CELL
C0346182|T047||CCS_10|IMMATURE GERM CELL TERATOMA OF OVARY
C0346182|T047||CCS_10|IMMATURE GERM CELL TERATOMA OF THE OVARY
C0346182|T047||CCS_10|IMMATURE OVARIAN TERATOMA
C0346182|T047||CCS_10|IMMATURE TERATOMA OF THE OVARY
C0346182|T047||CCS_10|MALIGNANT GERM CELL TERATOMA OF OVARY
C0346182|T047||CCS_10|MALIGNANT GERM CELL TERATOMA OF THE OVARY
C0346182|T047||CCS_10|MALIGNANT OVARIAN GERM CELL TERATOMA
C0346182|T047||CCS_10|MALIGNANT OVARIAN TERATOMA
C0346182|T047||CCS_10|MALIGNANT TERATOMA OF THE OVARY
C0346182|T047||CCS_10|OVARIAN IMMATURE GERM CELL TERATOMA
C0346182|T047||CCS_10|OVARIAN IMMATURE TERATOMA
C2842146|T047||CCS_10|MALIGNANT NEOPLASM OF RIGHT OVARY
C2842147|T047||CCS_10|MALIGNANT NEOPLASM OF UNSPECIFIED OVARY
C2016058|T047||CCS_10|CARCINOMA SIMPLEX OF OVARY 
C2016058|T047||CCS_10|CARCINOMA SIMPLEX OF OVARY
C2212041|T047||CCS_10|ADENOCARCINOID TUMOR OF OVARY
C2212041|T047||CCS_10|ADENOCARCINOID TUMOR OF OVARY 
C0392998|T047||CCS_10|CARCINOSARCOMA OF OVARY
C0392998|T047||CCS_10|CARCINOSARCOMA OF OVARY 
C0392998|T047||CCS_10|CARCINOSARCOMA OF OVARY 
C0392998|T047||CCS_10|OVARIAN CARCINOSARCOMA
C0392998|T047||CCS_10|MALIGNANT MIXED MESODERMAL MÜLLERIAN NEOPLASM OF OVARY
C0392998|T047||CCS_10|OVARIAN MALIGNANT MIXED MÜLLERIAN TUMOR
C0392998|T047||CCS_10|MALIGNANT MIXED MESODERMAL MÜLLERIAN TUMOR OF THE OVARY
C0392998|T047||CCS_10|OVARIAN MALIGNANT MIXED MÜLLERIAN NEOPLASM
C0392998|T047||CCS_10|MALIGNANT MIXED MESODERMAL MÜLLERIAN NEOPLASM OF THE OVARY
C0392998|T047||CCS_10|OVARIAN MALIGNANT MIXED MESODERMAL MÜLLERIAN TUMOR
C0392998|T047||CCS_10|MALIGNANT MIXED MESODERMAL MÜLLERIAN TUMOR OF OVARY
C0392998|T047||CCS_10|OVARIAN MALIGNANT MIXED MESODERMAL MÜLLERIAN NEOPLASM
C0392998|T047||CCS_10|OVARIAN MALIGNANT MIXED MESODERMAL (MÜLLERIAN) TUMOR
C0392998|T047||CCS_10|OVARIAN MALIGNANT MESODERMAL (MÜLLERIAN) MIXED TUMOR
C0392998|T047||CCS_10|MULLERIAN SARCOMA, OVARIAN MALIGNANT MIXED MESODERMAL
C0392998|T047||CCS_10|MULLERIAN TUMOR, OVARIAN MALIGNANT MIXED MESODERMAL
C0392998|T047||CCS_10|CARCINOSARCOMA, OVARIAN
C0392998|T047||CCS_10|MALIGNANT MIXED MESODERMAL MULLERIAN TUMOR, OVARIAN
C0392998|T047||CCS_10|OVARIAN MMMT
C0392998|T047||CCS_10|CARCINOSARCOMA OF THE OVARY
C2212004|T047||CCS_10|MALIGNANT SMALL CELL NEOPLASM OF OVARY 
C2212004|T047||CCS_10|OVARIAN NEOPLASM MALIGNANT SMALL CELL TYPE
C2212004|T047||CCS_10|MALIGNANT SMALL CELL NEOPLASM OF OVARY
C2011392|T047||CCS_10|GIANT CELL TYPE NEOPLASM OF OVARY 
C2011392|T047||CCS_10|OVARIAN NEOPLASM MALIGNANT GIANT CELL TYPE
C2011392|T047||CCS_10|GIANT CELL TYPE NEOPLASM OF OVARY
C2018675|T047||CCS_10|SPINDLE CELL TYPE NEOPLASM OF OVARY 
C2018675|T047||CCS_10|SPINDLE CELL TYPE NEOPLASM OF OVARY
C2018675|T047||CCS_10|OVARIAN NEOPLASM MALIGNANT SPINDLE CELL TYPE
C2075635|T047||CCS_10|OVARIAN NEOPLASM MALIGNANT CLEAR CELL TYPE
C2075635|T047||CCS_10|MALIGNANT CLEAR CELL TYPE NEOPLASM OF THE OVARY 
C2075635|T047||CCS_10|MALIGNANT CLEAR CELL TYPE NEOPLASM OF THE OVARY
C2075635|T047||CCS_10|CLEAR CELL TYPE NEOPLASM OF OVARY
C0029925|T047||CCS_10|OVARIAN CARCINOMA
C0029925|T047||CCS_10|CARCINOMA OF OVARY 
C0029925|T047||CCS_10|CARCINOMA OF OVARY
C2212016|T047||CCS_10|MALIGNANT EPITHELIOID TROPHOBLASTIC TUMOR OF OVARY
C2212016|T047||CCS_10|MALIGNANT EPITHELIOID TROPHOBLASTIC TUMOR OF OVARY 
C0334525|T047||CCS_10|MALIGNANT STRUMA OVARII
C0334525|T047||CCS_10|MALIGNANT STRUMA OVARII 
C0334525|T047||CCS_10|STRUMA OVARII, MALIGNANT
C0334525|T047||CCS_10|STRUMA OVARII, MALIGNANT (MORPHOLOGIC ABNORMALITY)
C0334525|T047||CCS_10|STRUMA; OVARII, MALIGNANT
C0280746|T047||CCS_10|SARCOMA OF OVARY
C0280746|T047||CCS_10|SARCOMA OF OVARY 
C0280746|T047||CCS_10|SARCOMA OF OVARY 
C0280746|T047||CCS_10|OVARIAN SARCOMA
C0280746|T047||CCS_10|SARCOMA OF THE OVARY
C0280746|T047||CCS_10|SARCOMA, OVARIAN
C1335161|T047||CCS_10|FIBROSARCOMA OF OVARY 
C1335161|T047||CCS_10|FIBROSARCOMA OF OVARY
C1335161|T047||CCS_10|FIBROSARCOMA OF THE OVARY
C1335161|T047||CCS_10|OVARIAN FIBROSARCOMA
C2212040|T047||CCS_10|MYOSARCOMA OF OVARY 
C2212040|T047||CCS_10|MYOSARCOMA OF OVARY
C2212048|T047||CCS_10|MALIGNANT GONADAL NEOPLASM OF OVARY 
C2212048|T047||CCS_10|MALIGNANT GONADAL NEOPLASM OF OVARY
C2212049|T047||CCS_10|MALIGNANT MESONEPHROMA OF OVARY 
C2212049|T047||CCS_10|MALIGNANT MESONEPHROMA OF OVARY
C2212050|T047||CCS_10|MALIGNANT LYMPHOMA OF OVARY
C2212050|T047||CCS_10|MALIGNANT LYMPHOMA OF OVARY 
C2212053|T047||CCS_10|MALIGNANT PLASMACYTOMA OF OVARY
C2212053|T047||CCS_10|MALIGNANT PLASMACYTOMA OF OVARY 
C2212055|T047||CCS_10|MALIGNANT MASTOCYTOSIS OF OVARY 
C2212055|T047||CCS_10|MALIGNANT MASTOCYTOSIS OF OVARY
C2212056|T047||CCS_10|MULLERIAN MIXED TUMOR OF OVARY 
C2212056|T047||CCS_10|MULLERIAN MIXED TUMOR OF OVARY
C2212057|T047||CCS_10|MALIGNANT MESODERMAL MIXED TUMOR OF OVARY 
C2212057|T047||CCS_10|MALIGNANT MESODERMAL MIXED TUMOR OF OVARY
C2212058|T047||CCS_10|ADENOCARCINOFIBROMA OF OVARY
C2212058|T047||CCS_10|ADENOCARCINOFIBROMA OF OVARY 
C2217304|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGING
C2217304|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGING 
C2217304|T047||CCS_10|MALIGNANT OVARIAN NEOPLASM STAGING
C2217304|T047||CCS_10|MALIGNANT TUMOR OF OVARY STAGING
C2217304|T047||CCS_10|OVARIAN CANCER STAGING
C0346181|T047||CCS_10|CHORIOCARCINOMA OF OVARY 
C0346181|T047||CCS_10|CHORIOCARCINOMA OF OVARY
C0346181|T047||CCS_10|OVARIAN GERM CELL CHORIOCARCINOMA
C0346181|T047||CCS_10|CHORIOCARCINOMA OF OVARY 
C0346181|T047||CCS_10|CHORIOCARCINOMA, OVARIAN GERM CELL
C0346181|T047||CCS_10|CHORIOCARCINOMA OF THE OVARY
C0346181|T047||CCS_10|GERM CELL CHORIOCARCINOMA OF OVARY
C0346181|T047||CCS_10|GERM CELL CHORIOCARCINOMA OF THE OVARY
C0346181|T047||CCS_10|OVARIAN CHORIOCARCINOMA
C2062541|T047||CCS_10|MALIGNANT CARCINOID TUMOR OF OVARY 
C2062541|T047||CCS_10|MALIGNANT CARCINOID TUMOR OF OVARY
C2011182|T047||CCS_10|GERMINOMA OF OVARY
C2011182|T047||CCS_10|GERMINOMA OF OVARY 
C2212020|T047||CCS_10|OVARIAN ADENOCARCINOMA SCIRRHOUS
C2212020|T047||CCS_10|SCIRRHOUS ADENOCARCINOMA OF OVARY 
C2212020|T047||CCS_10|SCIRRHOUS ADENOCARCINOMA OF OVARY
C2037342|T047||CCS_10|OVARIAN ADENOCARCINOMA SUPERFICIAL SPREADING
C2037342|T047||CCS_10|SUPERFICIAL SPREADING ADENOCARCINOMA OF OVARY 
C2037342|T047||CCS_10|SUPERFICIAL SPREADING ADENOCARCINOMA OF OVARY
C2212021|T047||CCS_10|BASAL CELL ADENOCARCINOMA OF OVARY
C2212021|T047||CCS_10|BASAL CELL ADENOCARCINOMA OF OVARY 
C2033126|T047||CCS_10|PAPILLARY ADENOCARCINOMA OF OVARY 
C2033126|T047||CCS_10|PAPILLARY ADENOCARCINOMA OF OVARY
C2189642|T047||CCS_10|VILLOUS ADENOCARCINOMA OF OVARY 
C2189642|T047||CCS_10|VILLOUS ADENOCARCINOMA OF OVARY
C2016016|T047||CCS_10|ADENOCARCINOMA IN VILLOUS ADENOMA OF OVARY 
C2016016|T047||CCS_10|ADENOCARCINOMA IN VILLOUS ADENOMA OF OVARY
C2016015|T047||CCS_10|ADENOCARCINOMA IN TUBULOVILLOUS ADENOMA OF OVARY
C2016015|T047||CCS_10|ADENOCARCINOMA IN TUBULOVILLOUS ADENOMA OF OVARY 
C2212022|T047||CCS_10|MIXED CELL ADENOCARCINOMA OF OVARY
C2212022|T047||CCS_10|MIXED CELL ADENOCARCINOMA OF OVARY 
C2212026|T047||CCS_10|ENDOCERVICAL TYPE MUCINOUS ADENOCARCINOMA OF OVARY 
C2212026|T047||CCS_10|ENDOCERVICAL TYPE MUCINOUS ADENOCARCINOMA OF OVARY
C2212027|T047||CCS_10|MUCIN-PRODUCING ADENOCARCINOMA OF OVARY 
C2212027|T047||CCS_10|MUCIN-PRODUCING ADENOCARCINOMA OF OVARY
C2212028|T047||CCS_10|ADENOCARCINOMA OF OVARY WITH METAPLASIA
C2212028|T047||CCS_10|ADENOCARCINOMA OF OVARY WITH METAPLASIA 
C2212028|T047||CCS_10|OVARIAN ADENOCARCINOMA WITH METAPLASIA
C2212029|T047||CCS_10|ADENOCARCINOMA OF OVARY WITH SQUAMOUS METAPLASIA
C2212029|T047||CCS_10|OVARIAN ADENOCARCINOMA WITH SQUAMOUS METAPLASIA
C2212029|T047||CCS_10|ADENOCARCINOMA OF OVARY WITH SQUAMOUS METAPLASIA 
C2016017|T047||CCS_10|ADENOCARCINOMA WITH CARTILAGINOUS OR OSSEOUS METAPLASIA OF OVARY
C2016017|T047||CCS_10|ADENOCARCINOMA OF OVARY WITH CARTILAGINOUS AND OSSEOUS METAPLASIA 
C2016017|T047||CCS_10|ADENOCARCINOMA OF OVARY WITH CARTILAGINOUS AND OSSEOUS METAPLASIA
C2016017|T047||CCS_10|OVARIAN ADENOCARCINOMA WITH CARTILAGINOUS OR OSSEOUS METAPLASIA
C2016017|T047||CCS_10|OVARIAN ADENOCARCINOMA WITH CARTILAGINOUS AND OSSEOUS METAPLASIA
C2212030|T047||CCS_10|OVARIAN ADENOCARCINOMA WITH SPINDLE CELL METAPLASIA
C2212030|T047||CCS_10|ADENOCARCINOMA OF OVARY WITH SPINDLE CELL METAPLASIA
C2212030|T047||CCS_10|ADENOCARCINOMA OF OVARY WITH SPINDLE CELL METAPLASIA 
C2212031|T047||CCS_10|ADENOCARCINOMA OF OVARY WITH APOCRINE METAPLASIA
C2212031|T047||CCS_10|OVARIAN ADENOCARCINOMA WITH APOCRINE METAPLASIA
C2212031|T047||CCS_10|ADENOCARCINOMA OF OVARY WITH APOCRINE METAPLASIA 
C2016018|T047||CCS_10|ADENOCARCINOMA OF OVARY WITH NEUROENDOCRINE DIFFERENTIATION
C2016018|T047||CCS_10|ADENOCARCINOMA OF OVARY WITH NEUROENDOCRINE DIFFERENTIATION 
C2016018|T047||CCS_10|OVARIAN ADENOCARCINOMA WITH NEUROENDOCRINE DIFFERENTIATION
C1335167|T047||CCS_10|MUCINOUS ADENOCARCINOMA OF OVARY 
C1335167|T047||CCS_10|MUCINOUS ADENOCARCINOMA OF OVARY
C1335167|T047||CCS_10|MUCINOUS ADENOCARCINOMA OF THE OVARY
C1335167|T047||CCS_10|MUCINOUS CARCINOMA OF OVARY
C1335167|T047||CCS_10|MUCINOUS CARCINOMA OF THE OVARY
C1335167|T047||CCS_10|OVARIAN MUCINOUS ADENOCARCINOMA
C1335167|T047||CCS_10|OVARIAN MUCINOUS CARCINOMA
C0346163|T047||CCS_10|OVARIAN ENDOMETRIOID ADENOCARCINOMA NOS
C0346163|T047||CCS_10|ENDOMETRIOID ADENOCARCINOMA OF OVARY 
C0346163|T047||CCS_10|ENDOMETRIOID ADENOCARCINOMA OF OVARY
C0346163|T047||CCS_10|OVARIAN ENDOMETRIOID CARCINOMA
C0346163|T047||CCS_10|OVARIAN MALIGNANT CARCINOMA ENDOMETRIOID
C0346163|T047||CCS_10|ENDOMETRIOID CARCINOMA OF OVARY
C0346163|T047||CCS_10|ENDOMETRIOID CARCINOMA OF OVARY 
C0346163|T047||CCS_10|OVARIAN ENDOMETRIOID ADENOCARCINOMA NOT OTHERWISE SPECIFIED
C0346163|T047||CCS_10|ENDOMETRIOID CARCINOMA OVARY
C0346163|T047||CCS_10|ENDOMETRIOID CARCINOMA OVARY 
C0346163|T047||CCS_10|OVARIAN ENDOMETRIOID ADENOCARCINOMA
C0346163|T047||CCS_10|ADENOCARCINOMA OF THE OVARY, ENDOMETRIOID
C0346163|T047||CCS_10|ENDOMETRIOID ADENOCARCINOMA OF THE OVARY
C0346163|T047||CCS_10|OVARIAN CANCER, ENDOMETRIOID ADENOCARCINOMA
C0346163|T047||CCS_10|OVARY CANCER, ENDOMETRIOID ADENOCARCINOMA
C0346163|T047||CCS_10|ENDOMETRIOID CANCER OF OVARY
C0346163|T047||CCS_10|ENDOMETRIOID CANCER OF THE OVARY
C0346163|T047||CCS_10|ENDOMETRIOID CARCINOMA OF THE OVARY
C0346163|T047||CCS_10|OVARIAN ENDOMETRIOID CANCER
C1518693|T047||CCS_10|CLEAR CELL ADENOCARCINOMA OF OVARY 
C1518693|T047||CCS_10|CLEAR CELL ADENOCARCINOMA OF OVARY
C1518693|T047||CCS_10|OVARIAN CLEAR CELL ADENOCARCINOMA
C2977928|T047||CCS_10|MALIGNANT NEOPLASM OF LEFT OVARY
C2212005|T047||CCS_10|MALIGNANT EPITHELIOMA OF OVARY
C2212005|T047||CCS_10|MALIGNANT EPITHELIOMA OF OVARY 
C2111648|T047||CCS_10|LARGE CELL CARCINOMA OF OVARY 
C2111648|T047||CCS_10|LARGE CELL CARCINOMA OF OVARY
C1335174|T047||CCS_10|LARGE CELL NEUROENDOCRINE CARCINOMA OF OVARY 
C1335174|T047||CCS_10|LARGE CELL NEUROENDOCRINE CARCINOMA OF OVARY
C1335174|T047||CCS_10|OVARIAN LARGE CELL NEC
C1335174|T047||CCS_10|LARGE CELL NEUROENDOCRINE CARCINOMA OF THE OVARY
C1335174|T047||CCS_10|LARGE-CELL NEUROENDOCRINE CARCINOMA OF OVARY
C1335174|T047||CCS_10|LARGE-CELL NEUROENDOCRINE CARCINOMA OF THE OVARY
C1335174|T047||CCS_10|NON-SMALL-CELL TYPE NEUROENDOCRINE CARCINOMA OF OVARY
C1335174|T047||CCS_10|NON-SMALL-CELL TYPE NEUROENDOCRINE CARCINOMA OF THE OVARY
C1335174|T047||CCS_10|OVARIAN NON-SMALL-CELL TYPE NEUROENDOCRINE CARCINOMA
C1335174|T047||CCS_10|OVARIAN LARGE CELL NEUROENDOCRINE CARCINOMA
C2111649|T047||CCS_10|OVARIAN MALIGNANT CARCINOMA LARGE CELL WITH RHABDOID PHENOTYPE
C2111649|T047||CCS_10|LARGE CELL CARCINOMA OF OVARY WITH RHABDOID PHENOTYPE
C2111649|T047||CCS_10|LARGE CELL CARCINOMA OF OVARY WITH RHABDOID PHENOTYPE 
C2012100|T047||CCS_10|GLASSY CELL CARCINOMA OF OVARY 
C2012100|T047||CCS_10|GLASSY CELL CARCINOMA OF OVARY
C0334398|T047||CCS_10|MALIGNANT THECOMA OF OVARY 
C0334398|T047||CCS_10|MALIGNANT THECOMA OF OVARY
C0334398|T047||CCS_10|THECOMA, OVARIAN, MALIGNANT
C0334398|T047||CCS_10|MALIGNANT OVARIAN THECAL CELL NEOPLASM
C0334398|T047||CCS_10|THECOMA, MALIGNANT
C0334398|T047||CCS_10|MALIGNANT THECAL CELL TUMOR OF THE OVARY
C0334398|T047||CCS_10|MALIGNANT THECAL CELL NEOPLASM OF OVARY
C0334398|T047||CCS_10|MALIGNANT THECAL CELL TUMOR OF OVARY
C0334398|T047||CCS_10|MALIGNANT THECOMA OF THE OVARY
C0334398|T047||CCS_10|MALIGNANT OVARIAN THECAL CELL TUMOR
C0334398|T047||CCS_10|MALIGNANT THECAL CELL NEOPLASM OF THE OVARY
C0334398|T047||CCS_10|MALIGNANT THECOMA
C0334398|T047||CCS_10|THECOMA, MALIGNANT (MORPHOLOGIC ABNORMALITY)
C0334398|T047||CCS_10|MALIGNANT; THECOMA
C0334398|T047||CCS_10|THECOMA; MALIGNANT
C0334398|T047||CCS_10|MALIGNANT OVARIAN THECOMA
C0346167|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF OVARY
C0346167|T047||CCS_10|ANAPLASTIC CARCINOMA OF OVARY
C0346167|T047||CCS_10|ANAPLASTIC CARCINOMA OF OVARY 
C0346167|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF OVARY 
C0346167|T047||CCS_10|UNDIFFERENTIATED OVARIAN CANCER
C0346167|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF OVARY 
C0346167|T047||CCS_10|ANAPLASTIC CARCINOMA OF THE OVARY
C0346167|T047||CCS_10|ANAPLASTIC OVARIAN CARCINOMA
C0346167|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF THE OVARY
C0346167|T047||CCS_10|UNDIFFERENTIATED OVARIAN CARCINOMA
C2082449|T047||CCS_10|PLEOMORPHIC CARCINOMA OF OVARY
C2082449|T047||CCS_10|PLEOMORPHIC CARCINOMA OF OVARY 
C2011259|T047||CCS_10|GIANT CELL CARCINOMA OF OVARY 
C2011259|T047||CCS_10|GIANT CELL CARCINOMA OF OVARY
C2018399|T047||CCS_10|SPINDLE CELL CARCINOMA OF OVARY
C2018399|T047||CCS_10|SPINDLE CELL CARCINOMA OF OVARY 
C2011224|T047||CCS_10|GIANT CELL AND SPINDLE CELL CARCINOMA OF OVARY
C2011224|T047||CCS_10|GIANT CELL AND SPINDLE CELL CARCINOMA OF OVARY 
C2142929|T047||CCS_10|PSEUDOSARCOMATOUS CARCINOMA OF OVARY 
C2142929|T047||CCS_10|PSEUDOSARCOMATOUS CARCINOMA OF OVARY
C2111811|T047||CCS_10|POLYGONAL CELL CARCINOMA OF OVARY 
C2111811|T047||CCS_10|POLYGONAL CELL CARCINOMA OF OVARY
C2016059|T047||CCS_10|CARCINOMA OF OVARY WITH OSTEOCLAST-LIKE GIANT CELLS 
C2016059|T047||CCS_10|CARCINOMA OF OVARY WITH OSTEOCLAST-LIKE GIANT CELLS
C2212006|T047||CCS_10|SMALL CELL CARCINOMA OF OVARY 
C2212006|T047||CCS_10|SMALL CELL CARCINOMA OF OVARY
C2212006|T047||CCS_10|OVARIAN SMALL CELL NEUROENDOCRINE CARCINOMA
C2212006|T047||CCS_10|OVARIAN SMALL CELL NEC
C2212006|T047||CCS_10|OVARIAN SMALL CELL CARCINOMA
C2033226|T047||CCS_10|PAPILLARY CARCINOMA OF OVARY
C2033226|T047||CCS_10|PAPILLARY CARCINOMA OF OVARY 
C2033303|T047||CCS_10|PAPILLARY SQUAMOUS CELL CARCINOMA OF OVARY 
C2033303|T047||CCS_10|PAPILLARY SQUAMOUS CELL CARCINOMA OF OVARY
C2189355|T047||CCS_10|VERRUCOUS CARCINOMA OF OVARY 
C2189355|T047||CCS_10|VERRUCOUS CARCINOMA OF OVARY
C2019443|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF OVARY 
C2019443|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF OVARY
C2019443|T047||CCS_10|OVARIAN SQUAMOUS CELL CARCINOMA
C2109313|T047||CCS_10|KERATINIZING SQUAMOUS CELL CARCINOMA OF OVARY
C2109313|T047||CCS_10|KERATINIZING SQUAMOUS CELL CARCINOMA OF OVARY 
C2212007|T047||CCS_10|NONKERATINIZING LARGE CELL SQUAMOUS CARCINOMA CELL OF OVARY 
C2212007|T047||CCS_10|NONKERATINIZING LARGE CELL SQUAMOUS CARCINOMA CELL OF OVARY
C2212007|T047||CCS_10|OVARIAN MALIGNANT CARCINOMA SQUAMOUS CELL LARGE CELL NONKERATINIZING
C2212008|T047||CCS_10|OVARIAN MALIGNANT CARCINOMA SQUAMOUS CELL SMALL CELL NONKERATINIZING
C2212008|T047||CCS_10|NONKERATINIZING SMALL CELL SQUAMOUS CELL CARCINOMA OF OVARY 
C2212008|T047||CCS_10|NONKERATINIZING SMALL CELL SQUAMOUS CELL CARCINOMA OF OVARY
C2018560|T047||CCS_10|SPINDLE CELL SQUAMOUS CELL CARCINOMA OF OVARY 
C2018560|T047||CCS_10|SPINDLE CELL SQUAMOUS CELL CARCINOMA OF OVARY
C2212009|T047||CCS_10|ADENOID SQUAMOUS CELL CARCINOMA OF OVARY
C2212009|T047||CCS_10|ADENOID SQUAMOUS CELL CARCINOMA OF OVARY 
C2212010|T047||CCS_10|MICROINVASIVE SQUAMOUS CELL CARCINOMA OF OVARY 
C2212010|T047||CCS_10|MICROINVASIVE SQUAMOUS CELL CARCINOMA OF OVARY
C2019488|T047||CCS_10|OVARIAN MALIGNANT CARCINOMA SQUAMOUS CELL WITH HORN FORMATION
C2019488|T047||CCS_10|SQUAMOUS CELL CARCINOMA WITH HORN FORMATION OF OVARY
C2019488|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF OVARY WITH HORN FORMATION 
C2019488|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF OVARY WITH HORN FORMATION
C2212012|T047||CCS_10|MYXOSARCOMA OF OVARY
C2212012|T047||CCS_10|MYXOSARCOMA OF OVARY 
C2212013|T047||CCS_10|OVARIAN SEROUS ADENOCARCINOFIBROMA
C2212013|T047||CCS_10|SEROUS ADENOCARCINOFIBROMA OF OVARY
C2212013|T047||CCS_10|SEROUS ADENOCARCINOFIBROMA OF OVARY 
C2212014|T047||CCS_10|MUCINOUS ADENOCARCINOFIBROMA OF OVARY
C2212014|T047||CCS_10|MUCINOUS ADENOCARCINOFIBROMA OF OVARY 
C2212014|T047||CCS_10|OVARIAN MUCINOUS ADENOCARCINOFIBROMA
C2212014|T047||CCS_10|OVARIAN MUCINOUS MALIGNANT ADENOFIBROMA
C2212017|T047||CCS_10|ADENOSQUAMOUS CARCINOMA OF OVARY 
C2212017|T047||CCS_10|ADENOSQUAMOUS CARCINOMA OF OVARY
C2212017|T047||CCS_10|OVARIAN ADENOACANTHOMA
C2212017|T047||CCS_10|OVARIAN ADENOSQUAMOUS CARCINOMA
C2212017|T047||CCS_10|OVARIAN ENDOMETRIOID ADENOCARCINOMA WITH SQUAMOUS DIFFERENTIATION
C2212018|T047||CCS_10|EPITHELIAL-MYOEPITHELIAL CARCINOMA OF OVARY
C2212018|T047||CCS_10|EPITHELIAL-MYOEPITHELIAL CARCINOMA OF OVARY 
C2017451|T047||CCS_10|SOLID CARCINOMA OF OVARY 
C2017451|T047||CCS_10|SOLID CARCINOMA OF OVARY
C2012542|T047||CCS_10|GRANULAR CELL CARCINOMA OF OVARY 
C2012542|T047||CCS_10|GRANULAR CELL CARCINOMA OF OVARY
C2212019|T047||CCS_10|MEDULLARY CARCINOMA OF OVARY
C2212019|T047||CCS_10|MEDULLARY CARCINOMA OF OVARY 
C2212023|T047||CCS_10|SECRETORY VARIANT ENDOMETRIOID ADENOCARCINOMA OF OVARY 
C2212023|T047||CCS_10|SECRETORY VARIANT ENDOMETRIOID ADENOCARCINOMA OF OVARY
C2075006|T047||CCS_10|CILIATED CELL VARIANT ENDOMETRIOID ADENOCARCINOMA OF OVARY 
C2075006|T047||CCS_10|CILIATED CELL VARIANT ENDOMETRIOID ADENOCARCINOMA OF OVARY
C2212024|T047||CCS_10|ENDOMETRIOID ADENOFIBROMA OF OVARY 
C2212024|T047||CCS_10|ENDOMETRIOID ADENOFIBROMA OF OVARY
C2212024|T047||CCS_10|OVARIAN ENDOMETRIOID ADENOFIBROMA
C2018502|T047||CCS_10|SPINDLE CELL SARCOMA OF OVARY 
C2018502|T047||CCS_10|SPINDLE CELL SARCOMA OF OVARY
C2011316|T047||CCS_10|GIANT CELL SARCOMA OF OVARY 
C2011316|T047||CCS_10|GIANT CELL SARCOMA OF OVARY
C2212032|T047||CCS_10|SMALL CELL SARCOMA OF OVARY 
C2212032|T047||CCS_10|SMALL CELL SARCOMA OF OVARY
C2212033|T047||CCS_10|EPITHELIOID SARCOMA OF OVARY
C2212033|T047||CCS_10|EPITHELIOID SARCOMA OF OVARY 
C2188139|T047||CCS_10|UNDIFFERENTIATED SARCOMA OF OVARY 
C2188139|T047||CCS_10|UNDIFFERENTIATED SARCOMA OF OVARY
C2188139|T047||CCS_10|HIGH GRADE OVARIAN ENDOMETRIOID STROMAL SARCOMA
C2188139|T047||CCS_10|UNDIFFERENTIATED OVARIAN SARCOMA
C2016060|T047||CCS_10|DESMOPLASTIC SMALL ROUND CELL TUMOR OF OVARY
C2016060|T047||CCS_10|DESMOPLASTIC SMALL ROUND CELL TUMOR OF OVARY 
C2212034|T047||CCS_10|MALIGNANT ENTEROCHROMAFFIN CELL CARCINOID TUMOR OF OVARY 
C2212034|T047||CCS_10|MALIGNANT ENTEROCHROMAFFIN CELL CARCINOID TUMOR OF OVARY
C2046334|T047||CCS_10|HISTIOCYTIC SARCOMA OF OVARY
C2046334|T047||CCS_10|HISTIOCYTIC SARCOMA OF OVARY 
C2111171|T047||CCS_10|LANGERHANS CELL SARCOMA OF OVARY 
C2111171|T047||CCS_10|LANGERHANS CELL SARCOMA OF OVARY
C2077757|T047||CCS_10|INTERDIGITATING DENDRITIC CELL SARCOMA OF OVARY
C2077757|T047||CCS_10|INTERDIGITATING DENDRITIC CELL SARCOMA OF OVARY 
C2212036|T047||CCS_10|FOLLICULAR DENDRITIC CELL SARCOMA OF OVARY
C2212036|T047||CCS_10|FOLLICULAR DENDRITIC CELL SARCOMA OF OVARY 
C2212037|T047||CCS_10|MALIGNANT ENTEROCHROMAFFIN-LIKE CELL CARCINOID TUMOR OF OVARY
C2212037|T047||CCS_10|MALIGNANT ENTEROCHROMAFFIN-LIKE CELL CARCINOID TUMOR OF OVARY 
C2212038|T047||CCS_10|FIBROMYXOSARCOMA OF OVARY 
C2212038|T047||CCS_10|FIBROMYXOSARCOMA OF OVARY
C2212039|T047||CCS_10|FASCIAL FIBROSARCOMA OF OVARY 
C2212039|T047||CCS_10|FASCIAL FIBROSARCOMA OF OVARY
C2016039|T047||CCS_10|INFANTILE FIBROSARCOMA OF OVARY 
C2016039|T047||CCS_10|INFANTILE FIBROSARCOMA OF OVARY
C2016081|T047||CCS_10|MALIGNANT SOLITARY FIBROUS TUMOR OF OVARY
C2016081|T047||CCS_10|MALIGNANT SOLITARY FIBROUS TUMOR OF OVARY 
C2016056|T047||CCS_10|GOBLET CELL CARCINOID OF OVARY
C2016056|T047||CCS_10|GOBLET CELL CARCINOID OF OVARY 
C2106919|T047||CCS_10|COMPOSITE CARCINOID TUMOR OF OVARY 
C2106919|T047||CCS_10|COMPOSITE CARCINOID TUMOR OF OVARY
C2016057|T047||CCS_10|NEUROENDOCRINE CARCINOMA OF OVARY
C2016057|T047||CCS_10|NEUROENDOCRINE CARCINOMA OF OVARY 
C2212042|T047||CCS_10|ATYPICAL CARCINOID TUMOR OF OVARY 
C2212042|T047||CCS_10|ATYPICAL CARCINOID TUMOR OF OVARY
C2212043|T047||CCS_10|ANGIOMYOSARCOMA OF OVARY
C2212043|T047||CCS_10|ANGIOMYOSARCOMA OF OVARY 
C2075522|T047||CCS_10|CLEAR CELL ADENOCARCINOFIBROMA OF OVARY 
C2075522|T047||CCS_10|CLEAR CELL ADENOCARCINOFIBROMA OF OVARY
C2075522|T047||CCS_10|OVARIAN CLEAR CELL ADENOCARCINOFIBROMA
C2075522|T047||CCS_10|OVARIAN CLEAR CELL MALIGNANT ADENOFIBROMA
C2212044|T047||CCS_10|EMBRYONAL CARCINOSARCOMA OF OVARY 
C2212044|T047||CCS_10|EMBRYONAL CARCINOSARCOMA OF OVARY
C2212045|T047||CCS_10|MALIGNANT MYOEPITHELIOMA OF OVARY
C2212045|T047||CCS_10|MALIGNANT MYOEPITHELIOMA OF OVARY 
C2033248|T047||CCS_10|PAPILLARY CYSTADENOCARCINOMA OF OVARY
C2033248|T047||CCS_10|PAPILLARY CYSTADENOCARCINOMA OF OVARY 
C2212047|T047||CCS_10|SIGNET RING CELL CARCINOMA OF OVARY 
C2212047|T047||CCS_10|SIGNET RING CELL CARCINOMA OF OVARY
C1335178|T047||CCS_10|SEROUS SURFACE PAPILLARY CARCINOMA OF OVARY 
C1335178|T047||CCS_10|SEROUS SURFACE PAPILLARY CARCINOMA OF OVARY
C1335178|T047||CCS_10|SEROUS SURFACE PAPILLARY CARCINOMA OF THE OVARY
C1335178|T047||CCS_10|OVARIAN SEROUS SURFACE PAPILLARY ADENOCARCINOMA
C2016082|T047||CCS_10|TERATOMA OF OVARY WITH MALIGNANT TRANSFORMATION
C2016082|T047||CCS_10|TERATOMA OF OVARY WITH MALIGNANT TRANSFORMATION 
C2217294|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGE IA
C2217294|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGE IA 
C2217294|T047||CCS_10|MALIGNANT OVARIAN NEOPLASM STAGE IA
C2217294|T047||CCS_10|MALIGNANT TUMOR OF OVARY STAGE IA
C2217294|T047||CCS_10|OVARIAN CANCER STAGE IA
C2217295|T047||CCS_10|MALIGNANT OVARIAN NEOPLASM STAGE IB
C2217295|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGE IB
C2217295|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGE IB 
C2217295|T047||CCS_10|MALIGNANT TUMOR OF OVARY STAGE IB
C2217295|T047||CCS_10|OVARIAN CANCER STAGE IB
C2217296|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGE IC
C2217296|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGE IC 
C2217296|T047||CCS_10|MALIGNANT OVARIAN NEOPLASM STAGE IC
C2217296|T047||CCS_10|OVARIAN CANCER STAGE IC
C2217296|T047||CCS_10|MALIGNANT TUMOR OF OVARY STAGE IC
C2217297|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGE IIA 
C2217297|T047||CCS_10|MALIGNANT OVARIAN NEOPLASM STAGE IIA
C2217297|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGE IIA
C2217297|T047||CCS_10|OVARIAN CANCER STAGE IIA
C2217297|T047||CCS_10|MALIGNANT TUMOR OF OVARY STAGE IIA
C2217298|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGE IIB 
C2217298|T047||CCS_10|MALIGNANT OVARIAN NEOPLASM STAGE IIB
C2217298|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGE IIB
C2217298|T047||CCS_10|MALIGNANT TUMOR OF OVARY STAGE IIB
C2217298|T047||CCS_10|OVARIAN CANCER STAGE IIB
C2217299|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGE IIC
C2217299|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGE IIC 
C2217299|T047||CCS_10|MALIGNANT OVARIAN NEOPLASM STAGE IIC
C2217299|T047||CCS_10|MALIGNANT TUMOR OF OVARY STAGE IIC
C2217299|T047||CCS_10|OVARIAN CANCER STAGE IIC
C2217300|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGE IIIA 
C2217300|T047||CCS_10|MALIGNANT OVARIAN NEOPLASM STAGE IIIA
C2217300|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGE IIIA
C2217300|T047||CCS_10|MALIGNANT TUMOR OF OVARY STAGE IIIA
C2217300|T047||CCS_10|OVARIAN CANCER STAGE IIIA
C2217301|T047||CCS_10|MALIGNANT OVARIAN NEOPLASM STAGE IIIB
C2217301|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGE IIIB
C2217301|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGE IIIB 
C2217301|T047||CCS_10|MALIGNANT TUMOR OF OVARY STAGE IIIB
C2217301|T047||CCS_10|OVARIAN CANCER STAGE IIIB
C2217302|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGE IIIC 
C2217302|T047||CCS_10|MALIGNANT OVARIAN NEOPLASM STAGE IIIC
C2217302|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGE IIIC
C2217302|T047||CCS_10|OVARIAN CANCER STAGE IIIC
C2217302|T047||CCS_10|MALIGNANT TUMOR OF OVARY STAGE IIIC
C2217303|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGE IV
C2217303|T047||CCS_10|MALIGNANT OVARIAN NEOPLASM STAGE IV
C2217303|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY STAGE IV 
C2217303|T047||CCS_10|MALIGNANT TUMOR OF OVARY STAGE IV
C2217303|T047||CCS_10|OVARIAN CANCER STAGE IV
C0346188|T047||CCS_10|YOLK SAC TUMOR OF OVARY 
C0346188|T047||CCS_10|YOLK SAC TUMOR OF OVARY
C0346188|T047||CCS_10|OVARIAN GERM CELL ENDODERMAL SINUS TUMOUR
C0346188|T047||CCS_10|ENDODERMAL SINUS TUMOR OF OVARY
C0346188|T047||CCS_10|ENDODERMAL SINUS TUMOR OF OVARY 
C0346188|T047||CCS_10|OVARIAN NEOPLASM MALIGNANT GERM CELL TUMOR ENDODERMAL SINUS
C0346188|T047||CCS_10|OVARIAN GERM CELL YOLK SAC TUMOR
C0346188|T047||CCS_10|OVARIAN GERM CELL ENDODERMAL SINUS TUMOR
C0346188|T047||CCS_10|OVARIAN GERM CELL YOLK SAC TUMOUR
C0346188|T047||CCS_10|ENDODERMAL SINUS TUMOUR OF OVARY
C0346188|T047||CCS_10|YOLK SAC TUMOUR OF OVARY
C0346188|T047||CCS_10|ENDODERMAL SINUS TUMOR OF OVARY 
C0346188|T047||CCS_10|ENDODERMAL SINUS TUMOR, OVARIAN GERM CELL
C0346188|T047||CCS_10|OVARIAN GERM CELL YOLK SAC CARCINOMA
C0346188|T047||CCS_10|YOLK SAC CARCINOMA, OVARIAN GERM CELL
C0346188|T047||CCS_10|ENDODERMAL SINUS NEOPLASM OF OVARY
C0346188|T047||CCS_10|ENDODERMAL SINUS NEOPLASM OF THE OVARY
C0346188|T047||CCS_10|ENDODERMAL SINUS TUMOR OF THE OVARY
C0346188|T047||CCS_10|GERM CELL ENDODERMAL SINUS NEOPLASM OF OVARY
C0346188|T047||CCS_10|GERM CELL ENDODERMAL SINUS NEOPLASM OF THE OVARY
C0346188|T047||CCS_10|GERM CELL ENDODERMAL SINUS TUMOR OF OVARY
C0346188|T047||CCS_10|GERM CELL ENDODERMAL SINUS TUMOR OF THE OVARY
C0346188|T047||CCS_10|OVARIAN ENDODERMAL SINUS NEOPLASM
C0346188|T047||CCS_10|OVARIAN ENDODERMAL SINUS TUMOR
C0346188|T047||CCS_10|OVARIAN GERM CELL ENDODERMAL SINUS NEOPLASM
C0346188|T047||CCS_10|OVARIAN YOLK SAC NEOPLASM
C0346188|T047||CCS_10|OVARIAN YOLK SAC TUMOR
C0346188|T047||CCS_10|YOLK SAC NEOPLASM OF OVARY
C0346188|T047||CCS_10|YOLK SAC NEOPLASM OF THE OVARY
C0346188|T047||CCS_10|YOLK SAC TUMOR OF THE OVARY
C0346161|T047||CCS_10|CARCINOMA OF OVARY
C0346161|T047||CCS_10|MALIGNANT EPITHELIAL TUMOR OF OVARY
C0346161|T047||CCS_10|MALIGNANT EPITHELIAL TUMOUR OF OVARY
C0346161|T047||CCS_10|MALIGNANT EPITHELIAL TUMOR OF OVARY 
C3469523|T047||CCS_10|OVARIAN CANCER SUSCEPTIBILITY 
C3469523|T047||CCS_10|OVARIAN CANCER SUSCEPTIBILITY
C3469523|T047||CCS_10|OVARIAN CANCER, SUSCEPTIBILITY TO
C0153577|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY AND OTHER UTERINE ADNEXA
C0153577|T047||CCS_10|CA OVARY/OTHER UTERINE ADNEXA
C0153577|T047||CCS_10|CA OVARY/OTHER UTERINE ADNEXA 
C0153577|T047||CCS_10|MALIGNANT NEOPLASM OF OVARY AND OTHER UTERINE ADNEXA 
C1299247|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF OVARY AND OTHER UTERINE ADNEXA 
C1299247|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF OVARY AND OTHER UTERINE ADNEXA
C1306468|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF OVARY
C1306468|T047||CCS_10|OVARIAN MALIGNANT NEOPLASM PRIMARY
C1306468|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF OVARY 
C1306468|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF OVARY 
C1299248|T047||CCS_10|CARCINOMA OF OVARY AND OTHER UTERINE ADNEXA 
C1299248|T047||CCS_10|CARCINOMA OF OVARY AND OTHER UTERINE ADNEXA
C3693886|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM FALLOPIAN TUBE 
C3693886|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM FALLOPIAN TUBE
C3693886|T047||CCS_10|OVARIAN NEOPLASM LEFT BY DIRECT EXTENSION FROM FALLOPIAN TUBE
C0346180|T047||CCS_10|OVARIAN GERM CELL CANCER
C0346180|T047||CCS_10|OVARIAN GERM CELL NEOPLASMS MALIGNANT
C0346180|T047||CCS_10|MALIGNANT GERM CELL TUMOR OF OVARY 
C0346180|T047||CCS_10|MALIGNANT GERM CELL TUMOR OF OVARY
C0346180|T047||CCS_10|OVARIAN NEOPLASM MALIGNANT GERM CELL TUMOR
C0346180|T047||CCS_10|OVARIAN GERM CELL CANCER NOS
C0346180|T047||CCS_10|MALIGNANT GERM CELL TUMOUR OF OVARY
C0346180|T047||CCS_10|MALIGNANT GERM CELL TUMOR OF OVARY 
C0346180|T047||CCS_10|MALIGNANT OVARIAN GERM CELL NEOPLASM
C0346180|T047||CCS_10|MALIGNANT GERM CELL NEOPLASM OF OVARY
C0346180|T047||CCS_10|MALIGNANT GERM CELL NEOPLASM OF THE OVARY
C0346180|T047||CCS_10|MALIGNANT GERM CELL TUMOR OF THE OVARY
C0346180|T047||CCS_10|MALIGNANT OVARIAN GERM CELL TUMOR
C3693885|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM RIGHT OVARY
C3693885|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM RIGHT OVARY 
C3693885|T047||CCS_10|OVARIAN NEOPLASM LEFT BY DIRECT EXTENSION FROM RIGHT OVARY
C3647143|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF OVARY
C3647143|T047||CCS_10|METASTASIS OF MALIGNANT NEOPLASM TO OVARY 
C3647143|T047||CCS_10|METASTASIS OF MALIGNANT NEOPLASM TO OVARY
C3647143|T047||CCS_10|METASTASES TO OVARY
C3647143|T047||CCS_10|SECOND MALIG NEO OVARY
C3647143|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF OVARY 
C3647143|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM GENITAL ORGANS OVARY
C3647143|T047||CCS_10|METASTASIS TO OVARY 
C3647143|T047||CCS_10|METASTASIS TO OVARY
C3647143|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO THE OVARY
C3647143|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM IN THE OVARY
C3647143|T047||CCS_10|OVARIAN METASTASES
C3647143|T047||CCS_10|METASTASIS TO OVARY [AMBIGUOUS]
C3647143|T047||CCS_10|METASTATIC MALIGNANT TUMOR TO THE OVARY
C3647143|T047||CCS_10|OVARIAN METASTASIS
C3693879|T047||CCS_10|OVARIAN NEOPLASM RIGHT BY DIRECT EXTENSION FROM VAGINA
C3693879|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM VAGINA 
C3693879|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM VAGINA
C3693881|T047||CCS_10|OVARIAN NEOPLASM RIGHT BY DIRECT EXTENSION FROM LEFT OVARY
C3693881|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM LEFT OVARY 
C3693881|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM LEFT OVARY
C0346175|T047||CCS_10|MALIGNANT GRANULOSA CELL TUMOR OF OVARY
C0346175|T047||CCS_10|MALIGNANT GRANULOSA CELL TUMOR OF OVARY 
C0346175|T047||CCS_10|OVARIAN NEOPLASM MALIGNANT GRANULOSA CELL
C0346175|T047||CCS_10|MALIGNANT GRANULOSA CELL NEOPLASM OF OVARY
C0346175|T047||CCS_10|MALIGNANT GRANULOSA CELL NEOPLASM OF OVARY 
C0346175|T047||CCS_10|MALIGNANT GRANULOSA CELL TUMOUR OF OVARY
C0346175|T047||CCS_10|MALIGNANT GRANULOSA CELL TUMOR OF OVARY 
C0346175|T047||CCS_10|MALIGNANT GRANULOSA CELL NEOPLASM OF THE OVARY
C0346175|T047||CCS_10|MALIGNANT GRANULOSA CELL TUMOR OF THE OVARY
C0346175|T047||CCS_10|MALIGNANT OVARIAN GRANULOSA CELL NEOPLASM
C0346175|T047||CCS_10|MALIGNANT OVARIAN GRANULOSA CELL TUMOR
C3693882|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM ENDOMETRIUM 
C3693882|T047||CCS_10|OVARIAN NEOPLASM RIGHT BY DIRECT EXTENSION FROM ENDOMETRIUM
C3693882|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM ENDOMETRIUM
C3693884|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM UTERINE CERVIX 
C3693884|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING LEFT OVARY BY DIRECT EXTENSION FROM UTERINE CERVIX
C3693884|T047||CCS_10|OVARIAN NEOPLASM LEFT BY DIRECT EXTENSION FROM UTERINE CERVIX
C3693880|T047||CCS_10|OVARIAN NEOPLASM RIGHT BY DIRECT EXTENSION FROM UTERUS
C3693880|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM UTERUS 
C3693880|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING RIGHT OVARY BY DIRECT EXTENSION FROM UTERUS
C3250633|T047||CCS_10|MALIG OVARIAN NEOPLASM TNM STAGING DISTANT METASTASIS (M) M0 
C3250633|T047||CCS_10|MALIG OVARIAN NEOPLASM TNM STAGING DISTANT METASTASIS (M) M0
C3250634|T047||CCS_10|MALIG OVARIAN NEOPLASM TNM STAGING DISTANT METASTASIS (M) M1
C3250634|T047||CCS_10|MALIG OVARIAN NEOPLASM TNM STAGING DISTANT METASTASIS (M) M1 
C3250632|T047||CCS_10|MALIG OVARIAN NEOPLASM TNM STAGING DISTANT METASTASIS (M) 
C3250632|T047||CCS_10|MALIG OVARIAN NEOPLASM TNM STAGING DISTANT METASTASIS (M)
C4030088|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM FIBROSARCOMA SOLITARY FIBROUS TUMOR
C4030088|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM FIBROSARCOMA SOLITARY FIBROUS TUMOR 
C4030115|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA PRECURSOR CELL LYMPHOBLASTIC 
C4030115|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA PRECURSOR CELL LYMPHOBLASTIC
C4030090|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM FIBROSARCOMA FIBROMYXOSARCOMA 
C4030090|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM FIBROSARCOMA FIBROMYXOSARCOMA
C4030122|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA MANTLE CELL
C4030122|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA MANTLE CELL 
C4030071|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM IMMATURE TERATOMA
C4030071|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM IMMATURE TERATOMA 
C4030060|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM PLASMACYTOMA
C4030060|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM PLASMACYTOMA 
C4030059|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM PLASMACYTOMA EXTRAMEDULLARY
C4030059|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM PLASMACYTOMA EXTRAMEDULLARY 
C4030166|T047||CCS_10|BIOPSY OVARY MALIGNANT CARCINOMA MEDULLARY 
C4030166|T047||CCS_10|BIOPSY OVARY MALIGNANT CARCINOMA MEDULLARY
C4030051|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM TERATOMA TERATOCARCINOMA
C4030051|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM TERATOMA TERATOCARCINOMA 
C4030045|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA HISTIOCYTIC
C4030045|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA HISTIOCYTIC 
C4030186|T047||CCS_10|BIOPSY OVARY MALIG LYMPHOMA PRECURSOR CELL LYMPHOBLASTIC T-CELL
C4030186|T047||CCS_10|BIOPSY OVARY MALIG LYMPHOMA PRECURSOR CELL LYMPHOBLASTIC T-CELL 
C4030114|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA SMALL B-CELL LYMPHOCYTIC
C4030114|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA SMALL B-CELL LYMPHOCYTIC 
C4030201|T047||CCS_10|BIOPSY OVARY MALIG ADENOCARCINOMA METAPLASTIC CARTILAGINOUS & OSSEOUS 
C4030201|T047||CCS_10|BIOPSY OVARY MALIG ADENOCARCINOMA METAPLASTIC CARTILAGINOUS & OSSEOUS
C4030104|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM CARCINOID TUMOR COMPOSITE 
C4030104|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM CARCINOID TUMOR COMPOSITE
C4030191|T047||CCS_10|BIOPSY OVARY MALIG LYMPHOMA HODGKIN'S LYMPHOCYT DEPLET RETICULAR
C4030191|T047||CCS_10|BIOPSY OVARY MALIG LYMPHOMA HODGKIN'S LYMPHOCYT DEPLET RETICULAR 
C4030058|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM SARCOMA 
C4030058|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM SARCOMA
C4030044|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA INTERDIGITATING DENDRITIC CELL 
C4030044|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA INTERDIGITATING DENDRITIC CELL
C4030040|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA SMALL CELL
C4030040|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA SMALL CELL 
C4030168|T047||CCS_10|BIOPSY OVARY MALIGNANT CARCINOMA LARGE CELL NEUROENDOCRINE 
C4030168|T047||CCS_10|BIOPSY OVARY MALIGNANT CARCINOMA LARGE CELL NEUROENDOCRINE
C4030160|T047||CCS_10|BIOPSY OVARY MALIGNANT CARCINOMA SEROUS SURFACE PAPILLARY 
C4030160|T047||CCS_10|BIOPSY OVARY MALIGNANT CARCINOMA SEROUS SURFACE PAPILLARY
C4030054|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM TERATOMA 
C4030054|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM TERATOMA
C4030102|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM CARCINOID TUMOR GOBLET CELL 
C4030102|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM CARCINOID TUMOR GOBLET CELL
C4030065|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM MYOSARCOMA
C4030065|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM MYOSARCOMA 
C4030134|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA FOLLICULAR GRADE 3 
C4030134|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA FOLLICULAR GRADE 3
C4030129|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA HODGKIN'S LYMPHOCYTIC DEPLETION
C4030129|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA HODGKIN'S LYMPHOCYTIC DEPLETION 
C4030083|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM GERMINOMA NONSEMINOMATOUS 
C4030083|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM GERMINOMA NONSEMINOMATOUS
C4030112|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM ADENOCARCINOFIBROMA CLEAR CELL 
C4030112|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM ADENOCARCINOFIBROMA CLEAR CELL
C4030049|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA DESMOPLASTIC SMALL ROUND CELL
C4030049|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA DESMOPLASTIC SMALL ROUND CELL 
C4030135|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA FOLLICULAR GRADE 2 
C4030135|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA FOLLICULAR GRADE 2
C4030177|T047||CCS_10|BIOPSY OVARY MALIGNANT CARCINOMA EMBRYONAL YOLK SAC TUMOR 
C4030177|T047||CCS_10|BIOPSY OVARY MALIGNANT CARCINOMA EMBRYONAL YOLK SAC TUMOR
C4030097|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM CARCINOSARCOMA MYOEPITHELIOMA
C4030097|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM CARCINOSARCOMA MYOEPITHELIOMA 
C4030111|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM ADENOCARCINOFIBROMA MUCINOUS
C4030111|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM ADENOCARCINOFIBROMA MUCINOUS 
C4030039|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA SPINDLE CELL
C4030039|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA SPINDLE CELL 
C4030064|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM MYOSARCOMA ANGIOMYOSARCOMA
C4030064|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM MYOSARCOMA ANGIOMYOSARCOMA 
C4030139|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA BURKITT'S 
C4030139|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA BURKITT'S
C4030120|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA MATURE T-CELL 
C4030120|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA MATURE T-CELL
C4030179|T047||CCS_10|BIOPSY OVARY MALIGNANT CARCINOMA EMBRYONAL
C4030179|T047||CCS_10|BIOPSY OVARY MALIGNANT CARCINOMA EMBRYONAL 
C4030178|T047||CCS_10|BIOPSY OVARY MALIGNANT CARCINOMA EMBRYONAL POLYEMBRYOMA
C4030178|T047||CCS_10|BIOPSY OVARY MALIGNANT CARCINOMA EMBRYONAL POLYEMBRYOMA 
C4030184|T047||CCS_10|BIOPSY OVARY MALIG NEOPLASM TERATOMA WITH MALIGNANT TRANSFORMATION 
C4030184|T047||CCS_10|BIOPSY OVARY MALIG NEOPLASM TERATOMA WITH MALIGNANT TRANSFORMATION
C4030062|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM MYOSARCOMA LEIOMYOSARCOMA EPITHELIOID
C4030062|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM MYOSARCOMA LEIOMYOSARCOMA EPITHELIOID 
C4030095|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM CLEAR CELL TYPE 
C4030095|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM CLEAR CELL TYPE
C4030069|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM MASTOCYTOSIS
C4030069|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM MASTOCYTOSIS 
C4030043|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA LANGERHANS CELL
C4030043|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA LANGERHANS CELL 
C4030038|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA UNDIFFERENTIATED 
C4030038|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA UNDIFFERENTIATED
C4030189|T047||CCS_10|BIOPSY OVARY MALIG LYMPHOMA HODGKIN'S NODULAR SCLEROSIS GRADE 2
C4030189|T047||CCS_10|BIOPSY OVARY MALIG LYMPHOMA HODGKIN'S NODULAR SCLEROSIS GRADE 2 
C4030132|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA HODGKIN'S 
C4030132|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA HODGKIN'S
C4030586|T047||CCS_10|BIOPSY OVARY MALIG LYMPHOMA HODGKIN'S NODULAR SCLEROSIS GRADE 1
C4030586|T047||CCS_10|BIOPSY OF OVARY SHOWED HODGKIN'S LYMPHOMA WITH GRADE 1 NODULAR SCLEROSIS 
C4030586|T047||CCS_10|BIOPSY OF OVARY SHOWED HODGKIN'S LYMPHOMA WITH GRADE 1 NODULAR SCLEROSIS
C4030066|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM MULLERIAN MIXED TUMOR 
C4030066|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM MULLERIAN MIXED TUMOR
C4030068|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM MESODERMAL MIXED TUMOR 
C4030068|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM MESODERMAL MIXED TUMOR
C4030101|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM CARCINOID TUMOR NEUROENDOCRINE
C4030101|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM CARCINOID TUMOR NEUROENDOCRINE 
C4030182|T047||CCS_10|BIOPSY OVARY MALIGNANT ADENOCARCINOMA VILLOUS 
C4030182|T047||CCS_10|BIOPSY OVARY MALIGNANT ADENOCARCINOMA VILLOUS
C4030061|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM MYOSARCOMA LEIOMYOSARCOMA MYXOID
C4030061|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM MYOSARCOMA LEIOMYOSARCOMA MYXOID 
C4030056|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM SPINDLE CELL TYPE
C4030056|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM SPINDLE CELL TYPE 
C4030192|T047||CCS_10|BIOPSY OVARY MALIG LYMPHOMA HODGKIN'S LYMPHOCYT DEPLET DIFFUSE FIBROSIS
C4030192|T047||CCS_10|BIOPSY OVARY MALIG LYMPHOMA HODGKIN'S LYMPHOCYT DEPLET DIFFUSE FIBROSIS 
C4030190|T047||CCS_10|BIOPSY OVARY MALIG LYMPHOMA HODGKIN'S NODULAR LYMPHOCYTE PREDOMINANCE 
C4030190|T047||CCS_10|BIOPSY OVARY MALIG LYMPHOMA HODGKIN'S NODULAR LYMPHOCYTE PREDOMINANCE
C4030048|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA EPITHELIOID
C4030048|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA EPITHELIOID 
C4030123|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA LYMPHOPLASMACYTIC 
C4030123|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA LYMPHOPLASMACYTIC
C4030583|T047||CCS_10|BIOPSY OF OVARY SHOWED MALIGNANT NEOPLASM
C4030583|T047||CCS_10|BIOPSY OF OVARY SHOWED MALIGNANT NEOPLASM 
C4030204|T047||CCS_10|BIOPSY OVARY MALIG ADENOCARC METAPLASTIC NEUROENDOCRINE DIFFERENTIATION 
C4030204|T047||CCS_10|BIOPSY OVARY MALIG ADENOCARC METAPLASTIC NEUROENDOCRINE DIFFERENTIATION
C4030047|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA FOLLICULAR DENDRITIC CELL 
C4030047|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA FOLLICULAR DENDRITIC CELL
C4030092|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM FIBROSARCOMA
C4030092|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM FIBROSARCOMA 
C4030187|T047||CCS_10|BIOPSY OVARY MALIG LYMPHOMA PRECURSOR CELL LYMPHOBLASTIC B-CELL
C4030187|T047||CCS_10|BIOPSY OVARY MALIG LYMPHOMA PRECURSOR CELL LYMPHOBLASTIC B-CELL 
C4030105|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM CARCINOID TUMOR ATYPICAL
C4030105|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM CARCINOID TUMOR ATYPICAL 
C4030202|T047||CCS_10|BIOPSY OVARY MALIG ADENOCARCINOMA ENDOMETRIOID SECRETORY VARIANT 
C4030202|T047||CCS_10|BIOPSY OVARY MALIG ADENOCARCINOMA ENDOMETRIOID SECRETORY VARIANT
C4030042|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA MAST CELL 
C4030042|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA MAST CELL
C4030138|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA COMPOSITE HODGKIN'S AND NON-HODGKIN'S
C4030138|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA COMPOSITE HODGKIN'S AND NON-HODGKIN'S 
C4030108|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM BRENNER TUMOR 
C4030108|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM BRENNER TUMOR
C4030110|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM ADENOCARCINOFIBROMA SEROUS
C4030110|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM ADENOCARCINOFIBROMA SEROUS 
C4030106|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM CARCINOID TUMOR ADENOCARCINOID 
C4030106|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM CARCINOID TUMOR ADENOCARCINOID
C4030103|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM CARCINOID TUMOR ENTEROCHROMAFFIN CELL 
C4030103|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM CARCINOID TUMOR ENTEROCHROMAFFIN CELL
C4030057|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM SMALL CELL TYPE
C4030057|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM SMALL CELL TYPE 
C4030137|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA FOLLICULAR
C4030137|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA FOLLICULAR 
C4030128|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA HODGKIN'S MIXED CELLULARITY
C4030128|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA HODGKIN'S MIXED CELLULARITY 
C4030127|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA HODGKIN'S NODULAR SCLEROSIS
C4030127|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA HODGKIN'S NODULAR SCLEROSIS 
C4030125|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA LARGE B-CELL DIFFUSE 
C4030125|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA LARGE B-CELL DIFFUSE
C4030119|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA MATURE T-CELL ANGIOIMMUNOBLASTIC 
C4030119|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA MATURE T-CELL ANGIOIMMUNOBLASTIC
C4030203|T047||CCS_10|BIOPSY OVARY MALIG ADENOCARCINOMA ENDOMETRIOID CILIATED CELL VARIANT
C4030203|T047||CCS_10|BIOPSY OVARY MALIG ADENOCARCINOMA ENDOMETRIOID CILIATED CELL VARIANT 
C4030113|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM ADENOCARCINOFIBROMA
C4030113|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM ADENOCARCINOFIBROMA 
C4030063|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM MYOSARCOMA LEIOMYOSARCOMA 
C4030063|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM MYOSARCOMA LEIOMYOSARCOMA
C4030126|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA HODGKIN'S SARCOMA
C4030126|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA HODGKIN'S SARCOMA 
C4030089|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM FIBROSARCOMA INFANTILE
C4030089|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM FIBROSARCOMA INFANTILE 
C4030133|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA HISTIOCYTOSIS
C4030133|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA HISTIOCYTOSIS 
C4030131|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA HODGKIN'S GRANULOMA
C4030131|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA HODGKIN'S GRANULOMA 
C4030093|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM EPITHELIOID TROPHOBLASTIC TUMOR 
C4030093|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM EPITHELIOID TROPHOBLASTIC TUMOR
C4030584|T047||CCS_10|BIOPSY OF OVARY SHOWED MALIGNANT ENDOMETRIOID ADENOFIBROMA 
C4030584|T047||CCS_10|BIOPSY OF OVARY SHOWED MALIGNANT ENDOMETRIOID ADENOFIBROMA
C4030584|T047||CCS_10|BIOPSY OVARY MALIGNANT ADENOCARCINOMA ENDOMETRIOID ADENOFIBROMA
C4030050|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM TERATOMA UNDIFFERENTIATED 
C4030050|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM TERATOMA UNDIFFERENTIATED
C4030052|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM TERATOMA MIXED GERM CELL TUMOR 
C4030052|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM TERATOMA MIXED GERM CELL TUMOR
C4030596|T047||CCS_10|BIOPSY OF OVARY SHOWED ADENOCARCINOMA WITH METAPLASIA
C4030596|T047||CCS_10|BIOPSY OF OVARY SHOWED ADENOCARCINOMA WITH METAPLASIA 
C4030596|T047||CCS_10|BIOPSY OVARY MALIGNANT ADENOCARCINOMA METAPLASTIC
C4030181|T047||CCS_10|BIOPSY OVARY MALIGNANT CARCINOMA ADENOSQUAMOUS 
C4030181|T047||CCS_10|BIOPSY OVARY MALIGNANT CARCINOMA ADENOSQUAMOUS
C4030121|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA MARGINAL ZONE B-CELL 
C4030121|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA MARGINAL ZONE B-CELL
C4030585|T047||CCS_10|BIOPSY OF OVARY SHOWED HODGKIN'S LYMPHOMA WITH NODULAR SCLEROSIS, CELLULAR PHASE 
C4030585|T047||CCS_10|BIOPSY OF OVARY SHOWED HODGKIN'S LYMPHOMA WITH NODULAR SCLEROSIS, CELLULAR PHASE
C4030585|T047||CCS_10|BIOPSY OVARY MALIG LYMPHOMA HODGKIN'S NODULAR SCLEROSIS CELLULAR PHASE
C4030053|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM TERATOMA INTERMEDIATE
C4030053|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM TERATOMA INTERMEDIATE 
C4030153|T047||CCS_10|BIOPSY OVARY MALIGNANT CARCINOMA SQUAMOUS CELL ADENOID
C4030153|T047||CCS_10|BIOPSY OVARY MALIGNANT CARCINOMA SQUAMOUS CELL ADENOID 
C4030107|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM CARCINOID TUMOR 
C4030107|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM CARCINOID TUMOR
C4030046|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA GIANT CELL 
C4030046|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA GIANT CELL
C4030041|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA MYXOSARCOMA 
C4030041|T047||CCS_10|BIOPSY OVARY MALIGNANT SARCOMA MYXOSARCOMA
C4030091|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM FIBROSARCOMA FASCIAL
C4030091|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM FIBROSARCOMA FASCIAL 
C4030188|T047||CCS_10|BIOPSY OVARY MALIG LYMPHOMA MIXED SMALL AND LARGE CELL, DIFFUSE
C4030188|T047||CCS_10|BIOPSY OVARY MALIG LYMPHOMA MIXED SMALL AND LARGE CELL, DIFFUSE 
C4030130|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA HODGKIN'S LYMPHOCYTE-RICH
C4030130|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA HODGKIN'S LYMPHOCYTE-RICH 
C4030124|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA LARGE B-CELL DIFFUSE IMMUNOBLASTIC
C4030124|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA LARGE B-CELL DIFFUSE IMMUNOBLASTIC 
C4030070|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM LYMPHOMA
C4030070|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM LYMPHOMA 
C4030067|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM MESONEPHROMA 
C4030067|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM MESONEPHROMA
C4030098|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM CARCINOSARCOMA EMBRYONAL 
C4030098|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM CARCINOSARCOMA EMBRYONAL
C4030159|T047||CCS_10|BIOPSY OVARY MALIGNANT CARCINOMA SIGNET RING CELL 
C4030159|T047||CCS_10|BIOPSY OVARY MALIGNANT CARCINOMA SIGNET RING CELL
C4030200|T047||CCS_10|BIOPSY OVARY MALIG CARCINOID TUMOR ENTEROCHROMAFFIN-LIKE CELL
C4030200|T047||CCS_10|BIOPSY OVARY MALIG CARCINOID TUMOR ENTEROCHROMAFFIN-LIKE CELL 
C4030082|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM GIANT CELL TYPE
C4030082|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM GIANT CELL TYPE 
C4030136|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA FOLLICULAR GRADE 1
C4030136|T047||CCS_10|BIOPSY OVARY MALIGNANT LYMPHOMA FOLLICULAR GRADE 1 
C4030055|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM STRUMA OVARII 
C4030055|T047||CCS_10|BIOPSY OVARY MALIGNANT NEOPLASM STRUMA OVARII
C4030196|T047||CCS_10|BIOPSY OVARY MALIG CHORIOCARCINOMA COMBINED W/ OTHER GERM CELL ELEMENTS
C4030196|T047||CCS_10|BIOPSY OVARY MALIG CHORIOCARCINOMA COMBINED W/ OTHER GERM CELL ELEMENTS 
C0022790|T047||CCS_10|KRUKENBERG TUMOR
C0022790|T047||CCS_10|KRUKENBERGS TUMOR
C0022790|T047||CCS_10|TUMOR, KRUKENBERG'S
C0022790|T047||CCS_10|TUMOR, KRUKENBERG
C0022790|T047||CCS_10|KRUKENBERG TUMOUR
C0022790|T047||CCS_10|KRUKENBURG TUMOUR
C0022790|T047||CCS_10|KRUKENBURG TUMOR
C0022790|T047||CCS_10|KRUKENBERG TUMOR 
C0022790|T047||CCS_10|KRUKENBURG TUMOR 
C0022790|T047||CCS_10|SIGNET RING CELL ADENOCARCINOMA METASTATIC TO OVARY 
C0022790|T047||CCS_10|SIGNET RING CELL ADENOCARCINOMA METASTATIC TO OVARY
C0022790|T047||CCS_10|METASTATIC CARCINOMA TO THE OVARY (KRUKENBERG TUMOR)
C0022790|T047||CCS_10|CARCINOMA, KRUKENBERG
C0022790|T047||CCS_10|KRUKENBERG TUMOR [DISEASE/FINDING]
C0022790|T047||CCS_10|KRUKENBERG'S TUMOR
C0022790|T047||CCS_10|KRUKENBERG CARCINOMA
C0022790|T047||CCS_10|CANCER METASTATIC TO OVARY
C0022790|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF OVARY
C0022790|T047||CCS_10|METASTASIS TO OVARY
C0022790|T047||CCS_10|OVARIAN METASTASIS
C0022790|T047||CCS_10|SECONDARY TUMOR TO OVARY
C0022790|T047||CCS_10|SECONDARY TUMOUR TO OVARY
C0022790|T047||CCS_10|SECONDARY CANCER OF OVARY
C0022790|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO OVARY
C0022790|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF OVARY 
C0022790|T047||CCS_10|KRUKENBERG; TUMOR
C0022790|T047||CCS_10|TUMOR; KRUKENBERG
C0022790|T047||CCS_10|KRUKENBERG NEOPLASM
C1386260|T047||CCS_10|ENDOMETRIOID; ADENOCARCINOMA, UNSPECIFIED SITE, FEMALE
C1386260|T047||CCS_10|ADENOCARCINOMA; ENDOMETRIOID, UNSPECIFIED SITE, FEMALE
C1386284|T047||CCS_10|ADENOCARCINOMA; PAPILLARY, SEROUS, UNSPECIFIED SITE
C1386284|T047||CCS_10|ADENOCARCINOMA; SEROUS PAPILLARY, UNSPECIFIED SITE
C1386284|T047||CCS_10|PAPILLARY; ADENOCARCINOMA, SEROUS, UNSPECIFIED SITE
C1386284|T047||CCS_10|SEROUS; ADENOCARCINOMA, PAPILLARY, UNSPECIFIED SITE
C1386285|T047||CCS_10|ADENOCARCINOMA; PAPILLOCYSTIC, UNSPECIFIED SITE
C1386285|T047||CCS_10|PAPILLOCYSTIC; ADENOCARCINOMA, UNSPECIFIED SITE
C1386286|T047||CCS_10|ADENOCARCINOMA; PSEUDOMUCINOUS, UNSPECIFIED SITE
C1386286|T047||CCS_10|PSEUDOMUCINOUS; ADENOCARCINOMA, UNSPECIFIED SITE
C0334341|T047||CCS_10|ENDOMETRIOID ADENOFIBROMA, MALIGNANT
C0334341|T047||CCS_10|ENDOMETRIOID CYSTADENOFIBROMA, MALIGNANT
C0334341|T047||CCS_10|MALIGNANT ENDOMETRIOID ADENOFIBROMA
C0334341|T047||CCS_10|MALIGNANT ENDOMETRIOID CYSTADENOFIBROMA
C0334341|T047||CCS_10|ENDOMETRIOID ADENOFIBROMA, MALIGNANT (MORPHOLOGIC ABNORMALITY)
C0334341|T047||CCS_10|CYSTADENOFIBROMA; ENDOMETRIOID, MALIGNANT
C0334341|T047||CCS_10|ENDOMETRIOID; ADENOFIBROMA, MALIGNANT
C0334341|T047||CCS_10|ENDOMETRIOID; CYSTADENOFIBROMA, MALIGNANT
C0334341|T047||CCS_10|ADENOFIBROMA; ENDOMETRIOID, MALIGNANT
C1388418|T047||CCS_10|MALIGNANT; ANDROBLASTOMA, UNSPECIFIED SITE, FEMALE
C1388418|T047||CCS_10|MALIGNANT; ARRHENOBLASTOMA, UNSPECIFIED SITE, FEMALE
C1388418|T047||CCS_10|ANDROBLASTOMA; MALIGNANT, UNSPECIFIED SITE, FEMALE
C1388418|T047||CCS_10|ARRHENOBLASTOMA; MALIGNANT, UNSPECIFIED SITE, FEMALE
C1390413|T047||CCS_10|BORDERLINE MALIGNANCY; MUCINOUS CYSTADENOMA, UNSPECIFIED SITE
C1390413|T047||CCS_10|CYSTADENOMA; MUCINOUS, BORDERLINE MALIGNANCY, UNSPECIFIED SITE
C1390413|T047||CCS_10|MUCINOUS; CYSTADENOMA, BORDERLINE MALIGNANCY, UNSPECIFIED SITE
C0851188|T047||CCS_10|BORDERLINE MALIGNANCY; MUCINOUS CYSTADENOMA, OVARY
C0851188|T047||CCS_10|CYSTADENOMA; MUCINOUS, BORDERLINE MALIGNANCY, OVARY
C0851188|T047||CCS_10|MUCINOUS; CYSTADENOMA, BORDERLINE MALIGNANCY, OVARY
C0851188|T047||CCS_10|OVARY; CYSTADENOMA, MUCINOUS, BORDERLINE MALIGNANCY
C0851188|T047||CCS_10|OVARY; MUCINOUS CYSTADENOMA, BORDERLINE MALIGNANCY
C1390414|T047||CCS_10|BORDERLINE MALIGNANCY; MUCINOUS PAPILLARY CYSTADENOMA, UNSPECIFIED SITE
C1390414|T047||CCS_10|BORDERLINE MALIGNANCY; PAPILLARY MUCINOUS CYSTADENOMA, UNSPECIFIED SITE
C1390414|T047||CCS_10|CYSTADENOMA; MUCINOUS, PAPILLARY, BORDERLINE MALIGNANCY, UNSPECIFIED SITE
C1390414|T047||CCS_10|CYSTADENOMA; PAPILLARY, MUCINOUS, BORDERLINE MALIGNANCY, UNSPECIFIED SITE
C1390414|T047||CCS_10|MUCINOUS; CYSTADENOMA, PAPILLARY, BORDERLINE MALIGNANCY, UNSPECIFIED SITE
C1390414|T047||CCS_10|PAPILLARY; CYSTADENOMA, MUCINOUS, BORDERLINE MALIGNANCY, UNSPECIFIED SITE
C0851177|T047||CCS_10|PAPILLARY MUCINOUS CYSTADENOMA OF OVARY OF BORDERLINE MALIGNANCY 
C0851177|T047||CCS_10|PAPILLARY MUCINOUS CYSTADENOMA OF OVARY OF BORDERLINE MALIGNANCY
C0851177|T047||CCS_10|PAPILLARY MUCINOUS OVARIAN CYSTADENOMA OF BORDERLINE MALIGNANCY
C0851177|T047||CCS_10|BORDERLINE MALIGNANCY; MUCINOUS PAPILLARY CYSTADENOMA, OVARY
C0851177|T047||CCS_10|BORDERLINE MALIGNANCY; PAPILLARY MUCINOUS CYSTADENOMA, OVARY
C0851177|T047||CCS_10|CYSTADENOMA; MUCINOUS, PAPILLARY, BORDERLINE MALIGNANCY, OVARY
C0851177|T047||CCS_10|CYSTADENOMA; PAPILLARY, MUCINOUS, BORDERLINE MALIGNANCY, OVARY
C0851177|T047||CCS_10|MUCINOUS; CYSTADENOMA, PAPILLARY, BORDERLINE MALIGNANCY, OVARY
C0851177|T047||CCS_10|OVARY; CYSTADENOMA, MUCINOUS PAPILLARY, BORDERLINE MALIGNANCY
C0851177|T047||CCS_10|OVARY; CYSTADENOMA, PAPILLARY MUCINOUS, BORDERLINE MALIGNANCY
C0851177|T047||CCS_10|OVARY; MUCINOUS PAPILLARY CYSTADENOMA, BORDERLINE MALIGNANCY
C0851177|T047||CCS_10|OVARY; PAPILLARY MUCINOUS CYSTADENOMA, BORDERLINE MALIGNANCY
C0851177|T047||CCS_10|PAPILLARY; CYSTADENOMA, MUCINOUS, BORDERLINE MALIGNANCY, OVARY
C0334356|T047||CCS_10|PAPILLARY CYSTADENOMA, BORDERLINE MALIGNANCY -RETIRED-
C0334356|T047||CCS_10|PAPILLARY CYSTADENOMA - BORDERLINE MALIGNANCY
C0334356|T047||CCS_10|PAPILLARY CYSTADENOMA - BORDERLINE MALIGNANCY 
C0334356|T047||CCS_10|PAPILLARY CYSTADENOMA, BORDERLINE MALIGNANCY
C0334356|T047||CCS_10|PAPILLARY CYSTADENOMA, BORDERLINE MALIGNANCY (MORPHOLOGIC ABNORMALITY)
C0334356|T047||CCS_10|[M] PAPILLARY CYSTADENOMA, BORDERLINE MALIGNANCY
C0334356|T047||CCS_10|[M]PAPILLARY CYSTADENOMA, BORDERLINE MALIGNANCY
C0334356|T047||CCS_10|BORDERLINE MALIGNANCY; PAPILLARY CYSTADENOMA, UNSPECIFIED SITE
C0334356|T047||CCS_10|CYSTADENOMA; PAPILLARY, BORDERLINE MALIGNANCY, UNSPECIFIED SITE
C0334356|T047||CCS_10|PAPILLARY; CYSTADENOMA, BORDERLINE MALIGNANCY, UNSPECIFIED SITE
C0334356|T047||CCS_10|LOW MALIGNANCY POTENTIAL PAPILLARY CYSTADENOMA
C0334356|T047||CCS_10|BORDERLINE MALIGNANCY PAPILLARY CYSTADENOMA
C0334356|T047||CCS_10|BORDERLINE PAPILLARY CYSTADENOMA
C0851186|T047||CCS_10|PAPILLARY CYSTADENOMA OF OVARY OF BORDERLINE MALIGNANCY 
C0851186|T047||CCS_10|PAPILLARY CYSTADENOMA OF OVARY OF BORDERLINE MALIGNANCY
C0851186|T047||CCS_10|PAPILLARY OVARIAN CYSTADENOMA OF BORDERLINE MALIGNANCY
C0851186|T047||CCS_10|BORDERLINE MALIGNANCY; PAPILLARY CYSTADENOMA, OVARY
C0851186|T047||CCS_10|CYSTADENOMA; PAPILLARY, BORDERLINE MALIGNANCY, OVARY
C0851186|T047||CCS_10|OVARY; CYSTADENOMA, PAPILLARY, BORDERLINE MALIGNANCY
C0851186|T047||CCS_10|OVARY; PAPILLARY CYSTADENOMA, BORDERLINE MALIGNANCY
C0851186|T047||CCS_10|PAPILLARY; CYSTADENOMA, BORDERLINE MALIGNANCY, OVARY
C1390415|T047||CCS_10|BORDERLINE MALIGNANCY; PAPILLARY PSEUDOMUCINOUS CYSTADENOMA, UNSPECIFIED SITE
C1390415|T047||CCS_10|BORDERLINE MALIGNANCY; PSEUDOMUCINOUS PAPILLARY CYSTADENOMA, UNSPECIFIED SITE
C1390415|T047||CCS_10|CYSTADENOMA; PAPILLARY, PSEUDOMUCINOUS, BORDERLINE MALIGNANCY, UNSPECIFIED SITE
C1390415|T047||CCS_10|CYSTADENOMA; PSEUDOMUCINOUS, PAPILLARY, BORDERLINE MALIGNANCY, UNSPECIFIED SITE
C1390415|T047||CCS_10|PAPILLARY; CYSTADENOMA, PSEUDOMUCINOUS, BORDERLINE MALIGNANCY, UNSPECIFIED SITE
C1390415|T047||CCS_10|PSEUDOMUCINOUS; CYSTADENOMA, PAPILLARY, BORDERLINE MALIGNANCY, UNSPECIFIED SITE
C1390416|T047||CCS_10|BORDERLINE MALIGNANCY; PAPILLARY PSEUDOMUCINOUS CYSTADENOMA, OVARY
C1390416|T047||CCS_10|BORDERLINE MALIGNANCY; PSEUDOMUCINOUS PAPILLARY CYSTADENOMA, OVARY
C1390416|T047||CCS_10|CYSTADENOMA; PAPILLARY, PSEUDOMUCINOUS, BORDERLINE MALIGNANCY, OVARY
C1390416|T047||CCS_10|CYSTADENOMA; PSEUDOMUCINOUS, PAPILLARY, BORDERLINE MALIGNANCY, OVARY
C1390416|T047||CCS_10|OVARY; CYSTADENOMA, PAPILLARY PSEUDOMUCINOUS, BORDERLINE MALIGNANCY
C1390416|T047||CCS_10|OVARY; CYSTADENOMA, PSEUDOMUCINOUS PAPILLARY, BORDERLINE MALIGNANCY
C1390416|T047||CCS_10|OVARY; PAPILLARY PSEUDOMUCINOUS CYSTADENOMA, BORDERLINE MALIGNANCY
C1390416|T047||CCS_10|OVARY; PSEUDOMUCINOUS PAPILLARY CYSTADENOMA, BORDERLINE MALIGNANCY
C1390416|T047||CCS_10|PAPILLARY; CYSTADENOMA, PSEUDOMUCINOUS, BORDERLINE MALIGNANCY, OVARY
C1390416|T047||CCS_10|PSEUDOMUCINOUS; CYSTADENOMA, PAPILLARY, BORDERLINE MALIGNANCY, OVARY
C1390417|T047||CCS_10|BORDERLINE MALIGNANCY; PAPILLARY SEROUS CYSTADENOMA, UNSPECIFIED SITE
C1390417|T047||CCS_10|BORDERLINE MALIGNANCY; SEROUS PAPILLARY CYSTADENOMA, UNSPECIFIED SITE
C1390417|T047||CCS_10|CYSTADENOMA; PAPILLARY, SEROUS, BORDERLINE MALIGNANCY, UNSPECIFIED SITE
C1390417|T047||CCS_10|CYSTADENOMA; SEROUS, PAPILLARY, BORDERLINE MALIGNANCY, UNSPECIFIED SITE
C1390417|T047||CCS_10|PAPILLARY; CYSTADENOMA, SEROUS, BORDERLINE MALIGNANCY, UNSPECIFIED SITE
C1390417|T047||CCS_10|SEROUS; CYSTADENOMA, PAPILLARY, BORDERLINE MALIGNANCY, UNSPECIFIED SITE
C0851187|T047||CCS_10|BORDERLINE MALIGNANCY; PAPILLARY SEROUS CYSTADENOMA, OVARY
C0851187|T047||CCS_10|BORDERLINE MALIGNANCY; SEROUS PAPILLARY CYSTADENOMA, OVARY
C0851187|T047||CCS_10|CYSTADENOMA; PAPILLARY, SEROUS, BORDERLINE MALIGNANCY, OVARY
C0851187|T047||CCS_10|CYSTADENOMA; SEROUS, PAPILLARY, BORDERLINE MALIGNANCY, OVARY
C0851187|T047||CCS_10|OVARY; CYSTADENOMA, PAPILLARY SEROUS, BORDERLINE MALIGNANCY
C0851187|T047||CCS_10|OVARY; CYSTADENOMA, SEROUS PAPILLARY, BORDERLINE MALIGNANCY
C0851187|T047||CCS_10|OVARY; PAPILLARY SEROUS CYSTADENOMA, BORDERLINE MALIGNANCY
C0851187|T047||CCS_10|OVARY; SEROUS PAPILLARY CYSTADENOMA, BORDERLINE MALIGNANCY
C0851187|T047||CCS_10|PAPILLARY; CYSTADENOMA, SEROUS, BORDERLINE MALIGNANCY, OVARY
C0851187|T047||CCS_10|SEROUS; CYSTADENOMA, PAPILLARY, BORDERLINE MALIGNANCY, OVARY
C1390418|T047||CCS_10|BORDERLINE MALIGNANCY; PSEUDOMUCINOUS CYSTADENOMA, UNSPECIFIED SITE
C1390418|T047||CCS_10|CYSTADENOMA; PSEUDOMUCINOUS, BORDERLINE MALIGNANCY, UNSPECIFIED SITE
C1390418|T047||CCS_10|PSEUDOMUCINOUS; CYSTADENOMA, BORDERLINE MALIGNANCY, UNSPECIFIED SITE
C1390419|T047||CCS_10|BORDERLINE MALIGNANCY; PSEUDOMUCINOUS CYSTADENOMA, OVARY
C1390419|T047||CCS_10|CYSTADENOMA; PSEUDOMUCINOUS, BORDERLINE MALIGNANCY, OVARY
C1390419|T047||CCS_10|OVARY; CYSTADENOMA, PSEUDOMUCINOUS, BORDERLINE MALIGNANCY
C1390419|T047||CCS_10|OVARY; PSEUDOMUCINOUS CYSTADENOMA, BORDERLINE MALIGNANCY
C1390419|T047||CCS_10|PSEUDOMUCINOUS; CYSTADENOMA, BORDERLINE MALIGNANCY, OVARY
C1390420|T047||CCS_10|BORDERLINE MALIGNANCY; SEROUS CYSTADENOMA, UNSPECIFIED SITE
C1390420|T047||CCS_10|CYSTADENOMA; SEROUS, BORDERLINE MALIGNANCY, UNSPECIFIED SITE
C1390420|T047||CCS_10|SEROUS; CYSTADENOMA, BORDERLINE MALIGNANCY, UNSPECIFIED SITE
C0851185|T047||CCS_10|SEROUS CYSTADENOMA OF BORDERLINE MALIGNANCY OF OVARY
C0851185|T047||CCS_10|SEROUS CYSTADENOMA OF BORDERLINE MALIGNANCY OF OVARY 
C0851185|T047||CCS_10|SEROUS OVARIAN CYSTADENOMA OF BORDERLINE MALIGNANCY
C0851185|T047||CCS_10|BORDERLINE MALIGNANCY; SEROUS CYSTADENOMA, OVARY
C0851185|T047||CCS_10|CYSTADENOMA; SEROUS, BORDERLINE MALIGNANCY, OVARY
C0851185|T047||CCS_10|OVARY; CYSTADENOMA, SEROUS, BORDERLINE MALIGNANCY
C0851185|T047||CCS_10|OVARY; SEROUS CYSTADENOMA, BORDERLINE MALIGNANCY
C0851185|T047||CCS_10|SEROUS; CYSTADENOMA, BORDERLINE MALIGNANCY, OVARY
C0206687|T047||CCS_10|CARCINOMA, ENDOMETRIOID
C0206687|T047||CCS_10|CARCINOMAS, ENDOMETRIOID
C0206687|T047||CCS_10|ENDOMETRIOID CARCINOMAS
C0206687|T047||CCS_10|ENDOMETRIOID CARCINOMA
C0206687|T047||CCS_10|ENDOMETRIOID CARCINOMA 
C0206687|T047||CCS_10|CARCINOMA, ENDOMETRIOID [DISEASE/FINDING]
C0206687|T047||CCS_10|ENDOMETRIOID ADENOCARCINOMA
C0206687|T047||CCS_10|ENDOMETRIOID CARCINOMA (MORPHOLOGIC ABNORMALITY)
C0206687|T047||CCS_10|CARCINOMA; ENDOMETRIOID, UNSPECIFIED SITE, FEMALE
C0206687|T047||CCS_10|ENDOMETRIOID; CARCINOMA, UNSPECIFIED SITE, FEMALE
C0206687|T047||CCS_10|ENDOMETRIOID CARCINOMA OF FEMALE REPRODUCTIVE SYSTEM
C0206687|T047||CCS_10|ENDOMETRIOID CARCINOMA OF THE FEMALE REPRODUCTIVE SYSTEM
C0206687|T047||CCS_10|FEMALE REPRODUCTIVE ENDOMETRIOID CARCINOMA
C0334401|T047||CCS_10|MALIGNANT GRANULOSA CELL TUMOR
C0334401|T047||CCS_10|GRANULOSA CELL TUMOR, MALIGNANT
C0334401|T047||CCS_10|GRANULOSA CELL CARCINOMA
C0334401|T047||CCS_10|MALIGNANT GRANULOSA CELL TUMOUR
C0334401|T047||CCS_10|GRANULOSA CELL TUMOUR, MALIGNANT
C0334401|T047||CCS_10|GRANULOSA CELL TUMOR, MALIGNANT (MORPHOLOGIC ABNORMALITY)
C0334401|T047||CCS_10|GRANULOSA CELL TUMOR, SARCOMATOID
C0334401|T047||CCS_10|GRANULOSA CELL TUMOUR, SARCOMATOID
C0334401|T047||CCS_10|CARCINOMA; GRANULOSA CELL
C0334401|T047||CCS_10|GRANULOSA CELL; CARCINOMA
C0334401|T047||CCS_10|GRANULOSA CELL; TUMOR, MALIGNANT
C0334401|T047||CCS_10|TUMOR; GRANULOSA CELL, MALIGNANT
C0334401|T047||CCS_10|MALIGNANT GRANULOSA CELL NEOPLASM
C1391921|T047||CCS_10|CARCINOMA; LEYDIG CELL, UNSPECIFIED SITE, FEMALE
C1391921|T047||CCS_10|LEYDIG CELL; CARCINOMA, UNSPECIFIED SITE, FEMALE
C1391935|T047||CCS_10|CARCINOMA; PAPILLARY, SEROUS, UNSPECIFIED SITE
C1391935|T047||CCS_10|CARCINOMA; SEROUS, PAPILLARY, UNSPECIFIED SITE
C1391935|T047||CCS_10|PAPILLARY; CARCINOMA, SEROUS, UNSPECIFIED SITE
C1391935|T047||CCS_10|SEROUS; CARCINOMA, PAPILLARY, UNSPECIFIED SITE
C1391936|T047||CCS_10|CARCINOMA; PAPILLARY, SEROUS, SUPERFICIAL, UNSPECIFIED SITE
C1391936|T047||CCS_10|CARCINOMA; SEROUS, SUPERFICIAL, PAPILLARY, UNSPECIFIED SITE
C1391936|T047||CCS_10|PAPILLARY; CARCINOMA, SEROUS, SUPERFICIAL, UNSPECIFIED SITE
C1391936|T047||CCS_10|SEROUS; CARCINOMA, SUPERFICIAL, PAPILLARY, UNSPECIFIED SITE
C1391937|T047||CCS_10|CARCINOMA; PAPILLOCYSTIC, UNSPECIFIED SITE
C1391937|T047||CCS_10|PAPILLOCYSTIC; CARCINOMA, UNSPECIFIED SITE
C1391941|T047||CCS_10|CARCINOMA; PSEUDOMUCINOUS, UNSPECIFIED SITE
C1391941|T047||CCS_10|PSEUDOMUCINOUS; CARCINOMA, UNSPECIFIED SITE
C1391945|T047||CCS_10|CARCINOMA; SERTOLI CELL, UNSPECIFIED SITE, FEMALE
C1391945|T047||CCS_10|SERTOLI CELL; CARCINOMA, UNSPECIFIED SITE, FEMALE
C0728814|T047||CCS_10|[M]THECA CELL CARCINOMA (MORPHOLOGIC ABNORMALITY)
C0728814|T047||CCS_10|[M]THECA CELL CARCINOMA
C0728814|T047||CCS_10|CARCINOMA; THECA CELL
C0728814|T047||CCS_10|THECA CELL; CARCINOMA
C1394299|T047||CCS_10|CYSTADENOCARCINOMA; ENDOMETRIOID, UNSPECIFIED SITE, FEMALE
C1394299|T047||CCS_10|ENDOMETRIOID; CYSTADENOCARCINOMA, UNSPECIFIED SITE, FEMALE
C0206699|T047||CCS_10|CYSTADENOCARCINOMA, MUCINOUS
C0206699|T047||CCS_10|CYSTADENOCARCINOMAS, MUCINOUS
C0206699|T047||CCS_10|MUCINOUS CYSTADENOCARCINOMAS
C0206699|T047||CCS_10|MUCINOUS CYSTADENOCARCINOMA
C0206699|T047||CCS_10|CYSTADENOCARCINOMA, MUCINOUS [DISEASE/FINDING]
C0206699|T047||CCS_10|[M]MUCINOUS CYSTADENOCARCINOMA NOS
C0206699|T047||CCS_10|[M]MUCINOUS CYSTADENOCARCINOMA NOS (MORPHOLOGIC ABNORMALITY)
C0206699|T047||CCS_10|PSEUDOMUCINOUS ADENOCARCINOMA
C0206699|T047||CCS_10|PSEUDOMUCINOUS CYSTADENOCARCINOMA
C0206699|T047||CCS_10|MUCINOUS CYSTADENOCARCINOMA (MORPHOLOGIC ABNORMALITY)
C0206699|T047||CCS_10|CYSTADENOCARCINOMA; MUCINOUS, UNSPECIFIED SITE
C0206699|T047||CCS_10|CYSTADENOCARCINOMA; PSEUDOMUCINOUS, UNSPECIFIED SITE
C0206699|T047||CCS_10|MUCINOUS; CYSTADENOCARCINOMA, UNSPECIFIED SITE
C0206699|T047||CCS_10|PSEUDOMUCINOUS; CYSTADENOCARCINOMA, UNSPECIFIED SITE
C0206699|T047||CCS_10|MUCINOUS CYSTADENOCARCINOMA, NOS
C0206699|T047||CCS_10|PSEUDOMUCINOUS CYSTADENOCARCINOMA, NOS
C0334364|T047||CCS_10|PAPILLARY MUCINOUS CYSTADENOCARCINOMA
C0334364|T047||CCS_10|PAPILLARY PSEUDOMUCINOUS ADENOCARCINOMA
C0334364|T047||CCS_10|PAPILLARY PSEUDOMUCINOUS CYSTADENOCARCINOMA
C0334364|T047||CCS_10|PAPILLARY MUCINOUS CYSTADENOCARCINOMA (MORPHOLOGIC ABNORMALITY)
C0334364|T047||CCS_10|CYSTADENOCARCINOMA; MUCINOUS, PAPILLARY, UNSPECIFIED SITE
C0334364|T047||CCS_10|CYSTADENOCARCINOMA; PAPILLARY, MUCINOUS, UNSPECIFIED SITE
C0334364|T047||CCS_10|MUCINOUS; CYSTADENOCARCINOMA, PAPILLARY, UNSPECIFIED SITE
C0334364|T047||CCS_10|PAPILLARY; CYSTADENOCARCINOMA, MUCINOUS, UNSPECIFIED SITE
C0206700|T047||CCS_10|CYSTADENOCARCINOMA, PAPILLARY
C0206700|T047||CCS_10|CYSTADENOCARCINOMAS, PAPILLARY
C0206700|T047||CCS_10|PAPILLARY CYSTADENOCARCINOMAS
C0206700|T047||CCS_10|PAPILLARY CYSTADENOCARCINOMA
C0206700|T047||CCS_10|CYSTADENOCARCINOMA, PAPILLARY [DISEASE/FINDING]
C0206700|T047||CCS_10|[M]PAPILLARY CYSTADENOCARCINOMA, NOS (MORPHOLOGIC ABNORMALITY)
C0206700|T047||CCS_10|[M]PAPILLARY CYSTADENOCARCINOMA, NOS
C0206700|T047||CCS_10|CYSTADENOCARCINOMA, PAPILLARY, MALIGNANT
C0206700|T047||CCS_10|PAPILLOCYSTIC ADENOCARCINOMA
C0206700|T047||CCS_10|PAPILLARY CYSTADENOCARCINOMA (MORPHOLOGIC ABNORMALITY)
C0206700|T047||CCS_10|CYSTADENOCARCINOMA; PAPILLARY, UNSPECIFIED SITE
C0206700|T047||CCS_10|PAPILLARY; CYSTADENOCARCINOMA, UNSPECIFIED SITE
C0206700|T047||CCS_10|PAPILLARY CYSTADENOCARCINOMA, NOS
C1394300|T047||CCS_10|CYSTADENOCARCINOMA; PAPILLARY, PSEUDOMUCINOUS, UNSPECIFIED SITE
C1394300|T047||CCS_10|CYSTADENOCARCINOMA; PSEUDOMUCINOUS, PAPILLARY, UNSPECIFIED SITE
C1394300|T047||CCS_10|PAPILLARY; CYSTADENOCARCINOMA, PSEUDOMUCINOUS, UNSPECIFIED SITE
C1394300|T047||CCS_10|PSEUDOMUCINOUS; CYSTADENOCARCINOMA, PAPILLARY, UNSPECIFIED SITE
C1394301|T047||CCS_10|CYSTADENOCARCINOMA; PAPILLARY, SEROUS, UNSPECIFIED SITE
C1394301|T047||CCS_10|CYSTADENOCARCINOMA; SEROUS, PAPILLARY, UNSPECIFIED SITE
C1394301|T047||CCS_10|PAPILLARY; CYSTADENOCARCINOMA, SEROUS, UNSPECIFIED SITE
C1394301|T047||CCS_10|SEROUS; CYSTADENOCARCINOMA, PAPILLARY, UNSPECIFIED SITE
C1394302|T047||CCS_10|CYSTADENOCARCINOMA; SEROUS, UNSPECIFIED SITE
C1394302|T047||CCS_10|SEROUS; CYSTADENOCARCINOMA, UNSPECIFIED SITE
C0334523|T047||CCS_10|TERATOMA WITH MALIGNANT TRANSFORMATION 
C0334523|T047||CCS_10|TERATOMA WITH MALIGNANT TRANSFORMATION
C0334523|T047||CCS_10|TERATOMA WITH MALIGNANT TRANSFORMATION (MORPHOLOGIC ABNORMALITY)
C0334523|T047||CCS_10|DERMOID CYST WITH MALIGNANT TRANSFORMATION
C0334523|T047||CCS_10|DERMOID CYST WITH MALIGNANT TRANSFORMATION (MORPHOLOGIC ABNORMALITY)
C0334523|T047||CCS_10|DERMOID CYST WITH SECONDARY TUMOR
C0334523|T047||CCS_10|DERMOID CYST WITH SECONDARY TUMOUR
C0334523|T047||CCS_10|DERMOID; CYST, WITH MALIGNANT TRANSFORMATION
C0334523|T047||CCS_10|MALIGNANT; TRANSFORMATION DERMOID CYST
C0334523|T047||CCS_10|TERATOMA WITH MALIGNANT TRANSFORMATION [DUP] (MORPHOLOGIC ABNORMALITY)
C0334523|T047||CCS_10|:: DERMOID CYST WITH MALIGNANT TRANSFORMATION
C1395294|T047||CCS_10|DERMOID; TUMOR, WITH MALIGNANT TRANSFORMATION
C1395294|T047||CCS_10|MALIGNANT; TRANSFORMATION DERMOID TUMOR
C1395294|T047||CCS_10|TUMOR; DERMOID, WITH MALIGNANT TRANSFORMATION
C1395294|T047||CCS_10|TRANSFORMATION; MALIGNANT, IN DERMOID TUMOR
C1395771|T047||CCS_10|TUMOR; YOLK SAC, UNSPECIFIED SITE, FEMALE
C1395771|T047||CCS_10|YOLK SAC; TUMOR, UNSPECIFIED SITE, FEMALE
C1395937|T047||CCS_10|DYSGERMINOMA; UNSPECIFIED SITE, FEMALE
C1396616|T047||CCS_10|ENDODERMAL; SINUS, TUMOR, UNSPECIFIED SITE, FEMALE
C1396616|T047||CCS_10|TUMOR; ENDODERMAL SINUS, UNSPECIFIED SITE, FEMALE
C1402882|T047||CCS_10|LEYDIG CELL; TUMOR, MALIGNANT, UNSPECIFIED SITE, FEMALE
C1402882|T047||CCS_10|TUMOR; LEYDIG CELL, MALIGNANT, UNSPECIFIED SITE, FEMALE
C1403527|T047||CCS_10|MALIGNANT; TRANSFORMATION DERMOID
C1334811|T047||CCS_10|MUCINOUS; TUMOR, UNSPECIFIED SITE
C1334811|T047||CCS_10|TUMOR; MUCINOUS, UNSPECIFIED SITE
C1334811|T047||CCS_10|MUCINOUS NEOPLASM
C1334811|T047||CCS_10|MUCINOUS TUMOR
C1408999|T047||CCS_10|OVARII; GOITER, MALIGNANT
C1406886|T047||CCS_10|OVARY; TERATOMA, EMBRYONAL, IMMATURE OR MALIGNANT
C1406886|T047||CCS_10|TERATOMA; OVARY, EMBRYONAL, IMMATURE OR MALIGNANT
C1407806|T047||CCS_10|PAPILLARY; TUMOR, MUCINOUS, UNSPECIFIED SITE
C1407806|T047||CCS_10|TUMOR; PAPILLARY MUCINOUS, UNSPECIFIED SITE
C0334366|T047||CCS_10|PAPILLARY MUCINOUS CYSTADENOMA, BORDERLINE MALIGNANCY -RETIRED-
C0334366|T047||CCS_10|PAPILLARY MUCINOUS CYSTADENOMA, BORDERLINE MALIGNANCY
C0334366|T047||CCS_10|PAPILLARY MUCINOUS CYSTADENOMA, BORDERLINE MALIGNANCY (MORPHOLOGIC ABNORMALITY)
C0334366|T047||CCS_10|PAPILLARY MUCINOUS CYSTADENOMA - BORDERLINE MALIGNANCY
C0334366|T047||CCS_10|PAPILLARY MUCINOUS TUMOR OF LOW MALIGNANT POTENTIAL
C0334366|T047||CCS_10|PAPILLARY MUCINOUS TUMOUR OF LOW MALIGNANT POTENTIAL
C0334366|T047||CCS_10|PAPILLARY PSEUDOMUCINOUS CYSTADENOMA, BORDERLINE MALIGNANCY
C0334366|T047||CCS_10|PAPILLARY; TUMOR, MUCINOUS, OF LOW MALIGNANT POTENTIAL
C0334366|T047||CCS_10|TUMOR; PAPILLARY, MUCINOUS, OF LOW MALIGNANT POTENTIAL
C0334366|T047||CCS_10|LOW MALIGNANCY POTENTIAL PAPILLARY MUCINOUS CYSTADENOMA
C0334366|T047||CCS_10|LOW MALIGNANCY POTENTIAL PAPILLARY PSEUDOMUCINOUS CYSTADENOMA
C0334366|T047||CCS_10|PAPILLARY MUCINOUS NEOPLASM OF LOW MALIGNANT POTENTIAL
C0334366|T047||CCS_10|BORDERLINE MALIGNANCY PAPILLARY MUCINOUS CYSTADENOMA
C0334366|T047||CCS_10|BORDERLINE MALIGNANCY PAPILLARY PSEUDOMUCINOUS CYSTADENOMA
C0334366|T047||CCS_10|BORDERLINE PAPILLARY MUCINOUS CYSTADENOMA
C0334366|T047||CCS_10|BORDERLINE PAPILLARY PSEUDOMUCINOUS CYSTADENOMA
C1407807|T047||CCS_10|PAPILLARY; TUMOR, SEROUS, LOW MALIGNANT POTENTIAL, UNSPECIFIED SITE
C1407807|T047||CCS_10|TUMOR; PAPILLARY SEROUS, LOW MALIGNANT POTENTIAL, UNSPECIFIED SITE
C1405367|T047||CCS_10|POLYVESICULAR; TUMOR, UNSPECIFIED SITE, FEMALE
C1405367|T047||CCS_10|TUMOR; POLYVESICULAR, UNSPECIFIED SITE, FEMALE
C1407812|T047||CCS_10|SEROUS; TUMOR, UNSPECIFIED SITE
C1407812|T047||CCS_10|TUMOR; SEROUS, UNSPECIFIED SITE
C1518236|T047||CCS_10|MALIGNANT OVARIAN SURFACE EPITHELIAL-STROMAL TUMOR
C1518236|T047||CCS_10|OVARIAN STROMAL CANCER
C1518236|T047||CCS_10|MALIGNANT OVARIAN EPITHELIAL TUMOR
C1518236|T047||CCS_10|CANCER, OVARIAN STROMAL
C1518236|T047||CCS_10|STROMAL CANCER, OVARIAN
C1518236|T047||CCS_10|MALIGNANT OVARIAN SURFACE EPITHELIAL-STROMAL NEOPLASM
C1518721|T047||CCS_10|OVARIAN MALIGNANT MESOTHELIOMA
C1335169|T047||CCS_10|OVARIAN MÜLLERIAN ADENOSARCOMA
C1335169|T047||CCS_10|OVARIAN MESODERMAL ADENOSARCOMA
C1335169|T047||CCS_10|OVARIAN ADENOSARCOMA
C1518720|T047||CCS_10|PRIMARY OVARIAN LYMPHOMA
C1518720|T047||CCS_10|OVARIAN LYMPHOMA
C0235770|T047||CCS_10|MALIGNANT OVARIAN CYST
C0235770|T047||CCS_10|OVARIAN CYST MALIGNANT
C1334609|T047||CCS_10|MALIGNANT OVARIAN SEX CORD-STROMAL NEOPLASM
C1334609|T047||CCS_10|MALIGNANT OVARIAN SEX CORD-STROMAL TUMOR
C1334609|T047||CCS_10|MALIGNANT SEX CORD-STROMAL TUMOR OF OVARY
C1334609|T047||CCS_10|MALIGNANT SEX CORD-STROMAL TUMOR OF THE OVARY
C1518746|T047||CCS_10|OVARIAN WILMS' TUMOR
C1518746|T047||CCS_10|OVARIAN WILMS TUMOR
C1827462|T047||CCS_10|CARCINOMA OF OVARY, STAGE 2 
C1827462|T047||CCS_10|CARCINOMA OF OVARY, STAGE 2
C1827462|T047||CCS_10|OVARIAN CANCER STAGE 2
C1827462|T047||CCS_10|CANCER OF OVARY, STAGE 2
C0346162|T047||CCS_10|SEROUS PAPILLARY CYSTADENOCARCINOMA OF OVARY
C0346162|T047||CCS_10|SEROUS PAPILLARY CYSTADENOCARCINOMA OF OVARY 
C0346162|T047||CCS_10|SEROUS PAPILLARY CYSTADENOCARCINOMA OVARY
C0346162|T047||CCS_10|SEROUS PAPILLARY CYSTADENOCARCINOMA OVARY 
C0279665|T047||CCS_10|MUCINOUS CYSTADENOCARCINOMA OF OVARY
C0279665|T047||CCS_10|MUCINOUS CYSTADENOCARCINOMA OF OVARY 
C0279665|T047||CCS_10|MUCINOUS CYSTADENOCARCINOMA OVARY
C0279665|T047||CCS_10|MUCINOUS CYSTADENOCARCINOMA OF OVARY 
C0279665|T047||CCS_10|OVARIAN MUCINOUS CYSTADENOCARCINOMA
C0279665|T047||CCS_10|CYSTADENOCARCINOMA OF THE OVARY, MUCINOUS
C0279665|T047||CCS_10|CYSTADENOCARCINOMA, MUCINOUS, OVARIAN
C0279665|T047||CCS_10|CYSTADENOCARCINOMA, OVARIAN MUCINOUS
C0279665|T047||CCS_10|MUCINOUS CYSTADENOCARCINOMA OF THE OVARY
C0279665|T047||CCS_10|OVARIAN CANCER, MUCINOUS CYSTADENOCARCINOMA
C0279665|T047||CCS_10|OVARY CANCER, MUCINOUS CYSTADENOCARCINOMA
C0521156|T047||CCS_10|EPITHELIAL OVARIAN TUMOR, INTERNATIONAL FEDERATION OF GYNECOLOGY AND OBSTETRICS STAGE IV 
C0521156|T047||CCS_10|EPITHELIAL OVARIAN TUMOR, FIGO STAGE IV 
C0521156|T047||CCS_10|EPITHELIAL OVARIAN TUMOR, INTERNATIONAL FEDERATION OF GYNECOLOGY AND OBSTETRICS STAGE IV
C0521156|T047||CCS_10|EPITHELIAL OVARIAN TUMOUR, INTERNATIONAL FEDERATION OF GYNECOLOGY AND OBSTETRICS STAGE IV
C0521156|T047||CCS_10|EPITHELIAL OVARIAN TUMOR, FIGO STAGE IV
C0521156|T047||CCS_10|EPITHELIAL OVARIAN TUMOUR, FIGO STAGE IV
C0521156|T047||CCS_10|EPITHELIAL OVARIAN TUMOR, FIGO STAGE IV (TUMOR STAGING)
C1096638|T047||CCS_10|CYSTADENOCARCINOMA OF OVARY 
C1096638|T047||CCS_10|CYSTADENOCARCINOMA OF OVARY
C1096638|T047||CCS_10|CYSTADENOCARCINOMA OVARY
C1096638|T047||CCS_10|CYSTADENOCARCINOMA OF OVARY 
C1096638|T047||CCS_10|CYSTADENOCARCINOMA OF THE OVARY
C1096638|T047||CCS_10|OVARIAN CYSTADENOCARCINOMA
C0346174|T047||CCS_10|OVARIAN NEOPLASM MALIGNANT GONADAL STROMAL TUMOR SEX CORD
C0346174|T047||CCS_10|MALIGNANT SEX CORD TUMOR OF OVARY
C0346174|T047||CCS_10|MALIGNANT SEX CORD TUMOR OF OVARY 
C0346174|T047||CCS_10|MALIGNANT SEX CORD TUMOUR OF OVARY
C0346174|T047||CCS_10|MALIGNANT SEX CORD TUMOR OF OVARY 
C1827620|T047||CCS_10|CARCINOMA OF OVARY, STAGE 4
C1827620|T047||CCS_10|CARCINOMA OF OVARY, STAGE 4 
C1827620|T047||CCS_10|OVARIAN CANCER STAGE 4
C1827620|T047||CCS_10|CANCER OF OVARY, STAGE 4
C0346183|T047||CCS_10|EMBRYONAL CARCINOMA OF OVARY
C0346183|T047||CCS_10|EMBRYONAL CARCINOMA OF OVARY 
C0346183|T047||CCS_10|OVARIAN EMBRYONAL CARCINOMA
C0346183|T047||CCS_10|EMBRYONAL CARCINOMA OF OVARY 
C0346183|T047||CCS_10|EMBRYONAL CARCINOMA OF THE OVARY
C0521152|T047||CCS_10|EPITHELIAL OVARIAN TUMOR, INTERNATIONAL FEDERATION OF GYNECOLOGY AND OBSTETRICS STAGE IIA 
C0521152|T047||CCS_10|EPITHELIAL OVARIAN TUMOR, FIGO STAGE IIA 
C0521152|T047||CCS_10|EPITHELIAL OVARIAN TUMOR, INTERNATIONAL FEDERATION OF GYNECOLOGY AND OBSTETRICS STAGE IIA
C0521152|T047||CCS_10|EPITHELIAL OVARIAN TUMOUR, INTERNATIONAL FEDERATION OF GYNAECOLOGY AND OBSTETRICS STAGE IIA
C0521152|T047||CCS_10|EPITHELIAL OVARIAN TUMOR, FIGO STAGE IIA
C0521152|T047||CCS_10|EPITHELIAL OVARIAN TUMOUR, FIGO STAGE IIA
C0521152|T047||CCS_10|EPITHELIAL OVARIAN TUMOR, FIGO STAGE IIA (TUMOR STAGING)
C1562619|T047||CCS_10|MALIGNANT MESONEPHROID TUMOR OF OVARY
C1562619|T047||CCS_10|MALIGNANT MESONEPHROID TUMOUR OF OVARY
C1562619|T047||CCS_10|PRIMARY MALIGNANT CLEAR CELL TUMOR OF OVARY 
C1562619|T047||CCS_10|PRIMARY MALIGNANT CLEAR CELL TUMOR OF OVARY
C1562619|T047||CCS_10|PRIMARY MALIGNANT CLEAR CELL TUMOUR OF OVARY
C0521154|T047||CCS_10|EPITHELIAL OVARIAN TUMOR, INTERNATIONAL FEDERATION OF GYNECOLOGY AND OBSTETRICS STAGE IIC
C0521154|T047||CCS_10|EPITHELIAL OVARIAN TUMOR, INTERNATIONAL FEDERATION OF GYNECOLOGY AND OBSTETRICS STAGE IIC 
C0521154|T047||CCS_10|EPITHELIAL OVARIAN TUMOR, FIGO STAGE IIC 
C0521154|T047||CCS_10|EPITHELIAL OVARIAN TUMOUR, INTERNATIONAL FEDERATION OF GYNECOLOGY AND OBSTETRICS STAGE IIC
C0521154|T047||CCS_10|EPITHELIAL OVARIAN TUMOR, FIGO STAGE IIC
C0521154|T047||CCS_10|EPITHELIAL OVARIAN TUMOUR, FIGO STAGE IIC
C0521154|T047||CCS_10|EPITHELIAL OVARIAN TUMOR, FIGO STAGE IIC (TUMOR STAGING)
C0346166|T047||CCS_10|OVARIAN NEOPLASM EPITHELIAL MIXED
C0346166|T047||CCS_10|MIXED EPITHELIAL NEOPLASM OF OVARY
C0346166|T047||CCS_10|MIXED EPITHELIAL NEOPLASM OF OVARY 
C0346166|T047||CCS_10|MIXED EPITHELIAL TUMOR OF OVARY
C0346166|T047||CCS_10|MIXED EPITHELIAL TUMOUR OF OVARY
C0346166|T047||CCS_10|MIXED EPITHELIAL TUMOR OF OVARY 
C0346166|T047||CCS_10|MIXED EPITHELIAL NEOPLASM OF THE OVARY
C0346166|T047||CCS_10|MIXED EPITHELIAL TUMOR OF THE OVARY
C0346166|T047||CCS_10|OVARIAN MIXED EPITHELIAL NEOPLASM
C0346166|T047||CCS_10|OVARIAN MIXED EPITHELIAL TUMOR
C1297996|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF RIGHT OVARY 
C1297996|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF RIGHT OVARY
C1297996|T047||CCS_10|OVARIAN MALIGNANT NEOPLASM PRIMARY RIGHT
C1297996|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF RIGHT OVARY 
C2016048|T047||CCS_10|MIXED CELLULARITY HODGKIN'S LYMPHOMA OF OVARY 
C2016048|T047||CCS_10|MIXED CELLULARITY HODGKIN'S LYMPHOMA OF OVARY
C2046511|T047||CCS_10|OVARIAN MALIGNANT LYMPHOMA HODGKIN'S AND NON-HODGKIN'S
C2046511|T047||CCS_10|COMPOSITE HODGKIN'S AND NON-HODGKIN'S LYMPHOMA OF OVARY 
C2046511|T047||CCS_10|COMPOSITE HODGKIN'S AND NON-HODGKIN'S LYMPHOMA OF OVARY
C2016073|T047||CCS_10|MANTLE CELL LYMPHOMA OF OVARY 
C2016073|T047||CCS_10|MANTLE CELL LYMPHOMA OF OVARY
C2016078|T047||CCS_10|NK/T-CELL LYMPHOMA OF OVARY 
C2016078|T047||CCS_10|NK/T-CELL LYMPHOMA OF OVARY
C2212025|T047||CCS_10|SEZARY SYNDROME OF OVARY 
C2212025|T047||CCS_10|SEZARY SYNDROME OF OVARY
C2016046|T047||CCS_10|OVARIAN HODGKIN LYMPHOMA LYMPHOCYTIC DEPLETION DIFFUSE FIBROSIS
C2016046|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION, DIFFUSE FIBROSIS OF OVARY
C2016046|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION, DIFFUSE FIBROSIS OF OVARY 
C2016049|T047||CCS_10|LYMPHOCYTE-RICH NODULAR HODGKIN'S LYMPHOMA OF OVARY 
C2016049|T047||CCS_10|LYMPHOCYTE-RICH NODULAR HODGKIN'S LYMPHOMA OF OVARY
C2016077|T047||CCS_10|MIXED SMALL AND LARGE CELL DIFFUSE LYMPHOMA OF OVARY 
C2016077|T047||CCS_10|MIXED SMALL AND LARGE CELL DIFFUSE LYMPHOMA OF OVARY
C2016071|T047||CCS_10|IMMUNOBLASTIC LARGE B-CELL DIFFUSE LYMPHOMA OF OVARY 
C2016071|T047||CCS_10|IMMUNOBLASTIC LARGE B-CELL DIFFUSE LYMPHOMA OF OVARY
C2016068|T047||CCS_10|GRADE 3 FOLLICULAR LYMPHOMA OF OVARY 
C2016068|T047||CCS_10|GRADE 3 FOLLICULAR LYMPHOMA OF OVARY
C2016070|T047||CCS_10|LARGE B-CELL DIFFUSE LYMPHOMA OF OVARY 
C2016070|T047||CCS_10|LARGE B-CELL DIFFUSE LYMPHOMA OF OVARY
C2016076|T047||CCS_10|ANGIOIMMUNOBLASTIC T-CELL LYMPHOMA OF OVARY 
C2016076|T047||CCS_10|ANGIOIMMUNOBLASTIC T-CELL LYMPHOMA OF OVARY
C2016076|T047||CCS_10|ANGIOIMMUNOBLASTIC LYMPHADENOPATHY WITH DYSPROTEINEMIA (AILD) OF OVARY
C2016044|T047||CCS_10|LYMPHOCYTE-RICH HODGKIN'S LYMPHOMA OF OVARY
C2016044|T047||CCS_10|LYMPHOCYTE-RICH HODGKIN'S LYMPHOMA OF OVARY 
C2016047|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION, RETICULAR OF OVARY
C2016047|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION, RETICULAR OF OVARY 
C2113645|T047||CCS_10|PRECURSOR B-CELL LYMPHOBLASTIC LYMPHOMA OF OVARY 
C2113645|T047||CCS_10|PRECURSOR B-CELL LYMPHOBLASTIC LYMPHOMA OF OVARY
C2212035|T047||CCS_10|MAST CELL SARCOMA OF OVARY 
C2212035|T047||CCS_10|MAST CELL SARCOMA OF OVARY
C2016067|T047||CCS_10|GRADE 2 FOLLICULAR LYMPHOMA OF OVARY 
C2016067|T047||CCS_10|GRADE 2 FOLLICULAR LYMPHOMA OF OVARY
C2016050|T047||CCS_10|NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF OVARY 
C2016050|T047||CCS_10|NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF OVARY
C2046584|T047||CCS_10|HODGKIN'S GRANULOMA OF OVARY
C2046584|T047||CCS_10|HODGKIN'S GRANULOMA OF OVARY 
C2016066|T047||CCS_10|GRADE 1 FOLLICULAR LYMPHOMA OF OVARY
C2016066|T047||CCS_10|GRADE 1 FOLLICULAR LYMPHOMA OF OVARY 
C2016075|T047||CCS_10|MATURE T-CELL LYMPHOMA OF OVARY
C2016075|T047||CCS_10|MATURE T-CELL LYMPHOMA OF OVARY 
C2113785|T047||CCS_10|PRECURSOR T-CELL LYMPHOBLASTIC LYMPHOMA OF OVARY
C2113785|T047||CCS_10|PRECURSOR T-CELL LYMPHOBLASTIC LYMPHOMA OF OVARY 
C2016045|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION OF OVARY 
C2016045|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION OF OVARY
C2016052|T047||CCS_10|GRADE 1 NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF OVARY
C2016052|T047||CCS_10|GRADE 1 NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF OVARY 
C2016053|T047||CCS_10|GRADE 2 NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF OVARY
C2016053|T047||CCS_10|GRADE 2 NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF OVARY 
C2016079|T047||CCS_10|SMALL B-CELL LYMPHOCYTIC LYMPHOMA OF OVARY 
C2016079|T047||CCS_10|SMALL B-CELL LYMPHOCYTIC LYMPHOMA OF OVARY
C2016074|T047||CCS_10|MARGINAL ZONE B-CELL LYMPHOMA OF OVARY 
C2016074|T047||CCS_10|MARGINAL ZONE B-CELL LYMPHOMA OF OVARY
C2113716|T047||CCS_10|PRECURSOR CELL LYMPHOBLASTIC LYMPHOMA OF OVARY 
C2113716|T047||CCS_10|PRECURSOR CELL LYMPHOBLASTIC LYMPHOMA OF OVARY
C2016051|T047||CCS_10|NODULAR SCLEROSING HODGKIN'S LYMPHOMA IN CELLULAR PHASE OF OVARY 
C2016051|T047||CCS_10|NODULAR SCLEROSING HODGKIN'S LYMPHOMA IN CELLULAR PHASE OF OVARY
C2046724|T047||CCS_10|HODGKIN'S SARCOMA OF OVARY 
C2046724|T047||CCS_10|HODGKIN'S SARCOMA OF OVARY
C2016072|T047||CCS_10|LYMPHOPLASMACYTIC LYMPHOMA OF OVARY 
C2016072|T047||CCS_10|LYMPHOPLASMACYTIC LYMPHOMA OF OVARY
C2016069|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF OVARY
C2016069|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF OVARY 
C0302592|T047||CCS_10|CARCINOMA OF CERVIX
C0302592|T047||CCS_10|CA CERVIX
C0302592|T047||CCS_10|CERVICAL CARCINOMA
C0302592|T047||CCS_10|CARCINOMA OF CERVIX 
C0302592|T047||CCS_10|CARCINOMA UTERINE CERIX
C0302592|T047||CCS_10|CARCINOMA;CERVIX
C0302592|T047||CCS_10|CA CERVIX UTERI NOS 
C0302592|T047||CCS_10|CANCER OF CERVIX
C0302592|T047||CCS_10|CERVICAL CARCINOMA (UTERUS)
C0302592|T047||CCS_10|CARCINOMA CERVIX UTERI
C0302592|T047||CCS_10|CA CERVIX UTERI NOS
C0302592|T047||CCS_10|CERVICAL CANCER
C0302592|T047||CCS_10|CERVICAL CANCER, NOS
C0302592|T047||CCS_10|CERVIX UTERI CANCER
C0302592|T047||CCS_10|CERVICAL CARCINOMA NOS
C0302592|T047||CCS_10|CERVIX CARCINOMA
C0302592|T047||CCS_10|CARCINOMA CERVIX
C0302592|T047||CCS_10|CARCINOMA UTERINE CERVIX
C0302592|T047||CCS_10|CARCINOMA OF CERVIX 
C0302592|T047||CCS_10|CANCER OF THE CERVIX
C0302592|T047||CCS_10|CERVIX CANCER
C0302592|T047||CCS_10|UTERINE CERVIX CANCER
C0302592|T047||CCS_10|UTERINE CERVIX CARCINOMA
C0302592|T047||CCS_10|CANCER OF UTERINE CERVIX
C0302592|T047||CCS_10|CANCER OF THE UTERINE CERVIX
C0302592|T047||CCS_10|CARCINOMA OF CERVIX UTERI
C0302592|T047||CCS_10|CARCINOMA OF UTERINE CERVIX
C0302592|T047||CCS_10|CARCINOMA OF THE CERVIX UTERI
C0302592|T047||CCS_10|CARCINOMA OF THE CERVIX
C0302592|T047||CCS_10|CARCINOMA OF THE UTERINE CERVIX
C0302592|T047||CCS_10|CERVIX UTERI CARCINOMA
C4048328|T047||CCS_10|CERVIX CANCER
C4048328|T047||CCS_10|CERVICAL CANCER
C4048328|T047||CCS_10|CANCER OF CERVIX
C4048328|T047||CCS_10|CERVICAL CANCER 
C4048328|T047||CCS_10|CANCERS, CERVIX
C4048328|T047||CCS_10|CANCER, CERVIX
C4048328|T047||CCS_10|CERVIX UTERI--CANCER
C4048328|T047||CCS_10|CA CERVIX
C4048328|T047||CCS_10|CANCER OF THE UTERINE CERVIX
C4048328|T047||CCS_10|CANCER OF THE CERVIX
C4048328|T047||CCS_10|UTERINE CERVICAL CANCER
C4048328|T047||CCS_10|UTERINE CERVIX CANCER
C4048328|T047||CCS_10|CANCER, UTERINE CERVICAL
C4048328|T047||CCS_10|CANCERS, UTERINE CERVICAL
C4048328|T047||CCS_10|CERVICAL CANCER, UTERINE
C4048328|T047||CCS_10|CERVICAL CANCERS, UTERINE
C4048328|T047||CCS_10|UTERINE CERVICAL CANCERS
C0279888|T047||CCS_10|CELLULAR DIAGNOSIS, CERVICAL CANCER
C0279888|T047||CCS_10|CERVICAL CANCER CELLULAR DIAGNOSIS
C0280232|T047||CCS_10|STAGE, CERVICAL CANCER
C0280232|T047||CCS_10|CERVICAL CANCER STAGE
C1280511|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF UTERINE CERVIX
C1280511|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF UTERINE CERVIX 
C4048331|T047|2.3|CCS_10|CANCER OF BRONCHUS; LUNG|CANCER OF BRONCHUS; LUNG
C0153615|T047||CCS_10|MALIGNANT NEOPLASM OF URACHUS
C0153615|T047||CCS_10|MALIGNANT NEOPLASM OF URACHUS 
C0153615|T047||CCS_10|MALIGNANT TUMOR OF URACHUS
C0153615|T047||CCS_10|MALIG NEO URACHUS
C0153615|T047||CCS_10|MALIGNANT TUMOUR OF URACHUS
C0153615|T047||CCS_10|MALIGNANT TUMOR OF URACHUS 
C0153611|T047||CCS_10|MALIGNANT NEOPLASM OF ANTERIOR WALL OF URINARY BLADDER
C0153611|T047||CCS_10|MALIGNANT NEOPLASM OF ANTERIOR WALL OF BLADDER
C0153611|T047||CCS_10|MALIGNANT NEOPLASM OF ANTERIOR WALL OF BLADDER 
C0153611|T047||CCS_10|MALIGNANT TUMOR OF ANTERIOR WALL OF BLADDER
C0153611|T047||CCS_10|MAL NEO BLADDER-ANTERIOR
C0153611|T047||CCS_10|MALIGNANT NEOPLASM OF ANTERIOR WALL OF URINARY BLADDER 
C0153613|T047||CCS_10|MALIGNANT NEOPLASM OF BLADDER NECK
C0153613|T047||CCS_10|MALIGNANT NEOPLASM OF URINARY BLADDER NECK
C0153613|T047||CCS_10|MALIGNANT NEOPLASM OF NECK OF BLADDER
C0153613|T047||CCS_10|MALIGNANT NEOPLASM OF NECK OF BLADDER 
C0153613|T047||CCS_10|MALIGNANT TUMOR OF NECK OF BLADDER
C0153613|T047||CCS_10|MAL NEO BLADDER NECK
C0153613|T047||CCS_10|MALIGNANT TUMOR OF BLADDER NECK
C0153613|T047||CCS_10|MALIGNANT TUMOUR OF BLADDER NECK
C0153613|T047||CCS_10|MALIGNANT TUMOR OF BLADDER NECK 
C0005684|T047||CCS_10|MALIGNANT NEOPLASM OF BLADDER
C0005684|T047||CCS_10|MALIGNANT NEOPLASM OF BLADDER, UNSPECIFIED
C0005684|T047||CCS_10|CANCER, URINARY BLADDER
C0005684|T047||CCS_10|BLADDER CANCER
C0005684|T047||CCS_10|MALIGNANT NEOPLASM OF BLADDER 
C0005684|T047||CCS_10|BLADDER CANCER 
C0005684|T047||CCS_10|CA BLADDER
C0005684|T047||CCS_10|BLADDER CANCERS
C0005684|T047||CCS_10|MALIGNANT TUMOR OF BLADDER
C0005684|T047||CCS_10|MALIG NEO BLADDER NOS
C0005684|T047||CCS_10|CANCER OF BLADDER
C0005684|T047||CCS_10|CANCER, BLADDER
C0005684|T047||CCS_10|BLADDER NEOPLASMS MALIGNANT
C0005684|T047||CCS_10|URINARY BLADDER CANCER
C0005684|T047||CCS_10|MALIGNANT TUMOUR OF URINARY BLADDER
C0005684|T047||CCS_10|MALIGNANT TUMOR OF URINARY BLADDER 
C0005684|T047||CCS_10|BLADDER CA
C0005684|T047||CCS_10|CA - BLADDER CANCER
C0005684|T047||CCS_10|MALIGNANT TUMOR OF URINARY BLADDER
C0005684|T047||CCS_10|MALIGNANT NEOPLASM OF URINARY BLADDER NOS
C0005684|T047||CCS_10|MALIGNANT NEOPLASM OF URINARY BLADDER NOS 
C0005684|T047||CCS_10|MALIGNANT NEOPLASM OF URINARY BLADDER
C0005684|T047||CCS_10|BLADDER--CANCER
C0005684|T047||CCS_10|BLADDER CANCER NOS
C0005684|T047||CCS_10|MALIGNANT NEOPLASM OF BLADDER, PART UNSPECIFIED
C0005684|T047||CCS_10|CANCER OF THE BLADDER
C0005684|T047||CCS_10|MALIGNANT NEOPLASM OF BLADDER, NOS
C0005684|T047||CCS_10|MALIGNANT BLADDER NEOPLASM
C0005684|T047||CCS_10|MALIGNANT BLADDER TUMOR
C0005684|T047||CCS_10|MALIGNANT NEOPLASM OF THE BLADDER
C0005684|T047||CCS_10|MALIGNANT NEOPLASM OF THE URINARY BLADDER
C0005684|T047||CCS_10|MALIGNANT NEOPLASM, BLADDER
C0005684|T047||CCS_10|MALIGNANT NEOPLASM, URINARY BLADDER
C0005684|T047||CCS_10|MALIGNANT TUMOR OF THE BLADDER
C0005684|T047||CCS_10|MALIGNANT TUMOR OF THE URINARY BLADDER
C0005684|T047||CCS_10|MALIGNANT TUMOR, URINARY BLADDER
C0005684|T047||CCS_10|MALIGNANT URINARY BLADDER NEOPLASM
C0005684|T047||CCS_10|MALIGNANT URINARY BLADDER TUMOR
C0005684|T047||CCS_10|URINARY BLADDER MALIGNANT NEOPLASM
C0005684|T047||CCS_10|URINARY BLADDER MALIGNANT TUMOR
C0005684|T047||CCS_10|NEOPLASM MALIG;BLADDER
C0005684|T047||CCS_10|MALIGNANT NEOSPLASM OF THE BLADDER
C0496827|T047||CCS_10|MALIGNANT NEOPLASM OF DOME OF BLADDER
C0496827|T047||CCS_10|MALIGNANT NEOPLASM OF APEX OF URINARY BLADDER
C0496827|T047||CCS_10|MALIGNANT NEOPLASM OF DOME OF BLADDER 
C0496827|T047||CCS_10|MALIGNANT TUMOR OF DOME OF BLADDER
C0496827|T047||CCS_10|MAL NEO BLADDER-DOME
C0496827|T047||CCS_10|MALIGNANT NEOPLASM OF DOME OF URINARY BLADDER
C0496827|T047||CCS_10|BLADDER, DOME
C0496827|T047||CCS_10|MALIGNANT TUMOR OF BLADDER DOME
C0496827|T047||CCS_10|MALIGNANT TUMOR OF VAULT OF BLADDER
C0496827|T047||CCS_10|MALIGNANT TUMOUR OF BLADDER DOME
C0496827|T047||CCS_10|MALIGNANT TUMOUR OF VAULT OF BLADDER
C0496827|T047||CCS_10|MALIGNANT NEOPLASM OF VAULT OF BLADDER
C0496827|T047||CCS_10|MALIGNANT TUMOR OF VAULT OF BLADDER 
C0496828|T047||CCS_10|MALIGNANT NEOPLASM OF LATERAL WALL OF BLADDER
C0496828|T047||CCS_10|MALIGNANT NEOPLASM OF LATERAL WALL OF URINARY BLADDER
C0496828|T047||CCS_10|MALIGNANT NEOPLASM OF LATERAL WALL OF BLADDER 
C0496828|T047||CCS_10|MALIGNANT TUMOR OF LATERAL WALL OF BLADDER
C0496828|T047||CCS_10|MAL NEO BLADDER-LATERAL
C0496828|T047||CCS_10|MALIGNANT NEOPLASM OF LATERAL WALL OF URINARY BLADDER 
C0349054|T047||CCS_10|MALIGNANT NEOPLASM OVERLAPPING BLADDER SITE
C0349054|T047||CCS_10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF BLADDER
C0349054|T047||CCS_10|MALIGNANT NEOPLASM BLADDER OVERLAPPING SITES
C0349054|T047||CCS_10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF BLADDER 
C0349054|T047||CCS_10|OVERLAPPING MALIGNANT NEOPLASM OF BLADDER
C0349054|T047||CCS_10|OVERLAPPING MALIGNANT NEOPLASM OF URINARY BLADDER 
C0349054|T047||CCS_10|OVERLAPPING MALIGNANT NEOPLASM OF URINARY BLADDER
C0349054|T047||CCS_10|MALIGNANT NEOPLASM, OVERLAPPING LESION OF BLADDER
C0349054|T047||CCS_10|MALIGNANT NEOPLASM, OVERLAPPING LESION OF BLADDER 
C0153612|T047||CCS_10|MALIGNANT NEOPLASM OF POSTERIOR WALL OF URINARY BLADDER
C0153612|T047||CCS_10|MALIGNANT NEOPLASM OF POSTERIOR WALL OF BLADDER
C0153612|T047||CCS_10|POSTERIOR WALL OF BLADDER
C0153612|T047||CCS_10|MALIGNANT NEOPLASM OF POSTERIOR WALL OF BLADDER 
C0153612|T047||CCS_10|MALIGNANT TUMOR OF POSTERIOR WALL OF BLADDER
C0153612|T047||CCS_10|MAL NEO BLADDER-POST
C0153612|T047||CCS_10|MALIGNANT NEOPLASM OF POSTERIOR WALL OF URINARY BLADDER 
C0496826|T047||CCS_10|MALIGNANT NEOPLASM OF TRIGONE OF BLADDER
C0496826|T047||CCS_10|MALIGNANT NEOPLASM OF TRIGONE OF URINARY BLADDER
C0496826|T047||CCS_10|MALIGNANT NEOPLASM OF TRIGONE OF BLADDER 
C0496826|T047||CCS_10|MALIGNANT TUMOR OF TRIGONE OF BLADDER
C0496826|T047||CCS_10|MAL NEO BLADDER-TRIGONE
C0496826|T047||CCS_10|MALIGNANT TUMOUR OF TRIGONE OF BLADDER
C0496826|T047||CCS_10|MALIGNANT TUMOR OF TRIGONE OF BLADDER 
C0496826|T047||CCS_10|MALIGNANT TUMOR OF TRIGONE OF URINARY BLADDER
C0496826|T047||CCS_10|MALIGNANT TUMOUR OF TRIGONE OF URINARY BLADDER
C0496826|T047||CCS_10|MALIGNANT TUMOR OF TRIGONE OF URINARY BLADDER 
C0153614|T047||CCS_10|MALIGNANT NEOPLASM OF URETERIC ORIFICE
C0153614|T047||CCS_10|MALIGNANT NEOPLASM OF URETERIC ORIFICE OF URINARY BLADDER
C0153614|T047||CCS_10|MALIGNANT NEOPLASM OF URETERIC ORIFICE 
C0153614|T047||CCS_10|MALIGNANT TUMOR OF URETERIC ORIFICE
C0153614|T047||CCS_10|MAL NEO URETERIC ORIFICE
C0153614|T047||CCS_10|CANCER OF URETERAL ORIFICE
C0153614|T047||CCS_10|CANCER OF URETERIC ORIFICE
C0153614|T047||CCS_10|MALIGNANT TUMOUR OF URETERIC ORIFICE
C0153614|T047||CCS_10|MALIGNANT TUMOR OF URETERIC ORIFICE 
C0855174|T047||CCS_10|BLADDER ADENOCARCINOMA RECURRENT
C0855174|T047||CCS_10|RECURRENT ADENOCARCINOMA OF BLADDER
C0855174|T047||CCS_10|RECURRENT ADENOCARCINOMA OF URINARY BLADDER
C0855174|T047||CCS_10|RECURRENT ADENOCARCINOMA OF THE BLADDER
C0855174|T047||CCS_10|RECURRENT ADENOCARCINOMA OF THE URINARY BLADDER
C0855174|T047||CCS_10|RECURRENT BLADDER ADENOCARCINOMA
C0855174|T047||CCS_10|RECURRENT URINARY BLADDER ADENOCARCINOMA
C0855174|T047||CCS_10|RELAPSED ADENOCARCINOMA OF BLADDER
C0855174|T047||CCS_10|RELAPSED ADENOCARCINOMA OF URINARY BLADDER
C0855174|T047||CCS_10|RELAPSED ADENOCARCINOMA OF THE BLADDER
C0855174|T047||CCS_10|RELAPSED ADENOCARCINOMA OF THE URINARY BLADDER
C0855174|T047||CCS_10|RELAPSED BLADDER ADENOCARCINOMA
C0855174|T047||CCS_10|RELAPSED URINARY BLADDER ADENOCARCINOMA
C0855174|T047||CCS_10|BLADDER ADENOCARCINOMA, RECURRENT
C0855175|T047||CCS_10|BLADDER ADENOCARCINOMA STAGE 0
C0855175|T047||CCS_10|STAGE 0 BLADDER ADENOCARCINOMA AJCC V7
C0855175|T047||CCS_10|STAGE 0 BLADDER ADENOCARCINOMA AJCC V6
C0855175|T047||CCS_10|STAGE 0 BLADDER ADENOCARCINOMA
C0855176|T047||CCS_10|BLADDER ADENOCARCINOMA STAGE I
C0855176|T047||CCS_10|STAGE I BLADDER ADENOCARCINOMA AJCC V7
C0855176|T047||CCS_10|STAGE I BLADDER ADENOCARCINOMA AJCC V6
C0855176|T047||CCS_10|STAGE I BLADDER ADENOCARCINOMA
C0855177|T047||CCS_10|BLADDER ADENOCARCINOMA STAGE II
C0855177|T047||CCS_10|STAGE II BLADDER ADENOCARCINOMA AJCC V6
C0855177|T047||CCS_10|STAGE II BLADDER ADENOCARCINOMA AJCC V7
C0855177|T047||CCS_10|STAGE II BLADDER ADENOCARCINOMA
C0855178|T047||CCS_10|BLADDER ADENOCARCINOMA STAGE III
C0855178|T047||CCS_10|STAGE III BLADDER ADENOCARCINOMA AJCC V7
C0855178|T047||CCS_10|STAGE III BLADDER ADENOCARCINOMA AJCC V6
C0855178|T047||CCS_10|STAGE III BLADDER ADENOCARCINOMA
C0855179|T047||CCS_10|BLADDER ADENOCARCINOMA STAGE IV
C0855179|T047||CCS_10|STAGE IV BLADDER ADENOCARCINOMA AJCC V7
C0855179|T047||CCS_10|STAGE IV BLADDER ADENOCARCINOMA
C0855180|T047||CCS_10|BLADDER ADENOCARCINOMA STAGE UNSPECIFIED
C0278827|T047||CCS_10|CA BLADDER RECURRENT
C0278827|T047||CCS_10|BLADDER CANCER RECURRENT
C0278827|T047||CCS_10|RECURRENT BLADDER CANCER
C0278827|T047||CCS_10|RECURRENT BLADDER CARCINOMA
C0278827|T047||CCS_10|CARCINOMA URINARY BLADDER RECURRENT
C0278827|T047||CCS_10|URINARY BLADDER CARCINOMA RECURRENT
C0278827|T047||CCS_10|CARCINOMA BLADDER RECURRENT
C0278827|T047||CCS_10|BLADDER CARCINOMA RECURRENT
C0278827|T047||CCS_10|BLADDER CANCER, RECURRENT
C0278827|T047||CCS_10|CANCER OF THE BLADDER, RECURRENT
C0278827|T047||CCS_10|CARCINOMA OF THE BLADDER, RECURRENT
C0278827|T047||CCS_10|RECURRENT CANCER OF THE BLADDER
C0278827|T047||CCS_10|RECURRENT CARCINOMA OF THE BLADDER
C0278827|T047||CCS_10|RECURRENT CANCER OF BLADDER
C0278827|T047||CCS_10|RECURRENT CANCER OF URINARY BLADDER
C0278827|T047||CCS_10|RECURRENT CANCER OF THE URINARY BLADDER
C0278827|T047||CCS_10|RECURRENT URINARY BLADDER CANCER
C0278827|T047||CCS_10|RELAPSED BLADDER CANCER
C0278827|T047||CCS_10|RELAPSED CANCER OF BLADDER
C0278827|T047||CCS_10|RELAPSED CANCER OF URINARY BLADDER
C0278827|T047||CCS_10|RELAPSED CANCER OF THE BLADDER
C0278827|T047||CCS_10|RELAPSED CANCER OF THE URINARY BLADDER
C0278827|T047||CCS_10|RELAPSED URINARY BLADDER CANCER
C0855181|T047||CCS_10|CA BLADDER STAGE 0, WITH CANCER IN SITU
C0855181|T047||CCS_10|BLADDER CANCER STAGE 0, WITH CANCER IN SITU
C0855181|T047||CCS_10|MALIGNANT NEOPLASM OF BLADDER STAGE 0, WITH CANCER IN SITU
C0855182|T047||CCS_10|CA BLADDER STAGE 0, WITHOUT CANCER IN SITU
C0855182|T047||CCS_10|BLADDER CANCER STAGE 0, WITHOUT CANCER IN SITU
C0855182|T047||CCS_10|MALIGNANT NEOPLASM OF BLADDER STAGE 0, WITHOUT CANCER IN SITU
C0855183|T047||CCS_10|CA BLADDER STAGE I, WITH CANCER IN SITU
C0855183|T047||CCS_10|BLADDER CANCER STAGE I, WITH CANCER IN SITU
C0855183|T047||CCS_10|MALIGNANT NEOPLASM OF BLADDER STAGE I, WITH CANCER IN SITU
C0855185|T047||CCS_10|CA BLADDER STAGE I, WITHOUT CANCER IN SITU
C0855185|T047||CCS_10|BLADDER CANCER STAGE I, WITHOUT CANCER IN SITU
C0855185|T047||CCS_10|MALIGNANT NEOPLASM OF BLADDER STAGE I, WITHOUT CANCER IN SITU
C0278823|T047||CCS_10|CA BLADDER STAGE II
C0278823|T047||CCS_10|BLADDER CANCER STAGE II
C0278823|T047||CCS_10|STAGE II BLADDER CARCINOMA AJCC V7
C0278823|T047||CCS_10|STAGE II BLADDER CANCER AJCC V7
C0278823|T047||CCS_10|STAGE II BLADDER CANCER AJCC V6
C0278823|T047||CCS_10|STAGE II BLADDER CARCINOMA AJCC V6
C0278823|T047||CCS_10|STAGE II BLADDER CANCER
C0278823|T047||CCS_10|CARCINOMA URINARY BLADDER STAGE II
C0278823|T047||CCS_10|CARCINOMA BLADDER STAGE II
C0278823|T047||CCS_10|BLADDER CARCINOMA STAGE II
C0278823|T047||CCS_10|URINARY BLADDER CARCINOMA STAGE II
C0278823|T047||CCS_10|BLADDER CANCER, STAGE B1
C0278823|T047||CCS_10|BLADDER CANCER, STAGE II
C0278823|T047||CCS_10|CANCER OF THE BLADDER, STAGE B1
C0278823|T047||CCS_10|CANCER OF THE BLADDER, STAGE II
C0278823|T047||CCS_10|CARCINOMA OF THE BLADDER, STAGE B1
C0278823|T047||CCS_10|CARCINOMA OF THE BLADDER, STAGE II
C0278823|T047||CCS_10|STAGE B1 CANCER OF THE BLADDER
C0278823|T047||CCS_10|STAGE B1 CARCINOMA OF THE BLADDER
C0278823|T047||CCS_10|STAGE II CANCER OF THE BLADDER
C0278823|T047||CCS_10|STAGE II CARCINOMA OF THE BLADDER
C0278823|T047||CCS_10|JEWETT-MARSHALL STAGE B BLADDER CANCER
C0278823|T047||CCS_10|JEWETT-MARSHALL STAGE B BLADDER CARCINOMA
C0278823|T047||CCS_10|JEWETT-MARSHALL STAGE B URINARY BLADDER CANCER
C0278823|T047||CCS_10|JEWETT-MARSHALL STAGE B URINARY BLADDER CARCINOMA
C0278823|T047||CCS_10|STAGE II BLADDER CARCINOMA
C0278823|T047||CCS_10|STAGE II CARCINOMA OF BLADDER
C0278823|T047||CCS_10|STAGE II CARCINOMA OF URINARY BLADDER
C0278823|T047||CCS_10|STAGE II CARCINOMA OF THE URINARY BLADDER
C0278823|T047||CCS_10|STAGE II URINARY BLADDER CARCINOMA
C0278823|T047||CCS_10|CANCER OF BLADDER STAGE II
C0278823|T047||CCS_10|CANCER OF THE BLADDER STAGE II
C0278824|T047||CCS_10|CA BLADDER STAGE III
C0278824|T047||CCS_10|BLADDER CANCER STAGE III
C0278824|T047||CCS_10|STAGE III BLADDER CANCER AJCC V6
C0278824|T047||CCS_10|STAGE III BLADDER CARCINOMA AJCC V7
C0278824|T047||CCS_10|STAGE III BLADDER CANCER AJCC V7
C0278824|T047||CCS_10|STAGE III BLADDER CARCINOMA AJCC V6
C0278824|T047||CCS_10|STAGE III BLADDER CANCER
C0278824|T047||CCS_10|CARCINOMA BLADDER STAGE III
C0278824|T047||CCS_10|CARCINOMA URINARY BLADDER STAGE III
C0278824|T047||CCS_10|BLADDER CARCINOMA STAGE III
C0278824|T047||CCS_10|URINARY BLADDER CARCINOMA STAGE III
C0278824|T047||CCS_10|BLADDER CANCER, STAGE III
C0278824|T047||CCS_10|CANCER OF THE BLADDER, STAGE III
C0278824|T047||CCS_10|CARCINOMA OF THE BLADDER, STAGE III
C0278824|T047||CCS_10|STAGE III CANCER OF THE BLADDER
C0278824|T047||CCS_10|STAGE III CARCINOMA OF THE BLADDER
C0278824|T047||CCS_10|JEWETT-MARSHALL STAGE C BLADDER CANCER
C0278824|T047||CCS_10|JEWETT-MARSHALL STAGE C URINARY BLADDER CANCER
C0278824|T047||CCS_10|JEWETT-MARSHALL STAGE C URINARY BLADDER CARCINOMA
C0278824|T047||CCS_10|STAGE III BLADDER CARCINOMA
C0278824|T047||CCS_10|STAGE III CARCINOMA OF BLADDER
C0278824|T047||CCS_10|STAGE III CARCINOMA OF URINARY BLADDER
C0278824|T047||CCS_10|STAGE III CARCINOMA OF THE URINARY BLADDER
C0278824|T047||CCS_10|STAGE III URINARY BLADDER CARCINOMA
C0278824|T047||CCS_10|CANCER OF BLADDER STAGE III
C0278824|T047||CCS_10|CANCER OF THE BLADDER STAGE III
C0278828|T047||CCS_10|CA BLADDER STAGE IV
C0278828|T047||CCS_10|BLADDER CANCER STAGE IV
C0278828|T047||CCS_10|CANCER OF BLADDER STAGE IV AJCC V6
C0278828|T047||CCS_10|STAGE IV CARCINOMA OF THE BLADDER AJCC V6
C0278828|T047||CCS_10|CANCER OF THE BLADDER STAGE IV AJCC V6
C0278828|T047||CCS_10|STAGE IV CARCINOMA OF URINARY BLADDER AJCC V6
C0278828|T047||CCS_10|STAGE IV CARCINOMA OF THE URINARY BLADDER AJCC V6
C0278828|T047||CCS_10|STAGE IV URINARY BLADDER CARCINOMA AJCC V6
C0278828|T047||CCS_10|STAGE IV CARCINOMA OF BLADDER AJCC V6
C0278828|T047||CCS_10|STAGE IV BLADDER CANCER AJCC V6
C0278828|T047||CCS_10|STAGE IV BLADDER CARCINOMA AJCC V6
C0278828|T047||CCS_10|METASTATIC CARCINOMA OF THE BLADDER
C0278828|T047||CCS_10|STAGE IV BLADDER CANCER
C0278828|T047||CCS_10|URINARY BLADDER CARCINOMA STAGE IV
C0278828|T047||CCS_10|CARCINOMA BLADDER STAGE IV
C0278828|T047||CCS_10|CARCINOMA URINARY BLADDER STAGE IV
C0278828|T047||CCS_10|BLADDER CARCINOMA STAGE IV
C0278828|T047||CCS_10|BLADDER CANCER, METASTATIC
C0278828|T047||CCS_10|BLADDER CANCER, STAGE IV
C0278828|T047||CCS_10|CANCER OF THE BLADDER, METASTATIC
C0278828|T047||CCS_10|CANCER OF THE BLADDER, STAGE IV
C0278828|T047||CCS_10|CARCINOMA OF THE BLADDER, METASTATIC
C0278828|T047||CCS_10|CARCINOMA OF THE BLADDER, STAGE IV
C0278828|T047||CCS_10|METASTATIC BLADDER CANCER
C0278828|T047||CCS_10|METASTATIC CANCER OF THE BLADDER
C0278828|T047||CCS_10|STAGE IV CANCER OF THE BLADDER
C0278828|T047||CCS_10|STAGE IV CARCINOMA OF THE BLADDER
C0278828|T047||CCS_10|JEWETT-MARSHALL STAGE D BLADDER CANCER
C0278828|T047||CCS_10|JEWETT-MARSHALL STAGE D BLADDER CARCINOMA
C0278828|T047||CCS_10|JEWETT-MARSHALL STAGE D URINARY BLADDER CANCER
C0278828|T047||CCS_10|JEWETT-MARSHALL STAGE D URINARY BLADDER CARCINOMA
C0855186|T047||CCS_10|BLADDER SQUAMOUS CELL CARCINOMA RECURRENT
C0855186|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE BLADDER RECURRENT
C0855186|T047||CCS_10|SQUAMOUS CELL BLADDER CARCINOMA RECURRENT
C0855186|T047||CCS_10|RECURRENT BLADDER EPIDERMOID CARCINOMA
C0855186|T047||CCS_10|RECURRENT BLADDER SQUAMOUS CELL CARCINOMA
C0855186|T047||CCS_10|RECURRENT EPIDERMOID CARCINOMA OF BLADDER
C0855186|T047||CCS_10|RECURRENT EPIDERMOID CARCINOMA OF URINARY BLADDER
C0855186|T047||CCS_10|RECURRENT EPIDERMOID CARCINOMA OF THE BLADDER
C0855186|T047||CCS_10|RECURRENT EPIDERMOID CARCINOMA OF THE URINARY BLADDER
C0855186|T047||CCS_10|RECURRENT SQUAMOUS CELL CARCINOMA OF BLADDER
C0855186|T047||CCS_10|RECURRENT SQUAMOUS CELL CARCINOMA OF URINARY BLADDER
C0855186|T047||CCS_10|RECURRENT SQUAMOUS CELL CARCINOMA OF THE BLADDER
C0855186|T047||CCS_10|RECURRENT SQUAMOUS CELL CARCINOMA OF THE URINARY BLADDER
C0855186|T047||CCS_10|RECURRENT URINARY BLADDER EPIDERMOID CARCINOMA
C0855186|T047||CCS_10|RECURRENT URINARY BLADDER SQUAMOUS CELL CARCINOMA
C0855186|T047||CCS_10|RELAPSED BLADDER EPIDERMOID CARCINOMA
C0855186|T047||CCS_10|RELAPSED BLADDER SQUAMOUS CELL CARCINOMA
C0855186|T047||CCS_10|RELAPSED EPIDERMOID CARCINOMA OF BLADDER
C0855186|T047||CCS_10|RELAPSED EPIDERMOID CARCINOMA OF URINARY BLADDER
C0855186|T047||CCS_10|RELAPSED EPIDERMOID CARCINOMA OF THE BLADDER
C0855186|T047||CCS_10|RELAPSED EPIDERMOID CARCINOMA OF THE URINARY BLADDER
C0855186|T047||CCS_10|RELAPSED SQUAMOUS CELL CARCINOMA OF BLADDER
C0855186|T047||CCS_10|RELAPSED SQUAMOUS CELL CARCINOMA OF URINARY BLADDER
C0855186|T047||CCS_10|RELAPSED SQUAMOUS CELL CARCINOMA OF THE BLADDER
C0855186|T047||CCS_10|RELAPSED SQUAMOUS CELL CARCINOMA OF THE URINARY BLADDER
C0855186|T047||CCS_10|RELAPSED URINARY BLADDER EPIDERMOID CARCINOMA
C0855186|T047||CCS_10|RELAPSED URINARY BLADDER SQUAMOUS CELL CARCINOMA
C0855186|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF BLADDER, RECURRENT
C0855186|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE BLADDER, RECURRENT
C0855187|T047||CCS_10|BLADDER SQUAMOUS CELL CARCINOMA STAGE 0
C0855187|T047||CCS_10|STAGE 0 BLADDER SQUAMOUS CELL CARCINOMA AJCC V6
C0855187|T047||CCS_10|STAGE 0 BLADDER SQUAMOUS CELL CARCINOMA AJCC V7
C0855187|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE BLADDER STAGE 0
C0855187|T047||CCS_10|SQUAMOUS CELL BLADDER CARCINOMA STAGE 0
C0855187|T047||CCS_10|STAGE 0 BLADDER SQUAMOUS CELL CARCINOMA
C0855187|T047||CCS_10|STAGE 0 SQUAMOUS CELL CARCINOMA OF BLADDER
C0855187|T047||CCS_10|STAGE 0 SQUAMOUS CELL CARCINOMA OF THE BLADDER
C0855188|T047||CCS_10|BLADDER SQUAMOUS CELL CARCINOMA STAGE I
C0855188|T047||CCS_10|STAGE I SQUAMOUS CELL CARCINOMA OF THE BLADDER AJCC V7
C0855188|T047||CCS_10|STAGE I SQUAMOUS CELL CARCINOMA OF THE BLADDER AJCC V6
C0855188|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE BLADDER STAGE I
C0855188|T047||CCS_10|SQUAMOUS CELL BLADDER CARCINOMA STAGE I
C0855188|T047||CCS_10|STAGE I SQUAMOUS CELL CARCINOMA OF BLADDER
C0855188|T047||CCS_10|STAGE I SQUAMOUS CELL CARCINOMA OF THE BLADDER
C0855189|T047||CCS_10|BLADDER SQUAMOUS CELL CARCINOMA STAGE II
C0855189|T047||CCS_10|STAGE II BLADDER SQUAMOUS CELL CARCINOMA AJCC V6
C0855189|T047||CCS_10|STAGE II BLADDER SQUAMOUS CELL CARCINOMA AJCC V7
C0855189|T047||CCS_10|SQUAMOUS CELL BLADDER CARCINOMA STAGE II
C0855189|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE BLADDER STAGE II
C0855189|T047||CCS_10|STAGE II BLADDER SQUAMOUS CELL CARCINOMA
C0855190|T047||CCS_10|BLADDER SQUAMOUS CELL CARCINOMA STAGE III
C0855190|T047||CCS_10|STAGE III BLADDER SQUAMOUS CELL CARCINOMA AJCC V6
C0855190|T047||CCS_10|STAGE III BLADDER SQUAMOUS CELL CARCINOMA AJCC V7
C0855190|T047||CCS_10|SQUAMOUS CELL BLADDER CARCINOMA STAGE III
C0855190|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE BLADDER STAGE III
C0855190|T047||CCS_10|STAGE III BLADDER SQUAMOUS CELL CARCINOMA
C0855191|T047||CCS_10|BLADDER SQUAMOUS CELL CARCINOMA STAGE IV
C0855191|T047||CCS_10|STAGE IV BLADDER SQUAMOUS CELL CARCINOMA AJCC V7
C0855191|T047||CCS_10|SQUAMOUS CELL BLADDER CARCINOMA STAGE IV
C0855191|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE BLADDER STAGE IV
C0855191|T047||CCS_10|STAGE IV BLADDER SQUAMOUS CELL CARCINOMA
C0855192|T047||CCS_10|BLADDER SQUAMOUS CELL CARCINOMA STAGE UNSPECIFIED
C0855192|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE BLADDER STAGE UNSPECIFIED
C0279680|T047||CCS_10|BLADDER TRANSITIONAL CELL CARCINOMA
C0279680|T047||CCS_10|TRANSITIONAL CELL CARCINOMA OF THE BLADDER
C0279680|T047||CCS_10|TRANSITIONAL CELL CARCINOMA OF BLADDER
C0279680|T047||CCS_10|TRANSITIONAL CELL CARCINOMA OF BLADDER 
C0279680|T047||CCS_10|TRANSITIONAL CELL CARCINOMA OF BLADDER 
C0279680|T047||CCS_10|BLADDER UROTHELIAL CARCINOMA
C0279680|T047||CCS_10|TRANSITIONAL CELL BLADDER CARCINOMA
C0279680|T047||CCS_10|UROTHELIAL CARCINOMA BLADDER
C0279680|T047||CCS_10|TCC - TRANSITIONAL CELL CARCINOMA OF BLADDER
C0279680|T047||CCS_10|BLADDER CANCER, TRANSITIONAL CELL CARCINOMA
C0279680|T047||CCS_10|CARCINOMA, TRANSITIONAL CELL, BLADDER
C0279680|T047||CCS_10|TRANSITIONAL CELL CARCINOMA OF THE URINARY BLADDER
C0279680|T047||CCS_10|URINARY BLADDER TRANSITIONAL CELL CARCINOMA
C0279680|T047||CCS_10|URINARY BLADDER UROTHELIAL CARCINOMA
C0279680|T047||CCS_10|UROTHELIAL CARCINOMA OF THE URINARY BLADDER
C1336089|T047||CCS_10|NON-INVASIVE BLADDER UROTHELIAL CARCINOMA
C1336089|T047||CCS_10|BLADDER TRANSITIONAL CELL CARCINOMA STAGE 0
C1336089|T047||CCS_10|STAGE 0 BLADDER UROTHELIAL CARCINOMA AJCC V7
C1336089|T047||CCS_10|STAGE 0 BLADDER UROTHELIAL CARCINOMA AJCC V6
C1336089|T047||CCS_10|STAGE 0 TRANSITIONAL CELL CARCINOMA OF BLADDER
C1336089|T047||CCS_10|STAGE 0 TRANSITIONAL CELL CARCINOMA OF URINARY BLADDER
C1336089|T047||CCS_10|STAGE 0 TRANSITIONAL CELL CARCINOMA OF THE BLADDER
C1336089|T047||CCS_10|STAGE 0 TRANSITIONAL CELL CARCINOMA OF THE URINARY BLADDER
C1336089|T047||CCS_10|STAGE 0 URINARY BLADDER TRANSITIONAL CELL CARCINOMA
C1336089|T047||CCS_10|STAGE 0 BLADDER UROTHELIAL CARCINOMA
C1739113|T047||CCS_10|BLADDER TRANSITIONAL CELL CARCINOMA RECURRENT
C1336450|T047||CCS_10|BLADDER TRANSITIONAL CELL CARCINOMA STAGE I
C1336450|T047||CCS_10|STAGE I BLADDER UROTHELIAL CARCINOMA AJCC V6
C1336450|T047||CCS_10|STAGE I BLADDER UROTHELIAL CARCINOMA AJCC V7
C1336450|T047||CCS_10|STAGE I TRANSITIONAL CELL CARCINOMA OF BLADDER
C1336450|T047||CCS_10|STAGE I TRANSITIONAL CELL CARCINOMA OF URINARY BLADDER
C1336450|T047||CCS_10|STAGE I TRANSITIONAL CELL CARCINOMA OF THE BLADDER
C1336450|T047||CCS_10|STAGE I TRANSITIONAL CELL CARCINOMA OF THE URINARY BLADDER
C1336450|T047||CCS_10|STAGE I URINARY BLADDER TRANSITIONAL CELL CARCINOMA
C1336450|T047||CCS_10|STAGE I BLADDER UROTHELIAL CARCINOMA
C0862432|T047||CCS_10|BLADDER TRANSITIONAL CELL CARCINOMA STAGE IV
C0862432|T047||CCS_10|STAGE IV BLADDER UROTHELIAL CARCINOMA AJCC V7
C0862432|T047||CCS_10|TRANSITIONAL CELL CARCINOMA OF THE BLADDER STAGE IV
C0862432|T047||CCS_10|UROTHELIAL CARCINOMA BLADDER STAGE IV
C0862432|T047||CCS_10|STAGE IV TRANSITIONAL CELL CARCINOMA OF BLADDER
C0862432|T047||CCS_10|STAGE IV TRANSITIONAL CELL CARCINOMA OF URINARY BLADDER
C0862432|T047||CCS_10|STAGE IV TRANSITIONAL CELL CARCINOMA OF THE BLADDER
C0862432|T047||CCS_10|STAGE IV TRANSITIONAL CELL CARCINOMA OF THE URINARY BLADDER
C0862432|T047||CCS_10|STAGE IV URINARY BLADDER TRANSITIONAL CELL CARCINOMA
C0862432|T047||CCS_10|STAGE IV BLADDER UROTHELIAL CARCINOMA
C0862402|T047||CCS_10|BLADDER TRANSITIONAL CELL CARCINOMA STAGE II
C0862402|T047||CCS_10|STAGE II BLADDER UROTHELIAL CARCINOMA AJCC V6
C0862402|T047||CCS_10|STAGE II BLADDER UROTHELIAL CARCINOMA AJCC V7
C0862402|T047||CCS_10|UROTHELIAL CARCINOMA BLADDER STAGE II
C0862402|T047||CCS_10|TRANSITIONAL CELL CARCINOMA OF THE BLADDER STAGE II
C0862402|T047||CCS_10|STAGE II TRANSITIONAL CELL CARCINOMA OF BLADDER
C0862402|T047||CCS_10|STAGE II TRANSITIONAL CELL CARCINOMA OF URINARY BLADDER
C0862402|T047||CCS_10|STAGE II TRANSITIONAL CELL CARCINOMA OF THE BLADDER
C0862402|T047||CCS_10|STAGE II TRANSITIONAL CELL CARCINOMA OF THE URINARY BLADDER
C0862402|T047||CCS_10|STAGE II URINARY BLADDER TRANSITIONAL CELL CARCINOMA
C0862402|T047||CCS_10|STAGE II BLADDER UROTHELIAL CARCINOMA
C0862417|T047||CCS_10|BLADDER TRANSITIONAL CELL CARCINOMA STAGE III
C0862417|T047||CCS_10|STAGE III BLADDER UROTHELIAL CARCINOMA AJCC V7
C0862417|T047||CCS_10|STAGE III BLADDER UROTHELIAL CARCINOMA AJCC V6
C0862417|T047||CCS_10|TRANSITIONAL CELL CARCINOMA OF THE BLADDER STAGE III
C0862417|T047||CCS_10|UROTHELIAL CARCINOMA BLADDER STAGE III
C0862417|T047||CCS_10|STAGE III TRANSITIONAL CELL CARCINOMA OF BLADDER
C0862417|T047||CCS_10|STAGE III TRANSITIONAL CELL CARCINOMA OF URINARY BLADDER
C0862417|T047||CCS_10|STAGE III TRANSITIONAL CELL CARCINOMA OF THE BLADDER
C0862417|T047||CCS_10|STAGE III TRANSITIONAL CELL CARCINOMA OF THE URINARY BLADDER
C0862417|T047||CCS_10|STAGE III URINARY BLADDER TRANSITIONAL CELL CARCINOMA
C0862417|T047||CCS_10|STAGE III BLADDER UROTHELIAL CARCINOMA
C1297936|T047||CCS_10|MALIGNANT NEOPLASM BLADDER BY DIRECT EXTENSION FROM ENDOMETRIUM
C1297936|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING BLADDER BY DIRECT EXTENSION FROM ENDOMETRIUM 
C1297936|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING BLADDER BY DIRECT EXTENSION FROM ENDOMETRIUM
C1297936|T047||CCS_10|MALIGNANT TUMOR INVOLVING BLADDER BY DIRECT EXTENSION FROM ENDOMETRIUM 
C1297936|T047||CCS_10|MALIGNANT TUMOR INVOLVING BLADDER BY DIRECT EXTENSION FROM ENDOMETRIUM
C1297936|T047||CCS_10|MALIGNANT TUMOUR INVOLVING BLADDER BY DIRECT EXTENSION FROM ENDOMETRIUM
C1297937|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING BLADDER BY DIRECT EXTENSION FROM FALLOPIAN TUBE
C1297937|T047||CCS_10|MALIGNANT NEOPLASM BLADDER BY DIRECT EXTENSION FROM FALLOPIAN TUBE
C1297937|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING BLADDER BY DIRECT EXTENSION FROM FALLOPIAN TUBE 
C1297937|T047||CCS_10|MALIGNANT TUMOR INVOLVING BLADDER BY DIRECT EXTENSION FROM FALLOPIAN TUBE 
C1297937|T047||CCS_10|MALIGNANT TUMOR INVOLVING BLADDER BY DIRECT EXTENSION FROM FALLOPIAN TUBE
C1297937|T047||CCS_10|MALIGNANT TUMOUR INVOLVING BLADDER BY DIRECT EXTENSION FROM FALLOPIAN TUBE
C1297938|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING BLADDER BY DIRECT EXTENSION FROM OVARY 
C1297938|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING BLADDER BY DIRECT EXTENSION FROM OVARY
C1297938|T047||CCS_10|MALIGNANT NEOPLASM BLADDER BY DIRECT EXTENSION FROM OVARY
C1297938|T047||CCS_10|MALIGNANT TUMOR INVOLVING BLADDER BY DIRECT EXTENSION FROM OVARY 
C1297938|T047||CCS_10|MALIGNANT TUMOR INVOLVING BLADDER BY DIRECT EXTENSION FROM OVARY
C1297938|T047||CCS_10|MALIGNANT TUMOUR INVOLVING BLADDER BY DIRECT EXTENSION FROM OVARY
C1297939|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING BLADDER BY DIRECT EXTENSION FROM PROSTATE
C1297939|T047||CCS_10|MALIGNANT NEOPLASM BLADDER BY DIRECT EXTENSION FROM PROSTATE
C1297939|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING BLADDER BY DIRECT EXTENSION FROM PROSTATE 
C1297939|T047||CCS_10|MALIGNANT TUMOR INVOLVING BLADDER BY DIRECT EXTENSION FROM PROSTATE 
C1297939|T047||CCS_10|MALIGNANT TUMOR INVOLVING BLADDER BY DIRECT EXTENSION FROM PROSTATE
C1297939|T047||CCS_10|MALIGNANT TUMOUR INVOLVING BLADDER BY DIRECT EXTENSION FROM PROSTATE
C1297940|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING BLADDER BY DIRECT EXTENSION FROM UTERINE CERVIX
C1297940|T047||CCS_10|MALIGNANT NEOPLASM BLADDER BY DIRECT EXTENSION FROM UTERINE CERVIX
C1297940|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING BLADDER BY DIRECT EXTENSION FROM UTERINE CERVIX 
C1297940|T047||CCS_10|MALIGNANT TUMOR INVOLVING BLADDER BY DIRECT EXTENSION FROM UTERINE CERVIX 
C1297940|T047||CCS_10|MALIGNANT TUMOR INVOLVING BLADDER BY DIRECT EXTENSION FROM UTERINE CERVIX
C1297940|T047||CCS_10|MALIGNANT TUMOUR INVOLVING BLADDER BY DIRECT EXTENSION FROM UTERINE CERVIX
C1297941|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING BLADDER BY DIRECT EXTENSION FROM UTERUS
C1297941|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING BLADDER BY DIRECT EXTENSION FROM UTERUS 
C1297941|T047||CCS_10|MALIGNANT NEOPLASM BLADDER BY DIRECT EXTENSION FROM UTERUS
C1297941|T047||CCS_10|MALIGNANT TUMOR INVOLVING BLADDER BY DIRECT EXTENSION FROM UTERUS 
C1297941|T047||CCS_10|MALIGNANT TUMOR INVOLVING BLADDER BY DIRECT EXTENSION FROM UTERUS
C1297941|T047||CCS_10|MALIGNANT TUMOUR INVOLVING BLADDER BY DIRECT EXTENSION FROM UTERUS
C1297942|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING BLADDER BY DIRECT EXTENSION FROM VAGINA
C1297942|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING BLADDER BY DIRECT EXTENSION FROM VAGINA 
C1297942|T047||CCS_10|MALIGNANT NEOPLASM BLADDER BY DIRECT EXTENSION FROM VAGINA
C1297942|T047||CCS_10|MALIGNANT TUMOR INVOLVING BLADDER BY DIRECT EXTENSION FROM VAGINA 
C1297942|T047||CCS_10|MALIGNANT TUMOR INVOLVING BLADDER BY DIRECT EXTENSION FROM VAGINA
C1297942|T047||CCS_10|MALIGNANT TUMOUR INVOLVING BLADDER BY DIRECT EXTENSION FROM VAGINA
C2033201|T047||CCS_10|PAPILLARY CARCINOMA OF BLADDER 
C2033201|T047||CCS_10|PAPILLARY CARCINOMA OF BLADDER
C2212520|T047||CCS_10|MULLERIAN MIXED TUMOR OF BLADDER
C2212520|T047||CCS_10|MULLERIAN MIXED TUMOR OF BLADDER 
C2212529|T047||CCS_10|MALIGNANT MESODERMAL MIXED TUMOR OF BLADDER
C2212529|T047||CCS_10|MALIGNANT MESODERMAL MIXED TUMOR OF BLADDER 
C2212590|T047||CCS_10|MALIGNANT SMALL CELL NEOPLASM OF BLADDER 
C2212590|T047||CCS_10|MALIGNANT SMALL CELL NEOPLASM OF BLADDER
C2011424|T047||CCS_10|GIANT CELL TYPE NEOPLASM OF BLADDER
C2011424|T047||CCS_10|GIANT CELL TYPE NEOPLASM OF BLADDER 
C2018634|T047||CCS_10|SPINDLE CELL TYPE NEOPLASM OF BLADDER 
C2018634|T047||CCS_10|SPINDLE CELL TYPE NEOPLASM OF BLADDER
C2075593|T047||CCS_10|CLEAR CELL TYPE NEOPLASM OF BLADDER 
C2075593|T047||CCS_10|CLEAR CELL TYPE NEOPLASM OF BLADDER
C1334563|T047||CCS_10|MALIGNANT PARAGANGLIOMA OF BLADDER 
C1334563|T047||CCS_10|MALIGNANT PARAGANGLIOMA OF BLADDER
C1334563|T047||CCS_10|MALIGNANT BLADDER PARAGANGLIOMA
C1334563|T047||CCS_10|MALIGNANT PARAGANGLIOMA OF URINARY BLADDER
C1334563|T047||CCS_10|MALIGNANT PARAGANGLIOMA OF THE BLADDER
C1334563|T047||CCS_10|MALIGNANT PARAGANGLIOMA OF THE URINARY BLADDER
C1334563|T047||CCS_10|MALIGNANT URINARY BLADDER PARAGANGLIOMA
C2212603|T047||CCS_10|MYOSARCOMA OF BLADDER
C2212603|T047||CCS_10|MYOSARCOMA OF BLADDER 
C2212605|T047||CCS_10|FIBROUS HISTIOCYTOMA OF BLADDER 
C2212605|T047||CCS_10|FIBROUS HISTIOCYTOMA OF BLADDER
C0279682|T047||CCS_10|ADENOCARCINOMA OF BLADDER
C0279682|T047||CCS_10|ADENOCARCINOMA OF BLADDER 
C0279682|T047||CCS_10|BLADDER ADENOCARCINOMA
C0279682|T047||CCS_10|ADENOCARCINOMA OF BLADDER 
C0279682|T047||CCS_10|ADENOCARCINOMA OF THE BLADDER
C0279682|T047||CCS_10|ADENOCARCINOMA, BLADDER
C0279682|T047||CCS_10|BLADDER CANCER, ADENOCARCINOMA
C0279682|T047||CCS_10|ADENOCARCINOMA OF URINARY BLADDER
C0279682|T047||CCS_10|ADENOCARCINOMA OF THE URINARY BLADDER
C0279682|T047||CCS_10|URINARY BLADDER ADENOCARCINOMA
C0279682|T047||CCS_10|BLADDER ADENOCARCINOMA NOS
C0279682|T047||CCS_10|BLADDER ADENOCARCINOMA, NOS
C0279682|T047||CCS_10|BLADDER ADENOCARCINOMA, NOT OTHERWISE SPECIFIED
C2007062|T047||CCS_10|CARCINOSARCOMA OF BLADDER 
C2007062|T047||CCS_10|CARCINOSARCOMA OF BLADDER
C0349666|T047||CCS_10|SARCOMA OF BLADDER
C0349666|T047||CCS_10|SARCOMA OF BLADDER 
C0349666|T047||CCS_10|URINARY BLADDER SARCOMA
C0349666|T047||CCS_10|SARCOMA OF BLADDER 
C0349666|T047||CCS_10|SARCOMA OF URINARY BLADDER
C0349666|T047||CCS_10|SARCOMA OF THE BLADDER
C0349666|T047||CCS_10|SARCOMA OF THE URINARY BLADDER
C0349666|T047||CCS_10|BLADDER SARCOMA
C2212616|T047||CCS_10|FIBROSARCOMA OF BLADDER 
C2212616|T047||CCS_10|FIBROSARCOMA OF BLADDER
C2212627|T047||CCS_10|MALIGNANT MESENCHYMOMA OF BLADDER 
C2212627|T047||CCS_10|MALIGNANT MESENCHYMOMA OF BLADDER
C2212628|T047||CCS_10|MALIGNANT LYMPHOMA OF BLADDER 
C2212628|T047||CCS_10|MALIGNANT LYMPHOMA OF BLADDER
C2212659|T047||CCS_10|MALIGNANT PLASMACYTOMA OF BLADDER
C2212659|T047||CCS_10|MALIGNANT PLASMACYTOMA OF BLADDER 
C2212661|T047||CCS_10|MALIGNANT MASTOCYTOSIS OF BLADDER
C2212661|T047||CCS_10|MALIGNANT MASTOCYTOSIS OF BLADDER 
C2216667|T047||CCS_10|STAGING OF BLADDER CANCER
C2216667|T047||CCS_10|STAGING OF MALIGNANT NEOPLASM OF BLADDER 
C2216667|T047||CCS_10|STAGING OF MALIGNANT NEOPLASM OF BLADDER
C2216667|T047||CCS_10|MALIGNANT NEOPLASM OF BLADDER STAGING
C0699885|T047||CCS_10|CARCINOMA OF BLADDER
C0699885|T047||CCS_10|BLADDER CARCINOMA
C0699885|T047||CCS_10|CARCINOMA OF BLADDER 
C0699885|T047||CCS_10|CARCINOMA;BLADDER
C0699885|T047||CCS_10|CARCINOMA BLADDER
C0699885|T047||CCS_10|BLADDER CANCER
C0699885|T047||CCS_10|BLADDER CARCINOMA NOS
C0699885|T047||CCS_10|CARCINOMA URINARY BLADDER
C0699885|T047||CCS_10|URINARY BLADDER CARCINOMA
C0699885|T047||CCS_10|CARCINOMA OF BLADDER 
C0699885|T047||CCS_10|CARCINOMA OF THE BLADDER
C0699885|T047||CCS_10|CANCER OF BLADDER
C0699885|T047||CCS_10|CANCER OF THE BLADDER
C0699885|T047||CCS_10|URINARY BLADDER CANCER
C0699885|T047||CCS_10|CANCER OF THE URINARY BLADDER
C0699885|T047||CCS_10|CARCINOMA OF URINARY BLADDER
C0699885|T047||CCS_10|CARCINOMA OF THE URINARY BLADDER
C0699885|T047||CCS_10|CANCER OF URINARY BLADDER
C2212587|T047||CCS_10|NONINVASIVE PAPILLARY TRANSITIONAL CELL CARCINOMA IN SITU OF BLADDER
C2212587|T047||CCS_10|NONINVASIVE PAPILLARY TRANSITIONAL CELL CARCINOMA IN SITU OF BLADDER 
C2212587|T047||CCS_10|BLADDER CARCINOMA IN SITU PAPILLARY TRANSITIONAL CELL NONINVASIVE
C2212591|T047||CCS_10|SIGNET RING CELL CARCINOMA OF BLADDER 
C2212591|T047||CCS_10|SIGNET RING CELL CARCINOMA OF BLADDER
C2212592|T047||CCS_10|MALIGNANT EPITHELIOMA OF BLADDER 
C2212592|T047||CCS_10|MALIGNANT EPITHELIOMA OF BLADDER
C2111591|T047||CCS_10|LARGE CELL CARCINOMA OF BLADDER
C2111591|T047||CCS_10|LARGE CELL CARCINOMA OF BLADDER 
C2111710|T047||CCS_10|LARGE CELL NEUROENDOCRINE CARCINOMA OF BLADDER 
C2111710|T047||CCS_10|LARGE CELL NEUROENDOCRINE CARCINOMA OF BLADDER
C2111592|T047||CCS_10|LARGE CELL CARCINOMA OF BLADDER WITH RHABDOID PHENOTYPE
C2111592|T047||CCS_10|BLADDER MALIGNANT CARCINOMA LARGE CELL WITH RHABDOID PHENOTYPE
C2111592|T047||CCS_10|LARGE CELL CARCINOMA OF BLADDER WITH RHABDOID PHENOTYPE 
C2012070|T047||CCS_10|GLASSY CELL CARCINOMA OF BLADDER
C2012070|T047||CCS_10|GLASSY CELL CARCINOMA OF BLADDER 
C2188054|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF BLADDER 
C2188054|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF BLADDER
C2212593|T047||CCS_10|ANAPLASTIC CARCINOMA OF BLADDER 
C2212593|T047||CCS_10|ANAPLASTIC CARCINOMA OF BLADDER
C2082422|T047||CCS_10|PLEOMORPHIC CARCINOMA OF BLADDER 
C2082422|T047||CCS_10|PLEOMORPHIC CARCINOMA OF BLADDER
C2011242|T047||CCS_10|GIANT CELL CARCINOMA OF BLADDER 
C2011242|T047||CCS_10|GIANT CELL CARCINOMA OF BLADDER
C2018384|T047||CCS_10|SPINDLE CELL CARCINOMA OF BLADDER 
C2018384|T047||CCS_10|SPINDLE CELL CARCINOMA OF BLADDER
C2011207|T047||CCS_10|GIANT CELL AND SPINDLE CELL CARCINOMA OF BLADDER 
C2011207|T047||CCS_10|GIANT CELL AND SPINDLE CELL CARCINOMA OF BLADDER
C2142912|T047||CCS_10|PSEUDOSARCOMATOUS CARCINOMA OF BLADDER
C2142912|T047||CCS_10|PSEUDOSARCOMATOUS CARCINOMA OF BLADDER 
C2111794|T047||CCS_10|POLYGONAL CELL CARCINOMA OF BLADDER
C2111794|T047||CCS_10|POLYGONAL CELL CARCINOMA OF BLADDER 
C2007057|T047||CCS_10|CARCINOMA OF BLADDER WITH OSTEOCLAST-LIKE GIANT CELLS 
C2007057|T047||CCS_10|CARCINOMA OF BLADDER WITH OSTEOCLAST-LIKE GIANT CELLS
C2007057|T047||CCS_10|BLADDER CARCINOMA WITH OSTEOCLAST-LIKE GIANT CELLS
C2212594|T047||CCS_10|SMALL CELL CARCINOMA OF BLADDER 
C2212594|T047||CCS_10|SMALL CELL CARCINOMA OF BLADDER
C2009873|T047||CCS_10|FUSIFORM TYPE SMALL CELL CARCINOMA OF BLADDER 
C2009873|T047||CCS_10|FUSIFORM TYPE SMALL CELL CARCINOMA OF BLADDER
C2212595|T047||CCS_10|MEDULLARY CARCINOMA OF BLADDER 
C2212595|T047||CCS_10|MEDULLARY CARCINOMA OF BLADDER
C2033276|T047||CCS_10|PAPILLARY SQUAMOUS CELL CARCINOMA OF BLADDER
C2033276|T047||CCS_10|PAPILLARY SQUAMOUS CELL CARCINOMA OF BLADDER 
C1511208|T047||CCS_10|VERRUCOUS CARCINOMA OF BLADDER 
C1511208|T047||CCS_10|VERRUCOUS CARCINOMA OF BLADDER
C1511208|T047||CCS_10|BLADDER VERRUCOUS CARCINOMA
C1511208|T047||CCS_10|BLADDER VERRUCOUS SQUAMOUS CELL CARCINOMA
C2018592|T047||CCS_10|SPINDLE CELL TRANSITIONAL CELL CARCINOMA OF BLADDER
C2018592|T047||CCS_10|SPINDLE CELL TRANSITIONAL CELL CARCINOMA OF BLADDER 
C1735888|T047||CCS_10|PAPILLARY TRANSITIONAL CELL CARCINOMA OF BLADDER 
C1735888|T047||CCS_10|PAPILLARY TRANSITIONAL CELL CARCINOMA OF BLADDER
C2212600|T047||CCS_10|MICROPAPILLARY TRANSITIONAL CELL CARCINOMA OF BLADDER
C2212600|T047||CCS_10|MICROPAPILLARY TRANSITIONAL CELL CARCINOMA OF BLADDER 
C2212601|T047||CCS_10|SCHNEIDERIAN CARCINOMA OF BLADDER
C2212601|T047||CCS_10|SCHNEIDERIAN CARCINOMA OF BLADDER 
C2212602|T047||CCS_10|BASALOID CARCINOMA OF BLADDER
C2212602|T047||CCS_10|BASALOID CARCINOMA OF BLADDER 
C2075828|T047||CCS_10|CLOACOGENIC CARCINOMA OF BLADDER 
C2075828|T047||CCS_10|CLOACOGENIC CARCINOMA OF BLADDER
C2007045|T047||CCS_10|CARCINOMA SIMPLEX OF BLADDER 
C2007045|T047||CCS_10|CARCINOMA SIMPLEX OF BLADDER
C2012537|T047||CCS_10|GRANULAR CELL CARCINOMA OF BLADDER 
C2012537|T047||CCS_10|GRANULAR CELL CARCINOMA OF BLADDER
C2017446|T047||CCS_10|SOLID CARCINOMA OF BLADDER 
C2017446|T047||CCS_10|SOLID CARCINOMA OF BLADDER
C3203710|T047||CCS_10|BLADDER TRANSITIONAL CELL CARCINOMA METASTATIC
C2033152|T047||CCS_10|PAPILLARY CARCINOMA IN SITU OF BLADDER 
C2033152|T047||CCS_10|PAPILLARY CARCINOMA IN SITU OF BLADDER
C2212585|T047||CCS_10|BLADDER CARCINOMA IN SITU PAPILLARY SQUAMOUS CELL NONINVASIVE
C2212585|T047||CCS_10|NONINVASIVE PAPILLARY SQUAMOUS CELL CARCINOMA IN SITU OF BLADDER
C2212585|T047||CCS_10|NONINVASIVE PAPILLARY SQUAMOUS CELL CARCINOMA IN SITU OF BLADDER 
C2019360|T047||CCS_10|SQUAMOUS CELL CARCINOMA IN SITU OF BLADDER 
C2019360|T047||CCS_10|SQUAMOUS CELL CARCINOMA IN SITU OF BLADDER
C2212586|T047||CCS_10|BLADDER CIS SQUAMOUS CELL WITH QUESTIONABLE STROMAL INVASION
C2212586|T047||CCS_10|BLADDER CARCINOMA IN SITU SQUAMOUS CELL WITH QUESTIONABLE STROMAL INVASION
C2212586|T047||CCS_10|SQUAMOUS CELL CARCINOMA IN SITU OF BLADDER WITH QUESTIONABLE STROMAL INVASION 
C2212586|T047||CCS_10|SQUAMOUS CELL CARCINOMA IN SITU OF BLADDER WITH QUESTIONABLE STROMAL INVASION
C2145423|T047||CCS_10|TRANSITIONAL CELL CARCINOMA IN SITU OF BLADDER
C2145423|T047||CCS_10|TRANSITIONAL CELL CARCINOMA IN SITU OF BLADDER 
C2212589|T047||CCS_10|BLADDER ADENOCARCINOMA IN SITU IN VILLOUS ADENOMA
C2212589|T047||CCS_10|ADENOCARCINOMA IN SITU IN VILLOUS ADENOMA OF BLADDER
C2212589|T047||CCS_10|ADENOCARCINOMA IN SITU IN VILLOUS ADENOMA OF BLADDER 
C2199211|T047||CCS_10|DUCTAL CARCINOMA IN SITU OF BLADDER
C2199211|T047||CCS_10|DUCTAL CARCINOMA IN SITU OF BLADDER 
C0346893|T047||CCS_10|MALIGNANT NEOPLASM OF OTHER SITE OF URINARY BLADDER 
C0346893|T047||CCS_10|MALIGNANT NEOPLASM OF OTHER SITE OF URINARY BLADDER
C1314699|T047||CCS_10|BLADDER MALIGNANT NEOPLASM PRIMARY
C1314699|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF BLADDER 
C1314699|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF BLADDER
C1314699|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF BLADDER 
C1282481|T047||CCS_10|MALIGNANT NEOPLASM BLADDER, LOCAL RECURRENCE
C1282481|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT NEOPLASM OF BLADDER
C1282481|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT NEOPLASM OF BLADDER 
C1282481|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOR OF URINARY BLADDER 
C1282481|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOR OF URINARY BLADDER
C1282481|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOUR OF URINARY BLADDER
C0347011|T047||CCS_10|METASTATIC NEOPLASM TO THE BLADDER
C0347011|T047||CCS_10|METASTASIS TO BLADDER 
C0347011|T047||CCS_10|METASTASIS TO BLADDER
C0347011|T047||CCS_10|METASTASIS TO THE BLADDER
C0347011|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BLADDER
C0347011|T047||CCS_10|METASTASES TO BLADDER
C0347011|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM URINARY BLADDER
C0347011|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BLADDER 
C0347011|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO THE BLADDER
C0347011|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM IN THE BLADDER
C0347011|T047||CCS_10|CANCER METASTATIC TO URINARY BLADDER
C0347011|T047||CCS_10|METASTATIC TUMOR TO BLADDER
C0347011|T047||CCS_10|METASTATIC TUMOUR TO BLADDER
C0347011|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO BLADDER
C0347011|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BLADDER 
C0347011|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO BLADDER, NOS
C0347011|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BLADDER, NOS
C0347011|T047||CCS_10|METASTATIC NEOPLASM TO THE URINARY BLADDER
C0347011|T047||CCS_10|METASTATIC TUMOR TO THE BLADDER
C0347011|T047||CCS_10|METASTATIC TUMOR TO THE URINARY BLADDER
C3694329|T047||CCS_10|MALIGNANT NEOPLASM OF APEX OF BLADDER 
C3694329|T047||CCS_10|MALIGNANT NEOPLASM OF APEX OF BLADDER
C3694329|T047||CCS_10|MALIGNANT NEOPLASM BLADDER APEX
C1282497|T047||CCS_10|METASTASIS FROM MALIGNANT NEOPLASM OF BLADDER
C1282497|T047||CCS_10|METASTASIS FROM MALIGNANT NEOPLASM OF BLADDER 
C1282497|T047||CCS_10|METASTASIS FROM MALIGNANT TUMOR OF BLADDER 
C1282497|T047||CCS_10|METASTASIS FROM MALIGNANT TUMOR OF BLADDER
C1282497|T047||CCS_10|METASTASIS FROM MALIGNANT TUMOUR OF BLADDER
C3839273|T047||CCS_10|MALIGNANT NEOPLASM OF AUGMENTED BLADDER 
C3839273|T047||CCS_10|MALIGNANT NEOPLASM OF AUGMENTED BLADDER
C3839273|T047||CCS_10|MALIGNANT TUMOR OF AUGMENTED BLADDER
C3839273|T047||CCS_10|MALIGNANT TUMOUR OF AUGMENTED BLADDER
C4031688|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA NODULAR LYMPHOCYTIC PREDOMINANCE
C4031688|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA NODULAR LYMPHOCYTIC PREDOMINANCE 
C4031667|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA MANTLE CELL
C4031667|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA MANTLE CELL 
C4031656|T047||CCS_10|BIOPSY OF BLADDER SHOWED MASTOCYTOSIS
C4031656|T047||CCS_10|BIOPSY OF BLADDER SHOWED MASTOCYTOSIS 
C4031722|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SQUAMOUS CELL KERATINIZING 
C4031722|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SQUAMOUS CELL KERATINIZING
C4031707|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOSARCOMA EMBRYONAL TYPE
C4031707|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOSARCOMA EMBRYONAL TYPE 
C4031671|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA HISTIOCYTOSIS
C4031671|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA HISTIOCYTOSIS 
C4031670|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA LARGE B-CELL DIFFUSE
C4031670|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA LARGE B-CELL DIFFUSE 
C4031648|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA LEIOMYOSARCOMA EPITHELIOID
C4031648|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA LEIOMYOSARCOMA EPITHELIOID 
C4031736|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA PAPILLARY
C4031736|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA PAPILLARY 
C4031735|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA PAPILLARY SQUAMOUS CELL
C4031735|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA PAPILLARY SQUAMOUS CELL 
C4031714|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA TRANSITIONAL CELL MICROPAPILLARY 
C4031714|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA TRANSITIONAL CELL MICROPAPILLARY
C4031661|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA PRECURSOR CELL LYMPHOBLASTIC
C4031661|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA PRECURSOR CELL LYMPHOBLASTIC 
C4031655|T047||CCS_10|BIOPSY OF BLADDER SHOWED MESENCHYMOMA 
C4031655|T047||CCS_10|BIOPSY OF BLADDER SHOWED MESENCHYMOMA
C4031641|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA RHABDOMYOSARCOMA SPINDLE CELL 
C4031641|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA RHABDOMYOSARCOMA SPINDLE CELL
C4031628|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA FOLLICULAR DENDRITIC CELL 
C4031628|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA FOLLICULAR DENDRITIC CELL
C4031749|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA BASALOID 
C4031749|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA BASALOID
C4031717|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SQUAMOUS CELL WITH HORN FORMATION
C4031717|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SQUAMOUS CELL WITH HORN FORMATION 
C4031706|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOSARCOMA MYOEPITHELIOMA
C4031706|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOSARCOMA MYOEPITHELIOMA 
C4031703|T047||CCS_10|BIOPSY OF BLADDER SHOWED CLEAR CELL TYPE
C4031703|T047||CCS_10|BIOPSY OF BLADDER SHOWED CLEAR CELL TYPE 
C4031702|T047||CCS_10|BIOPSY OF BLADDER SHOWED FIBROSARCOMA
C4031702|T047||CCS_10|BIOPSY OF BLADDER SHOWED FIBROSARCOMA 
C4031691|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA LYMPHOCYTIC DEPLETION
C4031691|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA LYMPHOCYTIC DEPLETION 
C4031672|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA FOLLICULAR GRADE 3 
C4031672|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA FOLLICULAR GRADE 3
C4031652|T047||CCS_10|BIOPSY OF BLADDER SHOWED MULLERIAN MIXED TUMOR
C4031652|T047||CCS_10|BIOPSY OF BLADDER SHOWED MULLERIAN MIXED TUMOR 
C4031644|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA RHABDOMYOSARCOMA EMBRYONAL
C4031644|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA RHABDOMYOSARCOMA EMBRYONAL 
C4031640|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA RHABDOMYOSARCOMA WITH GANGLIONIC DIFFERENTIATION
C4031640|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA RHABDOMYOSARCOMA WITH GANGLIONIC DIFFERENTIATION 
C4031746|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA GIANT CELL 
C4031746|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA GIANT CELL
C4031745|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA GIANT SELL AND SPINDLE CELL
C4031745|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA GIANT SELL AND SPINDLE CELL 
C4031726|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SOLID 
C4031726|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SOLID
C4031695|T047||CCS_10|BIOPSY OF BLADDER SHOWED HEPATOID ADENOCARCINOMA 
C4031695|T047||CCS_10|BIOPSY OF BLADDER SHOWED ADENOCARCINOMA HEPATOID
C4031695|T047||CCS_10|BIOPSY OF BLADDER SHOWED HEPATOID ADENOCARCINOMA
C4031687|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA NODULAR SCLEROSIS
C4031687|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA NODULAR SCLEROSIS 
C4031677|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA BURKITT'S
C4031677|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA BURKITT'S 
C4031659|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA PRECURSOR CELL LYMPHOBLASTIC T-CELL
C4031659|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA PRECURSOR CELL LYMPHOBLASTIC T-CELL 
C4031647|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA LEIOMYOSARCOMA MYXOID 
C4031647|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA LEIOMYOSARCOMA MYXOID
C4031645|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA RHABDOMYOSARCOMA ALVEOLAR 
C4031645|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA RHABDOMYOSARCOMA ALVEOLAR
C4031627|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA GIANT CELL 
C4031627|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA GIANT CELL
C4031623|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA MAST CELL 
C4031623|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA MAST CELL
C4031728|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SMALL CELL 
C4031728|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SMALL CELL
C4031690|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA LYMPHOCYTIC DEPLETION RETICULAR
C4031690|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA LYMPHOCYTIC DEPLETION RETICULAR 
C4031686|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA NODULAR SCLEROSIS CELLULAR PHASE
C4031686|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA NODULAR SCLEROSIS CELLULAR PHASE 
C4031683|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA SARCOMA
C4031683|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA SARCOMA 
C4031674|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA FOLLICULAR GRADE 1 
C4031674|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA FOLLICULAR GRADE 1
C4031669|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA LARGE B-CELL DIFFUSE IMMUNOBLASTIC 
C4031669|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA LARGE B-CELL DIFFUSE IMMUNOBLASTIC
C4031651|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA
C4031651|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA 
C4031634|T047||CCS_10|BIOPSY OF BLADDER SHOWED PLASMACYTOMA
C4031634|T047||CCS_10|BIOPSY OF BLADDER SHOWED PLASMACYTOMA 
C4031632|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA 
C4031632|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA
C4031625|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA INTERDIGITATING DENDRITIC CELL 
C4031625|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA INTERDIGITATING DENDRITIC CELL
C4031620|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA UNDIFFERENTIATED
C4031620|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA UNDIFFERENTIATED 
C4031730|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SIGNET RING CELL
C4031730|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SIGNET RING CELL 
C4031729|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SIMPLEX
C4031729|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SIMPLEX 
C4031701|T047||CCS_10|BIOPSY OF BLADDER SHOWED FIBROSARCOMA FASCIAL
C4031701|T047||CCS_10|BIOPSY OF BLADDER SHOWED FIBROSARCOMA FASCIAL 
C4031697|T047||CCS_10|BIOPSY OF BLADDER SHOWED FIBROUS HISTIOCYTOMA 
C4031697|T047||CCS_10|BIOPSY OF BLADDER SHOWED FIBROUS HISTIOCYTOMA
C4031668|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA LYMPHOPLASMACYTIC 
C4031668|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA LYMPHOPLASMACYTIC
C4031630|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA EMBRYONAL 
C4031630|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA EMBRYONAL
C4031626|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA HISTIOCYTIC
C4031626|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA HISTIOCYTIC 
C4031621|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA SPINDLE CELL 
C4031621|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA SPINDLE CELL
C4031750|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA ANAPLASTIC
C4031750|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA ANAPLASTIC 
C4031743|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA GRANULAR CELL 
C4031743|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA GRANULAR CELL
C4031739|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA LARGE CELL NEUROENDOCRINE
C4031739|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA LARGE CELL NEUROENDOCRINE 
C4031737|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA MEDULLARY
C4031737|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA MEDULLARY 
C4031732|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA PSEUDOSARCOMATOUS
C4031732|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA PSEUDOSARCOMATOUS 
C4031719|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SQUAMOUS CELL SMALL CELL, NONKERATINIZING 
C4031719|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SQUAMOUS CELL SMALL CELL, NONKERATINIZING
C4031698|T047||CCS_10|BIOPSY OF BLADDER SHOWED FIBROSARCOMA SOLITARY FIBROUS TUMOR
C4031698|T047||CCS_10|BIOPSY OF BLADDER SHOWED FIBROSARCOMA SOLITARY FIBROUS TUMOR 
C4031684|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA NODULAR SCLEROSIS GRADE 2 
C4031684|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA NODULAR SCLEROSIS GRADE 2
C4031675|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA FOLLICULAR
C4031675|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA FOLLICULAR 
C4031633|T047||CCS_10|BIOPSY OF BLADDER SHOWED PLASMACYTOMA EXTRAMEDULLARY
C4031633|T047||CCS_10|BIOPSY OF BLADDER SHOWED PLASMACYTOMA EXTRAMEDULLARY 
C4031624|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA LANGERHANS CELL 
C4031624|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA LANGERHANS CELL
C4031725|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SPINDLE CELL 
C4031725|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SPINDLE CELL
C4031700|T047||CCS_10|BIOPSY OF BLADDER SHOWED FIBROSARCOMA FIBROMYXOSARCOMA 
C4031700|T047||CCS_10|BIOPSY OF BLADDER SHOWED FIBROSARCOMA FIBROMYXOSARCOMA
C4031681|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA 
C4031681|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA
C4031666|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA MARGINAL ZONE B-CELL 
C4031666|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA MARGINAL ZONE B-CELL
C4031664|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA MATURE T-CELL ANGIOIMMUNOBLASTIC 
C4031664|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA MATURE T-CELL ANGIOIMMUNOBLASTIC
C4031657|T047||CCS_10|BIOPSY OF BLADDER SHOWED MALIGNANT NEOPLASM
C4031657|T047||CCS_10|BIOPSY OF BLADDER SHOWED MALIGNANT NEOPLASM 
C4031654|T047||CCS_10|BIOPSY OF BLADDER SHOWED MESODERMAL MIXED TUMOR
C4031654|T047||CCS_10|BIOPSY OF BLADDER SHOWED MESODERMAL MIXED TUMOR 
C4031619|T047||CCS_10|BIOPSY OF BLADDER SHOWED SMALL CELL TYPE 
C4031619|T047||CCS_10|BIOPSY OF BLADDER SHOWED SMALL CELL TYPE
C4031616|T047||CCS_10|BIOPSY OF BLADDER SHOWED SPINDLE CELL TYPE
C4031616|T047||CCS_10|BIOPSY OF BLADDER SHOWED SPINDLE CELL TYPE 
C4031738|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA LARGE CELL WITH RHABDOID PHENOTYPE
C4031738|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA LARGE CELL WITH RHABDOID PHENOTYPE 
C4031694|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA
C4031694|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA 
C4031660|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA PRECURSOR CELL LYMPHOBLASTIC B-CELL 
C4031660|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA PRECURSOR CELL LYMPHOBLASTIC B-CELL
C4031635|T047||CCS_10|BIOPSY OF BLADDER SHOWED PARAGANGLIOMA 
C4031635|T047||CCS_10|BIOPSY OF BLADDER SHOWED PARAGANGLIOMA
C4031631|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA DESMOPLASTIC SMALL ROUND CELL TUMOR 
C4031631|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA DESMOPLASTIC SMALL ROUND CELL TUMOR
C4031744|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA GLASSY CELL
C4031744|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA GLASSY CELL 
C4031740|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA LARGE CELL 
C4031740|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA LARGE CELL
C4031721|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SQUAMOUS CELL LARGE CELL, NONKERATINIZING 
C4031721|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SQUAMOUS CELL LARGE CELL, NONKERATINIZING
C4031720|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SQUAMOUS CELL MICROINVASIVE
C4031720|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SQUAMOUS CELL MICROINVASIVE 
C4031712|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA TRANSITIONAL CELL SPINDLE CELL
C4031712|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA TRANSITIONAL CELL SPINDLE CELL 
C4031710|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA VERRUCOUS
C4031710|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA VERRUCOUS 
C4031693|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA GRANULOMA 
C4031693|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA GRANULOMA
C4031692|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA LYMPHOCYTE-RICH 
C4031692|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA LYMPHOCYTE-RICH
C4031642|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA RHABDOMYOSARCOMA PLEOMORPHIC, ADULT TYPE 
C4031642|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA RHABDOMYOSARCOMA PLEOMORPHIC, ADULT TYPE
C4031639|T047||CCS_10|BIOPSY OF BLADDER SHOWED NON-HODGKIN'S LYMPHOMA 
C4031639|T047||CCS_10|BIOPSY OF BLADDER SHOWED NON-HODGKIN'S LYMPHOMA
C4031731|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SCHNEIDERIAN 
C4031731|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SCHNEIDERIAN
C4031727|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SMALL CELL FUSIFORM CELL 
C4031727|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SMALL CELL FUSIFORM CELL
C4031713|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA TRANSITIONAL CELL PAPILLARY
C4031713|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA TRANSITIONAL CELL PAPILLARY 
C4031699|T047||CCS_10|BIOPSY OF BLADDER SHOWED FIBROSARCOMA INFANTILE
C4031699|T047||CCS_10|BIOPSY OF BLADDER SHOWED FIBROSARCOMA INFANTILE 
C4031673|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA FOLLICULAR GRADE 2 
C4031673|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA FOLLICULAR GRADE 2
C4031665|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA MATURE T-CELL
C4031665|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA MATURE T-CELL 
C4031646|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA RHABDOMYOSARCOMA
C4031646|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA RHABDOMYOSARCOMA 
C4031748|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA CLOACOGENIC
C4031748|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA CLOACOGENIC 
C4031747|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA EPITHELIOMA
C4031747|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA EPITHELIOMA 
C4031724|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SQUAMOUS CELL 
C4031724|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SQUAMOUS CELL
C4031711|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA UNDIFFERENTIATED 
C4031711|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA UNDIFFERENTIATED
C4031709|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA WITH OSTEOCLAST-LIKE GIANT CELLS
C4031709|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA WITH OSTEOCLAST-LIKE GIANT CELLS 
C4031696|T047||CCS_10|BIOPSY OF BLADDER SHOWED GIANT CELL TYPE 
C4031696|T047||CCS_10|BIOPSY OF BLADDER SHOWED GIANT CELL TYPE
C4031663|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA MIXED SMALL AND LARGE CELL, DIFFUSE
C4031663|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA MIXED SMALL AND LARGE CELL, DIFFUSE 
C4031649|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA LEIOMYOSARCOMA
C4031649|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA LEIOMYOSARCOMA 
C4031658|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA SMALL B-CELL LYMPHOCYTIC
C4031658|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA SMALL B-CELL LYMPHOCYTIC 
C4031643|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA RHABDOMYOSARCOMA MIXED TYPE 
C4031643|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA RHABDOMYOSARCOMA MIXED TYPE
C4031734|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA PLEOMORPHIC
C4031734|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA PLEOMORPHIC 
C4031723|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SQUAMOUS CELL ADENOID 
C4031723|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SQUAMOUS CELL ADENOID
C4031685|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA NODULAR SCLEROSIS GRADE 1
C4031685|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA NODULAR SCLEROSIS GRADE 1 
C4031629|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA EPITHELIOID
C4031629|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA EPITHELIOID 
C4031733|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA POLYGONAL CELL
C4031733|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA POLYGONAL CELL 
C4031718|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SQUAMOUS CELL SPINDLE CELL
C4031718|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA SQUAMOUS CELL SPINDLE CELL 
C4031715|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA TRANSITIONAL CELL 
C4031715|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOMA TRANSITIONAL CELL
C4031708|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOSARCOMA
C4031708|T047||CCS_10|BIOPSY OF BLADDER SHOWED CARCINOSARCOMA 
C4031682|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA WITH LYMPHOCYTIC DEPLETION WITH DIFFUSE FIBROSIS 
C4031682|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA WITH LYMPHOCYTIC DEPLETION WITH DIFFUSE FIBROSIS
C4031689|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA MIXED CELLULARITY 
C4031689|T047||CCS_10|BIOPSY OF BLADDER SHOWED HODGKIN'S LYMPHOMA MIXED CELLULARITY
C4031676|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA COMPOSITE HODGKIN'S AND NON-HODGKIN'S 
C4031676|T047||CCS_10|BIOPSY OF BLADDER SHOWED LYMPHOMA COMPOSITE HODGKIN'S AND NON-HODGKIN'S
C4031650|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA ANGIOMYOSARCOMA 
C4031650|T047||CCS_10|BIOPSY OF BLADDER SHOWED MYOSARCOMA ANGIOMYOSARCOMA
C4031622|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA SMALL CELL
C4031622|T047||CCS_10|BIOPSY OF BLADDER SHOWED SARCOMA SMALL CELL 
C0279681|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF BLADDER 
C0279681|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF BLADDER
C0279681|T047||CCS_10|BLADDER SQUAMOUS CELL CARCINOMA
C0279681|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF BLADDER 
C0279681|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE BLADDER
C0279681|T047||CCS_10|BLADDER CANCER, SQUAMOUS CELL CARCINOMA
C0279681|T047||CCS_10|CARCINOMA, SQUAMOUS CELL, BLADDER
C0279681|T047||CCS_10|EPIDERMOID CARCINOMA OF BLADDER
C0279681|T047||CCS_10|EPIDERMOID CARCINOMA OF URINARY BLADDER
C0279681|T047||CCS_10|EPIDERMOID CARCINOMA OF THE BLADDER
C0279681|T047||CCS_10|EPIDERMOID CARCINOMA OF THE URINARY BLADDER
C0279681|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF URINARY BLADDER
C0279681|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE URINARY BLADDER
C0279681|T047||CCS_10|URINARY BLADDER EPIDERMOID CARCINOMA
C0279681|T047||CCS_10|URINARY BLADDER SQUAMOUS CELL CARCINOMA
C0279681|T047||CCS_10|BLADDER EPIDERMOID CARCINOMA
C1827293|T047||CCS_10|CARCINOMA OF URINARY BLADDER, INVASIVE 
C1827293|T047||CCS_10|CARCINOMA OF URINARY BLADDER, INVASIVE
C1827293|T047||CCS_10|CARCINOMA OF BLADDER, INVASIVE
C1827293|T047||CCS_10|CARCINOMA OF BLADDER, INVASIVE 
C1827293|T047||CCS_10|BLADDER MALIGNANT CARCINOMA INVASIVE
C1827293|T047||CCS_10|INVASIVE BLADDER CANCER
C0153616|T047||CCS_10|MALIGNANT NEOPLASM OF OTHER SPECIFIED SITES OF BLADDER
C0153616|T047||CCS_10|MALIG NEO BLADDER NEC
C0864967|T047||CCS_10|MALIGNANT NEOPLASM OF BLADDER WALL NOS
C1336527|T047||CCS_10|CARCINOMA OF URINARY BLADDER, SUPERFICIAL 
C1336527|T047||CCS_10|CARCINOMA OF URINARY BLADDER, SUPERFICIAL
C1336527|T047||CCS_10|CARCINOMA OF BLADDER, SUPERFICIAL 
C1336527|T047||CCS_10|BLADDER MALIGNANT CARCINOMA SUPERFICIAL
C1336527|T047||CCS_10|CARCINOMA OF BLADDER, SUPERFICIAL
C1336527|T047||CCS_10|SUPERFICIAL BLADDER CARCINOMA
C1336527|T047||CCS_10|SUPERFICIAL BLADDER CANCER
C1336527|T047||CCS_10|SUPERFICIAL URINARY BLADDER CANCER
C1336527|T047||CCS_10|SUPERFICIAL URINARY BLADDER CARCINOMA
C0280218|T047||CCS_10|STAGE, BLADDER CANCER
C0280218|T047||CCS_10|BLADDER CANCER STAGE
C0279879|T047||CCS_10|CELLULAR DIAGNOSIS, BLADDER CANCER
C0279879|T047||CCS_10|BLADDER CANCER CELLULAR DIAGNOSIS
C1332561|T047||CCS_10|PRIMARY BLADDER LYMPHOMA
C1332561|T047||CCS_10|LYMPHOMA OF BLADDER
C1332561|T047||CCS_10|LYMPHOMA OF URINARY BLADDER
C1332561|T047||CCS_10|LYMPHOMA OF THE BLADDER
C1332561|T047||CCS_10|LYMPHOMA OF THE URINARY BLADDER
C1332561|T047||CCS_10|URINARY BLADDER LYMPHOMA
C1332561|T047||CCS_10|BLADDER LYMPHOMA
C0862326|T047||CCS_10|MALIGNANT NEOPLASM OF BLADDER RECURRENT
C0862326|T047||CCS_10|RECURRENT MALIGNANT BLADDER NEOPLASM
C1276593|T047||CCS_10|T3B: BLADDER TUMOR INVADES PERIVESICAL TISSUE MACROSCOPICALLY (EXTRAVESICULAR MASS) 
C1276593|T047||CCS_10|T3B: BLADDER TUMOR INVADES PERIVESICAL TISSUE MACROSCOPICALLY (EXTRAVESICULAR MASS)
C1276593|T047||CCS_10|T3B: BLADDER TUMOUR INVADES PERIVESICAL TISSUE MACROSCOPICALLY (EXTRAVESICULAR MASS)
C1276593|T047||CCS_10|T3B: BLADDER TUMOR INVADES PERIVESICAL TISSUE MACROSCOPICALLY (EXTRAVESICULAR MASS) (TUMOR STAGING)
C1276588|T047||CCS_10|T2B: URINARY BLADDER TUMOR INVADES DEEP MUSCLE (OUTER HALF) 
C1276588|T047||CCS_10|T2B: URINARY BLADDER TUMOR INVADES DEEP MUSCLE (OUTER HALF)
C1276588|T047||CCS_10|T2B: URINARY BLADDER TUMOUR INVADES DEEP MUSCLE (OUTER HALF)
C1276588|T047||CCS_10|T2B: URINARY BLADDER TUMOR INVADES DEEP MUSCLE (OUTER HALF) (TUMOR STAGING)
C0349659|T047||CCS_10|RHABDOMYOSARCOMA OF BLADDER 
C0349659|T047||CCS_10|RHABDOMYOSARCOMA OF BLADDER
C0349659|T047||CCS_10|RHABDOMYOSARCOMA OF URINARY BLADDER
C0349659|T047||CCS_10|RHABDOMYOSARCOMA OF BLADDER 
C1276587|T047||CCS_10|T2A: URINARY BLADDER TUMOR INVADES SUPERFICIAL MUSCLE (INNER HALF) 
C1276587|T047||CCS_10|T2A: URINARY BLADDER TUMOR INVADES SUPERFICIAL MUSCLE (INNER HALF)
C1276587|T047||CCS_10|T2A: URINARY BLADDER TUMOUR INVADES SUPERFICIAL MUSCLE (INNER HALF)
C1276587|T047||CCS_10|T2A: URINARY BLADDER TUMOR INVADES SUPERFICIAL MUSCLE (INNER HALF) (TUMOR STAGING)
C1276592|T047||CCS_10|T3A: BLADDER TUMOR INVADES PERIVESICAL TISSUE MICROSCOPICALLY 
C1276592|T047||CCS_10|T3A: BLADDER TUMOR INVADES PERIVESICAL TISSUE MICROSCOPICALLY
C1276592|T047||CCS_10|T3A: BLADDER TUMOUR INVADES PERIVESICAL TISSUE MICROSCOPICALLY
C1276592|T047||CCS_10|T3A: BLADDER TUMOR INVADES PERIVESICAL TISSUE MICROSCOPICALLY (TUMOR STAGING)
C1276591|T047||CCS_10|T3: URINARY BLADDER TUMOR INVADES PERIVESICAL TISSUE 
C1276591|T047||CCS_10|T3: URINARY BLADDER TUMOR INVADES PERIVESICAL TISSUE
C1276591|T047||CCS_10|T3: URINARY BLADDER TUMOUR INVADES PERIVESICAL TISSUE
C1276591|T047||CCS_10|T3: URINARY BLADDER TUMOR INVADES PERIVESICAL TISSUE (TUMOR STAGING)
C2212650|T047||CCS_10|GRADE 3 FOLLICULAR LYMPHOMA OF BLADDER
C2212650|T047||CCS_10|GRADE 3 FOLLICULAR LYMPHOMA OF BLADDER 
C2212657|T047||CCS_10|NK/T-CELL LYMPHOMA OF BLADDER
C2212657|T047||CCS_10|NK/T-CELL LYMPHOMA OF BLADDER 
C2212631|T047||CCS_10|MIXED CELLULARITY HODGKIN'S LYMPHOMA OF BLADDER 
C2212631|T047||CCS_10|MIXED CELLULARITY HODGKIN'S LYMPHOMA OF BLADDER
C2046544|T047||CCS_10|HODGKIN'S GRANULOMA OF BLADDER 
C2046544|T047||CCS_10|HODGKIN'S GRANULOMA OF BLADDER
C2046684|T047||CCS_10|HODGKIN'S SARCOMA OF BLADDER 
C2046684|T047||CCS_10|HODGKIN'S SARCOMA OF BLADDER
C2212640|T047||CCS_10|SMALL B-CELL LYMPHOCYTIC LYMPHOMA OF BLADDER
C2212640|T047||CCS_10|SMALL B-CELL LYMPHOCYTIC LYMPHOMA OF BLADDER 
C2212649|T047||CCS_10|GRADE 2 FOLLICULAR LYMPHOMA OF BLADDER
C2212649|T047||CCS_10|GRADE 2 FOLLICULAR LYMPHOMA OF BLADDER 
C2212651|T047||CCS_10|MARGINAL ZONE B-CELL LYMPHOMA OF BLADDER
C2212651|T047||CCS_10|MARGINAL ZONE B-CELL LYMPHOMA OF BLADDER 
C2212653|T047||CCS_10|ANGIOIMMUNOBLASTIC T-CELL LYMPHOMA OF BLADDER 
C2212653|T047||CCS_10|ANGIOIMMUNOBLASTIC T-CELL LYMPHOMA OF BLADDER
C2212653|T047||CCS_10|ANGIOIMMUNOBLASTIC LYMPHADENOPATHY WITH DYSPROTEINEMIA (AILD) OF BLADDER
C2212662|T047||CCS_10|SEZARY SYNDROME OF BLADDER
C2212662|T047||CCS_10|SEZARY SYNDROME OF BLADDER 
C2046471|T047||CCS_10|BLADDER MALIGNANT LYMPHOMA HODGKIN'S AND NON-HODGKIN'S
C2046471|T047||CCS_10|COMPOSITE HODGKIN'S AND NON-HODGKIN'S LYMPHOMA OF BLADDER
C2046471|T047||CCS_10|COMPOSITE HODGKIN'S AND NON-HODGKIN'S LYMPHOMA OF BLADDER 
C2212644|T047||CCS_10|LARGE B-CELL DIFFUSE LYMPHOMA OF BLADDER 
C2212644|T047||CCS_10|LARGE B-CELL DIFFUSE LYMPHOMA OF BLADDER
C2113746|T047||CCS_10|PRECURSOR T-CELL LYMPHOBLASTIC LYMPHOMA OF BLADDER 
C2113746|T047||CCS_10|PRECURSOR T-CELL LYMPHOBLASTIC LYMPHOMA OF BLADDER
C2212614|T047||CCS_10|MAST CELL SARCOMA OF BLADDER 
C2212614|T047||CCS_10|MAST CELL SARCOMA OF BLADDER
C2212656|T047||CCS_10|ANAPLASTIC LARGE CELL LYMPHOMA, NULL CELL TYPE OF BLADDER
C2212656|T047||CCS_10|ANAPLASTIC LARGE CELL LYMPHOMA, NULL CELL TYPE OF BLADDER 
C2212641|T047||CCS_10|LYMPHOPLASMACYTIC LYMPHOMA OF BLADDER 
C2212641|T047||CCS_10|LYMPHOPLASMACYTIC LYMPHOMA OF BLADDER
C2212652|T047||CCS_10|MATURE T-CELL LYMPHOMA OF BLADDER 
C2212652|T047||CCS_10|MATURE T-CELL LYMPHOMA OF BLADDER
C2113675|T047||CCS_10|PRECURSOR CELL LYMPHOBLASTIC LYMPHOMA OF BLADDER
C2113675|T047||CCS_10|PRECURSOR CELL LYMPHOBLASTIC LYMPHOMA OF BLADDER 
C2212630|T047||CCS_10|LYMPHOCYTE-RICH HODGKIN'S LYMPHOMA OF BLADDER 
C2212630|T047||CCS_10|LYMPHOCYTE-RICH HODGKIN'S LYMPHOMA OF BLADDER
C2212642|T047||CCS_10|MANTLE CELL LYMPHOMA OF BLADDER
C2212642|T047||CCS_10|MANTLE CELL LYMPHOMA OF BLADDER 
C2212643|T047||CCS_10|MIXED SMALL AND LARGE CELL DIFFUSE LYMPHOMA OF BLADDER
C2212643|T047||CCS_10|MIXED SMALL AND LARGE CELL DIFFUSE LYMPHOMA OF BLADDER 
C2212647|T047||CCS_10|FOLLICULAR LYMPHOMA OF BLADDER 
C2212647|T047||CCS_10|FOLLICULAR LYMPHOMA OF BLADDER
C2212648|T047||CCS_10|GRADE 1 FOLLICULAR LYMPHOMA OF BLADDER
C2212648|T047||CCS_10|GRADE 1 FOLLICULAR LYMPHOMA OF BLADDER 
C2113606|T047||CCS_10|PRECURSOR B-CELL LYMPHOBLASTIC LYMPHOMA OF BLADDER
C2113606|T047||CCS_10|PRECURSOR B-CELL LYMPHOBLASTIC LYMPHOMA OF BLADDER 
C2212658|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF BLADDER 
C2212658|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF BLADDER
C0279565|T047||CCS_10|INVASIVE LOBULAR BREAST CARCINOMA
C0279565|T047||CCS_10|LOBULAR BREAST CARCINOMA INVASIVE
C0279565|T047||CCS_10|LOBULAR INVASIVE BREAST CARCINOMA
C0279565|T047||CCS_10|CARCINOMA; INFILTRATING LOBULAR, UNSPECIFIED SITE
C0279565|T047||CCS_10|INFILTRATING; LOBULAR CARCINOMA, UNSPECIFIED SITE
C0279565|T047||CCS_10|CLASSIC INVASIVE LOBULAR CARCINOMA
C0279565|T047||CCS_10|INFILTRATING LOBULAR ADENOCARCINOMA
C0279565|T047||CCS_10|INFILTRATING LOBULAR BREAST CARCINOMA
C0279565|T047||CCS_10|INFILTRATING LOBULAR CARCINOMA OF BREAST
C0279565|T047||CCS_10|INFILTRATING LOBULAR CARCINOMA OF THE BREAST
C0279565|T047||CCS_10|INVASIVE LOBULAR ADENOCARCINOMA
C0279565|T047||CCS_10|INVASIVE LOBULAR CARCINOMA OF BREAST
C0279565|T047||CCS_10|INVASIVE LOBULAR CARCINOMA OF THE BREAST
C0279565|T047||CCS_10|INVASIVE LOBULAR CARCINOMA, CLASSIC TYPE
C0279565|T047||CCS_10|INVASIVE LOBULAR CARCINOMA
C0281267|T047||CCS_10|BILATERAL BREAST CANCER
C0281267|T047||CCS_10|BILATERAL BREAST CARCINOMA
C0242787|T047||CCS_10|MALIGNANT NEOPLASM OF MALE BREAST
C0242787|T047||CCS_10|MALIGNANT NEOPLASM OF MALE BREAST 
C0242787|T047||CCS_10|MALIGNANT MALE BREAST NEOPLASM
C0242787|T047||CCS_10|MALIGNANT TUMOR OF MALE BREAST
C0242787|T047||CCS_10|MALIGNANT NEOPLASM OF MALE BREAST 
C0242787|T047||CCS_10|MALIGNANT NEOPLASM OF MALE BREAST NOS
C0242787|T047||CCS_10|MALIGNANT NEOPLASM OF MALE BREAST NOS 
C0242787|T047||CCS_10|BREAST NEOPLASM MALIGNANT MALE
C0242787|T047||CCS_10|MALIGNANT BREAST NEOPLASM MALE
C0242787|T047||CCS_10|MALIGNANT NEOPLASM OF MALE BREAST, NOS
C0242787|T047||CCS_10|NEOPLASM MALIG;BREAST:M
C0242787|T047||CCS_10|MALIGNANT NEOSPLASM OF THE MALE BREAST
C0496812|T047||CCS_10|AXILLARY TAIL OF BREAST
C0496812|T047||CCS_10|MALIGNANT NEOPLASM OF AXILLARY TAIL OF BREAST
C0496812|T047||CCS_10|BREAST NEOPLASM MALIGNANT AXILLARY TAIL
C0496812|T047||CCS_10|MALIGNANT NEOPLASM OF AXILLARY TAIL OF BREAST 
C0496812|T047||CCS_10|CA BREAST - AXILLARY TAIL 
C0496812|T047||CCS_10|CA BREAST - AXILLARY TAIL
C0496812|T047||CCS_10|MALIGNANT NEOPLASM OF AXILLARY TAIL OF BREAST 
C0496807|T047||CCS_10|MALIGNANT NEOPLASM OF CENTRAL PORTION OF BREAST
C0496807|T047||CCS_10|MALIGNANT NEOPLASM OF CENTRAL PORTION OF BREAST 
C0496807|T047||CCS_10|BREAST NEOPLASM MALIGNANT CENTRAL PORTION
C0006142|T047||CCS_10|CANCER, BREAST
C0006142|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST
C0006142|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST, UNSPECIFIED
C0006142|T047||CCS_10|BREAST CANCER
C0006142|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST 
C0006142|T047||CCS_10|BREAST CANCER 
C0006142|T047||CCS_10|MALIGNANT BREAST NEOPLASM
C0006142|T047||CCS_10|CA BREAST
C0006142|T047||CCS_10|CANCER OF BREAST
C0006142|T047||CCS_10|MALIGNANT TUMOR OF BREAST
C0006142|T047||CCS_10|MALIGNANT NEOPLASMS OF BREAST (C50)
C0006142|T047||CCS_10|CA BREAST - NOS
C0006142|T047||CCS_10|CA BREAST - NOS 
C0006142|T047||CCS_10|[X]MALIGNANT NEOPLASM OF BREAST 
C0006142|T047||CCS_10|[X]MALIGNANT NEOPLASM OF BREAST
C0006142|T047||CCS_10|BREAST--CANCER
C0006142|T047||CCS_10|-- BREAST CANCER
C0006142|T047||CCS_10|BREAST CANCER STAGE UNSPECIFIED
C0006142|T047||CCS_10|BREAST CANCER NOS
C0006142|T047||CCS_10|BREAST TUMOR MALIGNANT
C0006142|T047||CCS_10|BREAST TUMOUR MALIGNANT
C0006142|T047||CCS_10|MAMMARY CANCER
C0006142|T047||CCS_10|CANCER OF THE BREAST
C0006142|T047||CCS_10|BREAST CARCINOMA
C0006142|T047||CCS_10|CA - BREAST CANCER
C0006142|T047||CCS_10|MALIGNANT TUMOUR OF BREAST
C0006142|T047||CCS_10|MALIGNANT TUMOR OF BREAST 
C0006142|T047||CCS_10|MALIGNANT BREAST TUMOR
C0006142|T047||CCS_10|MALIGNANT NEOPLASM OF THE BREAST
C0006142|T047||CCS_10|MALIGNANT TUMOR OF THE BREAST
C0496809|T047||CCS_10|MALIGNANT NEOPLASM OF LOWER-INNER QUADRANT OF BREAST
C0496809|T047||CCS_10|MALIGNANT NEOPLASM OF LOWER INNER QUADRANT OF BREAST 
C0496809|T047||CCS_10|BREAST NEOPLASM MALIGNANT LOWER INNER QUADRANT
C0496809|T047||CCS_10|MALIGNANT NEOPLASM OF LOWER INNER QUADRANT OF BREAST
C0496809|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST LOWER INNER QUADRANT 
C0496809|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST LOWER INNER QUADRANT
C0496811|T047||CCS_10|MALIGNANT NEOPLASM OF LOWER-OUTER QUADRANT OF BREAST
C0496811|T047||CCS_10|MALIGNANT NEOPLASM OF LOWER OUTER QUADRANT OF BREAST
C0496811|T047||CCS_10|MALIGNANT NEOPLASM OF LOWER OUTER QUADRANT OF BREAST 
C0496811|T047||CCS_10|BREAST NEOPLASM MALIGNANT LOWER OUTER QUADRANT
C0496811|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST LOWER OUTER QUADRANT 
C0496811|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST LOWER OUTER QUADRANT
C0496806|T047||CCS_10|MALIGNANT NEOPLASM OF NIPPLE AND AREOLA
C0496806|T047||CCS_10|MALIGNANT NEOPLASM OF NIPPLE AND AREOLA 
C0496806|T047||CCS_10|BREAST NEOPLASM MALIGNANT NIPPLE / AREOLA
C0348912|T047||CCS_10|MALIGNANT NEOPLASM OVERLAPPING BREAST SITE
C0348912|T047||CCS_10|OVERLAPPING LESION OF BREAST
C0348912|T047||CCS_10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF BREAST
C0348912|T047||CCS_10|BREAST NEOPLASM MALIGNANT OVERLAPPING SITES
C0348912|T047||CCS_10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF BREAST 
C0348912|T047||CCS_10|MALIGNANT NEOPLASM, OVERLAPPING LESION OF BREAST
C0348912|T047||CCS_10|MALIGNANT NEOPLASM, OVERLAPPING LESION OF BREAST 
C0496808|T047||CCS_10|MALIGNANT NEOPLASM OF UPPER-INNER QUADRANT OF BREAST
C0496808|T047||CCS_10|BREAST NEOPLASM MALIGNANT UPPER INNER QUADRANT
C0496808|T047||CCS_10|MALIGNANT NEOPLASM OF UPPER INNER QUADRANT OF BREAST
C0496808|T047||CCS_10|MALIGNANT NEOPLASM OF UPPER INNER QUADRANT OF BREAST 
C0496808|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST UPPER INNER QUADRANT 
C0496808|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST UPPER INNER QUADRANT
C0496810|T047||CCS_10|MALIGNANT NEOPLASM OF UPPER-OUTER QUADRANT OF BREAST
C0496810|T047||CCS_10|MALIGNANT NEOPLASM OF UPPER OUTER QUADRANT OF BREAST 
C0496810|T047||CCS_10|BREAST NEOPLASM MALIGNANT UPPER OUTER QUADRANT
C0496810|T047||CCS_10|MALIGNANT NEOPLASM OF UPPER OUTER QUADRANT OF BREAST
C0496810|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST UPPER OUTER QUADRANT 
C0496810|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST UPPER OUTER QUADRANT
C0678222|T047||CCS_10|CARCINOMA OF BREAST
C0678222|T047||CCS_10|BREAST CARCINOMA
C0678222|T047||CCS_10|CARCINOMA OF BREAST 
C0678222|T047||CCS_10|BREAST CANCER DIAGNOSIS
C0678222|T047||CCS_10|CARCINOMA OF BREAST NOS 
C0678222|T047||CCS_10|CARCINOMA OF BREAST 
C0678222|T047||CCS_10|CARCINOMA OF BREAST NOS
C0678222|T047||CCS_10|BREAST CANCER, NOS
C0678222|T047||CCS_10|BREAST CANCER
C0678222|T047||CCS_10|CANCER, BREAST
C0678222|T047||CCS_10|BREAST CARCINOMA NOS
C0678222|T047||CCS_10|CARCINOMA BREAST
C0678222|T047||CCS_10|CA - CARCINOMA OF BREAST
C0678222|T047||CCS_10|CANCER OF BREAST
C0678222|T047||CCS_10|CANCER OF THE BREAST
C0678222|T047||CCS_10|MAMMARY CARCINOMA
C0678222|T047||CCS_10|CARCINOMA OF THE BREAST
C2842134|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST OF UNSPECIFIED SITE
C0030185|T047||CCS_10|PAGET'S DISEASE, MAMMARY
C0030185|T047||CCS_10|PAGETS DISEASE, BREAST
C0030185|T047||CCS_10|DISEASE, MAMMARY PAGET
C0030185|T047||CCS_10|DISEASE, MAMMARY PAGET'S
C0030185|T047||CCS_10|MAMMARY PAGETS DISEASE
C0030185|T047||CCS_10|PAGETS DISEASE, MAMMARY
C0030185|T047||CCS_10|PAGET'S DISEASE OF BREAST
C0030185|T047||CCS_10|MAMMARY PAGET'S DISEASE
C0030185|T047||CCS_10|PAGETS DIS BREAST
C0030185|T047||CCS_10|PAGET DIS MAMMARY
C0030185|T047||CCS_10|PAGETS DIS MAMMARY
C0030185|T047||CCS_10|MAMMARY PAGETS DIS
C0030185|T047||CCS_10|PAGET DIS BREAST
C0030185|T047||CCS_10|MAMMARY PAGET DIS
C0030185|T047||CCS_10|PAGET DISEASE OF THE BREAST
C0030185|T047||CCS_10|PAGET'S DISEASE OF THE BREAST
C0030185|T047||CCS_10|PAGET'S DISEASE (MAMMARY)
C0030185|T047||CCS_10|PAGET'S DISEASE OF BREAST 
C0030185|T047||CCS_10|PAGET DISEASE, MAMMARY
C0030185|T047||CCS_10|PAGET'S DISEASE, MAMMARY [DISEASE/FINDING]
C0030185|T047||CCS_10|MAMMARY PAGET DISEASE
C0030185|T047||CCS_10|PAGET DISEASE OF BREAST
C0030185|T047||CCS_10|PAGET'S DISEASE OF THE NIPPLE AND AREOLA
C0030185|T047||CCS_10|PAGET'S DISEASE OF THE NIPPLE
C0030185|T047||CCS_10|PAGET DISEASE, BREAST
C0030185|T047||CCS_10|PAGET'S DISEASE, MAMMARY (MORPHOLOGIC ABNORMALITY)
C0030185|T047||CCS_10|BREAST; PAGET
C0030185|T047||CCS_10|BREAST; DISORDER, PAGET
C0030185|T047||CCS_10|PAGET; BREAST
C2211687|T047||CCS_10|BREAST NEOPLASM MALIGNANT SMALL CELL TYPE
C2211687|T047||CCS_10|MALIGNANT SMALL CELL NEOPLASM OF BREAST 
C2211687|T047||CCS_10|MALIGNANT SMALL CELL NEOPLASM OF BREAST
C2011353|T047||CCS_10|GIANT CELL TYPE NEOPLASM OF BREAST
C2011353|T047||CCS_10|GIANT CELL TYPE NEOPLASM OF BREAST 
C2011353|T047||CCS_10|BREAST NEOPLASM MALIGNANT GIANT CELL TYPE
C2018637|T047||CCS_10|BREAST NEOPLASM MALIGNANT SPINDLE CELL TYPE
C2018637|T047||CCS_10|SPINDLE CELL TYPE NEOPLASM OF BREAST
C2018637|T047||CCS_10|SPINDLE CELL TYPE NEOPLASM OF BREAST 
C2075596|T047||CCS_10|BREAST NEOPLASM MALIGNANT CLEAR CELL TYPE
C2075596|T047||CCS_10|CLEAR CELL TYPE NEOPLASM OF BREAST 
C2075596|T047||CCS_10|CLEAR CELL TYPE NEOPLASM OF BREAST
C0349667|T047||CCS_10|SARCOMA OF BREAST
C0349667|T047||CCS_10|SARCOMA OF BREAST 
C0349667|T047||CCS_10|BREAST SARCOMA
C0349667|T047||CCS_10|SARCOMA OF BREAST 
C0349667|T047||CCS_10|SARCOMA OF THE BREAST
C2211725|T047||CCS_10|MYOSARCOMA OF BREAST 
C2211725|T047||CCS_10|MYOSARCOMA OF BREAST
C2211725|T047||CCS_10|BREAST NEOPLASM MALIGNANT MYOSARCOMA
C2007063|T047||CCS_10|CARCINOSARCOMA OF BREAST
C2007063|T047||CCS_10|CARCINOSARCOMA OF BREAST 
C2211730|T047||CCS_10|MALIGNANT MESENCHYMOMA OF BREAST
C2211730|T047||CCS_10|MALIGNANT MESENCHYMOMA OF BREAST 
C2211731|T047||CCS_10|MALIGNANT HEMANGIOENDOTHELIOMA OF BREAST
C2211731|T047||CCS_10|MALIGNANT HEMANGIOENDOTHELIOMA OF BREAST 
C0346154|T047||CCS_10|MALIGNANT CYSTOSARCOMA PHYLLODES OF THE BREAST
C0346154|T047||CCS_10|MALIGNANT PHYLLODES TUMOR OF BREAST
C0346154|T047||CCS_10|MALIGNANT PHYLLODES TUMOR OF BREAST 
C0346154|T047||CCS_10|MALIGNANT CYSTOSARCOMA PHYLLODES OF BREAST
C0346154|T047||CCS_10|MALIGNANT PHYLLODES TUMOUR OF BREAST
C0346154|T047||CCS_10|MALIGNANT PHYLLODES TUMOR OF BREAST 
C0346154|T047||CCS_10|MALIGNANT BREAST PHYLLODES NEOPLASM
C0346154|T047||CCS_10|MALIGNANT MAMMARY PHYLLODES NEOPLASM
C0346154|T047||CCS_10|MALIGNANT MAMMARY PHYLLODES TUMOR
C0346154|T047||CCS_10|MALIGNANT PHYLLODES BREAST NEOPLASM
C0346154|T047||CCS_10|MALIGNANT PHYLLODES NEOPLASM OF BREAST
C0346154|T047||CCS_10|MALIGNANT PHYLLODES NEOPLASM OF THE BREAST
C0346154|T047||CCS_10|MALIGNANT PHYLLODES TUMOR OF THE BREAST
C0346154|T047||CCS_10|MALIGNANT BREAST PHYLLODES TUMOR
C2211733|T047||CCS_10|MALIGNANT GRANULAR CELL TUMOR OF BREAST
C2211733|T047||CCS_10|MALIGNANT GRANULAR CELL TUMOR OF BREAST 
C2211755|T047||CCS_10|MALIGNANT PLASMACYTOMA OF BREAST 
C2211755|T047||CCS_10|MALIGNANT PLASMACYTOMA OF BREAST
C2211757|T047||CCS_10|MALIGNANT MASTOCYTOSIS OF BREAST
C2211757|T047||CCS_10|MALIGNANT MASTOCYTOSIS OF BREAST 
C2216702|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST STAGING 
C2216702|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST STAGING
C2216702|T047||CCS_10|MALIGNANT BREAST NEOPLASM STAGING
C2216702|T047||CCS_10|MALIGNANT TUMOR OF BREAST STAGING
C2216702|T047||CCS_10|BREAST CANCER STAGING
C2216702|T047||CCS_10|STAGE, BREAST CANCER
C2216702|T047||CCS_10|BREAST CANCER STAGE
C0858252|T047||CCS_10|ADENOCARCINOMA OF BREAST 
C0858252|T047||CCS_10|ADENOCARCINOMA OF BREAST
C0858252|T047||CCS_10|BREAST ADENOCARCINOMA
C0858252|T047||CCS_10|ADENOCARCINOMA OF THE BREAST
C1332630|T047||CCS_10|FIBROSARCOMA OF BREAST 
C1332630|T047||CCS_10|FIBROSARCOMA OF BREAST
C1332630|T047||CCS_10|FIBROSARCOMA OF THE BREAST
C1332630|T047||CCS_10|BREAST FIBROSARCOMA
C2062549|T047||CCS_10|BREAST NIPPLE EPITHELIOMA
C1332632|T047||CCS_10|LIPOSARCOMA OF BREAST 
C1332632|T047||CCS_10|LIPOSARCOMA OF BREAST
C1332632|T047||CCS_10|LIPOSARCOMA OF THE BREAST
C1332632|T047||CCS_10|BREAST LIPOSARCOMA
C0235653|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST (FEMALE), UNSPECIFIED
C0235653|T047||CCS_10|MALIGNANT NEOPLASM OF FEMALE BREAST
C0235653|T047||CCS_10|MALIGNANT NEOPLASM OF FEMALE BREAST 
C0235653|T047||CCS_10|CANCER OF FEMALE BREAST
C0235653|T047||CCS_10|MALIGNANT FEMALE BREAST NEOPLASM
C0235653|T047||CCS_10|MALIGNANT TUMOR OF FEMALE BREAST
C0235653|T047||CCS_10|MALIGN NEOPL BREAST NOS
C0235653|T047||CCS_10|MALIGNANT NEOPLASM OF FEMALE BREAST 
C0235653|T047||CCS_10|MALIGNANT NEOPLASM OF FEMALE BREAST NOS
C0235653|T047||CCS_10|MALIGNANT NEOPLASM OF FEMALE BREAST NOS 
C0235653|T047||CCS_10|BREAST CANCER FEMALE
C0235653|T047||CCS_10|FEMALE BREAST CANCER
C0235653|T047||CCS_10|MALIGNANT NEOPLASM OF FEMALE BREAST, UNSPECIFIED
C0235653|T047||CCS_10|BREAST NEOPLASM MALIGNANT FEMALE
C0235653|T047||CCS_10|BREAST CANCER FEMALE NOS
C0235653|T047||CCS_10|BREAST CANCER, FEMALE
C0235653|T047||CCS_10|MALIGNANT NEOPLASM OF FEMALE BREAST, NOS
C0235653|T047||CCS_10|NEOPLASM MALIG;BREAST;F
C0235653|T047||CCS_10|MALIGNANT NEOSPLASM OF THE FEMALE BREAST
C2211688|T047||CCS_10|MALIGNANT EPITHELIOMA OF BREAST
C2211688|T047||CCS_10|MALIGNANT EPITHELIOMA OF BREAST 
C2111593|T047||CCS_10|LARGE CELL CARCINOMA OF BREAST
C2111593|T047||CCS_10|LARGE CELL CARCINOMA OF BREAST 
C1511316|T047||CCS_10|LARGE CELL NEUROENDOCRINE CARCINOMA OF BREAST
C1511316|T047||CCS_10|LARGE CELL NEUROENDOCRINE CARCINOMA OF BREAST 
C1511316|T047||CCS_10|BREAST LARGE CELL NEUROENDOCRINE CARCINOMA
C2111594|T047||CCS_10|LARGE CELL CARCINOMA OF BREAST WITH RHABDOID PHENOTYPE 
C2111594|T047||CCS_10|BREAST MALIGNANT CARCINOMA LARGE CELL W/ RHABDOID PHENOTYPE
C2111594|T047||CCS_10|LARGE CELL CARCINOMA OF BREAST WITH RHABDOID PHENOTYPE
C2012071|T047||CCS_10|GLASSY CELL CARCINOMA OF BREAST
C2012071|T047||CCS_10|GLASSY CELL CARCINOMA OF BREAST 
C1336854|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF BREAST
C1336854|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF BREAST 
C2211689|T047||CCS_10|ANAPLASTIC CARCINOMA OF BREAST 
C2211689|T047||CCS_10|ANAPLASTIC CARCINOMA OF BREAST
C2211689|T047||CCS_10|ANAPLASTIC BREAST CARCINOMA
C1514169|T047||CCS_10|PLEOMORPHIC CARCINOMA OF BREAST
C1514169|T047||CCS_10|PLEOMORPHIC CARCINOMA OF BREAST 
C1514169|T047||CCS_10|PLEOMORPHIC BREAST CARCINOMA
C2011243|T047||CCS_10|GIANT CELL CARCINOMA OF BREAST 
C2011243|T047||CCS_10|GIANT CELL CARCINOMA OF BREAST
C2018385|T047||CCS_10|SPINDLE CELL CARCINOMA OF BREAST
C2018385|T047||CCS_10|SPINDLE CELL CARCINOMA OF BREAST 
C2011208|T047||CCS_10|GIANT CELL AND SPINDLE CELL CARCINOMA OF BREAST 
C2011208|T047||CCS_10|GIANT CELL AND SPINDLE CELL CARCINOMA OF BREAST
C2142913|T047||CCS_10|PSEUDOSARCOMATOUS CARCINOMA OF BREAST
C2142913|T047||CCS_10|PSEUDOSARCOMATOUS CARCINOMA OF BREAST 
C2111795|T047||CCS_10|POLYGONAL CELL CARCINOMA OF BREAST 
C2111795|T047||CCS_10|POLYGONAL CELL CARCINOMA OF BREAST
C2007022|T047||CCS_10|CARCINOMA OF BREAST WITH OSTEOCLAST-LIKE GIANT CELLS 
C2007022|T047||CCS_10|CARCINOMA OF BREAST WITH OSTEOCLAST-LIKE GIANT CELLS
C2007022|T047||CCS_10|BREAST CARCINOMA WITH OSTEOCLAST-LIKE GIANT CELLS
C3812899|T047||CCS_10|PAPILLARY CARCINOMA OF BREAST
C3812899|T047||CCS_10|PAPILLARY CARCINOMA OF BREAST 
C3812899|T047||CCS_10|PAPILLARY CARCINOMA OF THE BREAST (MORPHOLOGIC ABNORMALITY)
C3812899|T047||CCS_10|PAPILLARY CARCINOMA OF THE BREAST
C3812899|T047||CCS_10|PAPILLARY BREAST CARCINOMA
C2033277|T047||CCS_10|PAPILLARY SQUAMOUS CELL CARCINOMA OF BREAST 
C2033277|T047||CCS_10|PAPILLARY SQUAMOUS CELL CARCINOMA OF BREAST
C2189332|T047||CCS_10|VERRUCOUS CARCINOMA OF BREAST 
C2189332|T047||CCS_10|VERRUCOUS CARCINOMA OF BREAST
C1336079|T047||CCS_10|PRIMARY SQUAMOUS CELL CARCINOMA OF BREAST
C1336079|T047||CCS_10|PRIMARY SQUAMOUS CELL BREAST CARCINOMA
C1336079|T047||CCS_10|PRIMARY SQUAMOUS CELL CARCINOMA OF THE BREAST
C1336079|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF BREAST 
C1336079|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF BREAST
C1336079|T047||CCS_10|SCC OF BREAST
C1336079|T047||CCS_10|SCC OF THE BREAST
C1336079|T047||CCS_10|SQUAMOUS BREAST CARCINOMA
C1336079|T047||CCS_10|SQUAMOUS CARCINOMA OF BREAST
C1336079|T047||CCS_10|SQUAMOUS CARCINOMA OF THE BREAST
C1336079|T047||CCS_10|SQUAMOUS CELL BREAST CARCINOMA
C1336079|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE BREAST
C2109290|T047||CCS_10|KERATINIZING SQUAMOUS CELL CARCINOMA OF BREAST
C2109290|T047||CCS_10|KERATINIZING SQUAMOUS CELL CARCINOMA OF BREAST 
C2211690|T047||CCS_10|NONKERATINIZING LARGE CELL SQUAMOUS CARCINOMA CELL OF BREAST
C2211690|T047||CCS_10|NONKERATINIZING LARGE CELL SQUAMOUS CARCINOMA CELL OF BREAST 
C2211690|T047||CCS_10|BREAST MALIGNANT CARCINOMA SQUAMOUS CELL LARGE CELL NONKERATINIZING
C2018534|T047||CCS_10|SPINDLE CELL SQUAMOUS CELL CARCINOMA OF BREAST
C2018534|T047||CCS_10|SPINDLE CELL SQUAMOUS CELL CARCINOMA OF BREAST 
C2211692|T047||CCS_10|ADENOID SQUAMOUS CELL CARCINOMA OF BREAST 
C2211692|T047||CCS_10|ADENOID SQUAMOUS CELL CARCINOMA OF BREAST
C2211693|T047||CCS_10|MICROINVASIVE SQUAMOUS CELL CARCINOMA OF BREAST 
C2211693|T047||CCS_10|MICROINVASIVE SQUAMOUS CELL CARCINOMA OF BREAST
C2019466|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF BREAST WITH HORN FORMATION
C2019466|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF BREAST WITH HORN FORMATION 
C2019466|T047||CCS_10|SQUAMOUS CELL CARCINOMA WITH HORN FORMATION OF BREAST
C1332638|T047||CCS_10|OAT CELL CARCINOMA OF BREAST
C1332638|T047||CCS_10|SMALL CELL CARCINOMA OF BREAST
C1332638|T047||CCS_10|SMALL CELL CARCINOMA OF BREAST 
C1332638|T047||CCS_10|MAMMARY SMALL CELL CARCINOMA
C1332638|T047||CCS_10|OAT CELL CARCINOMA OF THE BREAST
C1332638|T047||CCS_10|SMALL CELL CARCINOMA OF THE BREAST
C1332638|T047||CCS_10|SMALL CELL NEUROENDOCRINE CARCINOMA OF BREAST
C1332638|T047||CCS_10|SMALL CELL NEUROENDOCRINE CARCINOMA OF THE BREAST
C1332638|T047||CCS_10|BREAST SMALL CELL CARCINOMA
C2009874|T047||CCS_10|FUSIFORM TYPE SMALL CELL CARCINOMA OF BREAST 
C2009874|T047||CCS_10|FUSIFORM TYPE SMALL CELL CARCINOMA OF BREAST
C1332167|T047||CCS_10|ADENOID CYSTIC CARCINOMA OF BREAST
C1332167|T047||CCS_10|ADENOID CYSTIC CARCINOMA OF BREAST 
C1332167|T047||CCS_10|ADENOID CYSTIC BREAST CARCINOMA
C1332167|T047||CCS_10|ADENOCYSTIC BREAST CARCINOMA
C1332167|T047||CCS_10|ADENOCYSTIC CARCINOMA OF BREAST
C1332167|T047||CCS_10|ADENOCYSTIC CARCINOMA OF THE BREAST
C1332167|T047||CCS_10|ADENOID CYSTIC CARCINOMA OF THE BREAST
C1332167|T047||CCS_10|MAMMARY ADENOCYSTIC CARCINOMA
C2007046|T047||CCS_10|CARCINOMA SIMPLEX OF BREAST
C2007046|T047||CCS_10|CARCINOMA SIMPLEX OF BREAST 
C1517894|T047||CCS_10|LIPID-RICH CARCINOMA OF BREAST
C1517894|T047||CCS_10|LIPID-RICH CARCINOMA OF BREAST 
C1517894|T047||CCS_10|LIPID SECRETING BREAST CARCINOMA
C1517894|T047||CCS_10|LIPID-RICH BREAST CARCINOMA
C2012538|T047||CCS_10|GRANULAR CELL CARCINOMA OF BREAST 
C2012538|T047||CCS_10|GRANULAR CELL CARCINOMA OF BREAST
C1335964|T047||CCS_10|SIGNET RING CELL CARCINOMA OF BREAST
C1335964|T047||CCS_10|SIGNET RING CELL CARCINOMA OF BREAST 
C1335964|T047||CCS_10|MAMMARY SIGNET RING CELL CARCINOMA
C1335964|T047||CCS_10|PRIMARY MAMMARY SIGNET RING CELL CARCINOMA
C1335964|T047||CCS_10|PRIMARY SRC BREAST CARCINOMA
C1335964|T047||CCS_10|PRIMARY SRC CARCINOMA OF BREAST
C1335964|T047||CCS_10|PRIMARY SRC CARCINOMA OF THE BREAST
C1335964|T047||CCS_10|PRIMARY SIGNET RING CELL BREAST CARCINOMA
C1335964|T047||CCS_10|PRIMARY SIGNET RING CELL CARCINOMA OF BREAST
C1335964|T047||CCS_10|PRIMARY SIGNET RING CELL CARCINOMA OF THE BREAST
C1335964|T047||CCS_10|SRC BREAST CARCINOMA
C1335964|T047||CCS_10|SRC CARCINOMA OF BREAST
C1335964|T047||CCS_10|SRC CARCINOMA OF THE BREAST
C1335964|T047||CCS_10|SIGNET RING CELL BREAST CARCINOMA
C1335964|T047||CCS_10|SIGNET RING CELL CARCINOMA OF THE BREAST
C1334002|T047||CCS_10|COMEDOCARCINOMA OF BREAST 
C1334002|T047||CCS_10|COMEDOCARCINOMA OF BREAST
C1334002|T047||CCS_10|HIGH GRADE DUCTAL BREAST CARCINOMA IN SITU
C1334002|T047||CCS_10|COMEDO CARCINOMA
C1334002|T047||CCS_10|DIN 3
C1334002|T047||CCS_10|DUCTAL INTRAEPITHELIAL NEOPLASIA 3
C1334002|T047||CCS_10|DCIS GRADE 3
C1334002|T047||CCS_10|DUCTAL INTRAEPITHELIAL NEOPLASIA, GRADE 3
C1334002|T047||CCS_10|HIGH-GRADE DCIS OF BREAST
C1334002|T047||CCS_10|HIGH-GRADE DCIS OF THE BREAST
C1334002|T047||CCS_10|HIGH-GRADE DUCTAL CARCINOMA IN SITU OF BREAST
C1334002|T047||CCS_10|BREAST COMEDOCARCINOMA
C0334371|T047||CCS_10|CYSTIC HYPERSECRETORY CARCINOMA OF BREAST
C0334371|T047||CCS_10|CYSTIC HYPERSECRETORY BREAST CARCINOMA
C0334371|T047||CCS_10|SECRETORY CARCINOMA
C0334371|T047||CCS_10|CYSTIC HYPERSECRETORY CARCINOMA OF THE BREAST
C0334371|T047||CCS_10|SECRETORY CARCINOMA OF BREAST 
C0334371|T047||CCS_10|SECRETORY CARCINOMA OF BREAST
C0334371|T047||CCS_10|HYPERSECRETORY CYSTIC CARCINOMA OF BREAST 
C0334371|T047||CCS_10|HYPERSECRETORY CYSTIC CARCINOMA OF BREAST
C0334371|T047||CCS_10|SECRETORY BREAST CARCINOMA
C0334371|T047||CCS_10|JUVENILE CARCINOMA OF THE BREAST
C0334371|T047||CCS_10|SECRETORY CARCINOMA OF THE BREAST
C0334371|T047||CCS_10|JUVENILE CARCINOMA OF THE BREAST (MORPHOLOGIC ABNORMALITY)
C0334371|T047||CCS_10|INFILTRATING CYSTIC HYPERSECRETORY DUCT BREAST CARCINOMA
C0334371|T047||CCS_10|INVASIVE CYSTIC HYPERSECRETORY DUCT BREAST CARCINOMA
C0334371|T047||CCS_10|JUVENILE BREAST CARCINOMA
C0334371|T047||CCS_10|JUVENILE CARCINOMA OF BREAST
C0334371|T047||CCS_10|JUVENILE SECRETORY BREAST CARCINOMA
C0334371|T047||CCS_10|JUVENILE SECRETORY CARCINOMA OF BREAST
C0334371|T047||CCS_10|JUVENILE SECRETORY CARCINOMA OF THE BREAST
C0334376|T047||CCS_10|INTRACYSTIC CARCINOMA OF BREAST 
C0334376|T047||CCS_10|INTRACYSTIC CARCINOMA OF BREAST
C0334376|T047||CCS_10|INTRACYSTIC PAPILLARY BREAST CARCINOMA
C0334376|T047||CCS_10|[M] INTRACYSTIC CARCINOMA NOS
C0334376|T047||CCS_10|[M] INTRACYSTIC CARCINOMA NOS (MORPHOLOGIC ABNORMALITY)
C0334376|T047||CCS_10|INTRACYSTIC CARCINOMA
C0334376|T047||CCS_10|INTRACYSTIC CARCINOMA (MORPHOLOGIC ABNORMALITY)
C0334376|T047||CCS_10|INTRACYSTIC PAPILLARY ADENOCARCINOMA
C0334376|T047||CCS_10|INTRACYSTIC CARCINOMA, NOS
C0334376|T047||CCS_10|INTRACYSTIC BREAST CARCINOMA
C0334376|T047||CCS_10|NONINFILTRATING INTRACYSTIC BREAST CARCINOMA
C0860580|T047||CCS_10|MEDULLARY CARCINOMA OF BREAST 
C0860580|T047||CCS_10|MEDULLARY CARCINOMA OF BREAST
C0860580|T047||CCS_10|MEDULLARY BREAST CARCINOMA
C0860580|T047||CCS_10|INFILTRATING MEDULLARY CARCINOMA OF BREAST
C0860580|T047||CCS_10|INFILTRATING MEDULLARY CARCINOMA OF THE BREAST
C0860580|T047||CCS_10|INVASIVE MEDULLARY BREAST CARCINOMA
C0860580|T047||CCS_10|INVASIVE MEDULLARY CARCINOMA OF BREAST
C0860580|T047||CCS_10|INVASIVE MEDULLARY CARCINOMA OF THE BREAST
C0860580|T047||CCS_10|MEDULLARY BREAST CARCINOMA WITH LYMPHOID STROMA
C0860580|T047||CCS_10|MEDULLARY CARCINOMA OF THE BREAST
C2211694|T047||CCS_10|MEDULLARY CARCINOMA WITH LYMPHOID STROMA OF BREAST 
C2211694|T047||CCS_10|MEDULLARY CARCINOMA WITH LYMPHOID STROMA OF BREAST
C1879758|T047||CCS_10|ATYPICAL MEDULLARY BREAST CARCINOMA
C1879758|T047||CCS_10|INFILTRATING DUCTAL BREAST CARCINOMA WITH MEDULLARY FEATURES
C1879758|T047||CCS_10|ATYPICAL MEDULLARY CARCINOMA OF BREAST 
C1879758|T047||CCS_10|ATYPICAL MEDULLARY CARCINOMA OF BREAST
C2182973|T047||CCS_10|DESMOPLASTIC TYPE DUCTAL CARCINOMA OF BREAST
C2182973|T047||CCS_10|DESMOPLASTIC TYPE DUCTAL CARCINOMA OF BREAST 
C2076522|T047||CCS_10|INFILTRATING DUCTAL AND LOBULAR CARCINOMA OF BREAST 
C2076522|T047||CCS_10|INFILTRATING DUCTAL AND LOBULAR CARCINOMA OF BREAST
C2146658|T047||CCS_10|ACINAR CELL CARCINOMA OF BREAST 
C2146658|T047||CCS_10|ACINAR CELL CARCINOMA OF BREAST
C2146670|T047||CCS_10|ACINAR CELL CYSTADENOCARCINOMA OF BREAST
C2146670|T047||CCS_10|ACINAR CELL CYSTADENOCARCINOMA OF BREAST 
C1510796|T047||CCS_10|ADENOSQUAMOUS CARCINOMA OF BREAST
C1510796|T047||CCS_10|ADENOSQUAMOUS CARCINOMA OF BREAST 
C1510796|T047||CCS_10|ADENOSQUAMOUS BREAST CARCINOMA
C2211695|T047||CCS_10|EPITHELIAL-MYOEPITHELIAL CARCINOMA OF BREAST 
C2211695|T047||CCS_10|EPITHELIAL-MYOEPITHELIAL CARCINOMA OF BREAST
C1334708|T047||CCS_10|METAPLASTIC CARCINOMA OF BREAST 
C1334708|T047||CCS_10|METAPLASTIC CARCINOMA OF BREAST
C1334708|T047||CCS_10|METAPLASTIC BREAST CARCINOMA
C1334708|T047||CCS_10|METAPLASTIC CARCINOMA OF THE BREAST
C2211696|T047||CCS_10|SCIRRHOUS ADENOCARCINOMA OF BREAST
C2211696|T047||CCS_10|SCIRRHOUS ADENOCARCINOMA OF BREAST 
C2037312|T047||CCS_10|SUPERFICIAL SPREADING ADENOCARCINOMA OF BREAST
C2037312|T047||CCS_10|SUPERFICIAL SPREADING ADENOCARCINOMA OF BREAST 
C2211697|T047||CCS_10|BASAL CELL ADENOCARCINOMA OF BREAST
C2211697|T047||CCS_10|BASAL CELL ADENOCARCINOMA OF BREAST 
C2145023|T047||CCS_10|TRABECULAR ADENOCARCINOMA OF BREAST 
C2145023|T047||CCS_10|TRABECULAR ADENOCARCINOMA OF BREAST
C2033109|T047||CCS_10|PAPILLARY ADENOCARCINOMA OF BREAST 
C2033109|T047||CCS_10|PAPILLARY ADENOCARCINOMA OF BREAST
C2211698|T047||CCS_10|APOCRINE ADENOCARCINOMA OF BREAST 
C2211698|T047||CCS_10|APOCRINE ADENOCARCINOMA OF BREAST
C2211699|T047||CCS_10|INTRADUCTAL PAPILLARY ADENOCARCINOMA OF BREAST WITH INVASION
C2211699|T047||CCS_10|INTRADUCTAL PAPILLARY ADENOCARCINOMA OF BREAST WITH INVASION 
C2211700|T047||CCS_10|MIXED CELL ADENOCARCINOMA OF BREAST 
C2211700|T047||CCS_10|MIXED CELL ADENOCARCINOMA OF BREAST
C2211701|T047||CCS_10|POLYMORPHOUS LOW GRADE ADENOCARCINOMA OF BREAST 
C2211701|T047||CCS_10|POLYMORPHOUS LOW GRADE ADENOCARCINOMA OF BREAST
C2075524|T047||CCS_10|CLEAR CELL ADENOCARCINOMA OF BREAST 
C2075524|T047||CCS_10|CLEAR CELL ADENOCARCINOMA OF BREAST
C2211702|T047||CCS_10|MUCINOUS ADENOCARCINOMA OF BREAST 
C2211702|T047||CCS_10|MUCINOUS ADENOCARCINOMA OF BREAST
C2211703|T047||CCS_10|MUCIN-PRODUCING ADENOCARCINOMA OF BREAST 
C2211703|T047||CCS_10|MUCIN-PRODUCING ADENOCARCINOMA OF BREAST
C2211704|T047||CCS_10|BREAST ADENOCARCINOMA WITH METAPLASIA
C2211704|T047||CCS_10|ADENOCARCINOMA OF BREAST WITH METAPLASIA 
C2211704|T047||CCS_10|ADENOCARCINOMA OF BREAST WITH METAPLASIA
C1332613|T047||CCS_10|ADENOCARCINOMA OF BREAST WITH SQUAMOUS METAPLASIA 
C1332613|T047||CCS_10|ADENOCARCINOMA OF BREAST WITH SQUAMOUS METAPLASIA
C1332613|T047||CCS_10|BREAST ADENOCARCINOMA WITH SQUAMOUS METAPLASIA
C1332613|T047||CCS_10|ADENOACANTHOMA OF BREAST
C1332613|T047||CCS_10|ADENOACANTHOMA OF THE BREAST
C1332613|T047||CCS_10|ADENOCARCINOMA OF THE BREAST WITH SQUAMOUS METAPLASIA
C1332613|T047||CCS_10|BREAST ADENOACANTHOMA
C2211705|T047||CCS_10|ADENOCARCINOMA WITH CARTILAGINOUS OR OSSEOUS METAPLASIA OF BREAST
C2211705|T047||CCS_10|ADENOCARCINOMA OF BREAST WITH CARTILAGINOUS AND OSSEOUS METAPLASIA
C2211705|T047||CCS_10|BREAST ADENOCARCINOMA WITH CARTILAGINOUS OR OSSEOUS METAPLASIA
C2211705|T047||CCS_10|ADENOCARCINOMA OF BREAST WITH CARTILAGINOUS AND OSSEOUS METAPLASIA 
C2211705|T047||CCS_10|BREAST ADENOCARCINOMA WITH CARTILAGINOUS AND OSSEOUS METAPLASIA
C1511281|T047||CCS_10|BREAST ADENOCARCINOMA WITH SPINDLE CELL METAPLASIA
C1511281|T047||CCS_10|ADENOCARCINOMA OF BREAST WITH SPINDLE CELL METAPLASIA
C1511281|T047||CCS_10|ADENOCARCINOMA OF BREAST WITH SPINDLE CELL METAPLASIA 
C2211706|T047||CCS_10|ADENOCARCINOMA OF BREAST WITH APOCRINE METAPLASIA
C2211706|T047||CCS_10|BREAST ADENOCARCINOMA WITH APOCRINE METAPLASIA
C2211706|T047||CCS_10|ADENOCARCINOMA OF BREAST WITH APOCRINE METAPLASIA 
C2211707|T047||CCS_10|ADENOCARCINOMA OF BREAST WITH NEUROENDOCRINE DIFFERENTIATION 
C2211707|T047||CCS_10|ADENOCARCINOMA OF BREAST WITH NEUROENDOCRINE DIFFERENTIATION
C2211707|T047||CCS_10|BREAST ADENOCARCINOMA WITH NEUROENDOCRINE DIFFERENTIATION
C2170817|T047||CCS_10|TUBULAR ADENOCARCINOMA OF BREAST 
C2170817|T047||CCS_10|TUBULAR ADENOCARCINOMA OF BREAST
C2211708|T047||CCS_10|ALVEOLAR ADENOCARCINOMA OF BREAST
C2211708|T047||CCS_10|ALVEOLAR ADENOCARCINOMA OF BREAST 
C2163806|T047||CCS_10|CYSTADENOCARCINOMA OF BREAST 
C2163806|T047||CCS_10|CYSTADENOCARCINOMA OF BREAST
C2211732|T047||CCS_10|MALIGNANT EPITHELIOID HEMANGIOENDOTHELIOMA OF BREAST
C2211732|T047||CCS_10|MALIGNANT EPITHELIOID HEMANGIOENDOTHELIOMA OF BREAST 
C0334386|T047||CCS_10|PAGET'S DISEASE AND INFILTRATING DUCT CARCINOMA OF BREAST
C0334386|T047||CCS_10|PAGET'S DISEASE AND INFILTRATING DUCT CARCINOMA OF BREAST 
C0334386|T047||CCS_10|PAGET DISEASE AND INFILTRATING DUCT CARCINOMA OF BREAST
C0334386|T047||CCS_10|PAGET'S DISEASE AND INFILTRATING DUCT CARCINOMA OF BREAST (MORPHOLOGIC ABNORMALITY)
C0279566|T047||CCS_10|PAGET DISEASE AND INTRADUCTAL CARCINOMA OF THE BREAST
C0279566|T047||CCS_10|PAGET'S DISEASE AND INTRADUCTAL CARCINOMA OF THE BREAST
C0279566|T047||CCS_10|PAGET'S DISEASE AND INTRADUCTAL CARCINOMA OF BREAST 
C0279566|T047||CCS_10|PAGET'S DISEASE AND INTRADUCTAL CARCINOMA OF BREAST
C0279566|T047||CCS_10|PAGET DISEASE AND INTRADUCTAL CARCINOMA OF BREAST
C0279566|T047||CCS_10|PAGET'S DISEASE AND INTRADUCTAL CARCINOMA OF BREAST 
C0279566|T047||CCS_10|[M]PAGET'S DISEASE AND INTRADUCTAL CARCINOMA OF BREAST
C0279566|T047||CCS_10|[M] PAGET'S DISEASE AND INTRADUCTAL CARCINOMA OF BREAST
C0279566|T047||CCS_10|PAGET'S DISEASE AND INTRADUCTAL CARCINOMA OF BREAST (MORPHOLOGIC ABNORMALITY)
C0279566|T047||CCS_10|PAGET'S DISEASE OF THE BREAST WITH INTRADUCTAL CARCINOMA
C0279566|T047||CCS_10|PAGET'S DISEASE OF BREAST WITH INTRADUCTAL CARCINOMA
C2211718|T047||CCS_10|MALIGNANT SOLITARY FIBROUS TUMOR OF BREAST
C2211718|T047||CCS_10|MALIGNANT SOLITARY FIBROUS TUMOR OF BREAST 
C2211729|T047||CCS_10|EMBRYONAL CARCINOSARCOMA OF BREAST
C2211729|T047||CCS_10|EMBRYONAL CARCINOSARCOMA OF BREAST 
C1518167|T047||CCS_10|MALIGNANT MYOEPITHELIOMA OF BREAST 
C1518167|T047||CCS_10|MALIGNANT MYOEPITHELIOMA OF BREAST
C1518167|T047||CCS_10|BREAST MYOEPITHELIAL CARCINOMA
C1518167|T047||CCS_10|MALIGNANT BREAST MYOEPITHELIOMA
C2216703|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING
C2216703|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING 
C2216703|T047||CCS_10|MALIGNANT BREAST NEOPLASM TNM STAGING
C2216703|T047||CCS_10|MALIGNANT TUMOR OF BREAST TNM STAGING
C2216703|T047||CCS_10|BREAST CANCER TNM STAGING
C2216694|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST STAGE 0
C2216694|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST STAGE 0 
C2216694|T047||CCS_10|MALIGNANT BREAST NEOPLASM STAGE 0
C2216694|T047||CCS_10|BREAST CANCER STAGE 0
C2216694|T047||CCS_10|MALIGNANT TUMOR OF BREAST STAGE 0
C2216695|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST STAGE I 
C2216695|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST STAGE I
C2216695|T047||CCS_10|MALIGNANT BREAST NEOPLASM STAGE I
C2216695|T047||CCS_10|MALIGNANT TUMOR OF BREAST STAGE I
C2216695|T047||CCS_10|BREAST CANCER STAGE I
C2216695|T047||CCS_10|STAGE I BREAST CANCER
C2216695|T047||CCS_10|STAGE I BREAST CANCER AJCC V7
C2216696|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST STAGE IIA 
C2216696|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST STAGE IIA
C2216696|T047||CCS_10|MALIGNANT BREAST NEOPLASM STAGE IIA
C2216696|T047||CCS_10|BREAST CANCER STAGE IIA
C2216696|T047||CCS_10|MALIGNANT TUMOR OF BREAST STAGE IIA
C2216697|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST STAGE IIB 
C2216697|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST STAGE IIB
C2216697|T047||CCS_10|MALIGNANT BREAST NEOPLASM STAGE IIB
C2216697|T047||CCS_10|MALIGNANT TUMOR OF BREAST STAGE IIB
C2216697|T047||CCS_10|BREAST CANCER STAGE IIB
C2216698|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST STAGE IIIA 
C2216698|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST STAGE IIIA
C2216698|T047||CCS_10|MALIGNANT BREAST NEOPLASM STAGE IIIA
C2216698|T047||CCS_10|MALIGNANT TUMOR OF BREAST STAGE IIIA
C2216698|T047||CCS_10|BREAST CANCER STAGE IIIA
C2216699|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST STAGE IIIB 
C2216699|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST STAGE IIIB
C2216699|T047||CCS_10|MALIGNANT BREAST NEOPLASM STAGE IIIB
C2216699|T047||CCS_10|BREAST CANCER STAGE IIIB
C2216699|T047||CCS_10|MALIGNANT TUMOR OF BREAST STAGE IIIB
C2216700|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST STAGE IIIC
C2216700|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST STAGE IIIC 
C2216700|T047||CCS_10|MALIGNANT BREAST NEOPLASM STAGE IIIC
C2216700|T047||CCS_10|MALIGNANT TUMOR OF BREAST STAGE IIIC
C2216700|T047||CCS_10|BREAST CANCER STAGE IIIC
C2216700|T047||CCS_10|STAGE IIIC BREAST CANCER AJCC V6
C2216700|T047||CCS_10|STAGE IIIC BREAST CARCINOMA AJCC V6
C2216700|T047||CCS_10|STAGE IIIC BREAST CANCER
C2216701|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST STAGE IV
C2216701|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST STAGE IV 
C2216701|T047||CCS_10|MALIGNANT BREAST NEOPLASM STAGE IV
C2216701|T047||CCS_10|BREAST CANCER STAGE IV
C2216701|T047||CCS_10|MALIGNANT TUMOR OF BREAST STAGE IV
C2062550|T047||CCS_10|NEUROSARCOMA OF BREAST 
C2062550|T047||CCS_10|NEUROSARCOMA OF BREAST
C2211754|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF BREAST 
C2211754|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF BREAST
C3665394|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF BREAST
C3665394|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF BREAST 
C3665394|T047||CCS_10|SKIN NEOPLASM MALIGNANT BREAST
C3665394|T047||CCS_10|MALIGNANT SKIN NEOPLASM OF BREAST
C3665394|T047||CCS_10|MALIGNANT SKIN NEOPLASM OF BREAST 
C3469450|T047||CCS_10|SUSCEPTIBILITY TO FAMILIAL BREAST-OVARIAN CANCER SYNDROME 
C3469450|T047||CCS_10|SUSCEPTIBILITY TO FAMILIAL BREAST-OVARIAN CANCER SYNDROME
C3469522|T047||CCS_10|BREAST CANCER SUSCEPTIBILITY 
C3469522|T047||CCS_10|BREAST CANCER SUSCEPTIBILITY
C3469522|T047||CCS_10|BREAST CANCER, SUSCEPTIBILITY TO
C1306469|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF MALE BREAST 
C1306469|T047||CCS_10|BREAST NEOPLASM MALIGNANT MALE PRIMARY
C1306469|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF MALE BREAST
C1306469|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF MALE BREAST 
C0559019|T047||CCS_10|CA BREAST-UPPER,INNER QUADRANT 
C0559019|T047||CCS_10|CA BREAST-UPPER,INNER QUADRANT
C0559020|T047||CCS_10|CA BREAST-UPPER,OUTER QUADRANT
C0559020|T047||CCS_10|CA BREAST-UPPER,OUTER QUADRANT 
C1304708|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF FEMALE BREAST
C1304708|T047||CCS_10|BREAST NEOPLASM MALIGNANT FEMALE PRIMARY
C1304708|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF FEMALE BREAST 
C1304708|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF FEMALE BREAST 
C0346860|T047||CCS_10|MALIGNANT MALE BREAST TISSUE NEOPLASM
C0346860|T047||CCS_10|MALIGNANT MALE BREAST ECTOPIC TISSUE NEOPLASM
C0346860|T047||CCS_10|MALIGNANT MALE BREAST NEOPLASM OF ECTOPIC BREAST TISSUE
C0346860|T047||CCS_10|MALIGNANT NEOPLASM OF ECTOPIC TISSUE OF MALE BREAST
C0346860|T047||CCS_10|MALIGNANT MALE BREAST NEOPLASM OF ECTOPIC BREAST TISSUE 
C0346860|T047||CCS_10|MALIGNANT NEOPLASM OF ECTOPIC SITE OF MALE BREAST
C0346860|T047||CCS_10|MALIGNANT NEOPLASM OF ECTOPIC SITE OF MALE BREAST 
C0559021|T047||CCS_10|CA BREAST-LOWER,OUTER QUADRANT
C0559021|T047||CCS_10|CA BREAST-LOWER,OUTER QUADRANT 
C0559062|T047||CCS_10|CA BREAST-LOWER,INNER QUADRANT
C0559062|T047||CCS_10|CA BREAST-LOWER,INNER QUADRANT 
C0948966|T047||CCS_10|MALIGNANT NIPPLE NEOPLASM FEMALE
C0948966|T047||CCS_10|BREAST NEOPLASM MALIGNANT FEMALE NIPPLE
C0948966|T047||CCS_10|MALIGNANT NEOPLASM OF FEMALE NIPPLE 
C0948966|T047||CCS_10|MALIGNANT NEOPLASM OF FEMALE NIPPLE
C0948966|T047||CCS_10|MALIGNANT NEOPLASM OF NIPPLE OF FEMALE BREAST
C0948966|T047||CCS_10|FEMALE MALIGNANT NIPPLE NEOPLASM
C0346858|T047||CCS_10|MALIGNANT NEOPLASM OF AREOLA OF MALE BREAST
C0346858|T047||CCS_10|MALIGNANT NEOPLASM OF AREOLA OF MALE BREAST 
C0346858|T047||CCS_10|BREAST NEOPLASM MALIGNANT MALE AREOLA PRIMARY
C0346858|T047||CCS_10|MALIGNANT NEOPLASM OF AREOLA OF MALE BREAST 
C0346858|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF AREOLA OF MALE BREAST 
C0346858|T047||CCS_10|BREAST NEOPLASM MALIGNANT MALE AREOLA
C0346858|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF AREOLA OF MALE BREAST
C0346858|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF AREOLA OF MALE BREAST 
C0346857|T047||CCS_10|MALIGNANT NEOPLASM OF NIPPLE OF MALE BREAST
C0346857|T047||CCS_10|MALIGNANT NEOPLASM OF NIPPLE OF MALE BREAST 
C0346857|T047||CCS_10|BREAST NEOPLASM MALIGNANT MALE NIPPLE
C0346857|T047||CCS_10|MALIGNANT NEOPLASM OF NIPPLE OF MALE BREAST 
C0346857|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF NIPPLE OF MALE BREAST 
C0346857|T047||CCS_10|BREAST NEOPLASM MALIGNANT MALE NIPPLE PRIMARY
C0346857|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF NIPPLE OF MALE BREAST
C0346857|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF NIPPLE OF MALE BREAST 
C0346862|T047||CCS_10|MALIGNANT NEOPLASM OF AREOLA OF FEMALE BREAST
C0346862|T047||CCS_10|MALIGNANT NEOPLASM OF AREOLA OF FEMALE BREAST 
C0346862|T047||CCS_10|BREAST NEOPLASM MALIGNANT FEMALE AREOLA
C0346862|T047||CCS_10|BREAST NEOPLASM MALIGNANT FEMALE AREOLA PRIMARY
C0346862|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF AREOLA OF FEMALE BREAST
C0346862|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF AREOLA OF FEMALE BREAST 
C0346862|T047||CCS_10|MALIGNANT NEOPLASM OF AREOLA OF FEMALE BREAST 
C0346862|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF AREOLA OF FEMALE BREAST 
C3649897|T047||CCS_10|MALIGNANT BREAST TISSUE NEOPLASM
C3649897|T047||CCS_10|MALIGNANT BREAST TISSUE NEOPLASM 
C3649897|T047||CCS_10|BREAST NEOPLASM MALIGNANT BREAST TISSUE
C1299258|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF BREAST
C1299258|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF BREAST 
C1299258|T047||CCS_10|BREAST NEOPLASM MALIGNANT PRIMARY
C1299258|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF BREAST 
C2216720|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING REGIONAL LYMPH NODE (N) NX 
C2216720|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING REGIONAL LYMPH NODE (N) NX
C2216720|T047||CCS_10|MALIGNANT BREAST NEOPLASM NX
C2216720|T047||CCS_10|BREAST CANCER TNM STAGING REGIONAL LYMPH NODE (N) NX
C2216720|T047||CCS_10|MALIGNANT TUMOR OF BREAST TNM STAGING REGIONAL LYMPH NODE (N) NX
C2216707|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING DISTANT METASTASIS (M) MX 
C2216707|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING DISTANT METASTASIS (M) MX
C2216707|T047||CCS_10|MALIGNANT BREAST NEOPLASM MX
C2216707|T047||CCS_10|MALIGNANT TUMOR OF BREAST TNM STAGING DISTANT METASTASIS (M) MX
C2216707|T047||CCS_10|BREAST CANCER TNM STAGING DISTANT METASTASIS (M) MX
C2216718|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING REGIONAL LYMPH NODE (N) N2
C2216718|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING REGIONAL LYMPH NODE (N) N2 
C2216718|T047||CCS_10|MALIGNANT BREAST NEOPLASM N2
C2216718|T047||CCS_10|MALIGNANT TUMOR OF BREAST TNM STAGING REGIONAL LYMPH NODE (N) N2
C2216718|T047||CCS_10|BREAST CANCER TNM STAGING REGIONAL LYMPH NODE (N) N2
C2216716|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING REGIONAL LYMPH NODE (N) N0 
C2216716|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING REGIONAL LYMPH NODE (N) N0
C2216716|T047||CCS_10|MALIGNANT BREAST NEOPLASM N0
C2216716|T047||CCS_10|MALIGNANT TUMOR OF BREAST TNM STAGING REGIONAL LYMPH NODE (N) N0
C2216716|T047||CCS_10|BREAST CANCER TNM STAGING REGIONAL LYMPH NODE (N) N0
C2216719|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING REGIONAL LYMPH NODE (N) N3
C2216719|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING REGIONAL LYMPH NODE (N) N3 
C2216719|T047||CCS_10|MALIGNANT BREAST NEOPLASM N3
C2216719|T047||CCS_10|BREAST CANCER TNM STAGING REGIONAL LYMPH NODE (N) N3
C2216719|T047||CCS_10|MALIGNANT TUMOR OF BREAST TNM STAGING REGIONAL LYMPH NODE (N) N3
C2216721|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING REGIONAL LYMPH NODES (N)
C2216721|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING REGIONAL LYMPH NODES (N) 
C2216721|T047||CCS_10|MALIGNANT BREAST NEOPLASM TNM STAGING OF REGIONAL LYMPH NODES (N)
C2216721|T047||CCS_10|BREAST CANCER TNM STAGING REGIONAL LYMPH NODES (N)
C2216721|T047||CCS_10|MALIGNANT TUMOR OF BREAST TNM STAGING REGIONAL LYMPH NODES (N)
C2216706|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING DISTANT METASTASIS (M) M1 
C2216706|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING DISTANT METASTASIS (M) M1
C2216706|T047||CCS_10|MALIGNANT BREAST NEOPLASM M1
C2216706|T047||CCS_10|BREAST CANCER TNM STAGING DISTANT METASTASIS (M) M1
C2216706|T047||CCS_10|MALIGNANT TUMOR OF BREAST TNM STAGING DISTANT METASTASIS (M) M1
C2216705|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING DISTANT METASTASIS (M) M0
C2216705|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING DISTANT METASTASIS (M) M0 
C2216705|T047||CCS_10|MALIGNANT BREAST NEOPLASM M0
C2216705|T047||CCS_10|BREAST CANCER TNM STAGING DISTANT METASTASIS (M) M0
C2216705|T047||CCS_10|MALIGNANT TUMOR OF BREAST TNM STAGING DISTANT METASTASIS (M) M0
C2216717|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING REGIONAL LYMPH NODE (N) N1 
C2216717|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING REGIONAL LYMPH NODE (N) N1
C2216717|T047||CCS_10|MALIGNANT BREAST NEOPLASM N1
C2216717|T047||CCS_10|MALIGNANT TUMOR OF BREAST TNM STAGING REGIONAL LYMPH NODE (N) N1
C2216717|T047||CCS_10|BREAST CANCER TNM STAGING REGIONAL LYMPH NODE (N) N1
C2216704|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING DISTANT METASTASIS (M)
C2216704|T047||CCS_10|MALIGNANT NEOPLASM OF BREAST TNM STAGING DISTANT METASTASIS (M) 
C2216704|T047||CCS_10|MALIGNANT BREAST NEOPLASM TNM STAGING OF DISTANT METASTASIS (M)
C2216704|T047||CCS_10|BREAST CANCER TNM STAGING DISTANT METASTASIS (M)
C2216704|T047||CCS_10|MALIGNANT TUMOR OF BREAST TNM STAGING DISTANT METASTASIS (M)
C3694291|T047||CCS_10|METASTASIS FROM MALIGNANT NEOPLASM OF BREAST
C3694291|T047||CCS_10|METASTASIS FROM MALIGNANT NEOPLASM OF BREAST 
C0346153|T047||CCS_10|BREAST CANCER, FAMILIAL
C0346153|T047||CCS_10|FAMILIAL BREAST CANCER
C0346153|T047||CCS_10|FAMILIAL BREAST CANCER 
C0346153|T047||CCS_10|FAMILIAL CANCER OF BREAST
C0346153|T047||CCS_10|FAMILIAL CANCER OF BREAST 
C0346153|T047||CCS_10|FAMILIAL CANCER OF THE BREAST
C0346153|T047||CCS_10|HEREDITARY BREAST CANCER
C0346153|T047||CCS_10|HEREDITARY BREAST CARCINOMA
C0346153|T047||CCS_10|FAMILIAL BREAST CARCINOMA
C1562029|T047||CCS_10|BREAST NEOPLASM MALIGNANT HORMONE RECEPTOR POSITIVE
C1562029|T047||CCS_10|HORMONE RECEPTOR POSITIVE MALIGNANT NEOPLASM OF BREAST
C1562029|T047||CCS_10|HORMONE RECEPTOR POSITIVE MALIGNANT NEOPLASM OF BREAST 
C1562029|T047||CCS_10|HORMONE RECEPTOR POSITIVE MALIGNANT NEOPLASM OF BREAST 
C3695123|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT BREAST NEOPLASM
C3695123|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT BREAST NEOPLASM 
C3695123|T047||CCS_10|BREAST NEOPLASM MALIGNANT LOCAL RECURRENCE
C3695122|T047||CCS_10|BREAST NEOPLASM MALIGNANT STAGING TNM PATHOLOGIC (PN)
C3695122|T047||CCS_10|MALIGNANT BREAST NEOPLASM PATHOLOGIC (PN) STAGING
C3695122|T047||CCS_10|MALIGNANT BREAST NEOPLASM PATHOLOGIC (PN) STAGING 
C0349669|T047||CCS_10|MALIGNANT LYMPHOMA OF BREAST
C0349669|T047||CCS_10|MALIGNANT LYMPHOMA OF BREAST 
C4031559|T047||CCS_10|BIOPSY OF BREAST SHOWED CARCINOMA MEDULLARY ATYPICAL
C4031559|T047||CCS_10|BIOPSY OF BREAST SHOWED ATYPICAL MEDULLARY CARCINOMA
C4031559|T047||CCS_10|BIOPSY OF BREAST SHOWED ATYPICAL MEDULLARY CARCINOMA 
C4031545|T047||CCS_10|BIOPSY OF BREAST SHOWED SIGNET RING CELL CARCINOMA 
C4031545|T047||CCS_10|BIOPSY OF BREAST SHOWED SIGNET RING CELL CARCINOMA
C4031545|T047||CCS_10|BIOPSY OF BREAST SHOWED CARCINOMA SIGNET RING CELL
C4031466|T047||CCS_10|BIOPSY OF BREAST SHOWED PRECURSOR CELL LYMPHOBLASTIC LYMPHOMA
C4031466|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA PRECURSOR CELL LYMPHOBLASTIC
C4031466|T047||CCS_10|BIOPSY OF BREAST SHOWED PRECURSOR CELL LYMPHOBLASTIC LYMPHOMA 
C4031512|T047||CCS_10|BIOPSY OF BREAST SHOWED EPITHELIOID HEMANGIOENDOTHELIOMA
C4031512|T047||CCS_10|BIOPSY OF BREAST SHOWED HEMANGIOENDOTHELIOMA EPITHELIOID
C4031512|T047||CCS_10|BIOPSY OF BREAST SHOWED EPITHELIOID HEMANGIOENDOTHELIOMA 
C4031503|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOMA WITH GRADE 1 NODULAR SCLEROSIS
C4031503|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOMA WITH GRADE 1 NODULAR SCLEROSIS 
C4031503|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOMA WITH NODULAR SCLEROSIS GRADE 1
C4031490|T047||CCS_10|BIOPSY OF BREAST SHOWED PLEOMORPHIC LIPOSARCOMA 
C4031490|T047||CCS_10|BIOPSY OF BREAST SHOWED LIPOSARCOMA PLEOMORPHIC
C4031490|T047||CCS_10|BIOPSY OF BREAST SHOWED PLEOMORPHIC LIPOSARCOMA
C4031482|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA COMPOSITE HODGKIN'S AND NON-HODGKIN'S
C4031482|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA COMPOSITE HODGKIN'S AND NON-HODGKIN'S 
C4031526|T047||CCS_10|BIOPSY OF BREAST SHOWED DUCT CARCINOMA, DESMOPLASTIC TYPE
C4031526|T047||CCS_10|BIOPSY OF BREAST SHOWED DUCT CARCINOMA, DESMOPLASTIC TYPE 
C4031526|T047||CCS_10|BIOPSY OF BREAST SHOWED CARCINOMA DUCT, DESMOPLASTIC TYPE
C4031523|T047||CCS_10|BIOPSY OF BREAST SHOWED FIBROSARCOMA 
C4031523|T047||CCS_10|BIOPSY OF BREAST SHOWED FIBROSARCOMA
C4031505|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOMA WITH LYMPHOCYTIC DEPLETION WITH DIFFUSE FIBROSIS
C4031505|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOMA WITH LYMPHOCYTIC DEPLETION WITH DIFFUSE FIBROSIS 
C4031494|T047||CCS_10|BIOPSY OF BREAST SHOWED LIPOSARCOMA DEDIFFERENTIATED
C4031494|T047||CCS_10|BIOPSY OF BREAST SHOWED DEDIFFERENTIATED LIPOSARCOMA
C4031494|T047||CCS_10|BIOPSY OF BREAST SHOWED DEDIFFERENTIATED LIPOSARCOMA 
C4031489|T047||CCS_10|BIOPSY OF BREAST SHOWED ROUND CELL LIPOSARCOMA
C4031489|T047||CCS_10|BIOPSY OF BREAST SHOWED LIPOSARCOMA ROUND CELL
C4031489|T047||CCS_10|BIOPSY OF BREAST SHOWED ROUND CELL LIPOSARCOMA 
C4031513|T047||CCS_10|BIOPSY OF BREAST SHOWED HEMANGIOENDOTHELIOMA
C4031513|T047||CCS_10|BIOPSY OF BREAST SHOWED HEMANGIOENDOTHELIOMA 
C4031488|T047||CCS_10|BIOPSY OF BREAST SHOWED WELL DIFFERENTIATED LIPOSARCOMA 
C4031488|T047||CCS_10|BIOPSY OF BREAST SHOWED WELL DIFFERENTIATED LIPOSARCOMA
C4031488|T047||CCS_10|BIOPSY OF BREAST SHOWED LIPOSARCOMA WELL DIFFERENTIATED
C4031479|T047||CCS_10|BIOPSY OF BREAST SHOWED GRADE 2 FOLLICULAR LYMPHOMA
C4031479|T047||CCS_10|BIOPSY OF BREAST SHOWED GRADE 2 FOLLICULAR LYMPHOMA 
C4031479|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA FOLLICULAR GRADE 2
C4031472|T047||CCS_10|BIOPSY OF BREAST SHOWED MANTLE CELL LYMPHOMA
C4031472|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA MANTLE CELL
C4031472|T047||CCS_10|BIOPSY OF BREAST SHOWED MANTLE CELL LYMPHOMA 
C4031465|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA PRECURSOR CELL LYMPHOBLASTIC B-CELL
C4031465|T047||CCS_10|BIOPSY OF BREAST SHOWED PRECURSOR B-CELL LYMPHOBLASTIC LYMPHOMA 
C4031465|T047||CCS_10|BIOPSY OF BREAST SHOWED PRECURSOR B-CELL LYMPHOBLASTIC LYMPHOMA
C4031464|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA PRECURSOR CELL LYMPHOBLASTIC T-CELL
C4031464|T047||CCS_10|BIOPSY OF BREAST SHOWED PRECURSOR T-CELL LYMPHOBLASTIC LYMPHOMA 
C4031464|T047||CCS_10|BIOPSY OF BREAST SHOWED PRECURSOR T-CELL LYMPHOBLASTIC LYMPHOMA
C4031529|T047||CCS_10|BIOPSY OF BREAST SHOWED EMBRYONAL CARCINOSARCOMA 
C4031529|T047||CCS_10|BIOPSY OF BREAST SHOWED CARCINOSARCOMA EMBRYONAL
C4031529|T047||CCS_10|BIOPSY OF BREAST SHOWED EMBRYONAL CARCINOSARCOMA
C4031521|T047||CCS_10|BIOPSY OF BREAST SHOWED FASCIAL FIBROSARCOMA
C4031521|T047||CCS_10|BIOPSY OF BREAST SHOWED FASCIAL FIBROSARCOMA 
C4031521|T047||CCS_10|BIOPSY OF BREAST SHOWED FIBROSARCOMA FASCIAL
C4031506|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOMA WITH LYMPHOCYTIC DEPLETION
C4031506|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOMA WITH LYMPHOCYTIC DEPLETION 
C4031493|T047||CCS_10|BIOPSY OF BREAST SHOWED FIBROBLASTIC LIPOSARCOMA 
C4031493|T047||CCS_10|BIOPSY OF BREAST SHOWED FIBROBLASTIC LIPOSARCOMA
C4031493|T047||CCS_10|BIOPSY OF BREAST SHOWED LIPOSARCOMA FIBROBLASTIC
C4031483|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA BURKITT'S
C4031483|T047||CCS_10|BIOPSY OF BREAST SHOWED BURKITT'S LYMPHOMA
C4031483|T047||CCS_10|BIOPSY OF BREAST SHOWED BURKITT'S LYMPHOMA 
C4031558|T047||CCS_10|BIOPSY OF BREAST SHOWED MEDULLARY CARCINOMA WITH LYMPHOID STROMA 
C4031558|T047||CCS_10|BIOPSY OF BREAST SHOWED CARCINOMA MEDULLARY WITH LYMPHOID STROMA
C4031558|T047||CCS_10|BIOPSY OF BREAST SHOWED MEDULLARY CARCINOMA WITH LYMPHOID STROMA
C4031502|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOMA WITH GRADE 2 NODULAR SCLEROSIS
C4031502|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOMA WITH GRADE 2 NODULAR SCLEROSIS 
C4031502|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOMA WITH NODULAR SCLEROSIS GRADE 2
C4031474|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOPLASMACYTIC LYMPHOMA
C4031474|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA LYMPHOPLASMACYTIC
C4031474|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOPLASMACYTIC LYMPHOMA 
C4031501|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOMA WITH NODULAR SCLEROSIS IN CELLULAR PHASE 
C4031501|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOMA WITH NODULAR SCLEROSIS IN CELLULAR PHASE
C4031467|T047||CCS_10|BIOPSY OF BREAST SHOWED NON-HODGKIN'S LYMPHOMA
C4031467|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA NON-HODGKIN'S
C4031467|T047||CCS_10|BIOPSY OF BREAST SHOWED NON-HODGKIN'S LYMPHOMA 
C4031455|T047||CCS_10|BIOPSY OF BREAST SHOWED MYXOID LEIOMYOSARCOMA 
C4031455|T047||CCS_10|BIOPSY OF BREAST SHOWED MYXOID LEIOMYOSARCOMA
C4031455|T047||CCS_10|BIOPSY OF BREAST SHOWED MYOSARCOMA LEIOMYOSARCOMA MYXOID
C4031580|T047||CCS_10|BIOPSY OF BREAST SHOWED COMEDOCARCINOMA 
C4031580|T047||CCS_10|BIOPSY OF BREAST SHOWED CARCINOMA COMEDOCARCINOMA
C4031580|T047||CCS_10|BIOPSY OF BREAST SHOWED COMEDOCARCINOMA
C4031560|T047||CCS_10|BIOPSY OF BREAST SHOWED MEDULLARY CARCINOMA 
C4031560|T047||CCS_10|BIOPSY OF BREAST SHOWED MEDULLARY CARCINOMA
C4031560|T047||CCS_10|BIOPSY OF BREAST SHOWED CARCINOMA MEDULLARY
C4031519|T047||CCS_10|BIOPSY OF BREAST SHOWED INFANTILE FIBROSARCOMA 
C4031519|T047||CCS_10|BIOPSY OF BREAST SHOWED INFANTILE FIBROSARCOMA
C4031519|T047||CCS_10|BIOPSY OF BREAST SHOWED FIBROSARCOMA INFANTILE
C4031511|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOMA 
C4031511|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOMA
C4031510|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOMA GRANULOMA
C4031510|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOMA GRANULOMA 
C4031463|T047||CCS_10|BIOPSY OF BREAST SHOWED SMALL B-CELL LYMPHOCYTIC LYMPHOMA
C4031463|T047||CCS_10|BIOPSY OF BREAST SHOWED SMALL B-CELL LYMPHOCYTIC LYMPHOMA 
C4031463|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA SMALL B-CELL LYMPHOCYTIC
C4031452|T047||CCS_10|BIOPSY OF BREAST SHOWED PLASMACYTOMA EXTRAMEDULLARY
C4031452|T047||CCS_10|BIOPSY OF BREAST SHOWED EXTRAMEDULLARY PLASMACYTOMA
C4031452|T047||CCS_10|BIOPSY OF BREAST SHOWED EXTRAMEDULLARY PLASMACYTOMA 
C4031567|T047||CCS_10|BIOPSY OF BREAST SHOWED INFILTRATING DUCTAL CARCINOMA MIXED WITH OTHER TYPES 
C4031567|T047||CCS_10|BIOPSY OF BREAST SHOWED CARCINOMA INFILTRATING DUCTAL MIXED WITH OTHER TYPES
C4031567|T047||CCS_10|BIOPSY OF BREAST SHOWED INFILTRATING DUCTAL CARCINOMA MIXED WITH OTHER TYPES
C4031518|T047||CCS_10|BIOPSY OF BREAST SHOWED FIBROSARCOMA, SOLITARY FIBROUS TUMOR 
C4031518|T047||CCS_10|BIOPSY OF BREAST SHOWED FIBROSARCOMA, SOLITARY FIBROUS TUMOR
C4031518|T047||CCS_10|BIOPSY OF BREAST SHOWED FIBROSARCOMA SOLITARY FIBROUS TUMOR
C4031456|T047||CCS_10|BIOPSY OF BREAST SHOWED EPITHELIOID LEIOMYOSARCOMA 
C4031456|T047||CCS_10|BIOPSY OF BREAST SHOWED MYOSARCOMA LEIOMYOSARCOMA EPITHELIOID
C4031456|T047||CCS_10|BIOPSY OF BREAST SHOWED EPITHELIOID LEIOMYOSARCOMA
C4031453|T047||CCS_10|BIOPSY OF BREAST SHOWED PLASMACYTOMA 
C4031453|T047||CCS_10|BIOPSY OF BREAST SHOWED PLASMACYTOMA
C4031602|T047||CCS_10|BIOPSY OF BREAST SHOWED ADENOCARCINOMA MUCIN-PRODUCING
C4031602|T047||CCS_10|BIOPSY OF BREAST SHOWED MUCIN-PRODUCING ADENOCARCINOMA
C4031602|T047||CCS_10|BIOPSY OF BREAST SHOWED MUCIN-PRODUCING ADENOCARCINOMA 
C4031527|T047||CCS_10|BIOPSY OF BREAST SHOWED CLEAR CELL TYPE NEOPLASM 
C4031527|T047||CCS_10|BIOPSY OF BREAST SHOWED CLEAR CELL TYPE NEOPLASM
C4031527|T047||CCS_10|BIOPSY OF BREAST SHOWED CLEAR CELL TYPE
C4031481|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA FOLLICULAR
C4031481|T047||CCS_10|BIOPSY OF BREAST SHOWED FOLLICULAR LYMPHOMA
C4031481|T047||CCS_10|BIOPSY OF BREAST SHOWED FOLLICULAR LYMPHOMA 
C4031480|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA FOLLICULAR GRADE 1
C4031480|T047||CCS_10|BIOPSY OF BREAST SHOWED GRADE 1 FOLLICULAR LYMPHOMA
C4031480|T047||CCS_10|BIOPSY OF BREAST SHOWED GRADE 1 FOLLICULAR LYMPHOMA 
C4031473|T047||CCS_10|BIOPSY OF BREAST SHOWED MALT LYMPHOMA
C4031473|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA MALT
C4031473|T047||CCS_10|BIOPSY OF BREAST SHOWED MALT LYMPHOMA 
C4031469|T047||CCS_10|BIOPSY OF BREAST SHOWED MATURE T-CELL ANGIOIMMUNOBLASTIC LYMPHOMA 
C4031469|T047||CCS_10|BIOPSY OF BREAST SHOWED MATURE T-CELL ANGIOIMMUNOBLASTIC LYMPHOMA
C4031469|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA MATURE T-CELL ANGIOIMMUNOBLASTIC
C4031460|T047||CCS_10|BIOPSY OF BREAST SHOWED MESENCHYMOMA
C4031460|T047||CCS_10|BIOPSY OF BREAST SHOWED MESENCHYMOMA 
C4031600|T047||CCS_10|BIOPSY OF BREAST SHOWED POLYMORPHOUS ADENOCARCINOMA, LOW GRADE
C4031600|T047||CCS_10|BIOPSY OF BREAST SHOWED POLYMORPHOUS ADENOCARCINOMA, LOW GRADE 
C4031600|T047||CCS_10|BIOPSY OF BREAST SHOWED ADENOCARCINOMA POLYMORPHOUS, LOW GRADE
C4031522|T047||CCS_10|BIOPSY OF BREAST SHOWED ADENOFIBROSARCOMA
C4031522|T047||CCS_10|BIOPSY OF BREAST SHOWED ADENOFIBROSARCOMA 
C4031522|T047||CCS_10|BIOPSY OF BREAST SHOWED FIBROSARCOMA ADENOFIBROSARCOMA
C4031492|T047||CCS_10|BIOPSY OF BREAST SHOWED MIXED TYPE LIPOSARCOMA 
C4031492|T047||CCS_10|BIOPSY OF BREAST SHOWED MIXED TYPE LIPOSARCOMA
C4031492|T047||CCS_10|BIOPSY OF BREAST SHOWED LIPOSARCOMA MIXED TYPE
C4031478|T047||CCS_10|BIOPSY OF BREAST SHOWED GRADE 3 FOLLICULAR LYMPHOMA 
C4031478|T047||CCS_10|BIOPSY OF BREAST SHOWED GRADE 3 FOLLICULAR LYMPHOMA
C4031478|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA FOLLICULAR GRADE 3
C4031487|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA
C4031487|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA 
C4031462|T047||CCS_10|BIOPSY OF BREAST SHOWED MALIGNANT NEOPLASM 
C4031462|T047||CCS_10|BIOPSY OF BREAST SHOWED MALIGNANT NEOPLASM
C4031423|T047||CCS_10|BIOPSY OF BREAST SHOWED SMALL CELL TYPE NEOPLASM 
C4031423|T047||CCS_10|BIOPSY OF BREAST SHOWED SMALL CELL TYPE
C4031423|T047||CCS_10|BIOPSY OF BREAST SHOWED SMALL CELL TYPE NEOPLASM
C4031421|T047||CCS_10|BIOPSY OF BREAST SHOWED SPINDLE CELL TYPE NEOPLASM
C4031421|T047||CCS_10|BIOPSY OF BREAST SHOWED SPINDLE CELL TYPE
C4031421|T047||CCS_10|BIOPSY OF BREAST SHOWED SPINDLE CELL TYPE NEOPLASM 
C4031561|T047||CCS_10|BIOPSY OF BREAST SHOWED LOBULAR CARCINOMA MIXED WITH OTHER TYPES OF CARCINOMA 
C4031561|T047||CCS_10|BIOPSY OF BREAST SHOWED CARCINOMA LOBULAR MIXED WITH OTHER TYPES OF CARCINOM
C4031561|T047||CCS_10|BIOPSY OF BREAST SHOWED LOBULAR CARCINOMA MIXED WITH OTHER TYPES OF CARCINOMA
C4031528|T047||CCS_10|BIOPSY OF BREAST SHOWED MYOEPITHELIOMA CARCINOSARCOMA
C4031528|T047||CCS_10|BIOPSY OF BREAST SHOWED MYOEPITHELIOMA CARCINOSARCOMA 
C4031528|T047||CCS_10|BIOPSY OF BREAST SHOWED CARCINOSARCOMA MYOEPITHELIOMA
C4031520|T047||CCS_10|BIOPSY OF BREAST SHOWED FIBROMYXOSARCOMA
C4031520|T047||CCS_10|BIOPSY OF BREAST SHOWED FIBROSARCOMA FIBROMYXOSARCOMA
C4031520|T047||CCS_10|BIOPSY OF BREAST SHOWED FIBROMYXOSARCOMA 
C4031509|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOMA LYMPHOCYTE-RICH
C4031509|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOCYTE-RICH LYMPHOMA 
C4031509|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOCYTE-RICH LYMPHOMA
C4031504|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOMA WITH NODULAR SCLEROSIS
C4031504|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOMA WITH NODULAR SCLEROSIS 
C4031471|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA MARGINAL ZONE B-CELL
C4031471|T047||CCS_10|BIOPSY OF BREAST SHOWED MARGINAL ZONE B-CELL LYMPHOMA
C4031471|T047||CCS_10|BIOPSY OF BREAST SHOWED MARGINAL ZONE B-CELL LYMPHOMA 
C4031470|T047||CCS_10|BIOPSY OF BREAST SHOWED MATURE T-CELL LYMPHOMA
C4031470|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA MATURE T-CELL
C4031470|T047||CCS_10|BIOPSY OF BREAST SHOWED MATURE T-CELL LYMPHOMA 
C4031459|T047||CCS_10|BIOPSY OF BREAST SHOWED MYOSARCOMA 
C4031459|T047||CCS_10|BIOPSY OF BREAST SHOWED MYOSARCOMA
C4031546|T047||CCS_10|BIOPSY OF BREAST SHOWED SECRETORY CARCINOMA
C4031546|T047||CCS_10|BIOPSY OF BREAST SHOWED CARCINOMA SECRETORY
C4031546|T047||CCS_10|BIOPSY OF BREAST SHOWED SECRETORY CARCINOMA 
C4031507|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOMA SARCOMA
C4031507|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN SARCOMA
C4031507|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN SARCOMA 
C4031475|T047||CCS_10|BIOPSY OF BREAST SHOWED DIFFUSE LARGE B-CELL IMMUNOBLASTIC LYMPHOMA
C4031475|T047||CCS_10|BIOPSY OF BREAST SHOWED DIFFUSE LARGE B-CELL IMMUNOBLASTIC LYMPHOMA 
C4031475|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA LARGE B-CELL, DIFFUSE IMMUNOBLASTIC
C4031461|T047||CCS_10|BIOPSY OF BREAST SHOWED MASTOCYTOSIS
C4031461|T047||CCS_10|BIOPSY OF BREAST SHOWED MASTOCYTOSIS 
C4031429|T047||CCS_10|BIOPSY OF BREAST SHOWED SARCOMA NEUROSARCOMA
C4031429|T047||CCS_10|BIOPSY OF BREAST SHOWED NEUROSARCOMA
C4031429|T047||CCS_10|BIOPSY OF BREAST SHOWED NEUROSARCOMA 
C4031586|T047||CCS_10|BIOPSY OF BREAST SHOWED ACINAR CELL CARCINOMA 
C4031586|T047||CCS_10|BIOPSY OF BREAST SHOWED ACINAR CELL CARCINOMA
C4031586|T047||CCS_10|BIOPSY OF BREAST SHOWED CARCINOMA ACINAR CELL
C4031496|T047||CCS_10|BIOPSY OF BREAST SHOWED LARGE CELL NEUROENDOCRINE CARCINOMA
C4031496|T047||CCS_10|BIOPSY OF BREAST SHOWED CARCINOMA LARGE CELL NEUROENDOCRINE
C4031496|T047||CCS_10|BIOPSY OF BREAST SHOWED LARGE CELL NEUROENDOCRINE CARCINOMA 
C4031530|T047||CCS_10|BIOPSY OF BREAST SHOWED CARCINOSARCOMA
C4031530|T047||CCS_10|BIOPSY OF BREAST SHOWED CARCINOSARCOMA 
C4031495|T047||CCS_10|BIOPSY OF BREAST SHOWED LIPOSARCOMA 
C4031495|T047||CCS_10|BIOPSY OF BREAST SHOWED LIPOSARCOMA
C4031477|T047||CCS_10|BIOPSY OF BREAST SHOWED HISTIOCYTOSIS LYMPHOMA
C4031477|T047||CCS_10|BIOPSY OF BREAST SHOWED HISTIOCYTOSIS LYMPHOMA 
C4031477|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA HISTIOCYTOSIS
C4031476|T047||CCS_10|BIOPSY OF BREAST SHOWED DIFFUSE LARGE B-CELL LYMPHOMA 
C4031476|T047||CCS_10|BIOPSY OF BREAST SHOWED DIFFUSE LARGE B-CELL LYMPHOMA
C4031476|T047||CCS_10|BIOPSY OF BREAST SHOWED LYMPHOMA LARGE B-CELL, DIFFUSE
C4031457|T047||CCS_10|BIOPSY OF BREAST SHOWED MYOSARCOMA LEIOMYOSARCOMA
C4031457|T047||CCS_10|BIOPSY OF BREAST SHOWED LEIOMYOSARCOMA 
C4031457|T047||CCS_10|BIOPSY OF BREAST SHOWED LEIOMYOSARCOMA
C4031585|T047||CCS_10|BIOPSY OF BREAST SHOWED ACINAR CELL CYSTADENOCARCINOMA
C4031585|T047||CCS_10|BIOPSY OF BREAST SHOWED ACINAR CELL CYSTADENOCARCINOMA 
C4031585|T047||CCS_10|BIOPSY OF BREAST SHOWED CARCINOMA ACINAR CELL CYSTADENOCARCINOMA
C4031515|T047||CCS_10|BIOPSY OF BREAST SHOWED GIANT CELL TYPE NEOPLASM 
C4031515|T047||CCS_10|BIOPSY OF BREAST SHOWED GIANT CELL TYPE NEOPLASM
C4031515|T047||CCS_10|BIOPSY OF BREAST SHOWED GIANT CELL TYPE
C4031508|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S MIXED CELLULARITY LYMPHOMA
C4031508|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S LYMPHOMA MIXED CELLULARITY
C4031508|T047||CCS_10|BIOPSY OF BREAST SHOWED HODGKIN'S MIXED CELLULARITY LYMPHOMA 
C4031491|T047||CCS_10|BIOPSY OF BREAST SHOWED MYXOID LIPOSARCOMA 
C4031491|T047||CCS_10|BIOPSY OF BREAST SHOWED MYXOID LIPOSARCOMA
C4031491|T047||CCS_10|BIOPSY OF BREAST SHOWED LIPOSARCOMA MYXOID
C4031458|T047||CCS_10|BIOPSY OF BREAST SHOWED ANGIOMYOSARCOMA
C4031458|T047||CCS_10|BIOPSY OF BREAST SHOWED MYOSARCOMA ANGIOMYOSARCOMA
C4031458|T047||CCS_10|BIOPSY OF BREAST SHOWED ANGIOMYOSARCOMA 
C0346787|T047||CCS_10|MALIGNANT MELANOMA OF BREAST
C0346787|T047||CCS_10|MALIGNANT MELANOMA OF BREAST 
C0346787|T047||CCS_10|BREAST; MELANOMA
C0346787|T047||CCS_10|MELANOMA; BREAST
C0346787|T047||CCS_10|MALIGNANT BREAST MELANOMA
C0346787|T047||CCS_10|MALIGNANT MELANOMA OF THE BREAST
C0346787|T047||CCS_10|BREAST MELANOMA
C0346986|T047||CCS_10|METASTASIS OF MALIGNANT NEOPLASM TO SKIN OF BREAST 
C0346986|T047||CCS_10|METASTASIS OF MALIGNANT NEOPLASM TO SKIN OF BREAST
C0346986|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SKIN OF BREAST 
C0346986|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SKIN OF BREAST
C0346986|T047||CCS_10|SKIN NEOPLASM MALIGNANT BREAST SECONDARY
C0346986|T047||CCS_10|SECONDARY MALIGNANT SKIN NEOPLASM OF BREAST 
C0346986|T047||CCS_10|SECONDARY MALIGNANT SKIN NEOPLASM OF BREAST
C0346986|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO SKIN OF BREAST
C1282471|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOR OF BREAST 
C1282471|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOR OF BREAST
C1282471|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOUR OF BREAST
C1134719|T047||CCS_10|CARCINOMAS, INFILTRATING DUCT
C1134719|T047||CCS_10|INVASIVE DUCTAL BREAST CARCINOMA
C1134719|T047||CCS_10|INFILTRATING DUCTAL CARCINOMA OF BREAST
C1134719|T047||CCS_10|INFILTRATING DUCTAL CARCINOMA OF BREAST 
C1134719|T047||CCS_10|CARCINOMA, DUCTAL, BREAST
C1134719|T047||CCS_10|CARCINOMA, INVASIVE DUCTAL, BREAST
C1134719|T047||CCS_10|INVASIVE DUCTAL CARCINOMA, BREAST
C1134719|T047||CCS_10|CARCINOMA, DUCTAL, BREAST [DISEASE/FINDING]
C1134719|T047||CCS_10|CARCINOMA, INFILTRATING DUCT
C1134719|T047||CCS_10|INFILTRATING DUCTAL CARCINOMA
C1134719|T047||CCS_10|INVASIVE DUCTAL CARCINOMA, NOT OTHERWISE SPECIFIED
C1134719|T047||CCS_10|BREAST CANCER, INVASIVE DUCTAL
C1134719|T047||CCS_10|BREAST DUCTAL CANCER INFILTRATING
C1134719|T047||CCS_10|INVASIVE DUCTAL BREAST CANCER
C1134719|T047||CCS_10|BREAST DUCTAL CANCER INVASIVE
C1134719|T047||CCS_10|INFILTRATING DUCTAL BREAST CANCER
C1134719|T047||CCS_10|INFILTRATING DUCTULAR CARCINOMA
C1134719|T047||CCS_10|INFILTRATING DUCTULAR CARCINOMA (MORPHOLOGIC ABNORMALITY)
C1134719|T047||CCS_10|INFILTRATING DUCT CARCINOMA OF BREAST 
C1134719|T047||CCS_10|INFILTRATING DUCT CARCINOMA OF BREAST
C1134719|T047||CCS_10|INVASIVE DUCT CARCINOMA OF BREAST
C1134719|T047||CCS_10|INVASIVE DUCTAL CARCINOMA OF BREAST
C1134719|T047||CCS_10|DUCTAL INVASIVE BREAST CARCINOMA
C1134719|T047||CCS_10|CARCINOMA; DUCTAL, INFILTRATING, UNSPECIFIED SITE
C1134719|T047||CCS_10|CARCINOMA; DUCTULAR, INFILTRATING, UNSPECIFIED SITE
C1134719|T047||CCS_10|CARCINOMA; INFILTRATING DUCT, UNSPECIFIED SITE
C1134719|T047||CCS_10|CARCINOMA; INFILTRATING DUCTULAR, UNSPECIFIED SITE
C1134719|T047||CCS_10|DUCTAL; CARCINOMA, INFILTRATING, UNSPECIFIED SITE
C1134719|T047||CCS_10|DUCTULAR; CARCINOMA, INFILTRATING, UNSPECIFIED SITE
C1134719|T047||CCS_10|INFILTRATING; DUCTAL ADENOCARCINOMA, UNSPECIFIED SITE
C1134719|T047||CCS_10|INFILTRATING; DUCTAL CARCINOMA, UNSPECIFIED SITE
C1134719|T047||CCS_10|INFILTRATING; DUCTULAR CARCINOMA, UNSPECIFIED SITE
C1134719|T047||CCS_10|INFILTRATING DUCTAL ADENOCARCINOMA
C1134719|T047||CCS_10|INFILTRATING DUCTAL BREAST CARCINOMA
C1134719|T047||CCS_10|INFILTRATING DUCTAL CARCINOMA OF THE BREAST
C1134719|T047||CCS_10|INVASIVE DUCTAL ADENOCARCINOMA
C1134719|T047||CCS_10|INVASIVE DUCTAL CARCINOMA OF THE BREAST
C1134719|T047||CCS_10|INVASIVE DUCTAL CARCINOMA, NOS
C1134719|T047||CCS_10|INVASIVE DUCTAL CARCINOMA, NST
C1134719|T047||CCS_10|INVASIVE DUCTAL CARCINOMA
C1134719|T047||CCS_10|INVASIVE DUCTAL CARCINOMA, NO SPECIFIC TYPE
C1386255|T047||CCS_10|DUCTAL; INFILTRATING ADENOCARCINOMA, UNSPECIFIED SITE, FEMALE
C1386255|T047||CCS_10|ADENOCARCINOMA; DUCTAL INFILTRATING, UNSPECIFIED SITE, FEMALE
C1386267|T047||CCS_10|ADENOCARCINOMA; INFILTRATING DUCT, UNSPECIFIED SITE
C1386268|T047||CCS_10|ADENOCARCINOMA; INFILTRATING DUCT, UNSPECIFIED SITE, FEMALE
C1386269|T047||CCS_10|INFLAMMATORY; ADENOCARCINOMA, UNSPECIFIED SITE
C1386269|T047||CCS_10|ADENOCARCINOMA; INFLAMMATORY, UNSPECIFIED SITE
C1386276|T047||CCS_10|ADENOCARCINOMA; INTRADUCTAL, NONINFILTRATING, PAPILLARY, WITH INVASION, UNSPECIFIED SITE
C1386278|T047||CCS_10|ADENOCARCINOMA; INTRADUCTAL, PAPILLARY, WITH INVASION, UNSPECIFIED SITE
C1386278|T047||CCS_10|ADENOCARCINOMA; PAPILLARY, INTRADUCTAL, WITH INVASION, UNSPECIFIED SITE
C1386278|T047||CCS_10|PAPILLARY; ADENOCARCINOMA, INTRADUCTAL, WITH INVASION, UNSPECIFIED SITE
C1386282|T047||CCS_10|LOBULAR; ADENOCARCINOMA, UNSPECIFIED SITE
C1386282|T047||CCS_10|ADENOCARCINOMA; LOBULAR, UNSPECIFIED SITE
C1391891|T047||CCS_10|BREAST; CARCINOMA IN SITU, LOBULAR WITH INFILTRATING DUCT
C1391891|T047||CCS_10|CARCINOMA IN SITU; LOBULAR WITH INFILTRATING DUCT, BREAST
C1391891|T047||CCS_10|LOBULAR; CARCINOMA IN SITU, WITH INFILTRATING DUCT, BREAST
C1391892|T047||CCS_10|CARCINOMA IN SITU; LOBULAR WITH INFILTRATING DUCT, UNSPECIFIED SITE
C1391892|T047||CCS_10|LOBULAR; CARCINOMA IN SITU, WITH INFILTRATING DUCT, UNSPECIFIED SITE
C1391902|T047||CCS_10|CARCINOMA; DUCTAL WITH LOBULAR (INFILTRATING), UNSPECIFIED SITE
C1391902|T047||CCS_10|DUCTAL; CARCINOMA WITH LOBULAR (INFILTRATING), UNSPECIFIED SITE
C1391903|T047||CCS_10|CARCINOMA; DUCTAL, INFILTRATING, WITH LOBULAR CARCINOMA IN SITU, UNSPECIFIED SITE
C1391903|T047||CCS_10|DUCTAL; CARCINOMA, INFILTRATING, WITH LOBULAR CARCINOMA IN SITU, UNSPECIFIED SITE
C1391904|T047||CCS_10|CARCINOMA; DUCTAL, INFILTRATING, WITH LOBULAR CARCINOMA, UNSPECIFIED SITE
C1391904|T047||CCS_10|DUCTAL; CARCINOMA, INFILTRATING, WITH LOBULAR CARCINOMA, UNSPECIFIED SITE
C1391904|T047||CCS_10|INFILTRATING; DUCTAL CARCINOMA, WITH LOBULAR CARCINOMA, UNSPECIFIED SITE
C0334384|T047||CCS_10|CARCINOMA OF BREAST WITH DUCTAL AND LOBULAR FEATURES 
C0334384|T047||CCS_10|CARCINOMA OF BREAST WITH DUCTAL AND LOBULAR FEATURES
C0334384|T047||CCS_10|MIXED DUCTAL AND LOBULAR CARCINOMA OF BREAST
C0334384|T047||CCS_10|INFILTRATING DUCT AND LOBULAR CARCINOMA
C0334384|T047||CCS_10|INFILTRATING DUCT AND LOBULAR CARCINOMA 
C0334384|T047||CCS_10|BREAST NEOPLASM MALIGNANT CARCINOMA WITH DUCTAL AND LOBULAR FEATURES
C0334384|T047||CCS_10|CARCINOMA OF BREAST WITH DUCTAL AND LOBULAR FEATURES 
C0334384|T047||CCS_10|[M] INFILTRATING DUCT AND LOBULAR CARCINOMA
C0334384|T047||CCS_10|[M]INFILTRATING DUCT AND LOBULAR CARCINOMA
C0334384|T047||CCS_10|MIXED DUCTAL LOBULAR BREAST CARCINOMA
C0334384|T047||CCS_10|INFILTRATING DUCT AND LOBULAR CARCINOMA IN SITU
C0334384|T047||CCS_10|INTRADUCTAL AND LOBULAR CARCINOMA
C0334384|T047||CCS_10|LOBULAR AND DUCTAL CARCINOMA
C0334384|T047||CCS_10|INFILTRATING DUCT AND LOBULAR CARCINOMA (MORPHOLOGIC ABNORMALITY)
C0334384|T047||CCS_10|INFILTRATING LOBULAR CARCINOMA AND DUCTAL CARCINOMA IN SITU
C0334384|T047||CCS_10|CARCINOMA; INFILTRATING DUCT WITH LOBULAR CA, UNSPECIFIED SITE
C0334384|T047||CCS_10|DCIS AND ILC
C0334384|T047||CCS_10|DCIS AND INFILTRATING LOBULAR CARCINOMA
C0334384|T047||CCS_10|DUCTAL CARCINOMA IN SITU AND INFILTRATING LOBULAR CARCINOMA
C0334384|T047||CCS_10|DUCTAL AND LOBULAR CARCINOMA
C0334384|T047||CCS_10|INFILTRATING DUCTAL AND LOBULAR CARCINOMA IN SITU
C0334384|T047||CCS_10|LCIS AND INFILTRATING DUCTAL CARCINOMA
C0334384|T047||CCS_10|LOBULAR CARCINOMA IN SITU AND INFILTRATING DUCTAL CARCINOMA
C0334384|T047||CCS_10|LOBULAR CARCINOMA IN SITU AND INVASIVE DUCTAL CARCINOMA
C0334384|T047||CCS_10|MIXED DUCTAL AND LOBULAR BREAST CARCINOMA
C0334384|T047||CCS_10|MIXED DUCTAL AND LOBULAR CARCINOMA OF THE BREAST
C0334384|T047||CCS_10|MIXED LOBULAR AND DUCTAL BREAST CARCINOMA
C0334384|T047||CCS_10|MIXED LOBULAR AND DUCTAL CARCINOMA OF BREAST
C0334384|T047||CCS_10|MIXED LOBULAR AND DUCTAL CARCINOMA OF THE BREAST
C0334384|T047||CCS_10|MIXED LOBULAR AND DUCTAL CARCINOMA
C0334384|T047||CCS_10|NON-INFILTRATING DUCTAL CARCINOMA AND ILC
C0334384|T047||CCS_10|NON-INFILTRATING DUCTAL CARCINOMA AND INFILTRATING LOBULAR CARCINOMA
C0334384|T047||CCS_10|DUCTAL BREAST CARCINOMA IN SITU AND INVASIVE LOBULAR CARCINOMA
C0334384|T047||CCS_10|INVASIVE DUCTAL AND LOBULAR CARCINOMA IN SITU
C0334385|T047||CCS_10|INFLAMMATORY ADENOCARCINOMA
C0334385|T047||CCS_10|INFLAMMATORY CARCINOMA
C0334385|T047||CCS_10|INFLAMMATORY CARCINOMA (MORPHOLOGIC ABNORMALITY)
C0334385|T047||CCS_10|CARCINOMA; INFLAMMATORY, UNSPECIFIED SITE
C0334385|T047||CCS_10|INFLAMMATORY; CARCINOMA, UNSPECIFIED SITE
C1391916|T047||CCS_10|CARCINOMA; INTRADUCTAL, PAPILLARY WITH INVASION, UNSPECIFIED SITE
C1391916|T047||CCS_10|INTRADUCTAL; CARCINOMA, PAPILLARY WITH INVASION, UNSPECIFIED SITE
C0334318|T047||CCS_10|LIPID-RICH CARCINOMA 
C0334318|T047||CCS_10|LIPID-RICH CARCINOMA
C0334318|T047||CCS_10|[M] LIPID-RICH CARCINOMA
C0334318|T047||CCS_10|[M]LIPID-RICH CARCINOMA
C0334318|T047||CCS_10|LIPID-RICH CARCINOMA (MORPHOLOGIC ABNORMALITY)
C0334318|T047||CCS_10|CARCINOMA; LIPID-RICH
C0334318|T047||CCS_10|LIPID-RICH; CARCINOMA
C1391922|T047||CCS_10|CARCINOMA; LOBULAR WITH INTRADUCTAL, UNSPECIFIED SITE
C1391923|T047||CCS_10|CARCINOMA; LOBULAR, UNSPECIFIED SITE
C1391923|T047||CCS_10|LOBULAR; CARCINOMA, UNSPECIFIED SITE
C0334380|T047||CCS_10|MEDULLARY CARCINOMA WITH LYMPHOID STROMA
C0334380|T047||CCS_10|MEDULLARY CARCINOMA WITH LYMPHOID STROMA (MORPHOLOGIC ABNORMALITY)
C0334380|T047||CCS_10|CARCINOMA; MEDULLARY WITH LYMPHOID STROMA, UNSPECIFIED SITE
C0334380|T047||CCS_10|MEDULLARY; CARCINOMA WITH LYMPHOID STROMA, UNSPECIFIED SITE
C1391934|T047||CCS_10|CARCINOMA; PAPILLARY, INTRADUCTAL (NONINFILTRATING), WITH INVASION, UNSPECIFIED SITE
C1391934|T047||CCS_10|PAPILLARY; CARCINOMA, INTRADUCTAL (NONINFILTRATING), WITH INVASION, UNSPECIFIED SITE
C1403125|T047||CCS_10|LOBULAR; CARCINOMA, WITH INTRADUCTAL CARCINOMA, UNSPECIFIED SITE
C0279855|T047||CCS_10|CELLULAR DIAGNOSIS, BREAST CANCER
C0279855|T047||CCS_10|BREAST CANCER CELLULAR DIAGNOSIS
C0281663|T047||CCS_10|BREAST CANCER AND PREGNANCY
C0281663|T047||CCS_10|PREGNANCY AND BREAST CANCER
C0238033|T047||CCS_10|CANCER, MALE BREAST
C0238033|T047||CCS_10|CARCINOMA OF MALE BREAST
C0238033|T047||CCS_10|BREAST CANCER, MALE
C0238033|T047||CCS_10|MALE BREAST CANCER
C0238033|T047||CCS_10|CA BREAST - MALE 
C0238033|T047||CCS_10|CA BREAST - MALE
C0238033|T047||CCS_10|CARCINOMA OF MALE BREAST 
C0238033|T047||CCS_10|BREAST NEOPLASM MALIGNANT MALE CARCINOMA
C0238033|T047||CCS_10|BREAST CANCER MALE NOS
C0238033|T047||CCS_10|CANCER OF MALE BREAST
C0238033|T047||CCS_10|BREAST CANCER MALE
C0238033|T047||CCS_10|BREAST CARCINOMA, MALE
C0238033|T047||CCS_10|CARCINOMA OF MALE BREAST 
C0238033|T047||CCS_10|MALE BREAST CARCINOMA
C0238033|T047||CCS_10|CARCINOMA, MALE BREAST
C0238033|T047||CCS_10|CARCINOMA OF THE MALE BREAST
C0238033|T047||CCS_10|CARCINOMA;BREAST;M
C0238033|T047||CCS_10|CARCINOMA OF THE BREAST
C0346993|T047||CCS_10|METASTATIC NEOPLASM TO THE BREAST
C0346993|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BREAST 
C0346993|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BREAST
C0346993|T047||CCS_10|METASTASES TO BREAST
C0346993|T047||CCS_10|SECOND MALIG NEO BREAST
C0346993|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF FEMALE BREAST 
C0346993|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF FEMALE BREAST
C0346993|T047||CCS_10|BREAST NEOPLASM MALIGNANT FEMALE SECONDARY
C0346993|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO THE BREAST
C0346993|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM IN THE BREAST
C0346993|T047||CCS_10|BREAST METASTASES
C0346993|T047||CCS_10|METASTASIS TO BREAST
C0346993|T047||CCS_10|SECONDARY MALIGNANT DEPOSIT TO BREAST
C0346993|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO FEMALE BREAST
C0346993|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF FEMALE BREAST 
C0346993|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO FEMALE BREAST, NOS
C0346993|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF FEMALE BREAST, NOS
C0346993|T047||CCS_10|METASTATIC CANCER TO THE BREAST
C0346993|T047||CCS_10|METASTATIC TUMOR TO THE BREAST
C0346993|T047||CCS_10|BREAST METASTASIS
C1334565|T047||CCS_10|MALIGNANT BREAST ECCRINE SPIRADENOMA
C1334565|T047||CCS_10|MALIGNANT ECCRINE SPIRADENOMA OF BREAST
C1334565|T047||CCS_10|MALIGNANT ECCRINE SPIRADENOMA OF THE BREAST
C1334564|T047||CCS_10|MALIGNANT ADENOMYOEPITHELIOMA OF BREAST
C1334564|T047||CCS_10|MALIGNANT ADENOMYOEPITHELIOMA OF THE BREAST
C1334564|T047||CCS_10|MALIGNANT BREAST ADENOMYOEPITHELIOMA
C1334564|T047||CCS_10|BREAST ADENOMYOEPITHELIOMA WITH MALIGNANT CHANGE
C1704251|T047||CCS_10|PRIMARY BREAST LYMPHOMA
C1704251|T047||CCS_10|BREAST LYMPHOMA
C1704251|T047||CCS_10|LYMPHOMA OF BREAST
C1704251|T047||CCS_10|LYMPHOMA OF THE BREAST
C0859086|T047||CCS_10|MALIGNANT NIPPLE NEOPLASM NOS
C0859086|T047||CCS_10|MALIGNANT NIPPLE NEOPLASM
C0859086|T047||CCS_10|MALIGNANT NEOPLASM OF NIPPLE
C0859086|T047||CCS_10|MALIGNANT NEOPLASM OF THE NIPPLE
C0859086|T047||CCS_10|MALIGNANT NIPPLE TUMOR
C0859086|T047||CCS_10|MALIGNANT TUMOR OF NIPPLE
C0859086|T047||CCS_10|MALIGNANT TUMOR OF THE NIPPLE
C2211713|T047||CCS_10|MAST CELL SARCOMA OF BREAST 
C2211713|T047||CCS_10|MAST CELL SARCOMA OF BREAST
C0345867|T047||CCS_10|CARCINOMA IN SITU OF DESCENDING COLON
C0345867|T047||CCS_10|CARCINOMA IN SITU OF DESCENDING COLON 
C0700315|T047||CCS_10|LARGE INTESTINE ADENOCARCINOMA - SPLENIC FLEXURE CARCINOMA
C0700315|T047||CCS_10|CARCINOMA OF SPLENIC FLEXURE
C0700315|T047||CCS_10|CARCINOMA OF SPLENIC FLEXURE 
C0700315|T047||CCS_10|CARCINOMA OF SPLENIC FLEXURE 
C0728951|T047||CCS_10|CARCINOMA OF APPENDIX
C0728951|T047||CCS_10|CARCINOMA OF APPENDIX 
C0728951|T047||CCS_10|APPENDIX CANCER
C0728951|T047||CCS_10|(CA APPENDIX) OR (APPENDIX CARCINOMA)
C0728951|T047||CCS_10|APPENDIX CARCINOMA
C0728951|T047||CCS_10|CA APPENDIX
C0728951|T047||CCS_10|(CA APPENDIX) OR (APPENDIX CARCINOMA) 
C0728951|T047||CCS_10|CARCINOMA OF THE APPENDIX
C0856355|T047||CCS_10|CANCER OF SIGMOID COLON (EXCLUDING RECTOSIGMOID)
C0856355|T047||CCS_10|CANCER OF SIGMOID COLON (EXCL RECTOSIGMOID)
C0153439|T047||CCS_10|MALIGNANT NEOPLASM OF ASCENDING COLON
C0153439|T047||CCS_10|ASCENDING COLON
C0153439|T047||CCS_10|MALIGNANT NEOPLASM OF ASCENDING COLON 
C0153439|T047||CCS_10|CANCER OF ASCENDING COLON
C0153439|T047||CCS_10|MALIGNANT TUMOR OF ASCENDING COLON
C0153439|T047||CCS_10|MALIG NEO ASCEND COLON
C0153439|T047||CCS_10|CA ASCENDING COLON 
C0153439|T047||CCS_10|CA ASCENDING COLON
C0153439|T047||CCS_10|ASCENDING COLON CANCER
C0153439|T047||CCS_10|MALIGNANT TUMOUR OF ASCENDING COLON
C0153439|T047||CCS_10|MALIGNANT TUMOR OF ASCENDING COLON 
C0153439|T047||CCS_10|MALIGNANT NEOPLASM OF RIGHT COLON
C0496779|T047||CCS_10|MALIGNANT NEOPLASM OF APPENDIX
C0496779|T047||CCS_10|MALIGNANT NEOPLASM OF APPENDIX 
C0496779|T047||CCS_10|MALIGNANT APPENDICEAL NEOPLASM
C0496779|T047||CCS_10|MALIGNANT TUMOR OF APPENDIX
C0496779|T047||CCS_10|MALIGNANT NEO APPENDIX
C0496779|T047||CCS_10|APPENDIX CANCER
C0496779|T047||CCS_10|MALIGNANT NEOPLASM OF APPENDIX VERMIFORMIS
C0496779|T047||CCS_10|CANCER, APPENDICEAL
C0496779|T047||CCS_10|CANCER OF THE APPENDIX
C0496779|T047||CCS_10|CANCER OF APPENDIX
C0496779|T047||CCS_10|CANCER, APPENDIX
C0496779|T047||CCS_10|MALIGNANT TUMOUR OF APPENDIX
C0496779|T047||CCS_10|MALIGNANT TUMOR OF APPENDIX 
C0496779|T047||CCS_10|MALIGNANT APPENDIX NEOPLASM
C0496779|T047||CCS_10|MALIGNANT APPENDIX TUMOR
C0496779|T047||CCS_10|MALIGNANT NEOPLASM OF THE APPENDIX
C0496779|T047||CCS_10|MALIGNANT TUMOR OF THE APPENDIX
C0496779|T047||CCS_10|APPENDICEAL CANCER
C0349051|T047||CCS_10|MALIGNANT NEOPLASM OVERLAPPING COLON SITE
C0349051|T047||CCS_10|OVERLAPPING LESION OF COLON
C0349051|T047||CCS_10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF COLON
C0349051|T047||CCS_10|MALIGNANT NEOPLASM, OVERLAPPING LESION OF COLON 
C0349051|T047||CCS_10|MALIGNANT NEOPLASM, OVERLAPPING LESION OF COLON
C0349051|T047||CCS_10|LARGE INTESTINE NEOPLASM MALIGNANT, OVERLAPPING LESION OF COLON
C0349051|T047||CCS_10|MALIGNANT NEOPLASM, OVERLAPPING LESION OF COLON 
C0153433|T047||CCS_10|MALIGNANT NEOPLASM OF HEPATIC FLEXURE
C0153433|T047||CCS_10|MALIGNANT NEOPLASM OF HEPATIC FLEXURE OF COLON
C0153433|T047||CCS_10|MALIGNANT NEOPLASM OF HEPATIC FLEXURE 
C0153433|T047||CCS_10|MALIGNANT TUMOR OF HEPATIC FLEXURE
C0153433|T047||CCS_10|MAL NEO HEPATIC FLEXURE
C0153433|T047||CCS_10|CA HEPATIC FLEXURE - COLON 
C0153433|T047||CCS_10|CA HEPATIC FLEXURE - COLON
C0153433|T047||CCS_10|HEPATIC FLEXURE COLON CANCER
C0153433|T047||CCS_10|MALIGNANT TUMOUR OF HEPATIC FLEXURE
C0153433|T047||CCS_10|MALIGNANT TUMOR OF HEPATIC FLEXURE 
C0153434|T047||CCS_10|MALIGNANT NEOPLASM OF TRANSVERSE COLON
C0153434|T047||CCS_10|MALIGNANT NEOPLASM OF TRANSVERSE COLON 
C0153434|T047||CCS_10|MALIGNANT TUMOR OF TRANSVERSE COLON
C0153434|T047||CCS_10|MAL NEO TRANSVERSE COLON
C0153434|T047||CCS_10|CA TRANSVERSE COLON
C0153434|T047||CCS_10|CA TRANSVERSE COLON 
C0153434|T047||CCS_10|CANCER OF TRANSVERSE COLON
C0153434|T047||CCS_10|TRANSVERSE COLON CANCER
C0153434|T047||CCS_10|MALIGNANT TUMOUR OF TRANSVERSE COLON
C0153434|T047||CCS_10|MALIGNANT TUMOR OF TRANSVERSE COLON 
C0153435|T047||CCS_10|MALIGNANT NEOPLASM OF DESCENDING COLON
C0153435|T047||CCS_10|MALIGNANT NEOPLASM OF DESCENDING COLON 
C0153435|T047||CCS_10|MALIGNANT TUMOR OF DESCENDING COLON
C0153435|T047||CCS_10|MAL NEO DESCEND COLON
C0153435|T047||CCS_10|CA DESCENDING COLON
C0153435|T047||CCS_10|CA DESCENDING COLON 
C0153435|T047||CCS_10|CANCER OF DESCENDING COLON
C0153435|T047||CCS_10|DESCENDING COLON CANCER
C0153435|T047||CCS_10|MALIGNANT TUMOUR OF DESCENDING COLON
C0153435|T047||CCS_10|MALIGNANT TUMOR OF DESCENDING COLON 
C0153435|T047||CCS_10|MALIGNANT NEOPLASM OF LEFT COLON
C0153436|T047||CCS_10|MALIGNANT NEOPLASM OF SIGMOID COLON
C0153436|T047||CCS_10|MALIGNANT NEOPLASM OF SIGMOID COLON 
C0153436|T047||CCS_10|MALIGNANT TUMOR OF SIGMOID COLON
C0153436|T047||CCS_10|MAL NEO SIGMOID COLON
C0153436|T047||CCS_10|CA SIGMOID COLON
C0153436|T047||CCS_10|CA SIGMOID COLON 
C0153436|T047||CCS_10|SIGMOID COLON CANCER
C0153436|T047||CCS_10|MALIGNANT TUMOUR OF SIGMOID COLON
C0153436|T047||CCS_10|MALIGNANT TUMOR OF SIGMOID COLON 
C0153443|T047||CCS_10|MALIGNANT NEOPLASM OF RECTOSIGMOID JUNCTION
C0153443|T047||CCS_10|MAL NEO RECTOSIGMOID JCT
C0153443|T047||CCS_10|MALIGNANT NEOPLASM OF RECTOSIGMOID (COLON)
C0153443|T047||CCS_10|RECTAL NEOPLASM MALIGNANT RECTOSIGMOID JUNCTION
C0153443|T047||CCS_10|MALIGNANT NEOPLASM OF RECTOSIGMOID JUNCTION 
C0153443|T047||CCS_10|RECTOSIGMOID COLON CANCER
C0153443|T047||CCS_10|CA RECTOSIGMOID JUNCTION
C0153443|T047||CCS_10|MALIGNANT TUMOR OF RECTOSIGMOID JUNCTION
C0153443|T047||CCS_10|MALIGNANT TUMOUR OF RECTOSIGMOID JUNCTION
C0153443|T047||CCS_10|MALIGNANT TUMOR OF RECTOSIGMOID JUNCTION 
C0153443|T047||CCS_10|MALIGNANT NEOPLASM OF THE RECTOSIGMOID JUNCTION
C0153443|T047||CCS_10|MALIGNANT RECTOSIGMOID NEOPLASM
C0153443|T047||CCS_10|MALIGNANT RECTOSIGMOID TUMOR
C0153443|T047||CCS_10|MALIGNANT TUMOR OF THE RECTOSIGMOID JUNCTION
C0153443|T047||CCS_10|MALIGNANT NEOPLASM OF RECTOSIGMOID COLON
C0153443|T047||CCS_10|MALIGNANT NEOPLASM OF RECTOSIGMOID
C1096639|T047||CCS_10|MUCINOUS CYSTADENOCARCINOMA OF APPENDIX 
C1096639|T047||CCS_10|MUCINOUS CYSTADENOCARCINOMA OF APPENDIX
C1096639|T047||CCS_10|MUCINOUS CYSTADENOCARCINOMA APPENDIX
C1096639|T047||CCS_10|COLLOID CYSTADENOCARCINOMA OF APPENDIX
C1096639|T047||CCS_10|COLLOID CYSTADENOCARCINOMA OF THE APPENDIX
C1096639|T047||CCS_10|COLLOIDAL CYSTADENOCARCINOMA OF APPENDIX
C1096639|T047||CCS_10|COLLOIDAL CYSTADENOCARCINOMA OF THE APPENDIX
C1096639|T047||CCS_10|MUCINOUS CYSTADENOCARCINOMA OF THE APPENDIX
C1096639|T047||CCS_10|APPENDICEAL COLLOID CYSTADENOCARCINOMA
C1096639|T047||CCS_10|APPENDICEAL COLLOIDAL CYSTADENOCARCINOMA
C1096639|T047||CCS_10|APPENDICEAL MUCINOUS CYSTADENOCARCINOMA
C1096639|T047||CCS_10|APPENDIX COLLOID CYSTADENOCARCINOMA
C1096639|T047||CCS_10|APPENDIX COLLOIDAL CYSTADENOCARCINOMA
C1096639|T047||CCS_10|APPENDIX MUCINOUS CYSTADENOCARCINOMA
C0153440|T047||CCS_10|MALIGNANT NEOPLASM OF SPLENIC FLEXURE
C0153440|T047||CCS_10|MALIGNANT NEOPLASM OF SPLENIC FLEXURE OF COLON
C0153440|T047||CCS_10|MALIGNANT NEOPLASM OF SPLENIC FLEXURE 
C0153440|T047||CCS_10|MALIGNANT TUMOR OF SPLENIC FLEXURE
C0153440|T047||CCS_10|MAL NEO SPLENIC FLEXURE
C0153440|T047||CCS_10|CA SPLENIC FLEXURE - COLON 
C0153440|T047||CCS_10|CA SPLENIC FLEXURE - COLON
C0153440|T047||CCS_10|CANCER OF SPLENIC FLEXURE
C0153440|T047||CCS_10|SPLENIC FLEXURE COLON CANCER
C0153440|T047||CCS_10|MALIGNANT TUMOUR OF SPLENIC FLEXURE
C0153440|T047||CCS_10|MALIGNANT TUMOR OF SPLENIC FLEXURE 
C0153437|T047||CCS_10|MALIGNANT NEOPLASM OF CECUM
C0153437|T047||CCS_10|MALIGNANT NEOPLASM OF CAECUM
C0153437|T047||CCS_10|MALIGNANT NEOPLASM OF CECUM 
C0153437|T047||CCS_10|MALIGNANT TUMOR OF CECUM
C0153437|T047||CCS_10|MALIGNANT NEOPLASM CECUM
C0153437|T047||CCS_10|CA CAECUM
C0153437|T047||CCS_10|CA CECUM
C0153437|T047||CCS_10|CECUM--CANCER
C0153437|T047||CCS_10|CECAL CANCER
C0153437|T047||CCS_10|CAECAL CANCER
C0153437|T047||CCS_10|CANCER OF THE CECUM
C0153437|T047||CCS_10|CANCER, CECAL
C0153437|T047||CCS_10|CA - CANCER OF CAECUM
C0153437|T047||CCS_10|CA - CANCER OF CECUM
C0153437|T047||CCS_10|CANCER OF CAECUM
C0153437|T047||CCS_10|CANCER OF CECUM
C0153437|T047||CCS_10|MALIGNANT TUMOUR OF CAECUM
C0153437|T047||CCS_10|MALIGNANT TUMOR OF CECUM 
C0153437|T047||CCS_10|MALIGNANT CECUM NEOPLASM
C0153437|T047||CCS_10|MALIGNANT CECUM TUMOR
C0153437|T047||CCS_10|MALIGNANT NEOPLASM OF THE CECUM
C0153437|T047||CCS_10|MALIGNANT TUMOR OF THE CECUM
C0007102|T047||CCS_10|MALIGNANT NEOPLASM OF COLON
C0007102|T047||CCS_10|COLON CANCER
C0007102|T047||CCS_10|CANCER OF COLON
C0007102|T047||CCS_10|MALIGNANT NEOPLASM OF COLON, UNSPECIFIED
C0007102|T047||CCS_10|MALIGNANT TUMOR OF COLON
C0007102|T047||CCS_10|CANCERS, COLON
C0007102|T047||CCS_10|COLON CANCERS
C0007102|T047||CCS_10|CANCER, COLONIC
C0007102|T047||CCS_10|CANCERS, COLONIC
C0007102|T047||CCS_10|COLONIC CANCERS
C0007102|T047||CCS_10|MALIGNANT NEO COLON NOS
C0007102|T047||CCS_10|CANCER, COLON
C0007102|T047||CCS_10|MALIGNANT NEOPLASM OF COLON, UNSPECIFIED SITE
C0007102|T047||CCS_10|COLONIC CANCER
C0007102|T047||CCS_10|CA COLON NOS 
C0007102|T047||CCS_10|MALIGNANT NEOPLASM OF COLON NOS
C0007102|T047||CCS_10|CA COLON NOS
C0007102|T047||CCS_10|MALIGNANT NEOPLASM OF COLON (& NOS) 
C0007102|T047||CCS_10|MALIGNANT NEOPLASM OF COLON (& NOS)
C0007102|T047||CCS_10|MALIGNANT NEOPLASM OF COLON NOS 
C0007102|T047||CCS_10|-- COLON CANCER
C0007102|T047||CCS_10|COLON CANCER NOS
C0007102|T047||CCS_10|COLONIC CANCER NOS
C0007102|T047||CCS_10|CANCER OF THE COLON
C0007102|T047||CCS_10|CA - CANCER OF COLON
C0007102|T047||CCS_10|MALIGNANT TUMOUR OF COLON
C0007102|T047||CCS_10|MALIGNANT TUMOR OF COLON 
C0007102|T047||CCS_10|MALIGNANT NEOPLASM OF COLON, NOS
C0007102|T047||CCS_10|COLON NEOPLASM, MALIGNANT
C0007102|T047||CCS_10|COLON TUMOR, MALIGNANT
C0007102|T047||CCS_10|MALIGNANT COLON NEOPLASM
C0007102|T047||CCS_10|MALIGNANT COLON TUMOR
C0007102|T047||CCS_10|MALIGNANT COLONIC NEOPLASM
C0007102|T047||CCS_10|MALIGNANT COLONIC TUMOR
C0007102|T047||CCS_10|MALIGNANT NEOPLASM OF THE COLON
C0007102|T047||CCS_10|MALIGNANT TUMOR OF THE COLON
C1333990|T047||CCS_10|INCLUDING THIS BECAUSE IT READS AS PRIMARY DX OF CANCER, SUBTYPE IS DUE TO LYNCH SYNDROME
C1333990|T047||CCS_10|COLORECTAL CANCER HEREDITARY NONPOLYPOSIS
C3472669|T047||CCS_10|PRIMARY ADENOCARCINOMA OF COLON
C3472669|T047||CCS_10|PRIMARY ADENOCARCINOMA OF COLON 
C0346630|T047||CCS_10|MALIGNANT NEOPLASM OF OTHER SPECIFIED SITES OF COLON 
C0346630|T047||CCS_10|MALIGNANT NEOPLASM OF OTHER SPECIFIED SITES OF COLON
C1304819|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF COLON
C1304819|T047||CCS_10|LARGE INTESTINE NEOPLASM MALIGNANT, COLON PRIMARY
C1304819|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF COLON 
C1304819|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF COLON 
C0519037|T047||CCS_10|PRIMARY COLON LYMPHOMA
C0519037|T047||CCS_10|COLONIC LYMPHOMA
C0519037|T047||CCS_10|LYMPHOMA OF COLON 
C0519037|T047||CCS_10|LYMPHOMA OF COLON
C0519037|T047||CCS_10|COLON LYMPHOMA
C0519037|T047||CCS_10|LYMPHOMA OF THE COLON
C0346974|T047||CCS_10|METASTATIC NEOPLASM TO THE COLON
C0346974|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF COLON
C0346974|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF COLON 
C0346974|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF COLON 
C0346974|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM IN THE COLON
C0346974|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO THE COLON
C0346974|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO COLON
C0346974|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO COLON, NOS
C0346974|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF COLON, NOS
C0346974|T047||CCS_10|METASTATIC TUMOR TO THE COLON
C1282478|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT NEOPLASM OF COLON 
C1282478|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT NEOPLASM OF COLON
C1282478|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOR OF COLON 
C1282478|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOR OF COLON
C1282478|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOUR OF COLON
C1386266|T047||CCS_10|ADENOCARCINOMA; IN POLYPOSIS COLI
C1391915|T047||CCS_10|CARCINOMA; IN POLYPOSIS COLI
C1391915|T047||CCS_10|POLYPOSIS COLI; WITH CARCINOMA
C1391940|T047||CCS_10|CARCINOMA; POLIPOSIS COLI
C1391940|T047||CCS_10|POLIPOSIS COLI; CARCINOMA
C0334293|T047||CCS_10|ADENOCARCINOMA IN ADENOMATOUS POLYPOSIS COLI
C0334293|T047||CCS_10|ADENOCARCINOMA IN ADENOMATOUS POLYPOSIS COLI (MORPHOLOGIC ABNORMALITY)
C0334293|T047||CCS_10|POLYPOSIS COLI; ADENOCARCINOMA, ADENOMATOUS (IN)
C0279880|T047||CCS_10|CELLULAR DIAGNOSIS, COLON CANCER
C0279880|T047||CCS_10|COLON CANCER CELLULAR DIAGNOSIS
C0280252|T047||CCS_10|STAGE, COLON CANCER
C0280252|T047||CCS_10|COLON CANCER STAGE
C0699790|T047||CCS_10|CARCINOMA OF COLON
C0699790|T047||CCS_10|COLON CARCINOMA
C0699790|T047||CCS_10|COLON CANCER
C0699790|T047||CCS_10|CARCINOMA;COLON
C0699790|T047||CCS_10|CARCINOMA OF COLON 
C0699790|T047||CCS_10|CARCINOMA COLON
C0699790|T047||CCS_10|COLONIC CARCINOMA
C0699790|T047||CCS_10|CARCINOMA OF THE COLON
C1333098|T047||CCS_10|COLON SARCOMA
C1333098|T047||CCS_10|COLONIC SARCOMA
C1333098|T047||CCS_10|SARCOMA OF COLON
C1333098|T047||CCS_10|SARCOMA OF THE COLON
C0153441|T047||CCS_10|MALIGNANT NEOPLASM OF OTHER SPECIFIED SITES OF LARGE INTESTINE
C0153441|T047||CCS_10|MALIGNANT NEO COLON NEC
C1319315|T047||CCS_10|ADENOCARCINOMA OF LARGE INTESTINE 
C1319315|T047||CCS_10|ADENOCARCINOMA OF LARGE INTESTINE
C1319315|T047||CCS_10|COLORECTAL ADENOCARCINOMA
C1319315|T047||CCS_10|LARGE INTESTINE ADENOCARCINOMA
C1319315|T047||CCS_10|ADENOCARCINOMA OF LARGE INTESTINE 
C1319315|T047||CCS_10|ADENOCARCINOMA OF LARGE BOWEL
C1319315|T047||CCS_10|ADENOCARCINOMA OF THE LARGE BOWEL
C1319315|T047||CCS_10|ADENOCARCINOMA OF THE LARGE INTESTINE
C1319315|T047||CCS_10|LARGE BOWEL ADENOCARCINOMA
C0809966|T047|23|CCS_10|OTHER NON-EPITHELIAL CANCER OF SKIN|OTHER NON-EPITHELIAL CANCER OF SKIN
C0151779|T047||CCS_10|MALIGNANT MELANOMA OF SKIN
C0151779|T047||CCS_10|MALIGNANT MELANOMA OF SKIN, UNSPECIFIED
C0151779|T047||CCS_10|MELANOMA OF SKIN, SITE UNSPECIFIED
C0151779|T047||CCS_10|CUTANEOUS MELANOMA
C0151779|T047||CCS_10|MALIGNANT MELANOMA OF SKIN 
C0151779|T047||CCS_10|MALIG MELANOMA SKIN NOS
C0151779|T047||CCS_10|MELANOMAS OF SKIN
C0151779|T047||CCS_10|MELANOMA (MALIGNANT) NOS
C0151779|T047||CCS_10|SKIN MELANOMA
C0151779|T047||CCS_10|MELANOMA, CUTANEOUS MALIGNANT
C0151779|T047||CCS_10|DYSPLASTIC NEVUS SYNDROME, HEREDITARY
C0151779|T047||CCS_10|MELANOMA, FAMILIAL
C0151779|T047||CCS_10|FAMMM
C0151779|T047||CCS_10|FAMILIAL ATYPICAL MOLE-MALIGNANT MELANOMA SYNDROME
C0151779|T047||CCS_10|[X]MALIGNANT MELANOMA OF SKIN, UNSPECIFIED
C0151779|T047||CCS_10|MELANOMA OF SKIN
C0151779|T047||CCS_10|[X]MALIGNANT MELANOMA OF SKIN, UNSPECIFIED 
C0151779|T047||CCS_10|MALIGNANT MELANOMA OF SKIN NOS 
C0151779|T047||CCS_10|MALIGNANT MELANOMA OF SKIN NOS
C0151779|T047||CCS_10|MELANOMA OF SKIN 
C0151779|T047||CCS_10|CUTANEOUS MALIGNANT MELANOMA
C0151779|T047||CCS_10|MELANOMA, MALIGNANT
C0151779|T047||CCS_10|MALIGNANT MELANOMA OF SKIN STAGE UNSPECIFIED
C0151779|T047||CCS_10|MELANOMA SKIN
C0151779|T047||CCS_10|MELANOMA OF SKIN (MALIGNANT)
C0151779|T047||CCS_10|MM - MALIGNANT MELANOMA OF SKIN
C0151779|T047||CCS_10|MALIGNANT MELANOMA OF SKIN 
C0151779|T047||CCS_10|MELANOMA, CUTANEOUS
C0151779|T047||CCS_10|SKIN CANCER, MELANOMA
C0151779|T047||CCS_10|MELANOMA; SKIN
C0151779|T047||CCS_10|SKIN; MELANOMA
C0151779|T047||CCS_10|MALIGNANT MELANOMA OF SKIN, NOS
C0151779|T047||CCS_10|MALIGNANT CUTANEOUS MELANOMA
C0151779|T047||CCS_10|MALIGNANT MELANOMA (OF SKIN), STAGE UNSPECIFIED
C0151779|T047||CCS_10|MELANOMA OF THE SKIN
C0151779|T047||CCS_10|SKIN, MELANOMA
C0852524|T047||CCS_10|SKIN MELANOMAS (EXCL OCULAR)
C0852524|T047||CCS_10|SKIN MELANOMAS (EXCLUDING OCULAR)
C0852525|T047||CCS_10|SKIN NEOPLASMS MALIGNANT AND UNSPECIFIED (EXCL MELANOMA)
C0852525|T047||CCS_10|SKIN NEOPLASMS MALIGNANT AND UNSPECIFIED (EXCLUDING MELANOMA)
C0007114|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN, UNSPECIFIED
C0007114|T047||CCS_10|SKIN CANCERS
C0007114|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN
C0007114|T047||CCS_10|SKIN CANCER 
C0007114|T047||CCS_10|SKIN CANCER
C0007114|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN 
C0007114|T047||CCS_10|MALIGNANT SKIN NEOPLASM
C0007114|T047||CCS_10|CANCER OF SKIN
C0007114|T047||CCS_10|SKIN NEOPLASMS MALIGNANT AND UNSPECIFIED
C0007114|T047||CCS_10|CANCERS, SKIN
C0007114|T047||CCS_10|MALIGNANT TUMOR OF SKIN
C0007114|T047||CCS_10|CANCER, SKIN
C0007114|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN NOS
C0007114|T047||CCS_10|SKIN NEOPLASM, MALIGNANT
C0007114|T047||CCS_10|MALIGNANT TUMOUR OF SKIN 
C0007114|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN NOS 
C0007114|T047||CCS_10|CA - SKIN CANCER
C0007114|T047||CCS_10|MALIGNANT TUMOUR OF SKIN
C0007114|T047||CCS_10|[X]MALIGNANT NEOPLASM OF SKIN, UNSPECIFIED
C0007114|T047||CCS_10|[X]MALIGNANT NEOPLASM OF SKIN, UNSPECIFIED 
C0007114|T047||CCS_10|SKIN--CANCER
C0007114|T047||CCS_10|SKIN CANCER, NOS
C0007114|T047||CCS_10|-- SKIN CANCER
C0007114|T047||CCS_10|SKIN MALIGNANT NEOPLASM NOS
C0007114|T047||CCS_10|SKIN NEOPLASM MALIGNANT
C0007114|T047||CCS_10|MALIGNANT SKIN NEOPLASM NOS
C0007114|T047||CCS_10|SKIN NEOPLASM MALIGNANT NOS
C0007114|T047||CCS_10|CANCER OF THE SKIN
C0007114|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN 
C0007114|T047||CCS_10|SKIN CANCER, NONMELANOMATOUS (SQUAMOUS AND BASAL CELL)
C0007114|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN, NOS
C0007114|T047||CCS_10|MALIGNANT NEOPLASM OF THE SKIN
C0007114|T047||CCS_10|MALIGNANT SKIN TUMOR
C0007114|T047||CCS_10|MALIGNANT TUMOR OF THE SKIN
C0007114|T047||CCS_10|MELANOMA AND NON-MELANOMA SKIN CANCER
C0007114|T047||CCS_10|SKIN CANCER, INCLUDING MELANOMA
C0007114|T047||CCS_10|NEOPLASM MALIG;SKIN
C0007114|T047||CCS_10|MALIGNANT NEOSPLASM OF THE SKIN
C2146257|T047||CCS_10|TRICHILEMMOCARCINOMA OF SKIN 
C2146257|T047||CCS_10|TRICHILEMMOCARCINOMA OF SKIN
C0699893|T047||CCS_10|CARCINOMA OF SKIN
C0699893|T047||CCS_10|SKIN CARCINOMA
C0699893|T047||CCS_10|CARCINOMA OF SKIN 
C0699893|T047||CCS_10|CARCINOMA;SKIN
C0699893|T047||CCS_10|NONMELANOMA SKIN CANCER
C0699893|T047||CCS_10|CARCINOMA SKIN
C0699893|T047||CCS_10|SKIN CARCINOMA NOS
C0699893|T047||CCS_10|CARCINOMA OF THE SKIN
C0699893|T047||CCS_10|NON-MELANOMA CANCER OF SKIN
C0699893|T047||CCS_10|NON-MELANOMA CANCER OF THE SKIN
C0699893|T047||CCS_10|NON-MELANOMA SKIN CANCER
C0699893|T047||CCS_10|SKIN CANCER, NON-MELANOMA
C2211421|T047||CCS_10|ADENOCARCINOMA OF SKIN 
C2211421|T047||CCS_10|ADENOCARCINOMA OF SKIN
C2163816|T047||CCS_10|CYSTADENOCARCINOMA OF SKIN
C2163816|T047||CCS_10|CYSTADENOCARCINOMA OF SKIN 
C0334447|T047||CCS_10|MELANOMA ARISING FROM BLUE NEVUS
C0334447|T047||CCS_10|BLUE NEVUS-LIKE MELANOMA
C0334447|T047||CCS_10|MALIGNANT BLUE NEVUS OF SKIN 
C0334447|T047||CCS_10|MALIGNANT BLUE NEVUS OF SKIN
C0334447|T047||CCS_10|MALIGNANT BLUE NAEVUS
C0334447|T047||CCS_10|[M]BLUE NAEVUS, MALIGNANT
C0334447|T047||CCS_10|[M]BLUE NEVUS, MALIGNANT
C0334447|T047||CCS_10|MALIGNANT MELANOMA IN BLUE NEVUS
C0334447|T047||CCS_10|MALIGNANT MELANOMA IN BLUE NAEVUS
C0334447|T047||CCS_10|BLUE NAEVUS-LIKE MELANOMA
C0334447|T047||CCS_10|MALIGNANT BLUE NEVUS
C0334447|T047||CCS_10|BLUE NEVUS, MALIGNANT
C0334447|T047||CCS_10|BLUE NAEVUS, MALIGNANT
C0334447|T047||CCS_10|MALIGNANT BLUE NAEVUS OF SKIN
C0334447|T047||CCS_10|BLUE NEVUS, MALIGNANT (MORPHOLOGIC ABNORMALITY)
C0334447|T047||CCS_10|MALIGNANT BLUE NEVUS OF SKIN 
C0334447|T047||CCS_10|MALIGNANT BLUE NEVUS OF THE SKIN
C0334447|T047||CCS_10|MALIGNANT CUTANEOUS BLUE NEVUS
C0334447|T047||CCS_10|MALIGNANT SKIN BLUE NEVUS
C0856900|T047||CCS_10|SARCOMA OF SKIN 
C0856900|T047||CCS_10|SARCOMA OF SKIN
C0856900|T047||CCS_10|CUTANEOUS SARCOMA
C0856900|T047||CCS_10|SARCOMA OF THE SKIN
C0856900|T047||CCS_10|SKIN SARCOMA
C2211446|T047||CCS_10|FIBROSARCOMA OF SKIN 
C2211446|T047||CCS_10|FIBROSARCOMA OF SKIN
C2182812|T047||CCS_10|DERMATOFIBROSARCOMA OF SKIN
C2182812|T047||CCS_10|DERMATOFIBROSARCOMA OF SKIN 
C1333175|T047||CCS_10|LIPOSARCOMA OF SKIN 
C1333175|T047||CCS_10|LIPOSARCOMA OF SKIN
C1333175|T047||CCS_10|CUTANEOUS LIPOSARCOMA
C1333175|T047||CCS_10|LIPOSARCOMA OF THE SKIN
C1333175|T047||CCS_10|SKIN LIPOSARCOMA
C2211457|T047||CCS_10|MYOSARCOMA OF SKIN
C2211457|T047||CCS_10|MYOSARCOMA OF SKIN 
C1275281|T047||CCS_10|CARCINOSARCOMA OF SKIN 
C1275281|T047||CCS_10|CARCINOSARCOMA OF SKIN
C1275281|T047||CCS_10|CARCINOSARCOMA OF SKIN 
C2242810|T047||CCS_10|MALIGNANT HEMANGIOENDOTHELIOMA OF SKIN 
C2242810|T047||CCS_10|MALIGNANT HEMANGIOENDOTHELIOMA OF SKIN
C0346085|T047||CCS_10|MALIGNANT HEMANGIOPERICYTOMA OF SKIN 
C0346085|T047||CCS_10|MALIGNANT HEMANGIOPERICYTOMA OF SKIN
C0346085|T047||CCS_10|MALIGNANT SKIN HEMANGIOPERICYTOMA
C0346085|T047||CCS_10|MALIGNANT HEMANGIOPERICYTOMA OF THE SKIN
C0346085|T047||CCS_10|MALIGNANT HAEMANGIOPERICYTOMA OF SKIN
C0346085|T047||CCS_10|MALIGNANT HEMANGIOPERICYTOMA OF SKIN 
C2211463|T047||CCS_10|MALIGNANT NEURILEMOMA OF SKIN 
C2211463|T047||CCS_10|MALIGNANT NEURILEMOMA OF SKIN
C2211464|T047||CCS_10|MALIGNANT PERIPHERAL NERVE SHEATH TUMOR (MPNST) OF SKIN
C2211464|T047||CCS_10|MALIGNANT PERIPHERAL NERVE SHEATH TUMOR (MPNST) OF SKIN 
C1321781|T047||CCS_10|MALIGNANT MIXED TUMOR OF SKIN
C1321781|T047||CCS_10|MALIGNANT MIXED TUMOR OF SKIN 
C1321781|T047||CCS_10|MALIGNANT CHONDROID SYRINGOMA
C1321781|T047||CCS_10|ECCRINE MIXED TUMOR, MALIGNANT
C1321781|T047||CCS_10|ECCRINE MIXED TUMOUR, MALIGNANT
C1321781|T047||CCS_10|MALIGNANT CHONDROID SYRINGOMA (MORPHOLOGIC ABNORMALITY)
C1321781|T047||CCS_10|MALIGNANT CHONDROID SYRINGOMA OF SKIN 
C1321781|T047||CCS_10|MALIGNANT CHONDROID SYRINGOMA OF SKIN
C1321781|T047||CCS_10|MALIGNANT MIXED TUMOR OF THE SKIN
C1321781|T047||CCS_10|MALIGNANT MIXED TUMOUR OF THE SKIN
C2211466|T047||CCS_10|MALIGNANT LYMPHOMA OF SKIN 
C2211466|T047||CCS_10|MALIGNANT LYMPHOMA OF SKIN
C1707551|T047||CCS_10|CUTANEOUS MATURE B-CELL LYMPHOCYTIC NEOPLASM
C1707551|T047||CCS_10|CUTANEOUS MATURE B-CELL NEOPLASM
C0948976|T047||CCS_10|LEUKEMIA CUTIS
C0948976|T047||CCS_10|LEUKAEMIA CUTIS
C0948976|T047||CCS_10|LEUKEMIC INFILTRATION OF SKIN
C0948976|T047||CCS_10|SKIN NEOPLASM MALIGNANT SECONDARY LEUKEMIC INFILTRATION
C0948976|T047||CCS_10|LEUKEMIC INFILTRATION OF SKIN 
C0948976|T047||CCS_10|LEUKAEMIC INFILTRATION OF SKIN
C0948976|T047||CCS_10|LEUKEMIC INFILTRATION OF SKIN 
C2211422|T047||CCS_10|SCIRRHOUS ADENOCARCINOMA OF SKIN
C2211422|T047||CCS_10|SCIRRHOUS ADENOCARCINOMA OF SKIN 
C2037356|T047||CCS_10|SUPERFICIAL SPREADING ADENOCARCINOMA OF SKIN
C2037356|T047||CCS_10|SUPERFICIAL SPREADING ADENOCARCINOMA OF SKIN 
C2145030|T047||CCS_10|TRABECULAR ADENOCARCINOMA OF SKIN 
C2145030|T047||CCS_10|TRABECULAR ADENOCARCINOMA OF SKIN
C0346017|T047||CCS_10|ADENOID CYSTIC CARCINOMA OF SKIN 
C0346017|T047||CCS_10|ADENOID CYSTIC CARCINOMA OF SKIN
C0346017|T047||CCS_10|ADENOID CYSTIC ECCRINE CARCINOMA OF SKIN
C0346017|T047||CCS_10|ADENOID CYSTIC ECCRINE CARCINOMA OF SKIN 
C0346017|T047||CCS_10|SKIN NEOP MALIGNANT ADNEXA W/ ECCRINE DIFFERENTIATION ADENOID CYSTIC CARCINOMA
C0346017|T047||CCS_10|ADENOID CYSTIC ECCRINE CARCINOMA
C0346017|T047||CCS_10|PRIMARY CUTANEOUS ADENOCYSTIC CARCINOMA
C0346017|T047||CCS_10|ADENOID CYSTIC ECCRINE CARCINOMA (MORPHOLOGIC ABNORMALITY)
C0346017|T047||CCS_10|ADENOID CYSTIC ECCRINE CARCINOMA OF SKIN 
C0346017|T047||CCS_10|ADENOID CYSTIC ECCRINE CARCINOMA 
C0346017|T047||CCS_10|ADENOID CYSTIC CARCINOMA OF THE SKIN
C0346017|T047||CCS_10|ADENOID CYSTIC CUTANEOUS CARCINOMA
C0346017|T047||CCS_10|ADENOID CYSTIC SKIN CARCINOMA
C2138462|T047||CCS_10|CRIBRIFORM CARCINOMA OF SKIN
C2138462|T047||CCS_10|CRIBRIFORM CARCINOMA OF SKIN 
C2017457|T047||CCS_10|SOLID CARCINOMA OF SKIN 
C2017457|T047||CCS_10|SOLID CARCINOMA OF SKIN
C2007050|T047||CCS_10|CARCINOMA SIMPLEX OF SKIN 
C2007050|T047||CCS_10|CARCINOMA SIMPLEX OF SKIN
C2033135|T047||CCS_10|PAPILLARY ADENOCARCINOMA OF SKIN 
C2033135|T047||CCS_10|PAPILLARY ADENOCARCINOMA OF SKIN
C2189650|T047||CCS_10|VILLOUS ADENOCARCINOMA OF SKIN
C2189650|T047||CCS_10|VILLOUS ADENOCARCINOMA OF SKIN 
C2211424|T047||CCS_10|ADENOCARCINOMA IN VILLOUS ADENOMA OF SKIN 
C2211424|T047||CCS_10|ADENOCARCINOMA IN VILLOUS ADENOMA OF SKIN
C2211425|T047||CCS_10|ADENOCARCINOMA IN TUBULOVILLOUS ADENOMA OF SKIN 
C2211425|T047||CCS_10|ADENOCARCINOMA IN TUBULOVILLOUS ADENOMA OF SKIN
C2075542|T047||CCS_10|CLEAR CELL ADENOCARCINOMA OF SKIN 
C2075542|T047||CCS_10|CLEAR CELL ADENOCARCINOMA OF SKIN
C0206697|T047||CCS_10|CARCINOMA, SKIN APPENDAGE
C0206697|T047||CCS_10|APPENDAGE CARCINOMA, SKIN
C0206697|T047||CCS_10|APPENDAGE CARCINOMAS, SKIN
C0206697|T047||CCS_10|CARCINOMAS, SKIN APPENDAGE
C0206697|T047||CCS_10|SKIN APPENDAGE CARCINOMAS
C0206697|T047||CCS_10|SKIN APPENDAGE CARCINOMA
C0206697|T047||CCS_10|SKIN APPENDAGE CARCINOMA 
C0206697|T047||CCS_10|CARCINOMA, SKIN APPENDAGE [DISEASE/FINDING]
C0206697|T047||CCS_10|[M]SKIN APPENDAGE CARCINOMA
C0206697|T047||CCS_10|[M]SKIN APPENDAGE CARCINOMA (MORPHOLOGIC ABNORMALITY)
C0206697|T047||CCS_10|CARCINOMA, ADNEXAL, MALIGNANT
C0206697|T047||CCS_10|CARCINOMA OF SKIN APPENDAGE
C0206697|T047||CCS_10|CARCINOMA OF ADNEXA
C0206697|T047||CCS_10|ADNEXAL CARCINOMA
C0206697|T047||CCS_10|SKIN APPENDAGE CARCINOMA (MORPHOLOGIC ABNORMALITY)
C2211430|T047||CCS_10|SEBACEOUS ADENOCARCINOMA OF SKIN 
C2211430|T047||CCS_10|SEBACEOUS ADENOCARCINOMA OF SKIN
C2026730|T047||CCS_10|CERUMINOUS ADENOCARCINOMA OF SKIN
C2026730|T047||CCS_10|CERUMINOUS ADENOCARCINOMA OF SKIN 
C2211431|T047||CCS_10|MUCINOUS ADENOCARCINOMA OF SKIN
C2211431|T047||CCS_10|MUCINOUS ADENOCARCINOMA OF SKIN 
C2211432|T047||CCS_10|MUCIN-PRODUCING ADENOCARCINOMA OF SKIN 
C2211432|T047||CCS_10|MUCIN-PRODUCING ADENOCARCINOMA OF SKIN
C1710103|T047||CCS_10|SKIN ADENOSQUAMOUS CARCINOMA
C1710103|T047||CCS_10|ADENOSQUAMOUS CARCINOMA OF SKIN
C1710103|T047||CCS_10|ADENOSQUAMOUS CARCINOMA OF SKIN 
C2211433|T047||CCS_10|EPITHELIAL-MYOEPITHELIAL CARCINOMA OF SKIN
C2211433|T047||CCS_10|EPITHELIAL-MYOEPITHELIAL CARCINOMA OF SKIN 
C2211434|T047||CCS_10|ADENOCARCINOMA OF SKIN WITH METAPLASIA
C2211434|T047||CCS_10|ADENOCARCINOMA OF SKIN WITH METAPLASIA 
C2211434|T047||CCS_10|SKIN ADENOCARCINOMA WITH METAPLASIA
C2211436|T047||CCS_10|ADENOCARCINOMA WITH CARTILAGINOUS OR OSSEOUS METAPLASIA OF SKIN
C2211436|T047||CCS_10|SKIN ADENOCARCINOMA WITH CARTILAGINOUS OR OSSEOUS METAPLASIA
C2211436|T047||CCS_10|ADENOCARCINOMA OF SKIN WITH CARTILAGINOUS AND OSSEOUS METAPLASIA 
C2211436|T047||CCS_10|ADENOCARCINOMA OF SKIN WITH CARTILAGINOUS AND OSSEOUS METAPLASIA
C2211437|T047||CCS_10|ADENOCARCINOMA OF SKIN WITH SPINDLE CELL METAPLASIA 
C2211437|T047||CCS_10|ADENOCARCINOMA OF SKIN WITH SPINDLE CELL METAPLASIA
C2211438|T047||CCS_10|ADENOCARCINOMA OF SKIN WITH APOCRINE METAPLASIA 
C2211438|T047||CCS_10|ADENOCARCINOMA OF SKIN WITH APOCRINE METAPLASIA
C2211439|T047||CCS_10|ADENOCARCINOMA OF SKIN WITH NEUROENDOCRINE DIFFERENTIATION
C2211439|T047||CCS_10|ADENOCARCINOMA OF SKIN WITH NEUROENDOCRINE DIFFERENTIATION 
C2018514|T047||CCS_10|SPINDLE CELL SARCOMA OF SKIN
C2018514|T047||CCS_10|SPINDLE CELL SARCOMA OF SKIN 
C2011328|T047||CCS_10|GIANT CELL SARCOMA OF SKIN
C2011328|T047||CCS_10|GIANT CELL SARCOMA OF SKIN 
C2211445|T047||CCS_10|SMALL CELL SARCOMA OF SKIN
C2211445|T047||CCS_10|SMALL CELL SARCOMA OF SKIN 
C2188151|T047||CCS_10|UNDIFFERENTIATED SARCOMA OF SKIN
C2188151|T047||CCS_10|UNDIFFERENTIATED SARCOMA OF SKIN 
C2182958|T047||CCS_10|DESMOPLASTIC SMALL ROUND CELL SARCOMA OF SKIN 
C2182958|T047||CCS_10|SKIN NEOPLASM MALIGNANT SARCOMA DESMOPLASTIC SMALL ROUND CELL
C2182958|T047||CCS_10|DESMOPLASTIC SMALL ROUND CELL SARCOMA OF SKIN
C2211447|T047||CCS_10|FIBROMYXOSARCOMA OF SKIN 
C2211447|T047||CCS_10|FIBROMYXOSARCOMA OF SKIN
C2211448|T047||CCS_10|FASCIAL FIBROSARCOMA OF SKIN
C2211448|T047||CCS_10|FASCIAL FIBROSARCOMA OF SKIN 
C2211449|T047||CCS_10|INFANTILE FIBROSARCOMA OF SKIN 
C2211449|T047||CCS_10|INFANTILE FIBROSARCOMA OF SKIN
C2211450|T047||CCS_10|MALIGNANT SOLITARY FIBROUS TUMOR OF SKIN
C2211450|T047||CCS_10|MALIGNANT SOLITARY FIBROUS TUMOR OF SKIN 
C2211451|T047||CCS_10|WELL DIFFERENTIATED LIPOSARCOMA OF SKIN
C2211451|T047||CCS_10|WELL DIFFERENTIATED LIPOSARCOMA OF SKIN 
C2211452|T047||CCS_10|MYXOID LIPOSARCOMA OF SKIN
C2211452|T047||CCS_10|MYXOID LIPOSARCOMA OF SKIN 
C2211453|T047||CCS_10|ROUND CELL LIPOSARCOMA OF SKIN
C2211453|T047||CCS_10|ROUND CELL LIPOSARCOMA OF SKIN 
C2211454|T047||CCS_10|PLEOMORPHIC LIPOSARCOMA OF SKIN
C2211454|T047||CCS_10|PLEOMORPHIC LIPOSARCOMA OF SKIN 
C2211455|T047||CCS_10|MIXED TYPE LIPOSARCOMA OF SKIN 
C2211455|T047||CCS_10|MIXED TYPE LIPOSARCOMA OF SKIN
C2211456|T047||CCS_10|FIBROBLASTIC LIPOSARCOMA OF SKIN 
C2211456|T047||CCS_10|FIBROBLASTIC LIPOSARCOMA OF SKIN
C2164525|T047||CCS_10|DEDIFFERENTIATED LIPOSARCOMA OF SKIN 
C2164525|T047||CCS_10|DEDIFFERENTIATED LIPOSARCOMA OF SKIN
C2200374|T047||CCS_10|RHABDOMYOSARCOMA OF SKIN 
C2200374|T047||CCS_10|RHABDOMYOSARCOMA OF SKIN
C2006989|T047||CCS_10|CARCINOMA EX PLEOMORPHIC ADENOMA OF SKIN 
C2006989|T047||CCS_10|CARCINOMA EX PLEOMORPHIC ADENOMA OF SKIN
C2211458|T047||CCS_10|EMBRYONAL RHABDOMYOSARCOMA OF SKIN
C2211458|T047||CCS_10|EMBRYONAL RHABDOMYOSARCOMA OF SKIN 
C2018456|T047||CCS_10|SPINDLE CELL RHABDOMYOSARCOMA OF SKIN
C2018456|T047||CCS_10|SPINDLE CELL RHABDOMYOSARCOMA OF SKIN 
C2211459|T047||CCS_10|ANGIOMYOSARCOMA OF SKIN 
C2211459|T047||CCS_10|ANGIOMYOSARCOMA OF SKIN
C2211460|T047||CCS_10|EMBRYONAL CARCINOSARCOMA OF SKIN 
C2211460|T047||CCS_10|EMBRYONAL CARCINOSARCOMA OF SKIN
C2211461|T047||CCS_10|MALIGNANT MYOEPITHELIOMA OF SKIN
C2211461|T047||CCS_10|MALIGNANT MYOEPITHELIOMA OF SKIN 
C0346081|T047||CCS_10|HEMANGIOSARCOMA OF SKIN 
C0346081|T047||CCS_10|HEMANGIOSARCOMA OF SKIN
C0346081|T047||CCS_10|SKIN ANGIOSARCOMA
C0346081|T047||CCS_10|CUTANEOUS HEMANGIOSARCOMA
C0346081|T047||CCS_10|HEMANGIOSARCOMA OF SKIN 
C0346081|T047||CCS_10|MALIGNANT NEOPLASM SARCOMA ANGIOSARCOMA OF SKIN
C0346081|T047||CCS_10|ANGIOSARCOMA OF SKIN 
C0346081|T047||CCS_10|ANGIOSARCOMA OF SKIN
C0346081|T047||CCS_10|ANGIOSARCOMA OF SKIN 
C0346081|T047||CCS_10|HEMANGIOSARCOMA OF THE SKIN
C0346081|T047||CCS_10|ANGIOSARCOMA OF THE SKIN
C0346081|T047||CCS_10|SKIN HEMANGIOSARCOMA
C0030186|T047||CCS_10|EXTRA MAMMARY PAGET DISEASE
C0030186|T047||CCS_10|EXTRA MAMMARY PAGET'S DISEASE
C0030186|T047||CCS_10|EXTRA-MAMMARY PAGETS DISEASE
C0030186|T047||CCS_10|EXTRAMAMMARY PAGETS DISEASE
C0030186|T047||CCS_10|PAGET DISEASE, EXTRA MAMMARY
C0030186|T047||CCS_10|PAGET'S DISEASE, EXTRA MAMMARY
C0030186|T047||CCS_10|PAGETS DISEASE, EXTRA-MAMMARY
C0030186|T047||CCS_10|PAGETS DISEASE, EXTRAMAMMARY
C0030186|T047||CCS_10|CUTANEOUS PAGET'S DISEASE
C0030186|T047||CCS_10|PAGET'S DISEASE OF SKIN
C0030186|T047||CCS_10|PAGET'S DISEASE OF THE SKIN
C0030186|T047||CCS_10|PAGET'S SKIN DISEASE
C0030186|T047||CCS_10|PAGET DISEASE, EXTRAMAMMARY
C0030186|T047||CCS_10|PAGETS DIS EXTRA MAMMARY
C0030186|T047||CCS_10|PAGETS DIS EXTRAMAMMARY
C0030186|T047||CCS_10|EXTRAMAMMARY PAGETS DIS
C0030186|T047||CCS_10|PAGET DIS EXTRA MAMMARY
C0030186|T047||CCS_10|EXTRA MAMMARY PAGET DIS
C0030186|T047||CCS_10|EXTRAMAMMARY PAGET DIS
C0030186|T047||CCS_10|PAGET DIS EXTRAMAMMARY
C0030186|T047||CCS_10|EXTRA MAMMARY PAGETS DIS
C0030186|T047||CCS_10|EXTRAMAMMARY PAGET'S DISEASE
C0030186|T047||CCS_10|EXTRAMAMMARY PAGET DISEASE
C0030186|T047||CCS_10|EXTRAMAMMARY PAGET'S DISEASE 
C0030186|T047||CCS_10|EXTRAMAMMARY, PAGET DISEASE
C0030186|T047||CCS_10|PAGET DISEASE EXTRAMAMMARY
C0030186|T047||CCS_10|PAGET DISEASE OF SKIN
C0030186|T047||CCS_10|PAGET DISEASE, EXTRAMAMMARY (EXCEPT PAGET DISEASE OF BONE)
C0030186|T047||CCS_10|EXTRA-MAMMARY PAGET DISEASE
C0030186|T047||CCS_10|EXTRA-MAMMARY PAGET'S DISEASE
C0030186|T047||CCS_10|PAGET DISEASE, EXTRA-MAMMARY
C0030186|T047||CCS_10|PAGET'S DISEASE, EXTRA-MAMMARY
C0030186|T047||CCS_10|PAGET'S DISEASE, EXTRAMAMMARY
C0030186|T047||CCS_10|PAGET DISEASE, EXTRAMAMMARY [DISEASE/FINDING]
C0030186|T047||CCS_10|EXTRAMAMMARY PAGET'S DISEASE (MORPHOLOGIC ABNORMALITY)
C0030186|T047||CCS_10|[M]PAGET'S DISEASE, EXTRAMAMMARY, EXCLUDING PAGET'S DISEASE OF BONE
C0030186|T047||CCS_10|PAGET'S DISEASE, EXTRAMAMMARY (EXCEPT PAGET'S DISEASE OF BONE)
C0030186|T047||CCS_10|PAGET'S DISEASE OF SKIN (MORPHOLOGIC ABNORMALITY)
C0030186|T047||CCS_10|PAGET'S DISEASE, EXTRAMAMMARY (EXCEPT PAGET'S DISEASE OF BONE) (MORPHOLOGIC ABNORMALITY)
C0030186|T047||CCS_10|[M]PAGET'S DISEASE, EXTRAMAMMARY, EXCLUDING PAGET'S DISEASE OF BONE (MORPHOLOGIC ABNORMALITY)
C3251593|T047||CCS_10|SKIN NEOPLASM LOCATION MALIGNANT 
C3251593|T047||CCS_10|SKIN NEOPLASM LOCATION MALIGNANT
C3251594|T047||CCS_10|SKIN NEOPLASM LOCATION MALIGNANT BASAL CELL CARCINOMA
C3251594|T047||CCS_10|SKIN NEOPLASM LOCATION MALIGNANT BASAL CELL CARCINOMA 
C3251595|T047||CCS_10|SKIN NEOPLASM LOCATION MALIGNANT SQUAMOUS CELL CARCINOMA
C3251595|T047||CCS_10|SKIN NEOPLASM LOCATION MALIGNANT SQUAMOUS CELL CARCINOMA 
C0375068|T047||CCS_10|OTHER MALIGNANT NEOPLASM OF SKIN, SITE UNSPECIFIED
C0553723|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF SKIN
C0553723|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE SKIN
C0553723|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF SKIN 
C0553723|T047||CCS_10|SQUAMOUS CELL CARCINOMA - SKIN
C0553723|T047||CCS_10|SQUAMOUS SKIN CARCINOMA
C0553723|T047||CCS_10|SPINOUS CELL CARCINOMA
C0553723|T047||CCS_10|CUTANEOUS SQUAMOUS CELL CARCINOMA
C0553723|T047||CCS_10|SCC - CUTANEOUS SQUAMOUS CELL CARCINOMA
C0553723|T047||CCS_10|SCC - SQUAMOUS CELL CARCINOMA OF SKIN
C0553723|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF SKIN 
C0553723|T047||CCS_10|CANCER OF THE SKIN, SQUAMOUS CELL
C0553723|T047||CCS_10|CARCINOMA OF THE SKIN, SQUAMOUS CELL
C0553723|T047||CCS_10|CARCINOMA, EPIDERMOID, SKIN
C0553723|T047||CCS_10|CARCINOMA, SQUAMOUS CELL, SKIN
C0553723|T047||CCS_10|EPIDERMOID CARCINOMA OF THE SKIN
C0553723|T047||CCS_10|SKIN CANCER, EPIDERMOID CARCINOMA
C0553723|T047||CCS_10|SKIN CANCER, SQUAMOUS CELL
C0553723|T047||CCS_10|EPIDERMOID CARCINOMA OF SKIN
C0553723|T047||CCS_10|EPIDERMOID SKIN CARCINOMA
C0553723|T047||CCS_10|SKIN SQUAMOUS CELL CARCINOMA
C0553723|T047||CCS_10|SQUAMOUS CELL SKIN CARCINOMA
C0007117|T047||CCS_10|BASAL CELL CARCINOMA
C0007117|T047||CCS_10|BASAL CELL CARCINOMA OF SKIN
C0007117|T047||CCS_10|BASAL CELL CARCINOMAS
C0007117|T047||CCS_10|BASAL CELL EPITHELIOMAS
C0007117|T047||CCS_10|CARCINOMA, BASAL CELL
C0007117|T047||CCS_10|CARCINOMAS, BASAL CELL
C0007117|T047||CCS_10|EPITHELIOMAS, BASAL CELL
C0007117|T047||CCS_10|BASAL CELL EPITHELIOMA
C0007117|T047||CCS_10|RODENT ULCERS
C0007117|T047||CCS_10|ULCERS, RODENT
C0007117|T047||CCS_10|BASAL CELL CARCINOMA OF SKIN 
C0007117|T047||CCS_10|CARCINOMA, BASAL CELL [DISEASE/FINDING]
C0007117|T047||CCS_10|EPITHELIOMA, BASAL CELL
C0007117|T047||CCS_10|RODENT ULCER
C0007117|T047||CCS_10|ULCER, RODENT
C0007117|T047||CCS_10|ULCER;RODENT
C0007117|T047||CCS_10|[M]BASAL CELL CARCINOMA NOS (MORPHOLOGIC ABNORMALITY)
C0007117|T047||CCS_10|[M]BASAL CELL CARCINOMA NOS
C0007117|T047||CCS_10|EPITHELIOMA BASAL CELL
C0007117|T047||CCS_10|BASAL CELL EPITHELIOMA 
C0007117|T047||CCS_10|MALIGNANT NEOPLASM CARCINOMA EPITHELIOMA BASAL CELL
C0007117|T047||CCS_10|BASAL CELL CANCER
C0007117|T047||CCS_10|BASALIOMA
C0007117|T047||CCS_10|CANCER OF SKIN, BASAL CELL
C0007117|T047||CCS_10|CARCINOMA BASAL CELL
C0007117|T047||CCS_10|BCC - BASAL CELL CARCINOMA
C0007117|T047||CCS_10|BCC - BASAL CELL CARCINOMA OF SKIN
C0007117|T047||CCS_10|BASILOMA
C0007117|T047||CCS_10|RU - RODENT ULCER
C0007117|T047||CCS_10|EPITHELIOMA BASAL CELL 
C0007117|T047||CCS_10|BASAL CELL CARCINOMA (MORPHOLOGIC ABNORMALITY)
C0007117|T047||CCS_10|BASAL CELL CARCINOMA OF SKIN 
C0007117|T047||CCS_10|BASAL CELL CARCINOMA OF THE SKIN
C0007117|T047||CCS_10|CARCINOMA OF THE SKIN, BASAL CELL
C0007117|T047||CCS_10|CARCINOMA, BASAL CELL, SKIN
C0007117|T047||CCS_10|BASAL CELL CARCINOMA, NOS
C0007117|T047||CCS_10|BCC
C0007117|T047||CCS_10|BASAL CELL SKIN CARCINOMA
C0007117|T047||CCS_10|SKIN BASAL CELL CARCINOMA
C1261513|T047||CCS_10|SKIN NEOPLASM NOSE MALIGNANT PRIMARY
C1261513|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF SKIN OF NOSE
C1261513|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF SKIN OF NOSE 
C1261513|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF SKIN OF NOSE 
C1314758|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF SKIN 
C1314758|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF SKIN
C1314758|T047||CCS_10|SKIN NEOPLASM MALIGNANT PRIMARY
C1314758|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF SKIN 
C0348363|T047||CCS_10|MALIGNANT NEOPLASM OVERLAPPING SKIN SITE
C0348363|T047||CCS_10|OVERLAPPING LESION OF SKIN
C0348363|T047||CCS_10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF SKIN 
C0348363|T047||CCS_10|SKIN NEOPLASM MALIGNANT OVERLAPPING SITES
C0348363|T047||CCS_10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF SKIN
C0348363|T047||CCS_10|[X]MALIGNANT NEOPLASM OVERLAPPING LESION OF SKIN
C0348363|T047||CCS_10|[X]MALIGNANT NEOPLASM OVERLAPPING LESION OF SKIN 
C0153346|T047||CCS_10|MALIGNANT NEOPLASM OF COMMISSURE OF LIP
C0153346|T047||CCS_10|LIP NEOPLASM MALIGNANT LABIAL COMMISSURE
C0153346|T047||CCS_10|MAL NEO LIP, COMMISSURE
C0153346|T047||CCS_10|MALIGNANT TUMOUR OF COMMISSURE OF LIP
C0153346|T047||CCS_10|MALIGNANT TUMOR OF COMMISSURE OF LIP
C0153346|T047||CCS_10|MALIGNANT TUMOR OF LABIAL COMMISSURE
C0153346|T047||CCS_10|MALIGNANT TUMOUR OF LABIAL COMMISSURE
C0153346|T047||CCS_10|MALIGNANT NEOPLASM OF LABIAL COMMISSURE
C0153346|T047||CCS_10|MALIGNANT NEOPLASM OF COMMISSURE OF LIP 
C0153346|T047||CCS_10|MALIGNANT TUMOR OF COMMISSURE OF LIP 
C0153346|T047||CCS_10|MALIGNANT NEOPLASM OF LABIAL COMMISSURE OF LIP
C0346735|T047||CCS_10|MALIGNANT SKIN NEOPLASM OF CHEEK (EXTERNAL)
C0346735|T047||CCS_10|MALIGNANT SKIN NEOPLASM OF CHEEK (EXTERNAL) 
C0346735|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF CHEEK, EXTERNAL 
C0346735|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF CHEEK, EXTERNAL
C0346026|T047||CCS_10|BENIGN MIXED TUMOR OF THE SKIN (CHONDROID SYRINGOMA)
C0346026|T047||CCS_10|MIXED TUMOR OF THE SKIN (CHONDROID SYRINGOMA)
C0346026|T047||CCS_10|ECCRINE MIXED TUMOR OF SKIN
C0346026|T047||CCS_10|ECCRINE MIXED TUMOUR OF SKIN
C0346026|T047||CCS_10|ECCRINE MIXED TUMOR
C0346026|T047||CCS_10|ECCRINE MIXED TUMOUR
C0346026|T047||CCS_10|MIXED TUMOR OF SKIN
C0346026|T047||CCS_10|MIXED TUMOUR OF SKIN
C0346026|T047||CCS_10|ECCRINE MIXED TUMOR (MORPHOLOGIC ABNORMALITY)
C0346026|T047||CCS_10|ECCRINE MIXED TUMOR OF SKIN 
C0346026|T047||CCS_10|ECCRINE MIXED TUMOR 
C0346026|T047||CCS_10|CHONDROID SYRINGOMA
C0346026|T047||CCS_10|BENIGN MIXED TUMOR OF SKIN (CHONDROID SYRINGOMA)
C0346026|T047||CCS_10|BENIGN MIXED TUMOR OF SKIN
C0346026|T047||CCS_10|BENIGN MIXED TUMOR OF THE SKIN
C1275323|T047||CCS_10|PRIMARY CUTANEOUS PLASMACYTOMA 
C1275323|T047||CCS_10|PRIMARY CUTANEOUS PLASMACYTOMA
C1275323|T047||CCS_10|SKIN MALIGNANT LYMPHOMA NON-HODGKIN'S PRIMARY CUTANEOUS PLASMACYTOMA
C1275323|T047||CCS_10|PRIMARY CUTANEOUS PLASMACYTIC B-CELL LYMPHOMA
C1275323|T047||CCS_10|PRIMARY CUTANEOUS PLASMACYTOMA 
C1275323|T047||CCS_10|PRIMARY CUTANEOUS PLASMACYTOMA (MORPHOLOGIC ABNORMALITY)
C1275318|T047||CCS_10|ANGIOCENTRIC NATURAL KILLER/T-CELL MALIGNANT LYMPHOMA INVOLVING SKIN
C1275318|T047||CCS_10|ANGIOCENTRIC NK/T-CELL MALIGNANT LYMPHOMA INVOLVING SKIN 
C1275318|T047||CCS_10|ANGIOCENTRIC NATURAL KILLER/T-CELL MALIGNANT LYMPHOMA INVOLVING SKIN 
C1275318|T047||CCS_10|ANGIOCENTRIC NK/T-CELL MALIGNANT LYMPHOMA INVOLVING SKIN
C1275318|T047||CCS_10|SKIN MALIGNANT LYMPHOMA NON-HODGKIN'S ANGIOCENTRIC NK/T-CELL
C1275318|T047||CCS_10|ANGIOCENTRIC NK/T-CELL MALIGNANT LYMPHOMA INVOLVING SKIN 
C1275318|T047||CCS_10|ANGIOCENTRIC LYMPHOMA INVOLVING SKIN
C3489398|T047||CCS_10|NEUROEPITHELIOMA, PERIPHERAL
C3489398|T047||CCS_10|PNE
C3489398|T047||CCS_10|SKIN NEOPLASM MALIGNANT PRIMARY PERIPHERAL NEUROEPITHELIOMA
C3489398|T047||CCS_10|PERIPHERAL NEUROEPITHELIOMA
C3489398|T047||CCS_10|PERIPHERAL NEUROEPITHELIOMA 
C3489398|T047||CCS_10|PNE - PERIPHERAL NEUROEPITHELIOMA
C3489398|T047||CCS_10|PERIPHERAL NEUROEPITHELIOMA 
C0346770|T047||CCS_10|MALIGNANT SKIN TUMOUR WITH ADNEXAL DIFFERENTIATION
C0346770|T047||CCS_10|MALIGNANT SKIN TUMOR WITH ADNEXAL DIFFERENTIATION
C0346770|T047||CCS_10|MALIGNANT TUMOR OF EPIDERMAL APPENDAGE
C0346770|T047||CCS_10|MALIGNANT TUMOUR OF EPIDERMAL APPENDAGE
C0346770|T047||CCS_10|MALIGNANT SKIN TUMOR WITH ADNEXAL DIFFERENTIATION 
C0346770|T047||CCS_10|MALIGNANT TUMOR OF EPIDERMAL APPENDAGE 
C0346770|T047||CCS_10|MALIGNANT CUTANEOUS ADNEXAL NEOPLASM
C0346770|T047||CCS_10|MALIGNANT EPIDERMAL APPENDAGE NEOPLASM
C0346770|T047||CCS_10|MALIGNANT EPIDERMAL APPENDAGE TUMOR
C0346770|T047||CCS_10|MALIGNANT NEOPLASM OF EPIDERMAL APPENDAGE
C0346770|T047||CCS_10|MALIGNANT NEOPLASM OF THE EPIDERMAL APPENDAGE
C0346770|T047||CCS_10|MALIGNANT SKIN ADNEXAL NEOPLASM
C0346770|T047||CCS_10|MALIGNANT SKIN ADNEXAL TUMOR
C0346770|T047||CCS_10|MALIGNANT SKIN APPENDAGE NEOPLASM
C0346770|T047||CCS_10|MALIGNANT TUMOR OF THE EPIDERMAL APPENDAGE
C0346728|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF EXTERNAL AUDITORY MEATUS
C0346728|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF EXTERNAL AUDITORY MEATUS 
C0346079|T047||CCS_10|PROLIFERATING ANGIOENDOTHELIOMATOSIS
C0346079|T047||CCS_10|NON-HODGKIN'S LYMPHOMA OF SKIN PROLIFERATING ANGIOENDOTHELIOMATOSIS
C0346079|T047||CCS_10|PROLIFERATING ANGIOENDOTHELIOMATOSIS 
C0346079|T047||CCS_10|PROLIFERATING ANGIOENDOTHELIOMATOSIS 
C0346024|T047||CCS_10|ECCRINE DERMAL DUCT NEOPLASM
C0346024|T047||CCS_10|DERMAL DUCT TUMOR
C0346024|T047||CCS_10|ECCRINE DERMAL DUCT TUMOUR OF SKIN
C0346024|T047||CCS_10|ECCRINE DERMAL DUCT TUMOR OF SKIN
C0346024|T047||CCS_10|DERMAL DUCT TUMOR (MORPHOLOGIC ABNORMALITY)
C0346024|T047||CCS_10|DERMAL DUCT TUMOUR
C0346024|T047||CCS_10|ECCRINE DERMAL DUCT TUMOR
C0346024|T047||CCS_10|ECCRINE DERMAL DUCT TUMOUR
C0346024|T047||CCS_10|ECCRINE DERMAL DUCT TUMOR OF SKIN 
C0346024|T047||CCS_10|ECCRINE DERMAL DUCT TUMOR 
C0346024|T047||CCS_10|DERMAL DUCT NEOPLASM
C0684352|T047||CCS_10|MALIGNANT NEOPLASM OF ADNEXA OF SKIN
C0684352|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF SKIN WITH ADNEXAL DIFFERENTIATION
C0684352|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF SKIN ADNEXA
C0684352|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF SKIN ADNEXA 
C0684352|T047||CCS_10|SKIN NEOPLASM MALIGNANT ADNEXA
C0684352|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN ADNEXA 
C0684352|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN ADNEXA
C0684352|T047||CCS_10|SKIN NEOPLASM MALIGNANT ADNEXA PRIMARY
C0684352|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF ADNEXA OF SKIN
C0684352|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF SKIN WITH ADNEXAL DIFFERENTIATION 
C0684352|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF ADNEXA OF SKIN 
C1304523|T047||CCS_10|AGGRESSIVE NATURAL KILLER-CELL LEUKEMIA INVOLVING SKIN
C1304523|T047||CCS_10|AGGRESSIVE NK-CELL LEUKEMIA INVOLVING SKIN 
C1304523|T047||CCS_10|AGGRESSIVE NATURAL KILLER-CELL LEUKEMIA INVOLVING SKIN 
C1304523|T047||CCS_10|AGGRESSIVE NK-CELL LEUKEMIA INVOLVING SKIN 
C1304523|T047||CCS_10|MALIGNANT NEOPLASM LYMPHOMA AGRESSIVE NK-CELL INVOLVING SKIN
C1304523|T047||CCS_10|AGGRESSIVE NK-CELL LEUKEMIA INVOLVING SKIN
C1304523|T047||CCS_10|AGGRESSIVE NATURAL KILLER-CELL LEUKAEMIA INVOLVING SKIN
C1304523|T047||CCS_10|AGGRESSIVE NK-CELL LEUKAEMIA INVOLVING SKIN
C2314897|T047||CCS_10|SKIN SQUAMOUS CELL CARCINOMA IN SITU
C2314897|T047||CCS_10|SQUAMOUS CELL CARCINOMA IN SITU OF SKIN
C2314897|T047||CCS_10|SQUAMOUS CELL CARCINOMA IN SITU OF SKIN 
C2314897|T047||CCS_10|CANCER IN SITU SKIN, SQUAMOUS CELL
C2314897|T047||CCS_10|INTRAEPIDERMAL SQUAMOUS CELL CARCINOMA
C2314897|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF SKIN IN SITU
C2314897|T047||CCS_10|IEC - INTRAEPIDERMAL CARCINOMA OF SKIN
C2314897|T047||CCS_10|INTRAEPIDERMAL CARCINOMA OF SKIN
C2314897|T047||CCS_10|SCC - SQUAMOUS CELL CARCINOMA IN SITU OF SKIN
C2314897|T047||CCS_10|SQUAMOUS CELL CARCINOMA IN SITU OF THE SKIN
C0346734|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF TEMPLE 
C0346734|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF TEMPLE
C0346734|T047||CCS_10|SKIN NEOPLASM TEMPLE MALIGNANT
C0346734|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF TEMPLE 
C0346082|T047||CCS_10|STEWART-TREVES SYNDROME
C0346082|T047||CCS_10|POSTMASTECTOMY EXTREMITY ANGIOSARCOMA
C0346082|T047||CCS_10|ANGIOSARCOMA ASSOCIATED WITH CHRONIC LYMPHEDEMA
C0346082|T047||CCS_10|LYMPHANGIOSARCOMA FOLLOWING MASTECTOMY
C0346082|T047||CCS_10|STEWART TREVES SYNDROME
C0346082|T047||CCS_10|STEWART-TREVES SYNDROME 
C0346082|T047||CCS_10|BENIGN NEOPLASM STEWART-TREVES SYNDROME
C0346082|T047||CCS_10|POSTMASTECTOMY LYMPHANGIOSARCOMA SYNDROME
C0346082|T047||CCS_10|LYMPHANGIOSARCOMA OF STEWART AND TREVES
C0346082|T047||CCS_10|LYMPHANGIOSARCOMA OF SKIN
C0346082|T047||CCS_10|STEWART-TREVES SYNDROME 
C0346082|T047||CCS_10|LYMPHANGIOSARCOMA OF THE SKIN
C0346082|T047||CCS_10|SKIN LYMPHANGIOSARCOMA
C0346769|T047||CCS_10|MALIGNANT NEOPLASM OF OTHER SPECIFIED SKIN SITES 
C0346769|T047||CCS_10|MALIGNANT NEOPLASM OF OTHER SPECIFIED SKIN SITES
C0559018|T047||CCS_10|CA SKIN - OTHER
C0559018|T047||CCS_10|CA SKIN - OTHER NOS 
C0559018|T047||CCS_10|CA SKIN - OTHER NOS
C3665499|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF ELBOW
C3665499|T047||CCS_10|SKIN NEOPLASM ELBOW MALIGNANT
C3665499|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF ELBOW 
C3665401|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF THIGH 
C3665401|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF THIGH
C3665401|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF THIGH 
C2210570|T047||CCS_10|SKIN BIOPSY SPECIMEN MALIGNANT NEOPLASM 
C2210570|T047||CCS_10|SKIN BIOPSY SPECIMEN MALIGNANT NEOPLASM
C3665399|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF HAND
C3665399|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF HAND 
C3665399|T047||CCS_10|SKIN NEOPLASM HAND MALIGNANT
C3665399|T047||CCS_10|MALIGNANT SKIN NEOPLASM OF HAND
C3665399|T047||CCS_10|MALIGNANT SKIN NEOPLASM OF HAND 
C1282486|T047||CCS_10|SKIN NEOPLASM MALIGNANT, LOCAL RECURRENCE
C1282486|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT SKIN NEOPLASM
C1282486|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT SKIN NEOPLASM 
C1282486|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOR OF SKIN 
C1282486|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOR OF SKIN
C1282486|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOUR OF SKIN
C1304404|T047||CCS_10|MALIGNANT VASCULAR NEOPLASM OF SKIN 
C1304404|T047||CCS_10|MALIGNANT VASCULAR NEOPLASM OF SKIN
C1304404|T047||CCS_10|SKIN MALIGNANT NEOPLASM VASCULAR
C1304404|T047||CCS_10|MALIGNANT VASCULAR TUMOR OF SKIN 
C1304404|T047||CCS_10|MALIGNANT VASCULAR TUMOR OF SKIN
C1304404|T047||CCS_10|MALIGNANT VASCULAR TUMOUR OF SKIN
C1304404|T047||CCS_10|MALIGNANT CUTANEOUS VASCULAR NEOPLASM
C1304404|T047||CCS_10|MALIGNANT CUTANEOUS VASCULAR TUMOR
C1304404|T047||CCS_10|MALIGNANT SKIN VASCULAR NEOPLASM
C1304404|T047||CCS_10|MALIGNANT SKIN VASCULAR TUMOR
C1282490|T047||CCS_10|METASTASIS FROM MALIGNANT NEOPLASM OF SKIN 
C1282490|T047||CCS_10|METASTASIS FROM MALIGNANT NEOPLASM OF SKIN
C1282490|T047||CCS_10|SKIN NEOPLASM MALIGNANT METASTASIS
C1282490|T047||CCS_10|METASTASIS FROM MALIGNANT TUMOR OF SKIN 
C1282490|T047||CCS_10|METASTASIS FROM MALIGNANT TUMOR OF SKIN
C1282490|T047||CCS_10|METASTASIS FROM MALIGNANT TUMOUR OF SKIN
C0346031|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN WITH APOCRINE DIFFERENTIATION
C0346031|T047||CCS_10|SKIN NEOPLASM MALIGNANT WITH APOCRINE DIFFERENTIATION
C0346031|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN WITH APOCRINE DIFFERENTIATION 
C0346031|T047||CCS_10|MALIGNANT SKIN TUMOR WITH APOCRINE DIFFERENTIATION
C0346031|T047||CCS_10|MALIGNANT SKIN TUMOUR WITH APOCRINE DIFFERENTIATION
C0346031|T047||CCS_10|MALIGNANT SKIN TUMOR WITH APOCRINE DIFFERENTIATION 
C1304452|T047||CCS_10|MALIGNANT FIBROHISTIOCYTIC NEOPLASM OF SKIN
C1304452|T047||CCS_10|MALIGNANT FIBROHISTIOCYTIC NEOPLASM OF SKIN 
C1304452|T047||CCS_10|SKIN NEOPLASM MALIGNANT FIBROHISTIOCYTIC
C1304452|T047||CCS_10|MALIGNANT FIBROHISTIOCYTIC TUMOR OF SKIN 
C1304452|T047||CCS_10|MALIGNANT FIBROHISTIOCYTIC TUMOR OF SKIN
C1304452|T047||CCS_10|MALIGNANT FIBROHISTIOCYTIC TUMOUR OF SKIN
C0346811|T047||CCS_10|SKIN NEOPLASM MALIGNANT DERMIS
C0346811|T047||CCS_10|MALIGNANT NEOPLASM OF DERMIS
C0346811|T047||CCS_10|MALIGNANT NEOPLASM OF DERMIS 
C0346811|T047||CCS_10|MALIGNANT TUMOR OF DERMIS
C0346811|T047||CCS_10|MALIGNANT TUMOUR OF DERMIS
C0346811|T047||CCS_10|MALIGNANT TUMOR OF DERMIS 
C0346811|T047||CCS_10|MALIGNANT DERMAL NEOPLASM
C0346811|T047||CCS_10|MALIGNANT DERMIS NEOPLASM
C0346811|T047||CCS_10|MALIGNANT DERMIS TUMOR
C0346811|T047||CCS_10|MALIGNANT NEOPLASM OF THE DERMIS
C0346811|T047||CCS_10|MALIGNANT TUMOR OF THE DERMIS
C1275031|T047||CCS_10|PUVA THERAPY-ASSOCIATED SKIN MALIGNANCY 
C1275031|T047||CCS_10|PSORALEN AND LONG-WAVE ULTRAVIOLET RADIATION (PUVA) THERAPY-ASSOCIATED SKIN MALIGNANCY
C1275031|T047||CCS_10|PSORALEN AND LONG-WAVE ULTRAVIOLET RADIATION (PUVA) THERAPY-ASSOCIATED SKIN MALIGNANCY 
C1275031|T047||CCS_10|PSORALEN AND LONG-WAVE ULTRAVIOLET RADIATION THERAPY-ASSOCIATED SKIN MALIGNANCY 
C1275031|T047||CCS_10|PSORALEN AND LONG-WAVE ULTRAVIOLET RADIATION THERAPY-ASSOCIATED SKIN MALIGNANCY
C1275031|T047||CCS_10|PSORALEN AND LONG-WAVE ULTRAVIOLET RADIATION THERAPY-ASSOCIATED SKIN MALIGNANCY 
C1275031|T047||CCS_10|SKIN NEOPLASM MALIGNANT PSORALEN/LONG-WAVE ULTRAVIOLET RADIATION THERAPY ASSOC
C1275031|T047||CCS_10|PUVA THERAPY-ASSOCIATED SKIN MALIGNANCY
C1275046|T047||CCS_10|RADIATION-INDUCED SKIN MALIGNANCY
C1275046|T047||CCS_10|SKIN NEOPLASM MALIGNANT RADIATION-INDUCED
C1275046|T047||CCS_10|RADIATION-INDUCED SKIN MALIGNANCY 
C1275046|T047||CCS_10|RADIATION-INDUCED SKIN MALIGNANCY 
C1275056|T047||CCS_10|ARSENIC-INDUCED MALIGNANCY
C1275056|T047||CCS_10|SKIN NEOPLASM MALIGNANT ARSENIC-INDUCED
C1275056|T047||CCS_10|ARSENIC-INDUCED MALIGNANCY 
C1275056|T047||CCS_10|ARSENIC-INDUCED SKIN MALIGNANCY 
C1275056|T047||CCS_10|ARSENIC-INDUCED SKIN MALIGNANCY
C1998037|T047||CCS_10|MALIGNANT BASAL CELL TUMOR OF SKIN
C1998037|T047||CCS_10|MALIGNANT BASAL CELL NEOPLASM OF SKIN
C1998037|T047||CCS_10|MALIGNANT BASAL CELL TUMOUR OF SKIN
C1998037|T047||CCS_10|MALIGNANT BASAL CELL NEOPLASM OF SKIN 
C1998037|T047||CCS_10|MALIGNANT BASAL CELL NEOPLASM OF SKIN 
C1998037|T047||CCS_10|SKIN MALIGNANT NEOPLASM BASAL CELL
C0153687|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SKIN
C0153687|T047||CCS_10|METASTATIC NEOPLASM TO THE SKIN
C0153687|T047||CCS_10|METASTASIS OF MALIGNANT NEOPLASM TO SKIN 
C0153687|T047||CCS_10|METASTASIS TO THE SKIN
C0153687|T047||CCS_10|METASTASIS OF MALIGNANT NEOPLASM TO SKIN
C0153687|T047||CCS_10|METASTASES TO SKIN
C0153687|T047||CCS_10|SECONDARY MALIG NEO SKIN
C0153687|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SKIN 
C0153687|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM SKIN
C0153687|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SKIN NOS 
C0153687|T047||CCS_10|METASTASIS TO SKIN 
C0153687|T047||CCS_10|SKIN CANCER METASTATIC
C0153687|T047||CCS_10|METASTASIS TO SKIN
C0153687|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SKIN NOS
C0153687|T047||CCS_10|METASTASES TO SKIN, NOS
C0153687|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO THE SKIN
C0153687|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM IN THE SKIN
C0153687|T047||CCS_10|CANCER METASTATIC TO SKIN
C0153687|T047||CCS_10|SKIN METASTASES
C0153687|T047||CCS_10|CUTANEOUS METASTASIS
C0153687|T047||CCS_10|DERMAL METASTASIS
C0153687|T047||CCS_10|MALIGNANT INFILTRATION OF SKIN
C0153687|T047||CCS_10|SKIN SECONDARIES
C0153687|T047||CCS_10|SECONDARY CANCER OF SKIN
C0153687|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO SKIN
C0153687|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SKIN 
C0153687|T047||CCS_10|CANCER, METASTATIC TO SKIN
C0153687|T047||CCS_10|METASTATIC CANCER TO SKIN
C0153687|T047||CCS_10|SKIN, METASTATIC CANCER TO
C0153687|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO SKIN, NOS
C0153687|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SKIN, NOS
C0153687|T047||CCS_10|METASTATIC TUMOR TO THE SKIN
C0153687|T047||CCS_10|SKIN METASTASIS
C0349513|T047||CCS_10|SKIN NEOPLASM MALIGNANT WITH PILAR DIFFERENTIATION 
C0349513|T047||CCS_10|SKIN NEOPLASM MALIGNANT WITH PILAR DIFFERENTIATION
C0349513|T047||CCS_10|MALIGNANT TUMOR OF SKIN WITH PILAR DIFFERENTIATION
C0349513|T047||CCS_10|MALIGNANT TUMOUR OF SKIN WITH PILAR DIFFERENTIATION
C0349513|T047||CCS_10|MALIGNANT TUMOR OF SKIN WITH PILAR DIFFERENTIATION 
C0547064|T047||CCS_10|MALIGNANT SKIN TUMOR WITH ECCRINE DIFFERENTIATION
C0547064|T047||CCS_10|MALIGNANT SKIN NEOPLASM WITH ECCRINE DIFFERENTIATION
C0547064|T047||CCS_10|SKIN NEOPLASM MALIGNANT ADNEXA WITH ECCRINE DIFFERENTIATION
C0547064|T047||CCS_10|MALIGNANT SKIN NEOPLASM WITH ECCRINE DIFFERENTIATION 
C0547064|T047||CCS_10|MALIGNANT SKIN TUMOUR WITH ECCRINE DIFFERENTIATION
C0547064|T047||CCS_10|MALIGNANT SWEAT GLAND TUMOR
C0547064|T047||CCS_10|MALIGNANT SWEAT GLAND TUMOUR
C0547064|T047||CCS_10|MALIGNANT SKIN TUMOR WITH ECCRINE DIFFERENTIATION 
C0496797|T047||CCS_10|SKIN OF TRUNK
C0496797|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF TRUNK
C0496797|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF TRUNK 
C0496797|T047||CCS_10|SKIN NEOPLASM TRUNK MALIGNANT
C0496797|T047||CCS_10|CA SKIN - TRUNK 
C0496797|T047||CCS_10|CA SKIN - TRUNK
C0496797|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF TRUNK 
C0496797|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF TRUNK, NOS
C0345977|T047||CCS_10|MALIGNANT TUMOR OF SURFACE EPITHELIUM
C0345977|T047||CCS_10|MALIGNANT TUMOUR OF SURFACE EPITHELIUM
C0345977|T047||CCS_10|MALIGNANT EPITHELIAL NEOPLASM OF SKIN 
C0345977|T047||CCS_10|MALIGNANT EPITHELIAL NEOPLASM OF SKIN
C0345977|T047||CCS_10|MALIGNANT TUMOR OF SURFACE EPITHELIUM 
C1269827|T047||CCS_10|MALIGNANT SKIN NEOPLASM OF HEAD AND NECK 
C1269827|T047||CCS_10|MALIGNANT SKIN NEOPLASM OF HEAD AND NECK
C1269827|T047||CCS_10|SKIN NEOPLASM HEAD AND NECK MALIGNANT
C1269827|T047||CCS_10|CA SKIN - HEAD/NECK
C1269827|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN HEAD AND NECK 
C1269827|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN HEAD AND NECK
C0559017|T047||CCS_10|SKIN NEOPLASM LOWER EXTREMITIES MALIGNANT
C0559017|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF LOWER EXTREMITIES 
C0559017|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF LOWER EXTREMITIES
C0559017|T047||CCS_10|CA SKIN - LOWER LIMB 
C0559017|T047||CCS_10|CA SKIN - LOWER LIMB
C0559017|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF LOWER LIMB 
C0559017|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF LOWER LIMB
C0684431|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF UPPER LIMB
C0684431|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF ARM
C0684431|T047||CCS_10|SKIN NEOPLASM UPPER EXTREMITIES MALIGNANT
C0684431|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF UPPER EXTREMITIES 
C0684431|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF UPPER EXTREMITIES
C0684431|T047||CCS_10|CA SKIN - UPPER LIMB
C0684431|T047||CCS_10|CA SKIN - UPPER LIMB 
C0684431|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF UPPER LIMB 
C0684431|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF UPPER LIMB, NOS
C1274311|T047||CCS_10|HODGKIN DISEASE AFFECTING SKIN
C1274311|T047||CCS_10|HODGKIN'S DISEASE AFFECTING SKIN 
C1274311|T047||CCS_10|HODGKIN'S DISEASE AFFECTING SKIN
C1274311|T047||CCS_10|HODGKIN'S DISEASE AFFECTING SKIN 
C1275320|T047||CCS_10|SMALL B-CELL LYMPHOCYTIC LYMPHOMA OF SKIN 
C1275320|T047||CCS_10|SMALL B-CELL LYMPHOCYTIC LYMPHOMA OF SKIN
C1275320|T047||CCS_10|SMALL LYMPHOCYTIC B-CELL LYMPHOMA INVOLVING SKIN 
C1275320|T047||CCS_10|SMALL LYMPHOCYTIC B-CELL LYMPHOMA INVOLVING SKIN
C0334346|T047||CCS_10|APOCRINE ADENOCARCINOMA
C0334346|T047||CCS_10|APOCRINE ADENOCARCINOMA 
C0334346|T047||CCS_10|APOCRINE ADENOCARCINOMA (MORPHOLOGIC ABNORMALITY)
C0334346|T047||CCS_10|ADENOCARCINOMA; APOCRINE, UNSPECIFIED SITE
C0334346|T047||CCS_10|APOCRINE; ADENOCARCINOMA, UNSPECIFIED SITE
C1388303|T047||CCS_10|CARCINOMA; APOCRINE, UNSPECIFIED SITE
C1388303|T047||CCS_10|APOCRINE; CARCINOMA, UNSPECIFIED SITE
C1395263|T047||CCS_10|DERMATOFIBROSARCOMA; (SITE OF SKIN NOT SPECIFIED)
C0392784|T047||CCS_10|DERMATOFIBROSARCOMA PROTUBERANS
C0392784|T047||CCS_10|DERMATOFIBROSARCOMA PROTUBERANS 
C0392784|T047||CCS_10|DERMATOFIBROSARCOMA
C0392784|T047||CCS_10|DERMATOFIBROSARCOMA PROTUBERANS 
C0392784|T047||CCS_10|SOFT TISSUE MALIGNANT NEOPLASM DERMATOFIBROSARCOMA PROTUBERANS
C0392784|T047||CCS_10|[M]DERMATOFIBROMA PROTUBERANS
C0392784|T047||CCS_10|DFSP - DERMATOFIBROSARCOMA PROTRUBERANS
C0392784|T047||CCS_10|DERMATOFIBROSARCOMA (MORPHOLOGIC ABNORMALITY)
C0392784|T047||CCS_10|DERMATOFIBROSARCOMA; PROTUBERANS
C0392784|T047||CCS_10|PROTUBERANS; DERMATOFIBROSARCOMA
C0392784|T047||CCS_10|DERMATOFIBROSARCOMA PROTUBERANS, NOS
C0392784|T047||CCS_10|DFSP
C0280247|T047||CCS_10|STAGE/CELL TYPE, SKIN CANCER
C0280247|T047||CCS_10|SKIN CANCER STAGE
C1302772|T047||CCS_10|PRIMARY CUTANEOUS LYMPHOMA
C1302772|T047||CCS_10|SKIN MALIGNANT LYMPHOMA PRIMARY CUTANEOUS
C1302772|T047||CCS_10|PRIMARY CUTANEOUS LYMPHOMA 
C1302772|T047||CCS_10|PRIMARY CUTANEOUS LYMPHOMA 
C1302772|T047||CCS_10|CUTANEOUS LYMPHOMA
C1302772|T047||CCS_10|SKIN LYMPHOMA
C1302772|T047||CCS_10|PRIMARY CUTANEOUS LYMPHOMA (MORPHOLOGIC ABNORMALITY)
C0153604|T047||CCS_10|MALIGNANT NEOPLASM OF SCROTUM
C0153604|T047||CCS_10|MALIGNANT NEOPLASM OF SCROTUM 
C0153604|T047||CCS_10|SCROTAL CANCER
C0153604|T047||CCS_10|MALIGNANT TUMOR OF SCROTUM
C0153604|T047||CCS_10|MALIGN NEOPL SCROTUM
C0153604|T047||CCS_10|MALIGNANT TUMOUR OF SCROTUM
C0153604|T047||CCS_10|MALIGNANT TUMOUR OF SCROTUM 
C0153604|T047||CCS_10|CA - CANCER OF SCROTUM
C0153604|T047||CCS_10|CANCER OF SCROTUM
C0153604|T047||CCS_10|SCROTAL CA
C0153604|T047||CCS_10|MALIGNANT SCROTAL TUMOR
C0153604|T047||CCS_10|MALIGNANT SCROTAL TUMOUR
C0153604|T047||CCS_10|MALIGNANT TUMOR OF SCROTUM 
C0153604|T047||CCS_10|MALIGNANT NEOPLASM OF THE SCROTUM
C0153604|T047||CCS_10|MALIGNANT SCROTAL NEOPLASM
C0153604|T047||CCS_10|MALIGNANT TUMOR OF THE SCROTUM
C1707590|T047||CCS_10|CUTANEOUS PRECURSOR LYMPHOBLASTIC LYMPHOMA/LEUKEMIA
C1707590|T047||CCS_10|CUTANEOUS PRECURSOR LYMPHOID NEOPLASM
C1301363|T047||CCS_10|BLASTIC NK-CELL LYMPHOMA
C1301363|T047||CCS_10|EARLY PLASMACYTOID DENDRITIC CELL LEUKEMIA/LYMPHOMA
C1301363|T047||CCS_10|PRIMARY CUTANEOUS CD4+/CD56+ HEMATOLYMPHOID NEOPLASM
C1301363|T047||CCS_10|BLASTIC NATURAL KILLER LEUKEMIA/LYMPHOMA
C1301363|T047||CCS_10|CD4+/CD56+ HEMATODERMIC NEOPLASM
C1301363|T047||CCS_10|AGRANULAR CD4+ CD56+ HEMATODERMIC NEOPLASM/TUMOR
C1301363|T047||CCS_10|BLASTIC PLASMACYTOID DENDRITIC CELL NEOPLASM
C1301363|T047||CCS_10|AGRANULAR CD4+ NATURAL KILLER CELL LEUKEMIA
C1301363|T047||CCS_10|BLASTIC PLASMACYTOID DENDRITIC CELL NEOPLASM (MORPHOLOGIC ABNORMALITY)
C1301363|T047||CCS_10|BLASTIC PLASMACYTOID DENDRITIC CELL NEOPLASM 
C1301363|T047||CCS_10|MALIGNANT NEOPLASM LYMPHOMA NK-CELL BLASTIC
C1301363|T047||CCS_10|BLASTIC NK-CELL LYMPHOMA 
C1301363|T047||CCS_10|BLASTIC NK-CELL LYMPHOMA (MORPHOLOGIC ABNORMALITY)
C1301363|T047||CCS_10|NEOPLASM OF HEMATOPOIETIC CELL TYPE BLASTIC PLASMACYTOID DENDRITIC CELL
C1301363|T047||CCS_10|BLASTIC PLASMACYTOID DENDRITIC CELL NEOPLASM 
C1301363|T047||CCS_10|MONOMORPHIC NK-CELL LYMPHOMA
C2211472|T047||CCS_10|NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF SKIN 
C2211472|T047||CCS_10|NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF SKIN
C2211475|T047||CCS_10|GRADE 2 NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF SKIN
C2211475|T047||CCS_10|GRADE 2 NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF SKIN 
C2046521|T047||CCS_10|SKIN MALIGNANT LYMPHOMA HODGKIN'S AND NON-HODGKIN'S
C2046521|T047||CCS_10|COMPOSITE HODGKIN'S AND NON-HODGKIN'S LYMPHOMA OF SKIN
C2046521|T047||CCS_10|COMPOSITE HODGKIN'S AND NON-HODGKIN'S LYMPHOMA OF SKIN 
C2211476|T047||CCS_10|LYMPHOPLASMACYTIC LYMPHOMA OF SKIN 
C2211476|T047||CCS_10|LYMPHOPLASMACYTIC LYMPHOMA OF SKIN
C2211477|T047||CCS_10|MANTLE CELL LYMPHOMA OF SKIN
C2211477|T047||CCS_10|MANTLE CELL LYMPHOMA OF SKIN 
C2211483|T047||CCS_10|GRADE 2 FOLLICULAR LYMPHOMA OF SKIN 
C2211483|T047||CCS_10|GRADE 2 FOLLICULAR LYMPHOMA OF SKIN
C2211486|T047||CCS_10|ANGIOIMMUNOBLASTIC T-CELL LYMPHOMA OF SKIN 
C2211486|T047||CCS_10|ANGIOIMMUNOBLASTIC T-CELL LYMPHOMA OF SKIN
C2211486|T047||CCS_10|ANGIOIMMUNOBLASTIC LYMPHADENOPATHY WITH DYSPROTEINEMIA (AILD) OF SKIN
C2211471|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION, DIFFUSE FIBROSIS OF SKIN 
C2211471|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION, DIFFUSE FIBROSIS OF SKIN
C2211474|T047||CCS_10|GRADE 1 NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF SKIN 
C2211474|T047||CCS_10|GRADE 1 NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF SKIN
C2211479|T047||CCS_10|IMMUNOBLASTIC LARGE B-CELL DIFFUSE LYMPHOMA OF SKIN 
C2211479|T047||CCS_10|IMMUNOBLASTIC LARGE B-CELL DIFFUSE LYMPHOMA OF SKIN
C2211484|T047||CCS_10|GRADE 3 FOLLICULAR LYMPHOMA OF SKIN
C2211484|T047||CCS_10|GRADE 3 FOLLICULAR LYMPHOMA OF SKIN 
C2046594|T047||CCS_10|HODGKIN'S GRANULOMA OF SKIN
C2046594|T047||CCS_10|HODGKIN'S GRANULOMA OF SKIN 
C1367653|T047||CCS_10|PRIMARY CUTANEOUS MARGINAL ZONE B CELL LYMPHOMA OF MUCOSA-ASSOCIATED LYMPHOID TISSUE
C1367653|T047||CCS_10|MARGINAL ZONE B-CELL LYMPHOMA OF SKIN 
C1367653|T047||CCS_10|MARGINAL ZONE B-CELL LYMPHOMA OF SKIN
C1367653|T047||CCS_10|PRIMARY CUTANEOUS MARGINAL ZONE LYMPHOMA OF MUCOSA-ASSOCIATED LYMPHOID TISSUE
C1367653|T047||CCS_10|PRIMARY CUTANEOUS MARGINAL ZONE B-CELL LYMPHOMA OF MUCOSA-ASSOCIATED LYMPHOID TISSUE
C1367653|T047||CCS_10|SALT LYMPHOMA
C1367653|T047||CCS_10|SKIN-ASSOCIATED LYMPHOID TISSUE LYMPHOMA
C1367653|T047||CCS_10|CUTANEOUS IMMUNOCYTOMA
C1367653|T047||CCS_10|MARGINAL ZONE B CELL LYMPHOMA OF SKIN
C1367653|T047||CCS_10|MARGINAL ZONE B CELL LYMPHOMA OF THE SKIN
C1367653|T047||CCS_10|C-MALT
C2211488|T047||CCS_10|SUBCUTANEOUS PANNICULITIS-LIKE T-CELL LYMPHOMA OF SKIN 
C2211488|T047||CCS_10|SUBCUTANEOUS PANNICULITIS-LIKE T-CELL LYMPHOMA OF SKIN
C2211469|T047||CCS_10|MIXED CELLULARITY HODGKIN'S LYMPHOMA OF SKIN
C2211469|T047||CCS_10|MIXED CELLULARITY HODGKIN'S LYMPHOMA OF SKIN 
C2211473|T047||CCS_10|NODULAR SCLEROSING HODGKIN'S LYMPHOMA IN CELLULAR PHASE OF SKIN
C2211473|T047||CCS_10|NODULAR SCLEROSING HODGKIN'S LYMPHOMA IN CELLULAR PHASE OF SKIN 
C2211485|T047||CCS_10|MATURE T-CELL LYMPHOMA OF SKIN 
C2211485|T047||CCS_10|MATURE T-CELL LYMPHOMA OF SKIN
C2211470|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION OF SKIN
C2211470|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION OF SKIN 
C2046734|T047||CCS_10|HODGKIN'S SARCOMA OF SKIN
C2046734|T047||CCS_10|HODGKIN'S SARCOMA OF SKIN 
C2211482|T047||CCS_10|GRADE 1 FOLLICULAR LYMPHOMA OF SKIN 
C2211482|T047||CCS_10|GRADE 1 FOLLICULAR LYMPHOMA OF SKIN
C2211468|T047||CCS_10|LYMPHOCYTE-RICH HODGKIN'S LYMPHOMA OF SKIN 
C2211468|T047||CCS_10|LYMPHOCYTE-RICH HODGKIN'S LYMPHOMA OF SKIN
C2211478|T047||CCS_10|LARGE B-CELL DIFFUSE LYMPHOMA OF SKIN 
C2211478|T047||CCS_10|LARGE B-CELL DIFFUSE LYMPHOMA OF SKIN
C0238461|T047||CCS_10|ANAPLASTIC THYROID CARCINOMA
C0238461|T047||CCS_10|THYROID GLAND CARCINOSARCOMA
C0238461|T047||CCS_10|THYROID GLAND UNDIFFERENTIATED (ANAPLASTIC) CARCINOMA
C0238461|T047||CCS_10|UNDIFFERENTIATED (ANAPLASTIC) THYROID GLAND CARCINOMA
C0238461|T047||CCS_10|DEDIFFERENTIATED THYROID GLAND CARCINOMA
C0238461|T047||CCS_10|METAPLASTIC THYROID GLAND CARCINOMA
C0238461|T047||CCS_10|PLEOMORPHIC THYROID GLAND CARCINOMA
C0238461|T047||CCS_10|SARCOMATOID THYROID GLAND CARCINOMA
C0238461|T047||CCS_10|CARCINOSARCOMA OF THYROID GLAND
C0238461|T047||CCS_10|CARCINOSARCOMA OF THYROID GLAND 
C0238461|T047||CCS_10|ANAPLASTIC THYROID CANCER
C0238461|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF THYROID GLAND
C0238461|T047||CCS_10|ANAPLASTIC CARCINOMA OF THYROID GLAND
C0238461|T047||CCS_10|ANAPLASTIC THYROID CARCINOMA 
C0238461|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF THE THYROID GLAND
C0238461|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF THE THYROID GLAND 
C0238461|T047||CCS_10|ANAPLASTIC THYROID CARCINOMAS
C0238461|T047||CCS_10|CANCERS, ANAPLASTIC THYROID
C0238461|T047||CCS_10|THYROID CANCERS, ANAPLASTIC
C0238461|T047||CCS_10|THYROID CARCINOMA, ANAPLASTIC
C0238461|T047||CCS_10|CARCINOMA, ANAPLASTIC THYROID
C0238461|T047||CCS_10|ANAPLASTIC THYROID CANCERS
C0238461|T047||CCS_10|THYROID CARCINOMAS, ANAPLASTIC
C0238461|T047||CCS_10|CANCER, ANAPLASTIC THYROID
C0238461|T047||CCS_10|CARCINOMAS, ANAPLASTIC THYROID
C0238461|T047||CCS_10|THYROID CARCINOMA, ANAPLASTIC [DISEASE/FINDING]
C0238461|T047||CCS_10|THYROID CANCER, ANAPLASTIC
C0238461|T047||CCS_10|ANAPLASTIC THYROID CARCINOMA 
C0238461|T047||CCS_10|ANAPLASTIC CARCINOMA OF THE THYROID
C0238461|T047||CCS_10|THYROID CANCER, ANAPLASTIC CARCINOMA
C0238461|T047||CCS_10|THYROID CANCER, UNDIFFERENTIATED CARCINOMA
C0238461|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF THE THYROID
C0238461|T047||CCS_10|UNDIFFERENTIATED THYROID CANCER
C0238461|T047||CCS_10|ANAPLASTIC CARCINOMA OF THYROID
C0238461|T047||CCS_10|ANAPLASTIC CARCINOMA OF THE THYROID GLAND
C0238461|T047||CCS_10|ANAPLASTIC THYROID GLAND CARCINOMA
C0238461|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF THYROID
C0238461|T047||CCS_10|UNDIFFERENTIATED THYROID CARCINOMA
C0238461|T047||CCS_10|UNDIFFERENTIATED THYROID GLAND CARCINOMA
C0206682|T047||CCS_10|ADENOCARCINOMA, FOLLICULAR
C0206682|T047||CCS_10|ADENOCARCINOMAS, FOLLICULAR
C0206682|T047||CCS_10|FOLLICULAR ADENOCARCINOMAS
C0206682|T047||CCS_10|FOLLICULAR ADENOCARCINOMA
C0206682|T047||CCS_10|FOLLICULAR THYROID CARCINOMA
C0206682|T047||CCS_10|THYROID GLAND FOLLICULAR CARCINOMA
C0206682|T047||CCS_10|FOLLICULAR THYROID GLAND CARCINOMA
C0206682|T047||CCS_10|THYROID CARCINOMA, FOLLICULAR
C0206682|T047||CCS_10|FTC
C0206682|T047||CCS_10|FOLLICULAR ADENOCARCINOMA OF THYROID GLAND
C0206682|T047||CCS_10|FOLLICULAR ADENOCARCINOMA OF THYROID GLAND 
C0206682|T047||CCS_10|FOLLICULAR THYROID CANCER
C0206682|T047||CCS_10|ADENOCARCINOMA, FOLLICULAR [DISEASE/FINDING]
C0206682|T047||CCS_10|CARCINOMA, FOLLICULAR THYROID
C0206682|T047||CCS_10|CARCINOMAS, FOLLICULAR THYROID
C0206682|T047||CCS_10|FOLLICULAR THYROID CARCINOMAS
C0206682|T047||CCS_10|THYROID CARCINOMAS, FOLLICULAR
C0206682|T047||CCS_10|[M]FOLLICULAR ADENOCARCINOMA NOS (MORPHOLOGIC ABNORMALITY)
C0206682|T047||CCS_10|[M]FOLLICULAR ADENOCARCINOMA NOS
C0206682|T047||CCS_10|[M]FOLLICULAR CARCINOMA
C0206682|T047||CCS_10|CARCINOMA, FOLLICULAR CELL, MALIGNANT
C0206682|T047||CCS_10|FOLLICULAR THYROID CARCINOMA 
C0206682|T047||CCS_10|THYROID MALIGNANT CARCINOMA FOLLICUALR
C0206682|T047||CCS_10|FOLLICULAR CARCINOMA OF THYROID GLAND
C0206682|T047||CCS_10|FOLLICULAR CANCER OF THYROID
C0206682|T047||CCS_10|FOLLICULAR CARCINOMA OF THE THYROID GLAND
C0206682|T047||CCS_10|FOLLICULAR CARCINOMA
C0206682|T047||CCS_10|FOLLICULAR CARCINOMA OF THE THYROID
C0206682|T047||CCS_10|WELL-DIFFERENTIATED FOLLICULAR ADENOCARCINOMA
C0206682|T047||CCS_10|WELL-DIFFERENTIATED FOLLICULAR CARCINOMA
C0206682|T047||CCS_10|FOLLICULAR CARCINOMA OF THYROID
C0206682|T047||CCS_10|FOLLICULAR CANCER OF THE THYROID
C0206682|T047||CCS_10|THYROID FOLLICULAR CARCINOMA
C0206682|T047||CCS_10|FOLLICULAR CANCER OF THYROID GLAND
C0206682|T047||CCS_10|FOLLICULAR CANCER OF THE THYROID GLAND
C0206682|T047||CCS_10|FOLLICULAR ADENOCARCINOMA - WELL DIFFERENTIATED
C0206682|T047||CCS_10|FOLLICULAR ADENOCARCINOMA, WELL DIFFERENTIATED
C0206682|T047||CCS_10|FOLLICULAR CARCINOMA - WELL DIFFERENTIATED
C0206682|T047||CCS_10|FOLLICULAR CARCINOMA, WELL DIFFERENTIATED
C0206682|T047||CCS_10|FTC - FOLLICULAR THYROID CARCINOMA
C0206682|T047||CCS_10|FOLLICULAR ADENOCARCINOMA (MORPHOLOGIC ABNORMALITY)
C0206682|T047||CCS_10|FOLLICULAR ADENOCARCINOMA, WELL DIFFERENTIATED (MORPHOLOGIC ABNORMALITY)
C0206682|T047||CCS_10|FOLLICULAR THYROID CARCINOMA 
C0206682|T047||CCS_10|THYROID CANCER, FOLLICULAR
C0206682|T047||CCS_10|CARCINOMA; FOLLICULAR, PURE
C0206682|T047||CCS_10|CARCINOMA; FOLLICULAR, WELL DIFFERENTIATED
C0206682|T047||CCS_10|FOLLICULAR; ADENOCARCINOMA, WELL DIFFERENTIATED
C0206682|T047||CCS_10|FOLLICULAR; CARCINOMA, WELL DIFFERENTIATED
C0206682|T047||CCS_10|ADENOCARCINOMA; FOLLICULAR, WELL DIFFERENTIATED
C0206682|T047||CCS_10|FOLLICULAR ADENOCARCINOMA, NOS
C0206682|T047||CCS_10|FOLLICULAR CARCINOMA, NOS
C0238462|T047||CCS_10|MEDULLARY THYROID CARCINOMA
C0238462|T047||CCS_10|THYROID GLAND MEDULLARY CARCINOMA
C0238462|T047||CCS_10|THYROID GLAND NEUROENDOCRINE CARCINOMA
C0238462|T047||CCS_10|MEDULLARY THYROID GLAND CARCINOMA
C0238462|T047||CCS_10|MEDULLARY CARCINOMA
C0238462|T047||CCS_10|MTC
C0238462|T047||CCS_10|MEDULLARY THYROID CANCER
C0238462|T047||CCS_10|THYROID CANCER, MEDULLARY
C0238462|T047||CCS_10|THYROID CARCINOMA, MEDULLARY
C0238462|T047||CCS_10|MEDULLARY THYROID CANCER (MTC)
C0238462|T047||CCS_10|CARCINOMA, C-CELL, MALIGNANT
C0238462|T047||CCS_10|SOLID CARCINOMA OF THE THYROID GLAND
C0238462|T047||CCS_10|SOLID CARCINOMA OF THYROID GLAND
C0238462|T047||CCS_10|MEDULLARY THYROID CARCINOMA 
C0238462|T047||CCS_10|SOLID CARCINOMA OF THE THYROID GLAND 
C0238462|T047||CCS_10|MEDULLARY CARCINOMA OF THYROID GLAND
C0238462|T047||CCS_10|MEDULLARY CARCINOMA OF THE THYROID
C0238462|T047||CCS_10|C CELL CARCINOMA
C0238462|T047||CCS_10|MEDULLARY CARCINOMA OF THYROID
C0238462|T047||CCS_10|MEDULLARY CARCINOMA OF THE THYROID GLAND
C0238462|T047||CCS_10|THYROID MEDULLARY CARCINOMA
C0238462|T047||CCS_10|PARAFOLLICULAR CELL CARCINOMA
C0238462|T047||CCS_10|ULTIMOBRANCHIAL THYROID TUMOR
C0238462|T047||CCS_10|ULTIMOBRANCHIAL THYROID TUMOUR
C0238462|T047||CCS_10|MTC - MEDULLARY THYROID CARCINOMA
C0238462|T047||CCS_10|MEDULLARY THYROID CARCINOMA 
C0238463|T047||CCS_10|PAPILLARY THYROID CARCINOMA
C0238463|T047||CCS_10|THYROID GLAND PAPILLARY CARCINOMA
C0238463|T047||CCS_10|PAPILLARY THYROID GLAND CARCINOMA
C0238463|T047||CCS_10|THYROID CARCINOMA, PAPILLARY
C0238463|T047||CCS_10|TPC
C0238463|T047||CCS_10|THYROID PAPILLARY CARCINOMA
C0238463|T047||CCS_10|PAPILLARY CARCINOMA OF THYROID
C0238463|T047||CCS_10|PAPILLARY THYROID CANCER
C0238463|T047||CCS_10|THYROID CANCER, PAPILLARY
C0238463|T047||CCS_10|PAPILLARY CARCINOMA OF THE THYROID GLAND 
C0238463|T047||CCS_10|PAPILLARY CARCINOMA OF THE THYROID GLAND
C0238463|T047||CCS_10|PAPILLARY CARCINOMA OF THYROID GLAND
C0238463|T047||CCS_10|CARCINOMA PAPILLARY THYROID
C0238463|T047||CCS_10|PTC - PAPILLARY THYROID CARCINOMA
C0238463|T047||CCS_10|PAPILLARY THYROID CARCINOMA 
C0238463|T047||CCS_10|PAPILLARY CANCER OF THYROID GLAND
C0238463|T047||CCS_10|PAPILLARY CANCER OF THYROID
C0238463|T047||CCS_10|PAPILLARY CANCER OF THE THYROID GLAND
C0238463|T047||CCS_10|PAPILLARY CANCER OF THE THYROID
C0238463|T047||CCS_10|PAPILLARY CARCINOMA OF THE THYROID
C1096666|T047||CCS_10|THYROID CANCER METASTATIC
C2116054|T047||CCS_10|CARCINOMA SIMPLEX OF THE THYROID GLAND 
C2116054|T047||CCS_10|CARCINOMA SIMPLEX OF THYROID GLAND
C2116054|T047||CCS_10|CARCINOMA SIMPLEX OF THE THYROID GLAND
C2213252|T047||CCS_10|MALIGNANT SMALL CELL NEOPLASM OF THYROID GLAND
C2213252|T047||CCS_10|MALIGNANT SMALL CELL NEOPLASM OF THYROID GLAND 
C2011415|T047||CCS_10|GIANT CELL TYPE NEOPLASM OF THYROID GLAND
C2011415|T047||CCS_10|GIANT CELL TYPE NEOPLASM OF THYROID GLAND 
C2018696|T047||CCS_10|SPINDLE CELL TYPE NEOPLASM OF THYROID GLAND 
C2018696|T047||CCS_10|SPINDLE CELL TYPE NEOPLASM OF THYROID GLAND
C2075656|T047||CCS_10|CLEAR CELL TYPE NEOPLASM OF THYROID GLAND 
C2075656|T047||CCS_10|CLEAR CELL TYPE NEOPLASM OF THYROID GLAND
C0549473|T047||CCS_10|THYROID CARCINOMA
C0549473|T047||CCS_10|THYROID GLAND CARCINOMA
C0549473|T047||CCS_10|THYROID CANCER
C0549473|T047||CCS_10|THYROID CANCER 
C0549473|T047||CCS_10|CANCERS, THYROID
C0549473|T047||CCS_10|THYROID CANCERS
C0549473|T047||CCS_10|THYROID GLAND CANCER
C0549473|T047||CCS_10|CARCINOMA;THYROID GLAND
C0549473|T047||CCS_10|CANCER, THYROID
C0549473|T047||CCS_10|THYROID GLAND--CANCER
C0549473|T047||CCS_10|THYROID CANCER, NOS
C0549473|T047||CCS_10|CARCINOMA OF THYROID GLAND
C0549473|T047||CCS_10|THYROID CARCINOMA 
C0549473|T047||CCS_10|THYROID CARCINOMAS
C0549473|T047||CCS_10|CARCINOMAS, THYROID
C0549473|T047||CCS_10|CARCINOMA THYROID
C0549473|T047||CCS_10|THYROID CARCINOMA NOS
C0549473|T047||CCS_10|CANCER OF THYROID
C0549473|T047||CCS_10|CANCER OF THE THYROID
C0549473|T047||CCS_10|HEAD AND NECK CANCER, THYROID
C0549473|T047||CCS_10|CARCINOMA OF THYROID
C0549473|T047||CCS_10|CARCINOMA OF THE THYROID GLAND
C0549473|T047||CCS_10|CARCINOMA OF THE THYROID
C0549473|T047||CCS_10|CARCINOMA, THYROID
C1704228|T047||CCS_10|THYROID ADENOCARCINOMA
C1704228|T047||CCS_10|THYROID GLAND ADENOCARCINOMA
C1704228|T047||CCS_10|ADENOCARCINOMA OF THYROID GLAND 
C1704228|T047||CCS_10|ADENOCARCINOMA OF THYROID GLAND
C1704228|T047||CCS_10|ADENOCARCINOMA OF THYROID
C1704228|T047||CCS_10|THYROID ADENOCARCINOMA 
C1704228|T047||CCS_10|ADENOCARCINOMA THYROID
C2213264|T047||CCS_10|MALIGNANT FIBROUS HISTIOCYTOMA OF THYROID GLAND
C2213264|T047||CCS_10|MALIGNANT FIBROUS HISTIOCYTOMA OF THYROID GLAND 
C1336756|T047||CCS_10|THYROID GLAND SARCOMA
C1336756|T047||CCS_10|THYROID SARCOMA
C1336756|T047||CCS_10|SARCOMA OF THYROID GLAND 
C1336756|T047||CCS_10|SARCOMA OF THYROID GLAND
C1336756|T047||CCS_10|SARCOMA OF THYROID
C1336756|T047||CCS_10|SARCOMA OF THE THYROID GLAND
C1336756|T047||CCS_10|SARCOMA OF THE THYROID
C0349668|T047||CCS_10|MALIGNANT LYMPHOMA OF THYROID GLAND 
C0349668|T047||CCS_10|MALIGNANT LYMPHOMA OF THYROID GLAND
C0349668|T047||CCS_10|MALIGNANT LYMPHOMA OF THYROID GLAND 
C2213268|T047||CCS_10|MALIGNANT PLASMACYTOMA OF THYROID GLAND 
C2213268|T047||CCS_10|MALIGNANT PLASMACYTOMA OF THYROID GLAND
C2213270|T047||CCS_10|MALIGNANT MASTOCYTOSIS OF THYROID GLAND 
C2213270|T047||CCS_10|MALIGNANT MASTOCYTOSIS OF THYROID GLAND
C2217675|T047||CCS_10|MALIGNANT NEOPLASM OF THYROID GLAND STAGING
C2217675|T047||CCS_10|MALIGNANT NEOPLASM OF THYROID GLAND STAGING 
C2217675|T047||CCS_10|MALIGNANT THYROID NEOPLASM STAGING
C2217675|T047||CCS_10|MALIGNANT TUMOR OF THYROID GLAND STAGING
C2217675|T047||CCS_10|THYROID CANCER STAGING
C0347023|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO THE THYROID
C0347023|T047||CCS_10|METASTASIS TO THYROID
C0347023|T047||CCS_10|METASTASIS TO THYROID 
C0347023|T047||CCS_10|METASTASES TO THYROID
C0347023|T047||CCS_10|THYROID MALIGNANT NEOPLASM SECONDARY
C0347023|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF THYROID GLAND
C0347023|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF THYROID GLAND 
C0347023|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM IN THE THYROID GLAND
C0347023|T047||CCS_10|CANCER METASTATIC TO THYROID
C0347023|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO THYROID GLAND
C0347023|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF THYROID GLAND 
C0347023|T047||CCS_10|METASTASIS TO THE THYROID GLAND
C0347023|T047||CCS_10|METASTASIS TO THE THYROID
C0347023|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO THE THYROID GLAND
C0347023|T047||CCS_10|METASTATIC MALIGNANT TUMOR TO THE THYROID GLAND
C0347023|T047||CCS_10|METASTATIC MALIGNANT TUMOR TO THE THYROID
C0347023|T047||CCS_10|METASTATIC NEOPLASM TO THE THYROID GLAND
C0347023|T047||CCS_10|METASTATIC NEOPLASM TO THE THYROID
C0347023|T047||CCS_10|METASTATIC TUMOR TO THE THYROID GLAND
C0347023|T047||CCS_10|METASTATIC TUMOR TO THE THYROID
C0347023|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM TO THE THYROID GLAND
C0347023|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM TO THE THYROID
C0347023|T047||CCS_10|SECONDARY MALIGNANT TUMOR TO THE THYROID GLAND
C0347023|T047||CCS_10|SECONDARY MALIGNANT TUMOR TO THE THYROID
C2062941|T047||CCS_10|DIFFERENTIATED MALIGNANT NEOPLASM OF THYROID RECURRENCE AFTER ABLATION
C2062941|T047||CCS_10|DIFFERENTIATED MALIGNANT NEOPLASM OF THYROID RECURRENCE AFTER ABLATION 
C2062941|T047||CCS_10|MALIGNANT THYROID NEOPLASM RECURRENCE AFTER ABLATION (DIFFERENTIATED)
C2938921|T047||CCS_10|THYROID CANCER STAGE 0
C2082467|T047||CCS_10|PLEOMORPHIC CARCINOMA OF THYROID GLAND
C2082467|T047||CCS_10|PLEOMORPHIC CARCINOMA OF THE THYROID GLAND
C2082467|T047||CCS_10|PLEOMORPHIC CARCINOMA OF THE THYROID GLAND 
C2011267|T047||CCS_10|GIANT CELL CARCINOMA OF THYROID GLAND
C2011267|T047||CCS_10|GIANT CELL CARCINOMA OF THE THYROID GLAND 
C2011267|T047||CCS_10|GIANT CELL CARCINOMA OF THE THYROID GLAND
C2142937|T047||CCS_10|PSEUDOSARCOMATOUS CARCINOMA OF THE THYROID GLAND 
C2142937|T047||CCS_10|PSEUDOSARCOMATOUS CARCINOMA OF THE THYROID GLAND
C2142937|T047||CCS_10|PSEUDOSARCOMATOUS CARCINOMA OF THYROID GLAND
C2111819|T047||CCS_10|POLYGONAL CELL CARCINOMA OF THYROID GLAND
C2111819|T047||CCS_10|POLYGONAL CELL CARCINOMA OF THE THYROID GLAND 
C2111819|T047||CCS_10|POLYGONAL CELL CARCINOMA OF THE THYROID GLAND
C2116055|T047||CCS_10|THYROID CARCINOMA WITH OSTEOCLAST-LIKE GIANT CELLS
C2116055|T047||CCS_10|CARCINOMA OF THE THYROID GLAND WITH OSTEOCLAST-LIKE GIANT CELLS 
C2116055|T047||CCS_10|CARCINOMA OF THE THYROID GLAND WITH OSTEOCLAST-LIKE GIANT CELLS
C2116055|T047||CCS_10|CARCINOMA OF THYROID GLAND WITH OSTEOCLAST-LIKE GIANT CELLS
C2213254|T047||CCS_10|SMALL CELL CARCINOMA OF THE THYROID GLAND 
C2213254|T047||CCS_10|SMALL CELL CARCINOMA OF THE THYROID GLAND
C2213254|T047||CCS_10|SMALL CELL CARCINOMA OF THYROID GLAND
C2009891|T047||CCS_10|SMALL CELL FUSIFORM CELL CARCINOMA OF THE THYROID GLAND
C2009891|T047||CCS_10|FUSIFORM TYPE SMALL CELL CARCINOMA OF THYROID GLAND
C2009891|T047||CCS_10|SMALL CELL FUSIFORM CELL CARCINOMA OF THE THYROID GLAND 
C2146668|T047||CCS_10|ACINAR CELL CARCINOMA OF THYROID
C2146668|T047||CCS_10|ACINAR CELL CARCINOMA OF THE THYROID GLAND
C2146668|T047||CCS_10|ACINAR CELL CARCINOMA OF THE THYROID GLAND 
C2146668|T047||CCS_10|ACINAR CELL CARCINOMA OF THYROID GLAND
C1710177|T047||CCS_10|THYROID GLAND SQUAMOUS CELL CARCINOMA
C1710177|T047||CCS_10|SQUAMOUS CELL THYROID GLAND CARCINOMA
C1710177|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THYROID GLAND
C1710177|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE THYROID GLAND 
C1710177|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE THYROID GLAND
C2109326|T047||CCS_10|KERATINIZING SQUAMOUS CELL CARCINOMA OF THYROID GLAND
C2109326|T047||CCS_10|KERATINIZING SQUAMOUS CELL CARCINOMA OF THE THYROID GLAND 
C2109326|T047||CCS_10|KERATINIZING SQUAMOUS CELL CARCINOMA OF THE THYROID GLAND
C2213255|T047||CCS_10|LARGE CELL, NONKERATINIZING SQUAMOUS CELL CARCINOMA OF THE THYROID GLAND
C2213255|T047||CCS_10|NONKERATINIZING LARGE CELL SQUAMOUS CARCINOMA CELL OF THYROID GLAND
C2213255|T047||CCS_10|LARGE CELL, NONKERATINIZING SQUAMOUS CELL CARCINOMA OF THE THYROID GLAND 
C2213256|T047||CCS_10|SMALL CELL, NONKERATINIZING SQUAMOUS CELL CARCINOMA OF THE THYROID GLAND 
C2213256|T047||CCS_10|NONKERATINIZING SMALL CELL SQUAMOUS CELL CARCINOMA OF THYROID GLAND
C2213256|T047||CCS_10|SMALL CELL, NONKERATINIZING SQUAMOUS CELL CARCINOMA OF THE THYROID GLAND
C2018573|T047||CCS_10|SPINDLE CELL SQUAMOUS CELL CARCINOMA OF THE THYROID GLAND
C2018573|T047||CCS_10|SPINDLE CELL SQUAMOUS CELL CARCINOMA OF THE THYROID GLAND 
C2018573|T047||CCS_10|SPINDLE CELL SQUAMOUS CELL CARCINOMA OF THYROID GLAND
C2213257|T047||CCS_10|ADENOID SQUAMOUS CELL CARCINOMA OF THYROID GLAND
C2213257|T047||CCS_10|ADENOID SQUAMOUS CELL CARCINOMA OF THE THYROID GLAND 
C2213257|T047||CCS_10|ADENOID SQUAMOUS CELL CARCINOMA OF THE THYROID GLAND
C2213258|T047||CCS_10|MICROINVASIVE SQUAMOUS CELL CARCINOMA OF THE THYROID GLAND 
C2213258|T047||CCS_10|MICROINVASIVE SQUAMOUS CELL CARCINOMA OF THYROID GLAND
C2213258|T047||CCS_10|MICROINVASIVE SQUAMOUS CELL CARCINOMA OF THE THYROID GLAND
C2019459|T047||CCS_10|SQUAMOUS CELL CARCINOMA WITH HORN FORMATION OF THYROID
C2019459|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE THYROID GLAND WITH HORN FORMATION 
C2019459|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE THYROID GLAND WITH HORN FORMATION
C2019459|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THYROID GLAND WITH HORN FORMATION
C1883338|T047||CCS_10|THYROID GLAND FOLLICULAR CARCINOMA, MINIMALLY INVASIVE
C1883338|T047||CCS_10|MINIMALLY INVASIVE FOLLICULAR CARCINOMA OF THYROID GLAND
C1883338|T047||CCS_10|MINIMALLY INVASIVE FOLLICULAR CARCINOMA OF THE THYROID GLAND
C1883338|T047||CCS_10|MINIMALLY INVASIVE FOLLICULAR CARCINOMA OF THE THYROID GLAND 
C2116051|T047||CCS_10|INSULAR CARCINOMA OF THE THYROID GLAND 
C2116051|T047||CCS_10|INSULAR CARCINOMA OF THYROID GLAND
C2116051|T047||CCS_10|INSULAR CARCINOMA OF THE THYROID GLAND
C0334379|T047||CCS_10|MEDULLARY CARCINOMA WITH AMYLOID STROMA
C0334379|T047||CCS_10|THYROID GLAND MEDULLARY CARCINOMA WITH AMYLOID STROMA
C0334379|T047||CCS_10|MEDULLARY THYROID GLAND CARCINOMA WITH AMYLOID STROMA
C0334379|T047||CCS_10|MEDULLARY CARCINOMA WITH AMYLOID STROMA -RETIRED-
C0334379|T047||CCS_10|MEDULLARY CARCINOMA WITH AMYLOID STROMA (MORPHOLOGIC ABNORMALITY)
C0334379|T047||CCS_10|MEDULLARY THYROID CARCINOMA WITH AMYLOID STROMA
C0334379|T047||CCS_10|MEDULLARY THYROID CARCINOMA WITH AMYLOID STROMA 
C0334379|T047||CCS_10|MEDULLARY CARCINOMA OF THYROID WITH AMYLOID STROMA
C0334379|T047||CCS_10|MEDULLARY CARCINOMA OF THYROID GLAND WITH AMYLOID STROMA
C0334379|T047||CCS_10|CARCINOMA; MEDULLARY WITH AMYLOID STROMA, UNSPECIFIED SITE
C0334379|T047||CCS_10|MEDULLARY; CARCINOMA WITH AMYLOID STROMA, UNSPECIFIED SITE
C0334379|T047||CCS_10|MEDULLARY ADENOCARCINOMA WITH AMYLOID STROMA
C0334379|T047||CCS_10|PARAFOLLICULAR CELL ADENOCARCINOMA WITH AMYLOID STROMA
C0334379|T047||CCS_10|PARAFOLLICULAR CELL CARCINOMA WITH AMYLOID STROMA
C0334379|T047||CCS_10|C CELL ADENOCARCINOMA WITH AMYLOID STROMA
C0334379|T047||CCS_10|C CELL CARCINOMA WITH AMYLOID STROMA
C2116052|T047||CCS_10|MIXED MEDULLARY-FOLLICULAR CARCINOMA OF THYROID GLAND
C2116052|T047||CCS_10|MIXED MEDULLARY-FOLLICULAR THYROID CARCINOMA
C2116052|T047||CCS_10|MIXED MEDULLARY-FOLLICULAR THYROID CARCINOMA 
C1710414|T047||CCS_10|THYROID GLAND MIXED MEDULLARY AND FOLLICULAR CELL CARCINOMA
C1710414|T047||CCS_10|THYROID GLAND MIXED MEDULLARY AND PAPILLARY CARCINOMA
C1710414|T047||CCS_10|MIXED MEDULLARY-PAPILLARY THYROID CARCINOMA
C1710414|T047||CCS_10|MIXED MEDULLARY-PAPILLARY CARCINOMA OF THYROID GLAND
C1710414|T047||CCS_10|MIXED MEDULLARY-PAPILLARY THYROID CARCINOMA 
C2116053|T047||CCS_10|NONENCAPSULATED SCLEROSING CARCINOMA OF THE THYROID GLAND
C2116053|T047||CCS_10|NONENCAPSULATED SCLEROSING CARCINOMA OF THYROID GLAND
C2116053|T047||CCS_10|NONENCAPSULATED SCLEROSING CARCINOMA OF THE THYROID GLAND 
C2033139|T047||CCS_10|PAPILLARY ADENOCARCINOMA OF THYROID GLAND
C2033139|T047||CCS_10|PAPILLARY ADENOCARCINOMA OF THYROID GLAND 
C2116009|T047||CCS_10|ADENOCARCINOMA IN VILLOUS ADENOMA OF THYROID GLAND 
C2116009|T047||CCS_10|ADENOCARCINOMA IN VILLOUS ADENOMA OF THYROID GLAND
C2116008|T047||CCS_10|ADENOCARCINOMA IN TUBULOVILLOUS ADENOMA OF THYROID GLAND 
C2116008|T047||CCS_10|ADENOCARCINOMA IN TUBULOVILLOUS ADENOMA OF THYROID GLAND
C2163817|T047||CCS_10|CYSTADENOCARCINOMA OF THYROID GLAND
C2163817|T047||CCS_10|CYSTADENOCARCINOMA OF THE THYROID GLAND
C2163817|T047||CCS_10|CYSTADENOCARCINOMA OF THE THYROID GLAND 
C2033251|T047||CCS_10|PAPILLARY CYSTADENOCARCINOMA OF THE THYROID GLAND
C2033251|T047||CCS_10|PAPILLARY CYSTADENOCARCINOMA OF THYROID GLAND
C2033251|T047||CCS_10|PAPILLARY CYSTADENOCARCINOMA OF THE THYROID GLAND 
C2146680|T047||CCS_10|ACINAR CELL CYSTADENOCARCINOMA OF THYROID
C2146680|T047||CCS_10|ACINAR CELL CYSTADENOCARCINOMA OF THYROID GLAND
C2146680|T047||CCS_10|ACINAR CELL CYSTADENOCARCINOMA OF THE THYROID GLAND
C2146680|T047||CCS_10|ACINAR CELL CYSTADENOCARCINOMA OF THE THYROID GLAND 
C3714651|T047||CCS_10|FOLLICULAR VARIANT PAPILLARY CARCINOMA
C3714651|T047||CCS_10|FOLLICULAR VARIANT PAPILLARY THYROID GLAND CARCINOMA
C3714651|T047||CCS_10|FOLLICULAR VARIANT THYROID GLAND PAPILLARY CARCINOMA
C3714651|T047||CCS_10|FOLLICULAR VARIANT PAPILLARY CARCINOMA OF THE THYROID GLAND
C3714651|T047||CCS_10|FOLLICULAR VARIANT PAPILLARY CARCINOMA OF THYROID GLAND
C3714651|T047||CCS_10|FOLLICULAR VARIANT PAPILLARY CARCINOMA OF THE THYROID GLAND 
C3714651|T047||CCS_10|FOLLICULAR VARIANT PAPILLARY ADENOCARCINOMA
C3714651|T047||CCS_10|PAPILLARY CARCINOMA FOLLICULAR VARIANT
C1709457|T047||CCS_10|THYROID GLAND PAPILLARY MICROCARCINOMA
C1709457|T047||CCS_10|PAPILLARY MICROCARCINOMA OF THE THYROID GLAND
C1709457|T047||CCS_10|PAPILLARY MICROCARCINOMA OF THE THYROID
C1709457|T047||CCS_10|PAPILLARY THYROID GLAND MICROCARCINOMA
C1709457|T047||CCS_10|PAPILLARY THYROID MICROCARCINOMA
C1709457|T047||CCS_10|PAPILLARY MICROCARCINOMA OF THYROID GLAND
C1709457|T047||CCS_10|PAPILLARY MICROCARCINOMA OF THE THYROID GLAND 
C2016175|T047||CCS_10|PAPILLARY OXYPHILIC CELL CARCINOMA OF THE THYROID GLAND
C2016175|T047||CCS_10|PAPILLARY OXYPHILIC CELL CARCINOMA OF THYROID GLAND
C2016175|T047||CCS_10|PAPILLARY OXYPHILIC CELL CARCINOMA OF THE THYROID GLAND 
C1880498|T047||CCS_10|ENCAPSULATED THYROID GLAND PAPILLARY CARCINOMA
C1880498|T047||CCS_10|ENCAPSULATED PAPILLARY CARCINOMA OF THE THYROID GLAND
C1880498|T047||CCS_10|ENCAPSULATED PAPILLARY CARCINOMA OF THYROID GLAND
C1880498|T047||CCS_10|ENCAPSULATED PAPILLARY CARCINOMA OF THE THYROID GLAND 
C2106521|T047||CCS_10|PAPILLARY COLUMNAR CELL CARCINOMA OF THE THYROID GLAND
C2106521|T047||CCS_10|COLUMNAR CELL PAPILLARY CARCINOMA OF THYROID GLAND
C2106521|T047||CCS_10|PAPILLARY COLUMNAR CELL CARCINOMA OF THE THYROID GLAND 
C2033239|T047||CCS_10|THYROID MALIGNANT CARCINOMA PAPILLARY METASTATIC TO REGIONAL LYMPH NODE
C2033239|T047||CCS_10|PAPILLARY CARCINOMA OF THYROID METASTATIC TO REGIONAL LYMPH NODE
C2033239|T047||CCS_10|PAPILLARY THYROID CARCINOMA WITH METASTASIS TO REGIONAL LYMPH NODES 
C2033239|T047||CCS_10|PAPILLARY THYROID CARCINOMA WITH METASTASIS TO REGIONAL LYMPH NODES
C2033240|T047||CCS_10|THYROID MALIGNANT CARCINOMA PAPILLARY METASTATIC TO SUPRACLAVICULAR LYMPH NODE
C2033240|T047||CCS_10|PAPILLARY THYROID CARCINOMA WITH METASTASIS TO SUPRACLAVICULAR LYMPH NODES
C2033240|T047||CCS_10|PAPILLARY THYROID CARCINOMA WITH METASTASIS TO SUPRACLAVICULAR LYMPH NODES 
C2033240|T047||CCS_10|PAPILLARY CARCINOMA OF THYROID METASTATIC TO SUPRACLAVICULAR LYMPH NODE
C2217676|T047||CCS_10|MALIGNANT NEOPLASM OF THYROID STAGE I
C2217676|T047||CCS_10|MALIGNANT NEOPLASM OF THYROID STAGE I 
C2217676|T047||CCS_10|MALIGNANT TUMOR OF THYROID STAGE I
C2217676|T047||CCS_10|THYROID CANCER STAGE I
C2217677|T047||CCS_10|MALIGNANT NEOPLASM OF THYROID STAGE II
C2217677|T047||CCS_10|MALIGNANT NEOPLASM OF THYROID STAGE II 
C2217677|T047||CCS_10|THYROID CANCER STAGE II
C2217677|T047||CCS_10|MALIGNANT TUMOR OF THYROID STAGE II
C2217678|T047||CCS_10|MALIGNANT NEOPLASM OF THYROID STAGE III
C2217678|T047||CCS_10|MALIGNANT NEOPLASM OF THYROID STAGE III 
C2217678|T047||CCS_10|THYROID CANCER STAGE III
C2217678|T047||CCS_10|MALIGNANT TUMOR OF THYROID STAGE III
C3160834|T047||CCS_10|THYROID CANCER STAGE IV
C2213253|T047||CCS_10|MALIGNANT EPITHELIOMA OF THE THYROID GLAND
C2213253|T047||CCS_10|MALIGNANT EPITHELIOMA OF THYROID GLAND
C2213253|T047||CCS_10|MALIGNANT EPITHELIOMA OF THE THYROID GLAND 
C2111684|T047||CCS_10|LARGE CELL CARCINOMA OF THE THYROID GLAND 
C2111684|T047||CCS_10|LARGE CELL CARCINOMA OF THYROID GLAND
C2111684|T047||CCS_10|LARGE CELL CARCINOMA OF THE THYROID GLAND
C2111754|T047||CCS_10|LARGE CELL NEUROENDOCRINE CARCINOMA OF THYROID GLAND
C2111754|T047||CCS_10|LARGE CELL NEUROENDOCRINE CARCINOMA OF THE THYROID GLAND 
C2111754|T047||CCS_10|LARGE CELL NEUROENDOCRINE CARCINOMA OF THE THYROID GLAND
C2111685|T047||CCS_10|THYROID MALIGNANT CARCINOMA LARGE CELL WITH RHABDOID PHENOTYPE
C2111685|T047||CCS_10|LARGE CELL CARCINOMA OF THE THYROID GLAND WITH RHABDOID PHENOTYPE
C2111685|T047||CCS_10|LARGE CELL CARCINOMA OF THE THYROID GLAND WITH RHABDOID PHENOTYPE 
C2111685|T047||CCS_10|LARGE CELL CARCINOMA OF THYROID GLAND WITH RHABDOID PHENOTYPE
C2012119|T047||CCS_10|GLASSY CELL CARCINOMA OF THYROID GLAND
C2012119|T047||CCS_10|GLASSY CELL CARCINOMA OF THE THYROID GLAND 
C2012119|T047||CCS_10|GLASSY CELL CARCINOMA OF THE THYROID GLAND
C2018407|T047||CCS_10|SPINDLE CELL CARCINOMA OF THYROID GLAND
C2018407|T047||CCS_10|SPINDLE CELL CARCINOMA OF THE THYROID GLAND 
C2018407|T047||CCS_10|SPINDLE CELL CARCINOMA OF THE THYROID GLAND
C2011232|T047||CCS_10|GIANT CELL AND SPINDLE CELL CARCINOMA OF THE THYROID GLAND
C2011232|T047||CCS_10|GIANT CELL AND SPINDLE CELL CARCINOMA OF THE THYROID GLAND 
C2011232|T047||CCS_10|GIANT CELL AND SPINDLE CELL CARCINOMA OF THYROID GLAND
C2213259|T047||CCS_10|SCIRRHOUS ADENOCARCINOMA OF THYROID GLAND 
C2213259|T047||CCS_10|SCIRRHOUS ADENOCARCINOMA OF THYROID GLAND
C2037361|T047||CCS_10|SUPERFICIAL SPREADING ADENOCARCINOMA OF THYROID GLAND 
C2037361|T047||CCS_10|SUPERFICIAL SPREADING ADENOCARCINOMA OF THYROID GLAND
C2213260|T047||CCS_10|BASAL CELL ADENOCARCINOMA OF THYROID GLAND
C2213260|T047||CCS_10|BASAL CELL ADENOCARCINOMA OF THYROID GLAND 
C2213260|T047||CCS_10|BASAL CELL ADENOCARCINOMA OF THYROID
C2145031|T047||CCS_10|TRABECULAR ADENOCARCINOMA OF THYROID GLAND 
C2145031|T047||CCS_10|TRABECULAR ADENOCARCINOMA OF THYROID GLAND
C2189655|T047||CCS_10|VILLOUS ADENOCARCINOMA OF THYROID GLAND
C2189655|T047||CCS_10|VILLOUS ADENOCARCINOMA OF THYROID GLAND 
C2016174|T047||CCS_10|OXYPHILIC ADENOCARCINOMA OF THYROID GLAND
C2016174|T047||CCS_10|OXYPHILIC ADENOCARCINOMA OF THYROID GLAND 
C2075544|T047||CCS_10|CLEAR CELL ADENOCARCINOMA OF THYROID GLAND
C2075544|T047||CCS_10|CLEAR CELL ADENOCARCINOMA OF THYROID GLAND 
C2116005|T047||CCS_10|ALVEOLAR ADENOCARCINOMA OF THYROID GLAND 
C2116005|T047||CCS_10|ALVEOLAR ADENOCARCINOMA OF THYROID GLAND
C2203046|T047||CCS_10|WELL DIFFERENTIATED FOLLICULAR ADENOCARCINOMA OF THYROID GLAND 
C2203046|T047||CCS_10|WELL DIFFERENTIATED FOLLICULAR ADENOCARCINOMA OF THYROID GLAND
C2213261|T047||CCS_10|FOLLICULAR TRABECULAR ADENOCARCINOMA OF THYROID GLAND 
C2213261|T047||CCS_10|FOLLICULAR TRABECULAR ADENOCARCINOMA OF THYROID GLAND
C2116050|T047||CCS_10|FETAL ADENOCARCINOMA OF THYROID GLAND
C2116050|T047||CCS_10|FETAL ADENOCARCINOMA OF THYROID GLAND 
C2213262|T047||CCS_10|EMBRYONAL CARCINOSARCOMA OF THYROID GLAND 
C2213262|T047||CCS_10|EMBRYONAL CARCINOSARCOMA OF THYROID GLAND
C2213263|T047||CCS_10|MALIGNANT MYOEPITHELIOMA OF THYROID GLAND
C2213263|T047||CCS_10|MALIGNANT MYOEPITHELIOMA OF THYROID GLAND 
C2046351|T047||CCS_10|HISTIOCYTIC SARCOMA OF THYROID GLAND 
C2046351|T047||CCS_10|HISTIOCYTIC SARCOMA OF THYROID GLAND
C2111188|T047||CCS_10|LANGERHANS CELL SARCOMA OF THYROID GLAND 
C2111188|T047||CCS_10|LANGERHANS CELL SARCOMA OF THYROID GLAND
C2077774|T047||CCS_10|INTERDIGITATING DENDRITIC CELL SARCOMA OF THYROID GLAND 
C2077774|T047||CCS_10|INTERDIGITATING DENDRITIC CELL SARCOMA OF THYROID GLAND
C2213266|T047||CCS_10|FOLLICULAR DENDRITIC CELL SARCOMA OF THYROID GLAND 
C2213266|T047||CCS_10|FOLLICULAR DENDRITIC CELL SARCOMA OF THYROID GLAND
C2033237|T047||CCS_10|THYROID MALIGNANT CARCINOMA PAPILLARY METASTATIC TO CERVICAL LYMPH NODE
C2033237|T047||CCS_10|PAPILLARY THYROID CARCINOMA WITH METASTASIS TO CERVICAL LYMPH NODES 
C2033237|T047||CCS_10|PAPILLARY THYROID CARCINOMA WITH METASTASIS TO CERVICAL LYMPH NODES
C2033237|T047||CCS_10|PAPILLARY CARCINOMA OF THYROID METASTATIC TO CERVICAL LYMPH NODE
C3163939|T047||CCS_10|CARCINOMA OF THYROID
C3163939|T047||CCS_10|MALIGNANT EPITHELIAL NEOPLASM OF THYROID
C3163939|T047||CCS_10|MALIGNANT EPITHELIAL NEOPLASM OF THYROID 
C2116063|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF THYROID GLAND 
C2116063|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF THYROID GLAND
C2098465|T047||CCS_10|THYROID BIOPSY SHOWING MALIGNANT NEOPLASM
C2098465|T047||CCS_10|THYROID BIOPSY MALIGNANT NEOPLASM 
C2098465|T047||CCS_10|THYROID BIOPSY MALIGNANT NEOPLASM
C0278861|T047||CCS_10|RECURRENT THYROID CARCINOMA
C0278861|T047||CCS_10|RECURRENT THYROID GLAND CARCINOMA
C0278861|T047||CCS_10|THYROID CANCER RECURRENT
C0278861|T047||CCS_10|RECURRENT THYROID CANCER
C0278861|T047||CCS_10|THYROID CANCER, RECURRENT
C0278861|T047||CCS_10|RECURRENT CANCER OF THYROID GLAND
C0278861|T047||CCS_10|RECURRENT CANCER OF THYROID
C0278861|T047||CCS_10|RECURRENT CANCER OF THE THYROID GLAND
C0278861|T047||CCS_10|RECURRENT CANCER OF THE THYROID
C0278861|T047||CCS_10|RELAPSED CANCER OF THYROID GLAND
C0278861|T047||CCS_10|RELAPSED CANCER OF THYROID
C0278861|T047||CCS_10|RELAPSED CANCER OF THE THYROID GLAND
C0278861|T047||CCS_10|RELAPSED CANCER OF THE THYROID
C0278861|T047||CCS_10|RELAPSED THYROID CANCER
C0278861|T047||CCS_10|RELAPSED THYROID GLAND CANCER
C0205642|T047||CCS_10|ADENOCARCINOMAS, OXYPHILIC
C0205642|T047||CCS_10|OXYPHILIC ADENOCARCINOMAS
C0205642|T047||CCS_10|OXYPHILIC ADENOCARCINOMA
C0205642|T047||CCS_10|OXYPHILIC ADENOCARCINOMA 
C0205642|T047||CCS_10|OXYPHILIC ADENOCARCINOMA 
C0205642|T047||CCS_10|HUERTHLE CELL CARCINOMA
C0205642|T047||CCS_10|ONCOCYTOMA, MALIGNANT
C0205642|T047||CCS_10|HURTHLE CELL ADENOCARCINOMA
C0205642|T047||CCS_10|ONCOCYTIC ADENOCARCINOMA
C0205642|T047||CCS_10|ONCOCYTIC CARCINOMA
C0205642|T047||CCS_10|HURTHLE CELL CARCINOMA
C0205642|T047||CCS_10|FOLLICULAR CARCINOMA, OXYPHILIC CELL
C0205642|T047||CCS_10|OXYPHILIC ADENOCARCINOMA (MORPHOLOGIC ABNORMALITY)
C0205642|T047||CCS_10|HURTHLE CELL; ADENOCARCINOMA
C0205642|T047||CCS_10|HURTHLE CELL; CARCINOMA
C0205642|T047||CCS_10|CARCINOMA; HURTHLE CELL
C0205642|T047||CCS_10|ADENOCARCINOMA; HURTHLE CELL
C0205642|T047||CCS_10|ADENOCARCINOMA, OXYPHILIC
C1306310|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF THYROID GLAND 
C1306310|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF THYROID GLAND
C1306310|T047||CCS_10|THYROID MALIGNANT NEOPLASM PRIMARY
C1306310|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF THYROID GLAND 
C1282509|T047||CCS_10|METASTASIS FROM MALIGNANT NEOPLASM OF THYROID
C1282509|T047||CCS_10|METASTASIS FROM MALIGNANT NEOPLASM OF THYROID 
C1282509|T047||CCS_10|METASTASIS FROM MALIGNANT TUMOR OF THYROID 
C1282509|T047||CCS_10|METASTASIS FROM MALIGNANT TUMOR OF THYROID
C1282509|T047||CCS_10|METASTASIS FROM MALIGNANT TUMOUR OF THYROID
C1282469|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT NEOPLASM OF THYROID GLAND
C1282469|T047||CCS_10|THYROID MALIGNANT NEOPLASM LOCAL RECURRENCE
C1282469|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT NEOPLASM OF THYROID GLAND 
C1282469|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOR OF THYROID GLAND 
C1282469|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOR OF THYROID GLAND
C1282469|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOUR OF THYROID GLAND
C4038608|T047||CCS_10|DIFFUSE SCLEROSING PAPILLARY THYROID CARCINOMA 
C4038608|T047||CCS_10|DIFFUSE SCLEROSING PAPILLARY THYROID CARCINOMA
C1266050|T047||CCS_10|POORLY DIFFERENTIATED THYROID CARCINOMA
C1266050|T047||CCS_10|THYROID GLAND POORLY DIFFERENTIATED CARCINOMA
C1266050|T047||CCS_10|POORLY DIFFERENTIATED THYROID GLAND CARCINOMA
C1266050|T047||CCS_10|INSULAR CARCINOMA (MORPHOLOGIC ABNORMALITY)
C1266050|T047||CCS_10|INSULAR CARCINOMA
C1266050|T047||CCS_10|POORLY DIFFERENTIATED CARCINOMA OF THYROID GLAND
C1266050|T047||CCS_10|POORLY DIFFERENTIATED CARCINOMA OF THE THYROID GLAND
C0206683|T047||CCS_10|CARCINOMA, PAPILLARY, FOLLICULAR
C0206683|T047||CCS_10|THYROID GLAND PAPILLARY AND FOLLICULAR CARCINOMA
C0206683|T047||CCS_10|CARCINOMA, PAPILLARY, FOLLICULAR [DISEASE/FINDING]
C0206683|T047||CCS_10|PAPILLARY AND FOLLICULAR ADENOCARCINOMA
C0206683|T047||CCS_10|PAPILLARY AND FOLLICULAR CARCINOMA
C0206683|T047||CCS_10|FOLLICULAR VARIANT THYROID GLAND PAPILLARY CARCINOMA
C0206683|T047||CCS_10|PAPILLARY ADENOCARCINOMA - FOLLICULAR VARIANT
C0206683|T047||CCS_10|PAPILLARY ADENOCARCINOMA, FOLLICULAR VARIANT
C0206683|T047||CCS_10|PAPILLARY CARCINOMA - FOLLICULAR VARIANT
C0206683|T047||CCS_10|PAPILLARY CARCINOMA, FOLLICULAR VARIANT
C0206683|T047||CCS_10|PAPILLARY AND FOLLICULAR ADENOCARCINOMA (MORPHOLOGIC ABNORMALITY)
C0206683|T047||CCS_10|PAPILLARY CARCINOMA, FOLLICULAR VARIANT (MORPHOLOGIC ABNORMALITY)
C0206683|T047||CCS_10|CARCINOMA; FOLLICULAR WITH PAPILLARY
C0206683|T047||CCS_10|CARCINOMA; PAPILLARY WITH FOLLICULAR
C0206683|T047||CCS_10|CARCINOMA; PAPILLARY, FOLLICULAR VARIANT
C0206683|T047||CCS_10|FOLLICULAR; ADENOCARCINOMA WITH PAPILLARY
C0206683|T047||CCS_10|FOLLICULAR; CARCINOMA, WITH PAPILLARY
C0206683|T047||CCS_10|ADENOCARCINOMA; FOLLICULAR WITH PAPILLARY
C0206683|T047||CCS_10|ADENOCARCINOMA; PAPILLARY WITH FOLLICULAR
C0206683|T047||CCS_10|ADENOCARCINOMA; PAPILLARY, FOLLICULAR VARIANT
C0206683|T047||CCS_10|PAPILLARY; ADENOCARCINOMA WITH FOLLICULAR
C0206683|T047||CCS_10|PAPILLARY; ADENOCARCINOMA, FOLLICULAR VARIANT
C0206683|T047||CCS_10|PAPILLARY; CARCINOMA, FOLLICULAR VARIANT
C0206683|T047||CCS_10|PAPILLARY; CARCINOMA, WITH FOLLICULAR
C1386262|T047||CCS_10|FOLLICULAR; ADENOCARCINOMA, INTERMEDIATE DIFFERENTIATION
C1386262|T047||CCS_10|ADENOCARCINOMA; FOLLICULAR, INTERMEDIATE DIFFERENTIATION
C1386263|T047||CCS_10|FOLLICULAR; ADENOCARCINOMA, UNSPECIFIED SITE
C1386263|T047||CCS_10|ADENOCARCINOMA; FOLLICULAR, UNSPECIFIED SITE
C0334327|T047||CCS_10|FOLLICULAR ADENOCARCINOMA - MODERATELY DIFFERENTIATED
C0334327|T047||CCS_10|FOLLICULAR ADENOCARCINOMA - TRABECULAR
C0334327|T047||CCS_10|FOLLICULAR ADENOCARCINOMA, MODERATELY DIFFERENTIATED
C0334327|T047||CCS_10|FOLLICULAR ADENOCARCINOMA, TRABECULAR
C0334327|T047||CCS_10|FOLLICULAR CARCINOMA - MODERATELY DIFFERENTIATED
C0334327|T047||CCS_10|FOLLICULAR CARCINOMA - TRABECULAR
C0334327|T047||CCS_10|FOLLICULAR CARCINOMA, MODERATELY DIFFERENTIATED
C0334327|T047||CCS_10|FOLLICULAR CARCINOMA, TRABECULAR
C0334327|T047||CCS_10|FOLLICULAR ADENOCARCINOMA, TRABECULAR (MORPHOLOGIC ABNORMALITY)
C0334327|T047||CCS_10|CARCINOMA; FOLLICULAR, TRABECULAR
C0334327|T047||CCS_10|CARCINOMA; TRABECULAR, FOLLICULAR
C0334327|T047||CCS_10|LANGHANS; WUCHERNDE STRUMAW
C0334327|T047||CCS_10|FOLLICULAR; ADENOCARCINOMA, TRABECULAR
C0334327|T047||CCS_10|FOLLICULAR; CARCINOMA, TRABECULAR
C0334327|T047||CCS_10|ADENOCARCINOMA; FOLLICULAR, TRABECULAR
C0334327|T047||CCS_10|ADENOCARCINOMA; TRABECULAR FOLLICULAR
C0334327|T047||CCS_10|TRABECULAR; FOLLICULAR ADENOCARCINOMA
C0334327|T047||CCS_10|WUCHERNDE STRUMA LANGHANS
C0334327|T047||CCS_10|TRABECULAR FOLLICULAR ADENOCARCINOMA
C0334330|T047||CCS_10|NONENCAPSULATED SCLEROSING ADENOCARCINOMA
C0334330|T047||CCS_10|NONENCAPSULATED SCLEROSING CARCINOMA
C0334330|T047||CCS_10|NONENCAPSULATED SCLEROSING CARCINOMA (MORPHOLOGIC ABNORMALITY)
C0334330|T047||CCS_10|PAPILLARY CARCINOMA, DIFFUSE SCLEROSING
C0334330|T047||CCS_10|CARCINOMA; NONENCAPSULATED SCLEROSING
C0334330|T047||CCS_10|ADENOCARCINOMA; NONENCAPSULATED SCLEROSING
C0334330|T047||CCS_10|NONENCAPSULATED SCLEROSING; CARCINOMA
C0334330|T047||CCS_10|NONENCAPSULATED; SCLEROSING ADENOCARCINOMA
C0334330|T047||CCS_10|NONENCAPSULATED SCLEROSING NEOPLASM
C1541839|T047||CCS_10|CARCINOMA; C-CELL, UNSPECIFIED SITE
C1541839|T047||CCS_10|C-CELL; CARCINOMA, UNSPECIFIED SITE
C1391909|T047||CCS_10|CARCINOMA; FOLLICULAR, INTERMEDIATE DIFFERENTIATION
C1391909|T047||CCS_10|FOLLICULAR; CARCINOMA, INTERMEDIATE DIFFERENTIATION
C1391910|T047||CCS_10|CARCINOMA; FOLLICULAR, UNSPECIFIED SITE
C1391910|T047||CCS_10|FOLLICULAR; CARCINOMA, UNSPECIFIED SITE
C1391938|T047||CCS_10|CARCINOMA; PARAFOLLICULAR CELL, UNSPECIFIED SITE
C1391938|T047||CCS_10|PARAFOLLICULAR CELL; CARCINOMA, UNSPECIFIED SITE
C1397650|T047||CCS_10|FOLLICULAR; CARCINOMA, PURE FOLLICLE
C1399823|T047||CCS_10|HURTHLE CELL; TUMOR, MALIGNANT
C1399823|T047||CCS_10|TUMOR; HURTHLE CELL, MALIGNANT
C1321862|T047||CCS_10|NONENCAPSULATED SCLEROSING PAPILLARY THYROID CARCINOMA
C1321862|T047||CCS_10|THYROID GLAND DIFFUSE SCLEROSING PAPILLARY CARCINOMA
C1321862|T047||CCS_10|NONENCAPSULATED SCLEROSING TUMOR
C1321862|T047||CCS_10|NONENCAPSULATED SCLEROSING TUMOUR
C1321862|T047||CCS_10|NONENCAPSULATED; SCLEROSING TUMOR
C1321862|T047||CCS_10|TUMOR; NONENCAPSULATED SCLEROSING
C1410366|T047||CCS_10|STRUMA; TOXIC, TUMOR, MALIGNANT
C1410366|T047||CCS_10|TOXIC; GOITER, TUMOR, MALIGNANT
C0280258|T047||CCS_10|STAGE/CELL TYPE, THYROID CANCER
C0280258|T047||CCS_10|THYROID CANCER STAGE
C1336753|T047||CCS_10|THYROID GLAND LYMPHOMA
C1336753|T047||CCS_10|THYROID LYMPHOMA
C1336753|T047||CCS_10|PRIMARY THYROID GLAND LYMPHOMA
C1336753|T047||CCS_10|LYMPHOMA OF THYROID GLAND
C1336753|T047||CCS_10|LYMPHOMA OF THYROID
C1336753|T047||CCS_10|LYMPHOMA OF THE THYROID GLAND
C1336753|T047||CCS_10|LYMPHOMA OF THE THYROID
C0686505|T047||CCS_10|MALIGNANT NEOPLASM OF THYROGLOSSAL DUCT
C0686505|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF THYROGLOSSAL DUCT
C0686505|T047||CCS_10|THYROID NEOPLASM LOCATION: ECTOPIC THYROGLOSSAL DUCT MALIGNANT PRIMARY
C0686505|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF THYROGLOSSAL DUCT 
C0686505|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF THYROGLOSSAL DUCT 
C1302463|T047||CCS_10|PT4B: EXTRATHYROIDAL ANAPLASTIC CARCINOMA - SURGICALLY UNRESECTABLE (ANAPLASTIC CARCINOMA) (THYROID) 
C1302463|T047||CCS_10|PT4B: EXTRATHYROIDAL ANAPLASTIC CARCINOMA - SURGICALLY UNRESECTABLE (ANAPLASTIC CARCINOMA) (THYROID)
C1276616|T047||CCS_10|T2: TUMOR > 1 CM BUT < 4 CM, LIMITED TO THYROID 
C1276616|T047||CCS_10|T2: TUMOR > 1 CM BUT < 4 CM, LIMITED TO THYROID
C1276616|T047||CCS_10|T2: TUMOUR > 1 CM BUT < 4 CM, LIMITED TO THYROID
C1276616|T047||CCS_10|T2: TUMOR > 1 CM BUT < 4 CM, LIMITED TO THYROID (TUMOR STAGING)
C1276617|T047||CCS_10|T3: THYROID TUMOR > 4 CM, LIMITED TO THYROID 
C1276617|T047||CCS_10|T3: THYROID TUMOR > 4 CM, LIMITED TO THYROID
C1276617|T047||CCS_10|T3: THYROID TUMOUR > 4 CM, LIMITED TO THYROID
C1276617|T047||CCS_10|T3: THYROID TUMOR > 4 CM, LIMITED TO THYROID (TUMOR STAGING)
C1276618|T047||CCS_10|T4: THYROID TUMOR OF ANY SIZE EXTENDING BEYOND THE THYROID CAPSULE 
C1276618|T047||CCS_10|T4: THYROID TUMOR OF ANY SIZE EXTENDING BEYOND THE THYROID CAPSULE
C1276618|T047||CCS_10|T4: THYROID TUMOUR OF ANY SIZE EXTENDING BEYOND THE THYROID CAPSULE
C1276618|T047||CCS_10|T4: THYROID TUMOR OF ANY SIZE EXTENDING BEYOND THE THYROID CAPSULE (TUMOR STAGING)
C0346398|T047||CCS_10|MIXED FOLLICULAR AND PAPILLARY THYROID CARCINOMA
C0346398|T047||CCS_10|THYROID MALIGNANT CARCINOMA MIXED FOLLICULAR AND PAPILLARY
C0346398|T047||CCS_10|MIXED FOLLICULAR AND PAPILLARY THYROID CARCINOMA 
C0346398|T047||CCS_10|MIXED FOLLICULAR AND PAPILLARY THYROID CARCINOMA 
C0749424|T047||CCS_10|THYROID HURTHLE CELL CARCINOMA
C0749424|T047||CCS_10|THYROID GLAND ONCOCYTIC FOLLICULAR CARCINOMA
C0749424|T047||CCS_10|HURTHLE CELL THYROID GLAND CARCINOMA
C0749424|T047||CCS_10|HURTHLE CELL CARCINOMA OF THYROID
C0749424|T047||CCS_10|HURTHLE CELL CARCINOMA OF THYROID 
C0749424|T047||CCS_10|THYROID CARCINOMA, HURTHLE CELL
C0749424|T047||CCS_10|THYROID CANCER, FOLLICULAR, HURTHLE CELL TYPE
C0749424|T047||CCS_10|FOLLICULAR THYROID CANCER, HURTHLE CELL TYPE
C0749424|T047||CCS_10|HURTHLE CELL CARCINOMA OF THE THYROID
C0749424|T047||CCS_10|THYROID CANCER, HURTHLE CELL
C0749424|T047||CCS_10|HURTHLE CELL CARCINOMA OF THYROID 
C0749424|T047||CCS_10|THYROID MALIGNANT CARCINOMA HURTHLE CELL
C0749424|T047||CCS_10|HURTHLE CELL THYROID NEOPLASIA
C0749424|T047||CCS_10|CANCER OF THYROID, HURTHLE CELL
C0749424|T047||CCS_10|HURTHLE CELL NEOPLASM OF THE THYROID
C0749424|T047||CCS_10|HURTHLE CELL CARCINOMA OF THYROID GLAND
C0749424|T047||CCS_10|HURTHLE CELL CARCINOMA OF THE THYROID GLAND
C0749424|T047||CCS_10|ONCOCYTIC CARCINOMA OF THYROID
C0749424|T047||CCS_10|ONCOCYTIC CARCINOMA OF THE THYROID
C0749424|T047||CCS_10|THYROID GLAND HURTHLE CELL CARCINOMA
C0749424|T047||CCS_10|THYROID ONCOCYTIC CARCINOMA
C1302519|T047||CCS_10|PT4A: INTRATHYROIDAL ANAPLASTIC CARCINOMA - SURGICALLY RESECTABLE (ANAPLASTIC CARCINOMA) (THYROID) 
C1302519|T047||CCS_10|PT4A: INTRATHYROIDAL ANAPLASTIC CARCINOMA - SURGICALLY RESECTABLE (ANAPLASTIC CARCINOMA) (THYROID)
C2213271|T047||CCS_10|SEZARY SYNDROME OF THYROID GLAND 
C2213271|T047||CCS_10|SEZARY SYNDROME OF THYROID GLAND
C2113733|T047||CCS_10|PRECURSOR CELL LYMPHOBLASTIC LYMPHOMA OF THYROID GLAND 
C2113733|T047||CCS_10|PRECURSOR CELL LYMPHOBLASTIC LYMPHOMA OF THYROID GLAND
C2213265|T047||CCS_10|MAST CELL SARCOMA OF THYROID GLAND
C2213265|T047||CCS_10|MAST CELL SARCOMA OF THYROID GLAND 
C0346643|T047||CCS_10|MALIGNANT NEOPLASM OF HEPATIC DUCT
C0346643|T047||CCS_10|MALIGNANT EXTRAHEPATIC NEOPLASM HEPATIC DUCT
C0346643|T047||CCS_10|MALIGNANT NEOPLASM OF HEPATIC DUCT 
C0346643|T047||CCS_10|MALIGNANT NEOPLASM OF HEPATIC DUCT 
C0546835|T047||CCS_10|MALIGNANT NEOPLASM OF INTRAHEPATIC BILIARY PASSAGES
C0546835|T047||CCS_10|MALIGNANT NEOPLASM OF INTRAHEPATIC BILE DUCTS
C0546835|T047||CCS_10|MALIGNANT NEOPLASM OF INTRAHEPATIC BILE DUCT 
C0546835|T047||CCS_10|MALIGNANT NEOPLASM OF INTRAHEPATIC BILE DUCT
C0546835|T047||CCS_10|MALIGNANT TUMOR OF INTRAHEPATIC BILE DUCT
C0546835|T047||CCS_10|MAL NEO INTRAHEPAT DUCTS
C0546835|T047||CCS_10|CA INTRAHEPATIC BILE DUCTS
C0546835|T047||CCS_10|MALIGNANT NEOPLASM OF INTRAHEPATIC BILE DUCTS NOS 
C0546835|T047||CCS_10|CA INTRAHEPATIC BILE DUCTS 
C0546835|T047||CCS_10|MALIGNANT NEOPLASM OF INTRAHEPATIC BILE DUCTS NOS
C0546835|T047||CCS_10|MALIGNANT NEOPLASM OF INTRAHEPATIC BILIARY PASSAGES 
C0546835|T047||CCS_10|MALIGNANT NEOPLASM OF INTRAHEPATIC BILE DUCTS 
C0546835|T047||CCS_10|INTRAHEPATIC BILE DUCT CANCER
C0546835|T047||CCS_10|INTRAHEPATIC BILE DUCT CANCER NOS
C0546835|T047||CCS_10|MALIGNANT NEOPLASM OF INTRAHEPATIC GALL DUCT
C0546835|T047||CCS_10|MALIGNANT NEOPLASM OF INTRAHEPATIC GALL DUCT 
C2239176|T047||CCS_10|LIVER CELL CARCINOMA
C2239176|T047||CCS_10|CARCINOMA, HEPATOCELLULAR
C2239176|T047||CCS_10|CARCINOMAS, HEPATOCELLULAR
C2239176|T047||CCS_10|HEPATOCELLULAR CARCINOMAS
C2239176|T047||CCS_10|HEPATOMA
C2239176|T047||CCS_10|HEPATOMAS
C2239176|T047||CCS_10|HEPATOCELLULAR CARCINOMA
C2239176|T047||CCS_10|THIS IS UNCOMMON AND I WOULD TYPICALLY ERE ON EXCLUDING SINCE IT COULD BE OTHER THINGS (LEFT COMMON CAROTID) HOWEVER ON A LIVER INTAKE FORM I WILL INCLUDE IT
C2239176|T047||CCS_10|CARCINOMA OF LIVER 
C2239176|T047||CCS_10|HEPATOCELLULAR CARCINOMA OF LIVER 
C2239176|T047||CCS_10|HEPATOCELLULAR CARCINOMA OF LIVER
C2239176|T047||CCS_10|LIVER NEOPLASM MALIGNANT CARCINOMA
C2239176|T047||CCS_10|CARCINOMA OF LIVER
C2239176|T047||CCS_10|LIVER CARCINOMA
C2239176|T047||CCS_10|LIVER CELL CANCER (HEPATOCELLULAR CARCINOMA)
C2239176|T047||CCS_10|CARCINOMA, HEPATOCELLULAR [DISEASE/FINDING]
C2239176|T047||CCS_10|CANCERS, ADULT LIVER
C2239176|T047||CCS_10|ADULT LIVER CANCER
C2239176|T047||CCS_10|CANCER, ADULT LIVER
C2239176|T047||CCS_10|ADULT LIVER CANCERS
C2239176|T047||CCS_10|LIVER CANCERS, ADULT
C2239176|T047||CCS_10|LIVER CANCER, ADULT
C2239176|T047||CCS_10|LIVER CELL CARCINOMA, ADULT
C2239176|T047||CCS_10|LIVER CELL CARCINOMAS
C2239176|T047||CCS_10|CELL CARCINOMA, LIVER
C2239176|T047||CCS_10|CELL CARCINOMAS, LIVER
C2239176|T047||CCS_10|CARCINOMA, LIVER CELL
C2239176|T047||CCS_10|CARCINOMAS, LIVER CELL
C2239176|T047||CCS_10|HEPATIC CELL CARCINOMA
C2239176|T047||CCS_10|PRIMARY CARCINOMA OF LIVER
C2239176|T047||CCS_10|LIVER NEOPLASM MALIGNANT CARCINOMA PRIMARY
C2239176|T047||CCS_10|PRIMARY CARCINOMA OF LIVER 
C2239176|T047||CCS_10|HCC
C2239176|T047||CCS_10|CARCINOMA, HEPATOCELLULAR, MALIGNANT
C2239176|T047||CCS_10|[M]HEPATOCELLULAR CARCINOMA NOS
C2239176|T047||CCS_10|CARCINOMA OF THE LIVER CELLS
C2239176|T047||CCS_10|PRIMARY CARCINOMA OF THE LIVER CELLS
C2239176|T047||CCS_10|CARCINOMA OF LIVER CELLS
C2239176|T047||CCS_10|PRIMARY CARCINOMA OF LIVER CELLS
C2239176|T047||CCS_10|LIVER CELL CARCINOMA (CLINICAL)
C2239176|T047||CCS_10|HEPATOCELLULAR CARCINOMA (CLINICAL)
C2239176|T047||CCS_10|CARCINOMA LIVER
C2239176|T047||CCS_10|CARCINOMA HEPATOCELLULAR
C2239176|T047||CCS_10|HEPATOCARCINOMA
C2239176|T047||CCS_10|HEPATOMA, MALIGNANT
C2239176|T047||CCS_10|MALIGNANT HEPATOMA
C2239176|T047||CCS_10|LCC - LIVER CELL CARCINOMA
C2239176|T047||CCS_10|HCC - HEPATOCELLULAR CARCINOMA
C2239176|T047||CCS_10|HEPATOCELLULAR CARCINOMA (MORPHOLOGIC ABNORMALITY)
C2239176|T047||CCS_10|LIVER CELL CARCINOMA 
C2239176|T047||CCS_10|PRIMARY CARCINOMA OF LIVER 
C2239176|T047||CCS_10|CARCINOMA; HEPATIC CELL
C2239176|T047||CCS_10|CARCINOMA; HEPATOCELLULAR
C2239176|T047||CCS_10|HEPATIC CELL; CARCINOMA
C2239176|T047||CCS_10|HEPATOCELLULAR; CARCINOMA
C2239176|T047||CCS_10|HEPATOCELLULAR CARCINOMA, NOS
C2239176|T047||CCS_10|HEPATOMA, NOS
C2239176|T047||CCS_10|CARCINOMA OF LIVER, SPECIFIED AS PRIMARY
C2239176|T047||CCS_10|CARCINOMA OF LIVER CELL
C0206624|T047||CCS_10|HEPATOBLASTOMA
C0206624|T047||CCS_10|HEPATOBLASTOMAS
C0206624|T047||CCS_10|HEPATOBLASTOMA OF LIVER
C0206624|T047||CCS_10|HEPATOBLASTOMA OF LIVER 
C0206624|T047||CCS_10|HEPATOBLASTOMA [DISEASE/FINDING]
C0206624|T047||CCS_10|HBL
C0206624|T047||CCS_10|HEPATOBLASTOMA, MALIGNANT
C0206624|T047||CCS_10|PEDIATRIC HEPATOBLASTOMA
C0206624|T047||CCS_10|PEDIATRIC EMBRYONAL HEPATOMA
C0206624|T047||CCS_10|HEPATOBLASTOMA NOS
C0206624|T047||CCS_10|EMBRYONAL HEPATOMA
C0206624|T047||CCS_10|HBL - HEPATOBLASTOMA
C0206624|T047||CCS_10|HEPATOBLASTOMA (CLINICAL)
C0206624|T047||CCS_10|HEPATOBLASTOMA 
C0206624|T047||CCS_10|HEPATOBLASTOMA (MORPHOLOGIC ABNORMALITY)
C0206624|T047||CCS_10|CHILDHOOD HEPATOBLASTOMA
C0206624|T047||CCS_10|HEPATOBLASTOMA, CHILDHOOD
C0206624|T047||CCS_10|EMBRYONAL; HEPATOMA
C0206624|T047||CCS_10|HEPATOMA; EMBRYONAL
C0345907|T047||CCS_10|ANGIOSARCOMA OF LIVER
C0345907|T047||CCS_10|HEPATIC ANGIOSARCOMA
C0345907|T047||CCS_10|HEMANGIOSARCOMA OF LIVER
C0345907|T047||CCS_10|HEMANGIOSARCOMA OF LIVER 
C0345907|T047||CCS_10|HEPATIC HEMANGIOSARCOMA
C0345907|T047||CCS_10|LIVER ANGIOSARCOMA
C0345907|T047||CCS_10|ANGIOSARCOMA OF LIVER 
C0345907|T047||CCS_10|HEMANGIOSARCOMA OF LIVER 
C0345907|T047||CCS_10|LIVER NEOPLASM MALIGNANT ANGIOSARCOMA
C0345907|T047||CCS_10|ANGIOSARCOMA OF LIVER 
C0345907|T047||CCS_10|PRIMARY ANGIOSARCOMA OF LIVER
C0345907|T047||CCS_10|LIVER; ANGIOSARCOMA
C0345907|T047||CCS_10|ANGIOSARCOMA; LIVER
C0345907|T047||CCS_10|HEMANGIOSARCOMA OF THE LIVER
C0345907|T047||CCS_10|LIVER HEMANGIOSARCOMA
C0345907|T047||CCS_10|ANGIOSARCOMA OF THE LIVER
C0345907|T047||CCS_10|PRIMARY ANGIOSARCOMA OF THE LIVER
C0345905|T047||CCS_10|INTRAHEPATIC BILE DUCT CARCINOMA
C0345905|T047||CCS_10|CHOLANGIOCARCINOMA OF INTRAHEPATIC BILE DUCT 
C0345905|T047||CCS_10|CHOLANGIOCARCINOMA OF INTRAHEPATIC BILE DUCT
C0345905|T047||CCS_10|CARCINOMA OF INTRAHEPATIC BILE DUCT
C0345905|T047||CCS_10|CARCINOMA OF INTRAHEPATIC BILE DUCT 
C0345905|T047||CCS_10|CHOLANGIOCARCINOMA, INTRAHEPATIC, MALIGNANT
C0345905|T047||CCS_10|INTRAHEPATIC CARCINOMA OF THE BILE DUCT
C0345905|T047||CCS_10|INTRAHEPATIC CARCINOMA OF BILE DUCT
C0345905|T047||CCS_10|CHOLANGIOCARCINOMAS, INTRAHEPATIC
C0345905|T047||CCS_10|INTRAHEPATIC CHOLANGIOCARCINOMAS
C0345905|T047||CCS_10|CHOLANGIOCARCINOMA, INTRAHEPATIC
C0345905|T047||CCS_10|INTRAHEPATIC CHOLANGIOCARCINOMA
C0345905|T047||CCS_10|INTRAHEPATIC BILE DUCT CARCINOMA 
C0345905|T047||CCS_10|INTRAHEPATIC CHOLANGIOCELLULAR CARCINOMA
C0348340|T047||CCS_10|OTHER SPECIFIED CARCINOMAS OF LIVER
C0348340|T047||CCS_10|[X]OTHER SPECIFIED CARCINOMAS OF LIVER
C0348340|T047||CCS_10|OTHER SPECIFIED CARCINOMA OF LIVER
C0348340|T047||CCS_10|OTHER SPECIFIED CARCINOMA OF LIVER 
C0348340|T047||CCS_10|[X]OTHER SPECIFIED CARCINOMAS OF LIVER 
C0345904|T047||CCS_10|LIVER, UNSPECIFIED
C0345904|T047||CCS_10|MALIGNANT NEOPLASM OF LIVER, UNSPECIFIED
C0345904|T047||CCS_10|MALIGNANT NEOPLASM OF LIVER
C0345904|T047||CCS_10|LIVER CANCER
C0345904|T047||CCS_10|LIVER CANCER 
C0345904|T047||CCS_10|LIVER NEOPLASM MALIGNANT
C0345904|T047||CCS_10|MALIGNANT NEOPLASM OF LIVER 
C0345904|T047||CCS_10|HEPATIC NEOPLASMS MALIGNANT
C0345904|T047||CCS_10|CANCER, HEPATIC
C0345904|T047||CCS_10|CANCERS, HEPATIC
C0345904|T047||CCS_10|HEPATIC CANCERS
C0345904|T047||CCS_10|CANCERS, LIVER
C0345904|T047||CCS_10|LIVER CANCERS
C0345904|T047||CCS_10|MALIGNANT TUMOR OF LIVER
C0345904|T047||CCS_10|MALIGNANT NEO LIVER NOS
C0345904|T047||CCS_10|MALIGNANT NEOPLASM OF LIVER, NOT SPECIFIED AS PRIMARY OR SECONDARY
C0345904|T047||CCS_10|HEPATIC CANCER
C0345904|T047||CCS_10|CANCER, LIVER
C0345904|T047||CCS_10|MALIG NEOPLASM OF LIVER, NOT SPECIFIED AS PRIMARY OR SEC
C0345904|T047||CCS_10|CANCERS, HEPATOCELLULAR
C0345904|T047||CCS_10|HEPATOCELLULAR CANCERS
C0345904|T047||CCS_10|MALIGNANT NEOPLASM OF LIVER UNSPECIFIED 
C0345904|T047||CCS_10|MALIGNANT TUMOR OF LIVER 
C0345904|T047||CCS_10|MALIGNANT NEOPLASM OF LIVER UNSPECIFIED
C0345904|T047||CCS_10|MALIGNANT TUMOUR OF LIVER
C0345904|T047||CCS_10|LIVER--CANCER
C0345904|T047||CCS_10|CANCER, HEPATOCELLULAR
C0345904|T047||CCS_10|HEPATIC NEOPLASM MALIGNANT NOS
C0345904|T047||CCS_10|MALIGNANT HEPATIC NEOPLASM
C0345904|T047||CCS_10|MALIGNANT LIVER TUMOR
C0345904|T047||CCS_10|HEPATIC TUMOUR MALIGNANT
C0345904|T047||CCS_10|LIVER, CANCER OF
C0345904|T047||CCS_10|MALIGNANT LIVER TUMOUR
C0345904|T047||CCS_10|HEPATIC NEOPLASM MALIGNANT
C0345904|T047||CCS_10|HEPATIC TUMOR MALIGNANT
C0345904|T047||CCS_10|HEPATOCELLULAR CANCER
C0345904|T047||CCS_10|CANCER OF THE LIVER
C0345904|T047||CCS_10|CA - LIVER CANCER
C0345904|T047||CCS_10|MALIGNANT NEOPLASM OF LIVER 
C0345904|T047||CCS_10|MALIGNANT NEOPLASM OF LIVER, NOS
C0345904|T047||CCS_10|CANCER OF LIVER
C0345904|T047||CCS_10|NEOPLASM MALIG;LIVER
C0345904|T047||CCS_10|MALIGNANT NEOSPLASM OF THE LIVER
C0348339|T047||CCS_10|OTHER SARCOMAS OF LIVER
C0348339|T047||CCS_10|OTHER SARCOMA OF LIVER
C0348339|T047||CCS_10|[X]OTHER SARCOMAS OF THE LIVER 
C0348339|T047||CCS_10|[X]OTHER SARCOMAS OF THE LIVER
C0348339|T047||CCS_10|OTHER SARCOMA OF LIVER 
C0153448|T047|16|CCS_10|MALIGNANT NEOPLASM OF LIVER AND INTRAHEPATIC BILE DUCTS|CANCER OF LIVER AND INTRAHEPATIC BILE DUCT
C0153448|T047|16|CCS_10|CANCER OF LIVER AND INTRAHEPATIC BILE DUCT|CANCER OF LIVER AND INTRAHEPATIC BILE DUCT
C0153448|T047|16|CCS_10|MALIGNANT NEOPLASM OF LIVER AND INTRAHEPATIC BILE DUCTS NOS|CANCER OF LIVER AND INTRAHEPATIC BILE DUCT
C0153448|T047|16|CCS_10|MALIGNANT NEOPLASM OF LIVER AND INTRAHEPATIC BILE DUCTS NOS |CANCER OF LIVER AND INTRAHEPATIC BILE DUCT
C0153448|T047|16|CCS_10|MALIGNANT NEOPLASM OF LIVER AND INTRAHEPATIC BILE DUCTS |CANCER OF LIVER AND INTRAHEPATIC BILE DUCT
C0153448|T047|16|CCS_10|MALIGNANT NEOPLASM OF LIVER AND INTRAHEPATIC BILE DUCTS |CANCER OF LIVER AND INTRAHEPATIC BILE DUCT
C2837938|T047||CCS_10|MALIGNANT NEOPLASM OF LIVER, PRIMARY, UNSPECIFIED AS TO TYPE
C2188066|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF INTRAHEPATIC BILE DUCT
C2188066|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF INTRAHEPATIC BILE DUCT 
C2078126|T047||CCS_10|UNDIFFERENTIATED SARCOMA OF INTRAHEPATIC BILE DUCT 
C2078126|T047||CCS_10|UNDIFFERENTIATED SARCOMA OF INTRAHEPATIC BILE DUCT
C0279000|T047||CCS_10|LIVER AND INTRAHEPATIC BILE DUCT CARCINOMA
C0279000|T047||CCS_10|LIVER AND INTRAHEPATIC BILIARY TRACT CARCINOMA
C0279000|T047||CCS_10|LIVER AND HEPATOBILIARY CANCER, NOS
C0279000|T047||CCS_10|LIVER/HEPATOBILIARY CANCER
C0279000|T047||CCS_10|LIVER CANCER
C0279000|T047||CCS_10|LIVER AND INTRAHEPATIC BILIARY TRACT CANCER
C0279000|T047||CCS_10|HEPATIC CANCER
C0279000|T047||CCS_10|CANCER OF LIVER
C0279000|T047||CCS_10|CANCER OF THE LIVER
C0279000|T047||CCS_10|LIVER AND INTRAHEPATIC BILE DUCT CANCER
C0279000|T047||CCS_10|PRIMARY LIVER CARCINOMA
C0279000|T047||CCS_10|CANCER OF LIVER AND INTRAHEPATIC BILIARY TRACT
C0279000|T047||CCS_10|CANCER OF THE LIVER AND INTRAHEPATIC BILIARY TRACT
C0024620|T047||CCS_10|PRIMARY LIVER CANCER
C0024620|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF LIVER
C0024620|T047||CCS_10|MAL NEO LIVER, PRIMARY
C0024620|T047||CCS_10|PRIMARY MALIGNANT LIVER NEOPLASM
C0024620|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF LIVER 
C0024620|T047||CCS_10|LIVER NEOPLASM MALIGNANT PRIMARY
C0024620|T047||CCS_10|CA LIVER - PRIMARY 
C0024620|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF LIVER NOS 
C0024620|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF LIVER 
C0024620|T047||CCS_10|CA LIVER - PRIMARY
C0024620|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF LIVER NOS
C0024620|T047||CCS_10|MALIGNANT NEOPLASM OF LIVER, PRIMARY
C0024620|T047||CCS_10|LIVER, CANCER OF, PRIMARY
C0024620|T047||CCS_10|PRIMARY CANCER OF LIVER
C0024620|T047||CCS_10|CANCER OF LIVER, PRIMARY
C0206630|T047||CCS_10|SARCOMA, ENDOMETRIAL STROMAL
C0206630|T047||CCS_10|ENDOMETRIAL STROMAL SARCOMAS
C0206630|T047||CCS_10|SARCOMAS, ENDOMETRIAL STROMAL
C0206630|T047||CCS_10|STROMAL SARCOMA, ENDOMETRIAL
C0206630|T047||CCS_10|STROMAL SARCOMAS, ENDOMETRIAL
C0206630|T047||CCS_10|SARCOMA, ENDOMETRIAL STROMAL [DISEASE/FINDING]
C0206630|T047||CCS_10|ENDOMETRIAL STROMAL SARCOMA
C0206630|T047||CCS_10|ENDOMETRIOID STROMAL SARCOMA
C0206630|T047||CCS_10|ENDOMETRIAL STROMAL SARCOMA 
C0206630|T047||CCS_10|STROMAL SARCOMA, ENDOMETRIAL, MALIGNANT
C0206630|T047||CCS_10|PRIMARY MALIGNANT STROMAL SARCOMA OF ENDOMETRIUM
C0206630|T047||CCS_10|ENDOMETRIAL SARCOMA
C0206630|T047||CCS_10|ENDOMETRIAL SARCOMA, NOS
C0206630|T047||CCS_10|STROMAL SARCOMA, NOS
C0346191|T047||CCS_10|CARCINOMA IN SITU OF ENDOMETRIUM
C0346191|T047||CCS_10|CA ENDOMETRIUM STAGE 0
C0346191|T047||CCS_10|ENDOMETRIAL CANCER STAGE 0
C0346191|T047||CCS_10|CARCINOMA IN SITU OF ENDOMETRIUM 
C0346191|T047||CCS_10|CANCER OF ENDOMETRIUM STAGE 0
C0346191|T047||CCS_10|ENDOMETRIAL CARCINOMA STAGE 0
C0346191|T047||CCS_10|CARCINOMA ENDOMETRIAL STAGE 0
C0346191|T047||CCS_10|STAGE 0 ENDOMETRIAL CANCER
C0346191|T047||CCS_10|CANCER OF THE ENDOMETRIUM, STAGE 0
C0346191|T047||CCS_10|CARCINOMA OF THE ENDOMETRIUM, STAGE 0
C0346191|T047||CCS_10|ENDOMETRIAL CANCER, STAGE 0
C0346191|T047||CCS_10|ENDOMETRIAL CARCINOMA, STAGE 0
C0346191|T047||CCS_10|STAGE 0 CANCER OF THE ENDOMETRIUM
C0346191|T047||CCS_10|STAGE 0 CARCINOMA OF THE ENDOMETRIUM
C0346191|T047||CCS_10|STAGE 0 UTERINE CANCER
C0346191|T047||CCS_10|UTERINE CANCER, STAGE 0
C0476089|T047||CCS_10|CARCINOMA OF ENDOMETRIUM
C0476089|T047||CCS_10|CANCER, ENDOMETRIAL
C0476089|T047||CCS_10|CANCERS, ENDOMETRIAL
C0476089|T047||CCS_10|ENDOMETRIAL CANCERS
C0476089|T047||CCS_10|ENDOMETRIAL CANCER
C0476089|T047||CCS_10|CA ENDOMETRIUM
C0476089|T047||CCS_10|ENDOMETRIAL CARCINOMA (NOS)
C0476089|T047||CCS_10|CANCERS, ENDOMETRIUM
C0476089|T047||CCS_10|ENDOMETRIUM CANCERS
C0476089|T047||CCS_10|CANCER, ENDOMETRIUM
C0476089|T047||CCS_10|ENDOMETRIAL CARCINOMA
C0476089|T047||CCS_10|ENDOMETRIAL CA
C0476089|T047||CCS_10|UTERINE NEOPLASM, MALIGNANT - OF ENDOMETRIUM CARCINOMA
C0476089|T047||CCS_10|ENDOMETRIAL CARCINOMA 
C0476089|T047||CCS_10|CARCINOMA, ENDOMETRIAL
C0476089|T047||CCS_10|CARCINOMAS, ENDOMETRIAL
C0476089|T047||CCS_10|ENDOMETRIAL CARCINOMAS
C0476089|T047||CCS_10|ENDOMETRIUM CARCINOMA
C0476089|T047||CCS_10|ENDOMETRIUM CARCINOMAS
C0476089|T047||CCS_10|ENDOMETRIUM--CANCER
C0476089|T047||CCS_10|CARCINOMA, ENDOMETRIAL, MALIGNANT
C0476089|T047||CCS_10|CARCINOMA OF THE ENDOMETRIUM
C0476089|T047||CCS_10|CANCER OF ENDOMETRIUM
C0476089|T047||CCS_10|CARCINOMA ENDOMETRIAL
C0476089|T047||CCS_10|ENDOMETRIAL CANCER NOS
C0476089|T047||CCS_10|ENDOMETRIUM CANCER
C0476089|T047||CCS_10|CANCER OF THE ENDOMETRIUM
C0476089|T047||CCS_10|ENDOMETRIAL CARCINOMA 
C0476089|T047||CCS_10|CARCINOMA;ENDOMETRIAL
C0813216|T047||CCS_10|CORPUS UTERI CARCINOMA
C0813216|T047||CCS_10|CARCINOMA OF CORPUS UTERI
C0813216|T047||CCS_10|MALIGNANT EPITHELIAL NEOPLASM OF BODY OF UTERUS 
C0813216|T047||CCS_10|MALIGNANT EPITHELIAL NEOPLASM OF BODY OF UTERUS
C0813216|T047||CCS_10|CARCINOMA BODY OF UTERUS
C0813216|T047||CCS_10|UTERINE NEOPLASM, MALIGNANT - OF CORPUS UTERI CARCINOMA
C0813216|T047||CCS_10|CARCINOMA OF CORPUS UTERI 
C0813216|T047||CCS_10|CARCINOMA CORPUS UTERI
C1153706|T047||CCS_10|UTERINE ADENOCARCINOMA
C1153706|T047||CCS_10|ADENOCARCINOMA OF UTERUS
C1153706|T047||CCS_10|ADENOCARCINOMA OF UTERUS 
C1153706|T047||CCS_10|ENDOMETRIAL ADENOCARCINOMA
C1153706|T047||CCS_10|[M]ENDOMETRIOID ADENOMAS AND CARCINOMAS
C1153706|T047||CCS_10|[M]ENDOMETRIOID ADENOMAS AND CARCINOMAS (MORPHOLOGIC ABNORMALITY)
C1153706|T047||CCS_10|[M]ENDOMETRIOID ADENOMA OR CARCINOMA NOS (MORPHOLOGIC ABNORMALITY)
C1153706|T047||CCS_10|[M]ENDOMETRIOID ADENOMA OR CARCINOMA NOS
C1153706|T047||CCS_10|ADENOCARCINOMA, ENDOMETRIAL, MALIGNANT
C1153706|T047||CCS_10|ADENOCARCINOMA OF ENDOMETRIUM 
C1153706|T047||CCS_10|ADENOCARCINOMA OF ENDOMETRIUM
C1153706|T047||CCS_10|UTERINE ADENOCARCINOMA ENDOMETRIUM
C1153706|T047||CCS_10|ADENOCARCINOMA OF THE ENDOMETRIUM
C1153706|T047||CCS_10|ADENOCARCINOMA ENDOMETRIAL
C1153706|T047||CCS_10|ADENOCARCINOMA OF ENDOMETRIUM 
C1153706|T047||CCS_10|ADENOCARCINOMA OF UTERUS 
C1153706|T047||CCS_10|ADENOCARCINOMA OF THE UTERUS
C1153706|T047||CCS_10|UTERINE CANCER, ADENOCARCINOMA
C1153706|T047||CCS_10|UTERUS CANCER, ADENOCARCINOMA
C0153574|T047||CCS_10|CORPUS UTERI, UNSPECIFIED
C0153574|T047||CCS_10|MALIGNANT NEOPLASM OF CORPUS UTERI
C0153574|T047||CCS_10|MALIGNANT NEOPLASM OF CORPUS UTERI, UNSPECIFIED
C0153574|T047||CCS_10|MALIGNANT NEOPLASM OF BODY OF UTERUS
C0153574|T047||CCS_10|MALIGNANT NEOPLASM OF CORPUS UTERI 
C0153574|T047||CCS_10|MALIGNANT TUMOR OF CORPUS UTERI
C0153574|T047||CCS_10|MALIGNANT NEOPLASM OF CORPUS UTERI NOS
C0153574|T047||CCS_10|MALIGNANT TUMOR OF BODY OF UTERUS
C0153574|T047||CCS_10|BODY OF UTERUS CA
C0153574|T047||CCS_10|MALIGNANT NEOPLASM OF BODY OF UTERUS NOS
C0153574|T047||CCS_10|UTERUS BODY CA
C0153574|T047||CCS_10|MALIGNANT NEOPLASM OF CORPUS UTERI NOS 
C0153574|T047||CCS_10|MALIGNANT TUMOUR OF BODY OF UTERUS
C0153574|T047||CCS_10|MALIGNANT TUMOUR OF BODY OF UTERUS 
C0153574|T047||CCS_10|MALIGNANT NEOPLASM OF BODY OF UTERUS NOS 
C0153574|T047||CCS_10|CANCER OF UTERINE BODY
C0153574|T047||CCS_10|UTERINE CANCER, BODY
C0153574|T047||CCS_10|CANCER OF BODY OF UTERUS
C0153574|T047||CCS_10|MALIGNANT NEOPLASM OF BODY OF UTERUS 
C0153574|T047||CCS_10|UTERINE CORPUS CANCER
C0153574|T047||CCS_10|MALIGNANT CORPUS UTERI NEOPLASM
C0153574|T047||CCS_10|MALIGNANT CORPUS UTERI TUMOR
C0153574|T047||CCS_10|MALIGNANT NEOPLASM OF UTERINE BODY
C0153574|T047||CCS_10|MALIGNANT NEOPLASM OF THE UTERINE BODY
C0153574|T047||CCS_10|MALIGNANT TUMOR OF UTERINE BODY
C0153574|T047||CCS_10|MALIGNANT TUMOR OF THE UTERINE BODY
C0153574|T047||CCS_10|MALIGNANT UTERINE BODY NEOPLASM
C0153574|T047||CCS_10|MALIGNANT UTERINE BODY TUMOR
C0153574|T047||CCS_10|MALIGNANT UTERINE CORPUS NEOPLASM
C0153574|T047||CCS_10|MALIGNANT UTERINE CORPUS TUMOR
C0338113|T047||CCS_10|SARCOMA OF UTERUS 
C0338113|T047||CCS_10|SARCOMA OF UTERUS
C0338113|T047||CCS_10|UTERINE SARCOMA
C0338113|T047||CCS_10|SARCOMA UTERUS
C0338113|T047||CCS_10|UTERINE SARCOMA NOS
C0338113|T047||CCS_10|SARCOMA OF UTERUS 
C0338113|T047||CCS_10|SARCOMA OF THE UTERUS
C0338113|T047||CCS_10|UTERINE CANCER, SARCOMA
C0338113|T047||CCS_10|UTERINE CORPUS CANCER, SARCOMA
C0338113|T047||CCS_10|UTERUS CANCER, SARCOMA
C0338113|T047||CCS_10|CORPUS UTERI SARCOMA
C0338113|T047||CCS_10|SARCOMA OF BODY OF UTERUS
C0338113|T047||CCS_10|SARCOMA OF CORPUS UTERI
C0338113|T047||CCS_10|SARCOMA OF UTERINE BODY
C0338113|T047||CCS_10|SARCOMA OF UTERINE CORPUS
C0338113|T047||CCS_10|SARCOMA OF THE BODY OF UTERUS
C0338113|T047||CCS_10|SARCOMA OF THE CORPUS UTERI
C0338113|T047||CCS_10|SARCOMA OF THE UTERINE BODY
C0338113|T047||CCS_10|SARCOMA OF THE UTERINE CORPUS
C0338113|T047||CCS_10|UTERINE BODY SARCOMA
C0338113|T047||CCS_10|UTERINE CORPUS SARCOMA
C0338113|T047||CCS_10|UTERUS SARCOMA
C0338113|T047||CCS_10|BODY OF UTERUS SARCOMA
C1297960|T047||CCS_10|UTERINE NEOPLASM, MALIGNANT CORPUS UTERI, BY DIRECT EXTENSION FROM BLADDER
C1297960|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM BLADDER 
C1297960|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM BLADDER
C1297960|T047||CCS_10|MALIGNANT TUMOR INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM BLADDER 
C1297960|T047||CCS_10|MALIGNANT TUMOR INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM BLADDER
C1297960|T047||CCS_10|MALIGNANT TUMOUR INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM BLADDER
C1297961|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM OVARY 
C1297961|T047||CCS_10|UTERINE NEOPLASM, MALIGNANT CORPUS UTERI, BY DIRECT EXTENSION FROM OVARY
C1297961|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM OVARY
C1297961|T047||CCS_10|MALIGNANT TUMOR INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM OVARY 
C1297961|T047||CCS_10|MALIGNANT TUMOR INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM OVARY
C1297961|T047||CCS_10|MALIGNANT TUMOUR INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM OVARY
C1297962|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM UTERINE CERVIX
C1297962|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM UTERINE CERVIX 
C1297962|T047||CCS_10|UTERINE NEOPLASM, MALIGNANT CORPUS UTERI BY DIRECT EXTENSION FROM UTERINE CERVIX
C1297962|T047||CCS_10|MALIGNANT TUMOR INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM UTERINE CERVIX 
C1297962|T047||CCS_10|MALIGNANT TUMOR INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM UTERINE CERVIX
C1297962|T047||CCS_10|MALIGNANT TUMOUR INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM UTERINE CERVIX
C1297963|T047||CCS_10|UTERINE NEOPLASM, MALIGNANT CORPUS UTERI, BY DIRECT EXTENSION FROM VAGINA
C1297963|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM VAGINA 
C1297963|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM VAGINA
C1297963|T047||CCS_10|MALIGNANT TUMOR INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM VAGINA 
C1297963|T047||CCS_10|MALIGNANT TUMOR INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM VAGINA
C1297963|T047||CCS_10|MALIGNANT TUMOUR INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM VAGINA
C1298046|T047||CCS_10|UTERINE NEOPLASM, MALIGNANT CORPUS UTERI BY DIRECT EXTENSION FROM FALLOPIAN TUBE
C1298046|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM FALLOPIAN TUBE 
C1298046|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM FALLOPIAN TUBE
C1298046|T047||CCS_10|MALIGNANT TUMOR INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM FALLOPIAN TUBE 
C1298046|T047||CCS_10|MALIGNANT TUMOR INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM FALLOPIAN TUBE
C1298046|T047||CCS_10|MALIGNANT TUMOUR INVOLVING UTERINE CORPUS BY DIRECT EXTENSION FROM FALLOPIAN TUBE
C0153567|T047||CCS_10|UTERINE CANCER
C0153567|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS, PART UNSPECIFIED
C0153567|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS 
C0153567|T047||CCS_10|CANCER OF UTERUS
C0153567|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS
C0153567|T047||CCS_10|UTERINE CANCER 
C0153567|T047||CCS_10|CANCER, UTERINE
C0153567|T047||CCS_10|CANCERS, UTERINE
C0153567|T047||CCS_10|UTERINE CANCERS
C0153567|T047||CCS_10|CANCERS, UTERUS
C0153567|T047||CCS_10|UTERUS CANCERS
C0153567|T047||CCS_10|MALIGNANT TUMOR OF UTERUS
C0153567|T047||CCS_10|MALIG NEOPL UTERUS NOS
C0153567|T047||CCS_10|CANCER, UTERUS
C0153567|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS, PART UNSPECIFIED 
C0153567|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS 
C0153567|T047||CCS_10|CA - CANCER OF UTERUS
C0153567|T047||CCS_10|MALIGNANT TUMOUR OF UTERUS
C0153567|T047||CCS_10|UTERINE CA NOS
C0153567|T047||CCS_10|CA UTERUS NOS
C0153567|T047||CCS_10|UTERUS--CANCER
C0153567|T047||CCS_10|UTERINE CANCER, NOS
C0153567|T047||CCS_10|-- UTERINE CANCER
C0153567|T047||CCS_10|UTERINE CANCER NOS
C0153567|T047||CCS_10|UTERUS CANCER
C0153567|T047||CCS_10|CANCER OF THE UTERUS
C0153567|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS, NOS
C0153567|T047||CCS_10|MALIGNANT NEOPLASM OF THE UTERUS
C0153567|T047||CCS_10|MALIGNANT TUMOR OF THE UTERUS
C0153567|T047||CCS_10|MALIGNANT UTERINE NEOPLASM
C0153567|T047||CCS_10|MALIGNANT UTERINE TUMOR
C0153567|T047||CCS_10|NEOPLASM MALIG;UTERUS
C0153567|T047||CCS_10|MALIGNANT NEOSPLASM OF THE UTERUS
C0153569|T047||CCS_10|MALIGNANT NEOPLASM OF ENDOCERVIX
C0153569|T047||CCS_10|MALIGNANT NEOPLASM OF CERVICAL CANAL 
C0153569|T047||CCS_10|MALIGNANT NEOPLASM OF ENDOCERVICAL CANAL
C0153569|T047||CCS_10|MALIGNANT NEOPLASM OF ENDOCERVICAL CANAL 
C0153569|T047||CCS_10|MALIGNANT NEOPLASM OF CERVICAL CANAL
C0153569|T047||CCS_10|MALIGNANT TUMOR OF ENDOCERVICAL CANAL
C0153569|T047||CCS_10|MALIGNANT TUMOR OF CERVICAL CANAL
C0153569|T047||CCS_10|MALIG NEO ENDOCERVIX
C0153569|T047||CCS_10|CERVICAL NEOPLASM MALIGNANT ENDOCERVIX
C0153569|T047||CCS_10|MALIGNANT NEOPLASM OF ENDOCERVIX 
C0153569|T047||CCS_10|MALIGNANT NEOPLASM OF ENDOCERVIX 
C0153569|T047||CCS_10|MALIGNANT NEOPLASM OF ENDOCERVIX NOS 
C0153569|T047||CCS_10|MALIGNANT NEOPLASM OF ENDOCERVIX NOS
C0153569|T047||CCS_10|MALIGNANT NEOPLASM OF ENDOCERVICAL CANAL 
C0153569|T047||CCS_10|MALIGNANT ENDOCERVICAL NEOPLASM
C0153569|T047||CCS_10|MALIGNANT ENDOCERVICAL TUMOR
C0153569|T047||CCS_10|MALIGNANT ENDOCERVIX NEOPLASM
C0153569|T047||CCS_10|MALIGNANT ENDOCERVIX TUMOR
C0153569|T047||CCS_10|MALIGNANT NEOPLASM OF UTERINE ENDOCERVIX
C0153569|T047||CCS_10|MALIGNANT NEOPLASM OF THE ENDOCERVIX
C0153569|T047||CCS_10|MALIGNANT NEOPLASM OF THE UTERINE ENDOCERVIX
C0153569|T047||CCS_10|MALIGNANT TUMOR OF ENDOCERVIX
C0153569|T047||CCS_10|MALIGNANT TUMOR OF UTERINE ENDOCERVIX
C0153569|T047||CCS_10|MALIGNANT TUMOR OF THE ENDOCERVIX
C0153569|T047||CCS_10|MALIGNANT TUMOR OF THE UTERINE ENDOCERVIX
C0153569|T047||CCS_10|MALIGNANT UTERINE ENDOCERVIX NEOPLASM
C0153569|T047||CCS_10|MALIGNANT UTERINE ENDOCERVIX TUMOR
C0153569|T047||CCS_10|MALIGNANT NEOPLASM OF CERVICAL CANAL NOS
C0153570|T047||CCS_10|MALIGNANT NEOPLASM OF EXOCERVIX
C0153570|T047||CCS_10|MALIGNANT NEOPLASM OF EXOCERVIX 
C0153570|T047||CCS_10|MALIGNANT TUMOR OF EXOCERVIX
C0153570|T047||CCS_10|MALIG NEO EXOCERVIX
C0153570|T047||CCS_10|MALIGNANT NEOPLASM OF EXOCERVIX 
C0153570|T047||CCS_10|CA CERVIX UTERI - EXOCERVIX 
C0153570|T047||CCS_10|CA CERVIX UTERI - EXOCERVIX
C0153570|T047||CCS_10|CANCER OF EXOCERVIX
C0153570|T047||CCS_10|MALIGNANT EXOCERVICAL NEOPLASM
C0153570|T047||CCS_10|MALIGNANT EXOCERVICAL TUMOR
C0153570|T047||CCS_10|MALIGNANT EXOCERVIX NEOPLASM
C0153570|T047||CCS_10|MALIGNANT EXOCERVIX TUMOR
C0153570|T047||CCS_10|MALIGNANT NEOPLASM OF UTERINE EXOCERVIX
C0153570|T047||CCS_10|MALIGNANT NEOPLASM OF THE EXOCERVIX
C0153570|T047||CCS_10|MALIGNANT NEOPLASM OF THE UTERINE EXOCERVIX
C0153570|T047||CCS_10|MALIGNANT TUMOR OF UTERINE EXOCERVIX
C0153570|T047||CCS_10|MALIGNANT TUMOR OF THE EXOCERVIX
C0153570|T047||CCS_10|MALIGNANT TUMOR OF THE UTERINE EXOCERVIX
C0153570|T047||CCS_10|MALIGNANT UTERINE EXOCERVIX NEOPLASM
C0153570|T047||CCS_10|MALIGNANT UTERINE EXOCERVIX TUMOR
C2211948|T047||CCS_10|MALIGNANT SMALL CELL NEOPLASM OF UTERUS
C2211948|T047||CCS_10|UTERINE NEOPLASM MALIGNANT SMALL CELL TYPE
C2211948|T047||CCS_10|MALIGNANT SMALL CELL NEOPLASM OF UTERUS 
C2011421|T047||CCS_10|UTERINE NEOPLASM MALIGNANT GIANT CELL TYPE
C2011421|T047||CCS_10|GIANT CELL TYPE NEOPLASM OF UTERUS 
C2011421|T047||CCS_10|GIANT CELL TYPE NEOPLASM OF UTERUS
C2018702|T047||CCS_10|UTERINE NEOPLASM MALIGNANT SPINDLE CELL TYPE
C2018702|T047||CCS_10|SPINDLE CELL TYPE NEOPLASM OF UTERUS 
C2018702|T047||CCS_10|SPINDLE CELL TYPE NEOPLASM OF UTERUS
C2075662|T047||CCS_10|CLEAR CELL TYPE NEOPLASM OF UTERUS
C2075662|T047||CCS_10|CLEAR CELL TYPE NEOPLASM OF UTERUS 
C2075662|T047||CCS_10|UTERINE NEOPLASM MALIGNANT CLEAR CELL TYPE
C0848454|T047||CCS_10|UTERINE CARCINOMA
C0848454|T047||CCS_10|CARCINOMA OF UTERUS 
C0848454|T047||CCS_10|CARCINOMA OF UTERUS
C0848454|T047||CCS_10|CARCINOMA;UTERUS
C0848454|T047||CCS_10|CARCINOMA OF THE UTERUS
C2211972|T047||CCS_10|MYOSARCOMA OF UTERUS 
C2211972|T047||CCS_10|MYOSARCOMA OF UTERUS
C2211981|T047||CCS_10|FIBROSARCOMA OF UTERUS 
C2211981|T047||CCS_10|FIBROSARCOMA OF UTERUS
C2211991|T047||CCS_10|MALIGNANT MESENCHYMOMA OF UTERUS 
C2211991|T047||CCS_10|MALIGNANT MESENCHYMOMA OF UTERUS
C2211992|T047||CCS_10|MALIGNANT MESONEPHROMA OF UTERUS 
C2211992|T047||CCS_10|MALIGNANT MESONEPHROMA OF UTERUS
C2211993|T047||CCS_10|MULLERIAN MIXED TUMOR OF UTERUS
C2211993|T047||CCS_10|MULLERIAN MIXED TUMOR OF UTERUS 
C1704376|T047||CCS_10|UTERINE CORPUS CARCINOSARCOMA
C1704376|T047||CCS_10|MALIGNANT MESODERMAL MIXED TUMOR OF UTERUS
C1704376|T047||CCS_10|MALIGNANT MESODERMAL MIXED TUMOR OF UTERUS 
C1704376|T047||CCS_10|MIXED MÜLLERIAN SARCOMA OF THE UTERUS
C1704376|T047||CCS_10|MIXED MÜLLERIAN SARCOMA OF UTERUS
C1704376|T047||CCS_10|UTERINE CORPUS MALIGNANT MIXED MESODERMAL (MÜLLERIAN) TUMOR
C1704376|T047||CCS_10|UTERINE CORPUS MALIGNANT MIXED MÜLLERIAN NEOPLASM
C1704376|T047||CCS_10|UTERINE MIXED MÜLLERIAN SARCOMA
C1704376|T047||CCS_10|UTERINE CORPUS MALIGNANT MIXED MÜLLERIAN TUMOR
C1704376|T047||CCS_10|CORPUS UTERI MALIGNANT MIXED MESODERMAL TUMOR
C1704376|T047||CCS_10|MALIGNANT MIXED MESODERMAL NEOPLASM OF UTERINE BODY
C1704376|T047||CCS_10|MALIGNANT MIXED MESODERMAL NEOPLASM OF UTERINE CORPUS
C1704376|T047||CCS_10|MALIGNANT MIXED MESODERMAL NEOPLASM OF UTERUS
C1704376|T047||CCS_10|MALIGNANT MIXED MESODERMAL NEOPLASM OF THE UTERINE BODY
C1704376|T047||CCS_10|MALIGNANT MIXED MESODERMAL NEOPLASM OF THE UTERINE CORPUS
C1704376|T047||CCS_10|MALIGNANT MIXED MESODERMAL NEOPLASM OF THE UTERUS
C1704376|T047||CCS_10|MALIGNANT MIXED MESODERMAL TUMOR OF UTERINE BODY
C1704376|T047||CCS_10|MALIGNANT MIXED MESODERMAL TUMOR OF UTERINE CORPUS
C1704376|T047||CCS_10|MALIGNANT MIXED MESODERMAL TUMOR OF UTERUS
C1704376|T047||CCS_10|MALIGNANT MIXED MESODERMAL TUMOR OF THE UTERINE BODY
C1704376|T047||CCS_10|MALIGNANT MIXED MESODERMAL TUMOR OF THE UTERINE CORPUS
C1704376|T047||CCS_10|MALIGNANT MIXED MESODERMAL TUMOR OF THE UTERUS
C1704376|T047||CCS_10|UTERINE BODY CARCINOSARCOMA
C1704376|T047||CCS_10|UTERINE BODY MALIGNANT MIXED MESODERMAL NEOPLASM
C1704376|T047||CCS_10|UTERINE BODY MALIGNANT MIXED MESODERMAL TUMOR
C1704376|T047||CCS_10|UTERINE CARCINOSARCOMA
C1704376|T047||CCS_10|UTERINE CORPUS MALIGNANT MIXED MESODERMAL NEOPLASM
C1704376|T047||CCS_10|UTERINE CORPUS MALIGNANT MIXED MESODERMAL TUMOR
C1704376|T047||CCS_10|UTERINE MALIGNANT MIXED MESODERMAL NEOPLASM
C1704376|T047||CCS_10|UTERINE MALIGNANT MIXED MESODERMAL TUMOR
C1704376|T047||CCS_10|CARCINOSARCOMA OF CORPUS UTERI
C1704376|T047||CCS_10|CARCINOSARCOMA OF UTERINE BODY
C1704376|T047||CCS_10|CARCINOSARCOMA OF UTERINE CORPUS
C1704376|T047||CCS_10|CARCINOSARCOMA OF UTERUS
C1704376|T047||CCS_10|CARCINOSARCOMA OF THE CORPUS UTERI
C1704376|T047||CCS_10|CARCINOSARCOMA OF THE UTERINE BODY
C1704376|T047||CCS_10|CARCINOSARCOMA OF THE UTERINE CORPUS
C1704376|T047||CCS_10|CARCINOSARCOMA OF THE UTERUS
C2211995|T047||CCS_10|MALIGNANT LYMPHOMA OF UTERUS
C2211995|T047||CCS_10|MALIGNANT LYMPHOMA OF UTERUS 
C2211998|T047||CCS_10|MALIGNANT PLASMACYTOMA OF UTERUS 
C2211998|T047||CCS_10|MALIGNANT PLASMACYTOMA OF UTERUS
C2212000|T047||CCS_10|MALIGNANT MASTOCYTOSIS OF UTERUS
C2212000|T047||CCS_10|MALIGNANT MASTOCYTOSIS OF UTERUS 
C2217776|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGING 
C2217776|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGING
C2217776|T047||CCS_10|UTERINE CANCER STAGING
C2217776|T047||CCS_10|MALIGNANT TUMOR OF UTERUS STAGING
C0496821|T047||CCS_10|MALIGNANT NEOPLASM OF FUNDUS UTERI
C0496821|T047||CCS_10|MALIGNANT NEOPLASM OF THE FUNDUS UTERI
C0496821|T047||CCS_10|MALIGNANT NEOPLASM OF FUNDUS OF UTERUS
C0496821|T047||CCS_10|MALIGNANT NEOPLASM OF FUNDUS OF UTERUS 
C0496821|T047||CCS_10|MALIGNANT TUMOR OF FUNDUS OF UTERUS
C0496821|T047||CCS_10|MALIGNANT NEOPLASM OF FUNDUS OF CORPUS UTERI
C0496821|T047||CCS_10|MALIGNANT NEOPLASM OF FUNDUS OF CORPUS UTERI 
C0496818|T047||CCS_10|MALIGNANT NEOPLASM OF ISTHMUS UTERI
C0496818|T047||CCS_10|MALIGNANT NEOPLASM OF ISTHMUS OF UTERUS
C0496818|T047||CCS_10|MALIGNANT NEOPLASM OF ISTHMUS OF UTERUS 
C0496818|T047||CCS_10|MALIGNANT TUMOR OF ISTHMUS OF UTERUS
C0496818|T047||CCS_10|MALIGNANT NEOPLASM OF ISTHMUS OF UTERINE BODY NOS 
C0496818|T047||CCS_10|MALIGNANT NEOPLASM OF ISTHMUS OF UTERINE BODY NOS
C0496818|T047||CCS_10|MALIGNANT NEOPLASM OF ISTHMUS OF UTERINE BODY
C0496818|T047||CCS_10|MALIGNANT NEOPLASM OF ISTHMUS OF UTERINE BODY 
C2103110|T047||CCS_10|ADENOSARCOMA OF UTERUS 
C2103110|T047||CCS_10|ADENOSARCOMA OF UTERUS
C2103110|T047||CCS_10|UTERINE ADENOSARCOMA
C2103110|T047||CCS_10|MULLERIAN ADENOSARCOMA OF THE UTERUS
C2103110|T047||CCS_10|ADENOSARCOMA OF THE UTERUS
C2103110|T047||CCS_10|ADENOSARCOMA OF UTERUS 
C2006983|T047||CCS_10|CARCINOFIBROMA OF UTERUS
C2006983|T047||CCS_10|CARCINOFIBROMA OF UTERUS 
C0280630|T047||CCS_10|UTERINE CARCINOSARCOMA
C0280630|T047||CCS_10|CARCINOSARCOMA OF THE UTERUS
C0280630|T047||CCS_10|UTERINE MALIGNANT MIXED MESODERMAL (MULLERIAN) TUMOR
C0280630|T047||CCS_10|MALIGNANT MIXED MESODERMAL (MULLERIAN) TUMOR OF THE UTERUS
C0280630|T047||CCS_10|CARCINOSARCOMA OF UTERUS 
C0280630|T047||CCS_10|CARCINOSARCOMA OF UTERUS
C0280630|T047||CCS_10|CARCINOSARCOMA OF UTERUS 
C0280630|T047||CCS_10|CARCINOSARCOMA UTERUS
C0280630|T047||CCS_10|CARCINO-SARCOMA UTERUS
C0280630|T047||CCS_10|CARCINOSARCOMA, UTERINE
C0280630|T047||CCS_10|MIXED MULLERIAN SARCOMA, UTERINE
C0280630|T047||CCS_10|UTERINE MIXED MULLERIAN SARCOMA
C0280630|T047||CCS_10|MULLERIAN SARCOMA, UTERINE MIXED
C0280630|T047||CCS_10|MULLERIAN TUMOR, UTERINE MIXED
C0153584|T047||CCS_10|MALIGNANT NEOPLASM OF UTERINE ADNEXA
C0153584|T047||CCS_10|MALIGNANT NEOPLASM OF UTERINE ADNEXA, UNSPECIFIED
C0153584|T047||CCS_10|UTERINE ADNEXA, UNSPECIFIED
C0153584|T047||CCS_10|MALIGNANT NEOPLASM OF UTERINE ADNEXA 
C0153584|T047||CCS_10|MALIGNANT NEOPLASM OF UTERINE ADNEXA 
C0153584|T047||CCS_10|MALIGNANT TUMOR OF UTERINE ADNEXA
C0153584|T047||CCS_10|MAL NEO ADNEXA NOS
C0153584|T047||CCS_10|MALIGNANT NEOPLASM OF UTERINE ADNEXA, UNSPECIFIED SITE
C0153584|T047||CCS_10|[X]MALIGNANT NEOPLASM OF UTERINE ADNEXA, UNSPECIFIED 
C0153584|T047||CCS_10|MALIGNANT NEOPLASM OF UTERINE ADNEXA NOS 
C0153584|T047||CCS_10|MALIGNANT NEOPLASM OF UTERINE ADNEXA NOS
C0153584|T047||CCS_10|[X]MALIGNANT NEOPLASM OF UTERINE ADNEXA, UNSPECIFIED
C0153584|T047||CCS_10|MALIGNANT NEOPLASM OF UTERINE ADNEXA, NOS
C2960452|T047||CCS_10|MALIGNANT EPITHELIAL NEOPLASM OF UTERUS 
C2960452|T047||CCS_10|MALIGNANT EPITHELIAL NEOPLASM OF UTERUS
C2960452|T047||CCS_10|CARCINOMA OF UTERUS
C0280631|T047||CCS_10|UTERINE LEIOMYOSARCOMA
C0280631|T047||CCS_10|LEIOMYOSARCOMA OF UTERUS
C0280631|T047||CCS_10|LEIOMYOSARCOMA OF UTERUS 
C0280631|T047||CCS_10|LEIOMYOSARCOMA OF UTERUS 
C0280631|T047||CCS_10|LEIOMYOSARCOMA OF THE UTERUS
C0280631|T047||CCS_10|LEIOMYOSARCOMA - UTERUS
C0280631|T047||CCS_10|LEIOMYOSARCOMA, UTERINE
C0280631|T047||CCS_10|CORPUS UTERI LEIOMYOSARCOMA
C0280631|T047||CCS_10|LEIOMYOSARCOMA OF BODY OF UTERUS
C0280631|T047||CCS_10|LEIOMYOSARCOMA OF CORPUS UTERI
C0280631|T047||CCS_10|LEIOMYOSARCOMA OF UTERINE BODY
C0280631|T047||CCS_10|LEIOMYOSARCOMA OF UTERINE CORPUS
C0280631|T047||CCS_10|LEIOMYOSARCOMA OF THE BODY OF UTERUS
C0280631|T047||CCS_10|LEIOMYOSARCOMA OF THE CORPUS UTERI
C0280631|T047||CCS_10|LEIOMYOSARCOMA OF THE UTERINE BODY
C0280631|T047||CCS_10|LEIOMYOSARCOMA OF THE UTERINE CORPUS
C0280631|T047||CCS_10|UTERINE BODY LEIOMYOSARCOMA
C0280631|T047||CCS_10|UTERINE CORPUS LEIOMYOSARCOMA
C0280631|T047||CCS_10|BODY OF UTERUS LEIOMYOSARCOMA
C3164916|T047||CCS_10|MALIGNANT MIXED MULLERIAN TUMOR OF UTERUS
C3164916|T047||CCS_10|MALIGNANT MIXED MULLERIAN TUMOUR OF UTERUS
C3164916|T047||CCS_10|MALIGNANT MIXED MULLERIAN TUMOR OF UTERUS 
C0153572|T047||CCS_10|MALIGNANT NEOPLASM OF PLACENTA
C0153572|T047||CCS_10|MALIGNANT NEOPLASM OF PLACENTA 
C0153572|T047||CCS_10|MALIGNANT TUMOR OF PLACENTA
C0153572|T047||CCS_10|MALIGNANT NEOPL PLACENTA
C0153572|T047||CCS_10|PLACENTAL CANCER
C0153572|T047||CCS_10|MALIGNANT NEOPLASM OF PLACENTA 
C0153572|T047||CCS_10|CANCER OF PLACENTA
C0153572|T047||CCS_10|DECIDUOMA, MALIGNANT
C0153572|T047||CCS_10|MALIGNANT PLACENTAL NEOPLASM
C0153572|T047||CCS_10|MALIGNANT TUMOR OF THE PLACENTA
C0153572|T047||CCS_10|MALIGNANT NEOPLASM OF THE PLACENTA
C0153572|T047||CCS_10|MALIGNANT PLACENTAL TUMOR
C0153572|T047||CCS_10|MALIGNANT PLACENTA NEOPLASM
C0153572|T047||CCS_10|MALIGNANT PLACENTA TUMOR
C0153572|T047||CCS_10|NEOPLASM MALIG;PLACENTA
C0153572|T047||CCS_10|MALIGNANT NEOSPLASM OF THE PLACENTA
C2211985|T047||CCS_10|ADULT TYPE PLEOMORPHIC RHABDOMYOSARCOMA OF UTERUS 
C2211985|T047||CCS_10|UTERINE RHABDOMYOSARCOMA PLEOMORPHIC, ADULT TYPE
C2211985|T047||CCS_10|ADULT TYPE PLEOMORPHIC RHABDOMYOSARCOMA OF UTERUS
C3468483|T047||CCS_10|ENDOMETRIAL CANCER SUSCEPTIBILITY 
C3468483|T047||CCS_10|ENDOMETRIAL CANCER SUSCEPTIBILITY
C0007103|T047||CCS_10|MALIGNANT NEOPLASM OF ENDOMETRIUM
C0007103|T047||CCS_10|ENDOMETRIAL NEOPLASMS MALIGNANT
C0007103|T047||CCS_10|MALIGNANT NEOPLASM OF ENDOMETRIUM 
C0007103|T047||CCS_10|UTERINE NEOPLASM, MALIGNANT - OF THE ENDOMETRIUM
C0007103|T047||CCS_10|ENDOMETRIAL CANCER
C0007103|T047||CCS_10|ENDOMETRIAL NEOPLASM MALIGNANT
C0007103|T047||CCS_10|MALIGNANT ENDOMETRIAL NEOPLASM
C0007103|T047||CCS_10|MALIGNANT NEOPLASM OF THE ENDOMETRIUM
C0007103|T047||CCS_10|NEOPLASM MALIG;ENDOMETRIAL
C1879358|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF ENDOMETRIUM
C1879358|T047||CCS_10|MALIGNANT NEOPLASM OF ENDOMETRIUM
C1879358|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF ENDOMETRIUM 
C1879358|T047||CCS_10|UTERINE NEOPLASM, MALIGNANT - OF THE ENDOMETRIUM PRIMARY
C1879358|T047||CCS_10|CANCER OF ENDOMETRIUM
C1879358|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF ENDOMETRIUM 
C0008493|T047||CCS_10|MALIGNANT HYDATIDIFORM MOLE
C0008493|T047||CCS_10|CHORIOADENOMAS
C0008493|T047||CCS_10|HYDATIDIFORM MOLE, INVASIVE
C0008493|T047||CCS_10|HYDATIDIFORM MOLES, INVASIVE
C0008493|T047||CCS_10|INVASIVE HYDATIDIFORM MOLES
C0008493|T047||CCS_10|INVASIVE MOLES
C0008493|T047||CCS_10|MOLES, INVASIVE
C0008493|T047||CCS_10|MOLES, INVASIVE HYDATIDIFORM
C0008493|T047||CCS_10|INVASIVE HYDATIDIFORM MOLE
C0008493|T047||CCS_10|MOLE, INVASIVE
C0008493|T047||CCS_10|MOLE, INVASIVE HYDATIDIFORM
C0008493|T047||CCS_10|INVASIVE HYDATIDIFORM MOLE 
C0008493|T047||CCS_10|MOLAR PREGNANCY, INVASIVE (NON-METASTATIC GTD)
C0008493|T047||CCS_10|CHORIOADENOMA DESTRUENS
C0008493|T047||CCS_10|CHORIOADENOMA
C0008493|T047||CCS_10|HYDATIDIFORM MOLE, INVASIVE [DISEASE/FINDING]
C0008493|T047||CCS_10|INVASIVE MOLE
C0008493|T047||CCS_10|MOLE;MALIGNANT
C0008493|T047||CCS_10|MOLAR PREGNANCY WITH INVASIVE HYDATIDIFORM MOLE
C0008493|T047||CCS_10|MALIGNANT HYDATIDIFORM MOLE 
C0008493|T047||CCS_10|MOLAR PREGNANCY WITH MALIGNANT HYDATIDIFORM MOLE
C0008493|T047||CCS_10|MOLAR PREGNANCY WITH CHORIOADENOMA DESTRUENS
C0008493|T047||CCS_10|INVASIVE MOLE - PLACENTA
C0008493|T047||CCS_10|MOLAR PREGNANCY WITH CHORIOADENOMA
C0008493|T047||CCS_10|IM - INVASIVE MOLE
C0008493|T047||CCS_10|CHORIADENOMA (DESTRUENS)
C0008493|T047||CCS_10|MOLAR PREGNANCY WITH INVASIVE MOLE
C0008493|T047||CCS_10|MOLAR PREGNANCY WITH INVASIVE HYDATIDIFORM MOLE 
C0008493|T047||CCS_10|[M]CHORIOADENOMA DESTRUENS
C0008493|T047||CCS_10|[M]INVASIVE HYDATIDIFORM MOLE
C0008493|T047||CCS_10|[M]CHORIOADENOMA
C0008493|T047||CCS_10|HYDATIDIFORM MOLE MALIGNANT
C0008493|T047||CCS_10|INVASIVE HYDATIDIFORM MOLE (MORPHOLOGIC ABNORMALITY)
C0008493|T047||CCS_10|GTT, INVASIVE MOLE
C0008493|T047||CCS_10|GESTATIONAL TROPHOBLASTIC TUMOR, INVASIVE MOLE
C0008493|T047||CCS_10|DESTRUCTIVE; MOLE
C0008493|T047||CCS_10|HYDATIDIFORM MOLE; INVASIVE
C0008493|T047||CCS_10|HYDATIDIFORM MOLE; MALIGNANT
C0008493|T047||CCS_10|INVASIVE; HYDATIDIFORM MOLE
C0008493|T047||CCS_10|INVASIVE; MOLE
C0008493|T047||CCS_10|MALIGNANT; HYDATIDIFORM MOLE
C0008493|T047||CCS_10|MALIGNANT; MOLE, HYDATIDIFORM
C0008493|T047||CCS_10|MOLE; HYDATIDIFORM, INVASIVE
C0008493|T047||CCS_10|MOLE; HYDATIDIFORM, MALIGNANT
C0008493|T047||CCS_10|MOLE; INVASIVE
C0008493|T047||CCS_10|MOLE; MALIGNANT, HYDATIDIFORM MOLE
C0008493|T047||CCS_10|INVASIVE MOLE, NOS
C0008493|T047||CCS_10|INVASIVE GESTATIONAL TROPHOBLASTIC NEOPLASM
C0008493|T047||CCS_10|MALIGNANT HYDATID MOLE
C0008493|T047||CCS_10|INVASIVE HYDATIDIFORM MOLE 
C0008493|T047||CCS_10|MALIGNANT MOLE
C1299275|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF BODY OF UTERUS
C1299275|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF BODY OF UTERUS 
C1299275|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF CORPUS UTERI
C1299275|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF CORPUS UTERI 
C1299275|T047||CCS_10|UTERINE NEOPLASM, MALIGNANT - CORPUS UTERI PRIMARY
C2703078|T047||CCS_10|MALIGNANT NEOPLASM OF PLACENTA
C2703078|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF PLACENTA
C2703078|T047||CCS_10|PLACENTAL NEOPLASM MALIGNANT PRIMARY
C2703078|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF PLACENTA 
C2703078|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF PLACENTA 
C1263776|T047||CCS_10|OVERLAPPING MALIGNANT NEOPLASM OF BODY OF UTERUS 
C1263776|T047||CCS_10|OVERLAPPING MALIGNANT NEOPLASM OF BODY OF UTERUS
C1263776|T047||CCS_10|OVERLAPPING MALIGNANT NEOPLASM OF CORPUS UTERI
C1306053|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF ISTHMUS OF UTERUS 
C1306053|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF ISTHMUS OF UTERUS
C1314886|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF PARAMETRIUM 
C1314886|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF PARAMETRIUM
C0007847|T047||CCS_10|MALIGNANT NEOPLASM OF CERVIX UTERI
C0007847|T047||CCS_10|MALIGNANT NEOPLASM OF CERVIX UTERI, UNSPECIFIED
C0007847|T047||CCS_10|MALIGNANT NEOPLASM OF UTERINE CERVIX
C0007847|T047||CCS_10|CANCER OF CERVIX
C0007847|T047||CCS_10|MALIGNANT NEOPLASM OF CERVIX
C0007847|T047||CCS_10|CERVICAL CANCER
C0007847|T047||CCS_10|MALIGNANT NEOPLASM OF CERVIX 
C0007847|T047||CCS_10|MALIGNANT CERVICAL NEOPLASM
C0007847|T047||CCS_10|MALIGNANT TUMOR OF CERVIX
C0007847|T047||CCS_10|MAL NEO CERVIX UTERI NOS
C0007847|T047||CCS_10|CERVIX NEOPLASMS MALIGNANT
C0007847|T047||CCS_10|MALIGNANT NEOPLASM OF CERVIX UTERI, UNSPECIFIED SITE
C0007847|T047||CCS_10|MALIGNANT NEOPLASM OF CERVIX UTERI 
C0007847|T047||CCS_10|CERVICAL NEOPLASM MALIGNANT CERVIX UTERI
C0007847|T047||CCS_10|MALIGNANT TUMOUR OF CERVIX 
C0007847|T047||CCS_10|MALIGNANT NEOPLASM OF CERVIX UTERI NOS 
C0007847|T047||CCS_10|MALIGNANT TUMOUR OF CERVIX
C0007847|T047||CCS_10|MALIGNANT NEOPLASM OF CERVIX UTERI NOS
C0007847|T047||CCS_10|CANCER OF THE UTERINE CERVIX
C0007847|T047||CCS_10|MALIGNANT TUMOR OF CERVIX 
C0007847|T047||CCS_10|MALIGNANT CERVICAL TUMOR
C0007847|T047||CCS_10|MALIGNANT CERVIX NEOPLASM
C0007847|T047||CCS_10|MALIGNANT CERVIX TUMOR
C0007847|T047||CCS_10|MALIGNANT CERVIX UTERI NEOPLASM
C0007847|T047||CCS_10|MALIGNANT CERVIX UTERI TUMOR
C0007847|T047||CCS_10|MALIGNANT NEOPLASM OF THE CERVIX UTERI
C0007847|T047||CCS_10|MALIGNANT NEOPLASM OF THE CERVIX
C0007847|T047||CCS_10|MALIGNANT NEOPLASM OF THE UTERINE CERVIX
C0007847|T047||CCS_10|MALIGNANT TUMOR OF CERVIX UTERI
C0007847|T047||CCS_10|MALIGNANT TUMOR OF UTERINE CERVIX
C0007847|T047||CCS_10|MALIGNANT TUMOR OF THE CERVIX UTERI
C0007847|T047||CCS_10|MALIGNANT TUMOR OF THE CERVIX
C0007847|T047||CCS_10|MALIGNANT TUMOR OF THE UTERINE CERVIX
C0007847|T047||CCS_10|MALIGNANT UTERINE CERVIX NEOPLASM
C0007847|T047||CCS_10|MALIGNANT UTERINE CERVIX TUMOR
C0007847|T047||CCS_10|NEOPLASM MALIG;CERVIX
C0007847|T047||CCS_10|MALIGNANT NEOSPLASM OF THE CERVIX
C0346995|T047||CCS_10|METASTASIS OF MALIGNANT NEOPLASM TO THE UTERUS
C0346995|T047||CCS_10|METASTASIS OF MALIGNANT NEOPLASM TO UTERUS 
C0346995|T047||CCS_10|METASTASIS OF MALIGNANT NEOPLASM TO UTERUS
C0346995|T047||CCS_10|METASTASES TO UTERUS
C0346995|T047||CCS_10|UTERINE NEOPLASM MALIGNANT SECONDARY
C0346995|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF UTERUS
C0346995|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF UTERUS 
C0346995|T047||CCS_10|CANCER METASTATIC TO UTERUS
C0346995|T047||CCS_10|METASTASIS TO UTERUS
C0346995|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO UTERUS
C0346995|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF UTERUS 
C0346995|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO UTERUS, NOS
C0346995|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF UTERUS, NOS
C1282495|T047||CCS_10|METASTASIS FROM MALIGNANT NEOPLASM OF UTERUS
C1282495|T047||CCS_10|METASTASIS FROM MALIGNANT NEOPLASM OF UTERUS 
C1282495|T047||CCS_10|METASTASIS FROM MALIGNANT TUMOR OF UTERUS 
C1282495|T047||CCS_10|METASTASIS FROM MALIGNANT TUMOR OF UTERUS
C1282495|T047||CCS_10|METASTASIS FROM MALIGNANT TUMOUR OF UTERUS
C3838720|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF UTERUS 
C3838720|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF UTERUS
C1336899|T047||CCS_10|HEMANGIOSARCOMA OF UTERUS
C1336899|T047||CCS_10|HEMANGIOSARCOMA OF THE UTERUS
C1336899|T047||CCS_10|ANGIOSARCOMA OF UTERUS
C1336899|T047||CCS_10|ANGIOSARCOMA OF THE UTERUS
C1336899|T047||CCS_10|UTERINE ANGIOSARCOMA
C1336899|T047||CCS_10|UTERINE HEMANGIOSARCOMA
C2217769|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGE IIA
C2217769|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGE IIA 
C2217769|T047||CCS_10|MALIGNANT TUMOR OF UTERUS STAGE IIA
C2217769|T047||CCS_10|UTERINE CANCER STAGE IIA
C2111694|T047||CCS_10|LARGE CELL CARCINOMA OF UTERUS WITH RHABDOID PHENOTYPE
C2111694|T047||CCS_10|LARGE CELL CARCINOMA OF UTERUS WITH RHABDOID PHENOTYPE 
C2111694|T047||CCS_10|UTERINE MALIGNANT CARCINOMA LARGE CELL WITH RHABDOID PHENOTYPE
C2018413|T047||CCS_10|SPINDLE CELL CARCINOMA OF UTERUS
C2018413|T047||CCS_10|SPINDLE CELL CARCINOMA OF UTERUS 
C2033322|T047||CCS_10|PAPILLARY SQUAMOUS CELL CARCINOMA OF UTERUS
C2033322|T047||CCS_10|PAPILLARY SQUAMOUS CELL CARCINOMA OF UTERUS 
C2211953|T047||CCS_10|NONKERATINIZING SQUAMOUS CELL CARCINOMA OF UTERUS
C2211953|T047||CCS_10|NONKERATINIZING SQUAMOUS CELL CARCINOMA OF UTERUS 
C2211953|T047||CCS_10|UTERINE MALIGNANT CARCINOMA SQUAMOUS CELL SMALL CELL NONKERATINIZING
C2211954|T047||CCS_10|ADENOID SQUAMOUS CELL CARCINOMA OF UTERUS
C2211954|T047||CCS_10|ADENOID SQUAMOUS CELL CARCINOMA OF UTERUS 
C2211956|T047||CCS_10|BASALOID SQUAMOUS CELL CARCINOMA OF UTERUS 
C2211956|T047||CCS_10|BASALOID SQUAMOUS CELL CARCINOMA OF UTERUS
C2075854|T047||CCS_10|CLOACOGENIC CARCINOMA OF UTERUS
C2075854|T047||CCS_10|CLOACOGENIC CARCINOMA OF UTERUS 
C2211979|T047||CCS_10|MAST CELL SARCOMA OF UTERUS
C2211979|T047||CCS_10|MAST CELL SARCOMA OF UTERUS 
C2188881|T047||CCS_10|LYMPHOCYTE-RICH NODULAR HODGKIN'S LYMPHOMA OF UTERUS 
C2188881|T047||CCS_10|LYMPHOCYTE-RICH NODULAR HODGKIN'S LYMPHOMA OF UTERUS
C2188883|T047||CCS_10|NODULAR SCLEROSING HODGKIN'S LYMPHOMA IN CELLULAR PHASE OF UTERUS 
C2188883|T047||CCS_10|NODULAR SCLEROSING HODGKIN'S LYMPHOMA IN CELLULAR PHASE OF UTERUS
C2188885|T047||CCS_10|GRADE 2 NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF UTERUS
C2188885|T047||CCS_10|GRADE 2 NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF UTERUS 
C2188897|T047||CCS_10|LYMPHOPLASMACYTIC LYMPHOMA OF UTERUS 
C2188897|T047||CCS_10|LYMPHOPLASMACYTIC LYMPHOMA OF UTERUS
C2188899|T047||CCS_10|MARGINAL ZONE B-CELL LYMPHOMA OF UTERUS
C2188899|T047||CCS_10|MARGINAL ZONE B-CELL LYMPHOMA OF UTERUS 
C2188900|T047||CCS_10|MATURE T-CELL LYMPHOMA OF UTERUS 
C2188900|T047||CCS_10|MATURE T-CELL LYMPHOMA OF UTERUS
C2188903|T047||CCS_10|NK/T-CELL LYMPHOMA OF UTERUS
C2188903|T047||CCS_10|NK/T-CELL LYMPHOMA OF UTERUS 
C2212001|T047||CCS_10|SEZARY SYNDROME OF UTERUS
C2212001|T047||CCS_10|SEZARY SYNDROME OF UTERUS 
C2111693|T047||CCS_10|LARGE CELL CARCINOMA OF UTERUS 
C2111693|T047||CCS_10|LARGE CELL CARCINOMA OF UTERUS
C2012125|T047||CCS_10|GLASSY CELL CARCINOMA OF UTERUS 
C2012125|T047||CCS_10|GLASSY CELL CARCINOMA OF UTERUS
C2033341|T047||CCS_10|PAPILLARY TRANSITIONAL CELL CARCINOMA OF UTERUS 
C2033341|T047||CCS_10|PAPILLARY TRANSITIONAL CELL CARCINOMA OF UTERUS
C2011238|T047||CCS_10|GIANT CELL AND SPINDLE CELL CARCINOMA OF UTERUS
C2011238|T047||CCS_10|GIANT CELL AND SPINDLE CELL CARCINOMA OF UTERUS 
C2007043|T047||CCS_10|CARCINOMA OF UTERUS WITH OSTEOCLAST-LIKE GIANT CELLS
C2007043|T047||CCS_10|CARCINOMA OF UTERUS WITH OSTEOCLAST-LIKE GIANT CELLS 
C2007043|T047||CCS_10|UTERINE CARCINOMA WITH OSTEOCLAST-LIKE GIANT CELLS
C0279764|T047||CCS_10|PAPILLARY CARCINOMA OF UTERUS
C0279764|T047||CCS_10|PAPILLARY CARCINOMA OF UTERUS 
C0279764|T047||CCS_10|ENDOMETRIAL PAPILLARY CARCINOMA
C0279764|T047||CCS_10|CARCINOMA OF THE UTERUS, PAPILLARY
C0279764|T047||CCS_10|CARCINOMA, PAPILLARY, ENDOMETRIAL
C0279764|T047||CCS_10|PAPILLARY CARCINOMA OF THE UTERUS
C0279764|T047||CCS_10|UTERINE CANCER, PAPILLARY CARCINOMA
C0279764|T047||CCS_10|UTERINE CORPUS CANCER, PAPILLARY CARCINOMA
C0279764|T047||CCS_10|UTERUS CANCER, PAPILLARY CARCINOMA
C2019462|T047||CCS_10|UTERINE MALIGNANT CARCINOMA SQUAMOUS CELL WITH HORN FORMATION
C2019462|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF UTERUS WITH HORN FORMATION 
C2019462|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF UTERUS WITH HORN FORMATION
C2019462|T047||CCS_10|SQUAMOUS CELL CARCINOMA WITH HORN FORMATION OF UTERUS
C2075582|T047||CCS_10|CLEAR CELL SQUAMOUS CELL CARCINOMA OF UTERUS
C2075582|T047||CCS_10|CLEAR CELL SQUAMOUS CELL CARCINOMA OF UTERUS 
C2211957|T047||CCS_10|SCHNEIDERIAN CARCINOMA OF UTERUS
C2211957|T047||CCS_10|SCHNEIDERIAN CARCINOMA OF UTERUS 
C2211957|T047||CCS_10|UTERINE MALIGNANT CARCINOMA SCHNEIDERIAN
C2211958|T047||CCS_10|BASALOID CARCINOMA OF UTERUS
C2211958|T047||CCS_10|BASALOID CARCINOMA OF UTERUS 
C2188891|T047||CCS_10|GRADE 1 FOLLICULAR LYMPHOMA OF UTERUS 
C2188891|T047||CCS_10|GRADE 1 FOLLICULAR LYMPHOMA OF UTERUS
C2188892|T047||CCS_10|GRADE 2 FOLLICULAR LYMPHOMA OF UTERUS
C2188892|T047||CCS_10|GRADE 2 FOLLICULAR LYMPHOMA OF UTERUS 
C2217767|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGE IB
C2217767|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGE IB 
C2217767|T047||CCS_10|MALIGNANT TUMOR OF UTERUS STAGE IB
C2217767|T047||CCS_10|UTERINE CANCER STAGE IB
C2217775|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGE IVB
C2217775|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGE IVB 
C2217775|T047||CCS_10|MALIGNANT TUMOR OF UTERUS STAGE IVB
C2217775|T047||CCS_10|UTERINE CANCER STAGE IVB
C2111825|T047||CCS_10|POLYGONAL CELL CARCINOMA OF UTERUS 
C2111825|T047||CCS_10|POLYGONAL CELL CARCINOMA OF UTERUS
C2018579|T047||CCS_10|SPINDLE CELL SQUAMOUS CELL CARCINOMA OF UTERUS 
C2018579|T047||CCS_10|SPINDLE CELL SQUAMOUS CELL CARCINOMA OF UTERUS
C2211960|T047||CCS_10|MUCOEPIDERMOID CARCINOMA OF UTERUS
C2211960|T047||CCS_10|MUCOEPIDERMOID CARCINOMA OF UTERUS 
C2017462|T047||CCS_10|SOLID CARCINOMA OF UTERUS 
C2017462|T047||CCS_10|SOLID CARCINOMA OF UTERUS
C2211984|T047||CCS_10|MALIGNANT SOLITARY FIBROUS TUMOR OF UTERUS 
C2211984|T047||CCS_10|MALIGNANT SOLITARY FIBROUS TUMOR OF UTERUS
C2188898|T047||CCS_10|MANTLE CELL LYMPHOMA OF UTERUS 
C2188898|T047||CCS_10|MANTLE CELL LYMPHOMA OF UTERUS
C2188895|T047||CCS_10|LARGE B-CELL DIFFUSE LYMPHOMA OF UTERUS
C2188895|T047||CCS_10|LARGE B-CELL DIFFUSE LYMPHOMA OF UTERUS 
C2113667|T047||CCS_10|PRECURSOR B-CELL LYMPHOBLASTIC LYMPHOMA OF UTERUS 
C2113667|T047||CCS_10|PRECURSOR B-CELL LYMPHOBLASTIC LYMPHOMA OF UTERUS
C2113807|T047||CCS_10|PRECURSOR T-CELL LYMPHOBLASTIC LYMPHOMA OF UTERUS 
C2113807|T047||CCS_10|PRECURSOR T-CELL LYMPHOBLASTIC LYMPHOMA OF UTERUS
C2103109|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF UTERUS 
C2103109|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF UTERUS
C2217766|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGE IA
C2217766|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGE IA 
C2217766|T047||CCS_10|MALIGNANT TUMOR OF UTERUS STAGE IA
C2217766|T047||CCS_10|UTERINE CANCER STAGE IA
C2111760|T047||CCS_10|LARGE CELL NEUROENDOCRINE CARCINOMA OF UTERUS
C2111760|T047||CCS_10|LARGE CELL NEUROENDOCRINE CARCINOMA OF UTERUS 
C2211950|T047||CCS_10|ANAPLASTIC CARCINOMA OF UTERUS
C2211950|T047||CCS_10|ANAPLASTIC CARCINOMA OF UTERUS 
C2211952|T047||CCS_10|MICROPAPILLARY TRANSITIONAL CELL CARCINOMA OF UTERUS
C2211952|T047||CCS_10|MICROPAPILLARY TRANSITIONAL CELL CARCINOMA OF UTERUS 
C2018619|T047||CCS_10|SPINDLE CELL TRANSITIONAL CELL CARCINOMA OF UTERUS 
C2018619|T047||CCS_10|SPINDLE CELL TRANSITIONAL CELL CARCINOMA OF UTERUS
C2211963|T047||CCS_10|MEDULLARY CARCINOMA OF UTERUS 
C2211963|T047||CCS_10|MEDULLARY CARCINOMA OF UTERUS
C2188880|T047||CCS_10|MIXED CELLULARITY HODGKIN'S LYMPHOMA OF UTERUS
C2188880|T047||CCS_10|MIXED CELLULARITY HODGKIN'S LYMPHOMA OF UTERUS 
C2188878|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION OF UTERUS
C2188878|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION OF UTERUS 
C2188896|T047||CCS_10|IMMUNOBLASTIC LARGE B-CELL DIFFUSE LYMPHOMA OF UTERUS 
C2188896|T047||CCS_10|IMMUNOBLASTIC LARGE B-CELL DIFFUSE LYMPHOMA OF UTERUS
C2188894|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF UTERUS 
C2188894|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF UTERUS
C2217773|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGE IIIC 
C2217773|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGE IIIC
C2217773|T047||CCS_10|UTERINE CANCER STAGE IIIC
C2217773|T047||CCS_10|MALIGNANT TUMOR OF UTERUS STAGE IIIC
C2109332|T047||CCS_10|KERATINIZING SQUAMOUS CELL CARCINOMA OF UTERUS 
C2109332|T047||CCS_10|KERATINIZING SQUAMOUS CELL CARCINOMA OF UTERUS
C2138886|T047||CCS_10|LARGE CELL NONKERATINIZING SQUAMOUS CELL CARCINOMA OF UTERUS 
C2138886|T047||CCS_10|UTERINE MALIGNANT CARCINOMA SQUAMOUS CELL LARGE CELL NONKERATINIZING
C2138886|T047||CCS_10|LARGE CELL NONKERATINIZING SQUAMOUS CELL CARCINOMA OF UTERUS
C2211955|T047||CCS_10|MICROINVASIVE SQUAMOUS CELL CARCINOMA OF UTERUS 
C2211955|T047||CCS_10|MICROINVASIVE SQUAMOUS CELL CARCINOMA OF UTERUS
C2188884|T047||CCS_10|GRADE 1 NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF UTERUS 
C2188884|T047||CCS_10|GRADE 1 NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF UTERUS
C2046746|T047||CCS_10|HODGKIN'S SARCOMA OF UTERUS
C2046746|T047||CCS_10|HODGKIN'S SARCOMA OF UTERUS 
C2188902|T047||CCS_10|MIXED SMALL AND LARGE CELL DIFFUSE LYMPHOMA OF UTERUS
C2188902|T047||CCS_10|MIXED SMALL AND LARGE CELL DIFFUSE LYMPHOMA OF UTERUS 
C2113738|T047||CCS_10|PRECURSOR CELL LYMPHOBLASTIC LYMPHOMA OF UTERUS 
C2113738|T047||CCS_10|PRECURSOR CELL LYMPHOBLASTIC LYMPHOMA OF UTERUS
C2009896|T047||CCS_10|FUSIFORM TYPE SMALL CELL CARCINOMA OF UTERUS
C2009896|T047||CCS_10|FUSIFORM TYPE SMALL CELL CARCINOMA OF UTERUS 
C2189372|T047||CCS_10|VERRUCOUS CARCINOMA OF UTERUS
C2189372|T047||CCS_10|VERRUCOUS CARCINOMA OF UTERUS 
C2145473|T047||CCS_10|TRANSITIONAL CELL CARCINOMA OF UTERUS 
C2145473|T047||CCS_10|TRANSITIONAL CELL CARCINOMA OF UTERUS
C2138465|T047||CCS_10|CRIBRIFORM CARCINOMA OF UTERUS 
C2138465|T047||CCS_10|CRIBRIFORM CARCINOMA OF UTERUS
C2211961|T047||CCS_10|ADENOSQUAMOUS CARCINOMA OF UTERUS 
C2211961|T047||CCS_10|ADENOSQUAMOUS CARCINOMA OF UTERUS
C2007053|T047||CCS_10|CARCINOMA SIMPLEX OF UTERUS
C2007053|T047||CCS_10|CARCINOMA SIMPLEX OF UTERUS 
C2007053|T047||CCS_10|CARCINOMA SIMPLEX OF URETHRA 
C2007053|T047||CCS_10|CARCINOMA SIMPLEX OF URETHRA
C2012551|T047||CCS_10|GRANULAR CELL CARCINOMA OF UTERUS 
C2012551|T047||CCS_10|GRANULAR CELL CARCINOMA OF UTERUS
C2182940|T047||CCS_10|DESMOPLASTIC SMALL ROUND CELL TUMOR OF UTERUS 
C2182940|T047||CCS_10|DESMOPLASTIC SMALL ROUND CELL TUMOR OF UTERUS
C2046534|T047||CCS_10|UTERINE MALIGNANT LYMPHOMA HODGKIN'S AND NON-HODGKIN'S
C2046534|T047||CCS_10|COMPOSITE HODGKIN'S AND NON-HODGKIN'S LYMPHOMA OF UTERUS 
C2046534|T047||CCS_10|COMPOSITE HODGKIN'S AND NON-HODGKIN'S LYMPHOMA OF UTERUS
C2188904|T047||CCS_10|SMALL B-CELL LYMPHOCYTIC LYMPHOMA OF UTERUS 
C2188904|T047||CCS_10|SMALL B-CELL LYMPHOCYTIC LYMPHOMA OF UTERUS
C2217770|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGE IIB
C2217770|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGE IIB 
C2217770|T047||CCS_10|UTERINE CANCER STAGE IIB
C2217770|T047||CCS_10|MALIGNANT TUMOR OF UTERUS STAGE IIB
C2217771|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGE IIIA 
C2217771|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGE IIIA
C2217771|T047||CCS_10|UTERINE CANCER STAGE IIIA
C2217771|T047||CCS_10|MALIGNANT TUMOR OF UTERUS STAGE IIIA
C2217772|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGE IIIB 
C2217772|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGE IIIB
C2217772|T047||CCS_10|MALIGNANT TUMOR OF UTERUS STAGE IIIB
C2217772|T047||CCS_10|UTERINE CANCER STAGE IIIB
C2211949|T047||CCS_10|MALIGNANT EPITHELIOMA OF UTERUS 
C2211949|T047||CCS_10|MALIGNANT EPITHELIOMA OF UTERUS
C2211951|T047||CCS_10|SMALL CELL CARCINOMA OF UTERUS 
C2211951|T047||CCS_10|SMALL CELL CARCINOMA OF UTERUS
C2211962|T047||CCS_10|EPITHELIAL-MYOEPITHELIAL CARCINOMA OF UTERUS 
C2211962|T047||CCS_10|EPITHELIAL-MYOEPITHELIAL CARCINOMA OF UTERUS
C2046606|T047||CCS_10|HODGKIN'S GRANULOMA OF UTERUS
C2046606|T047||CCS_10|HODGKIN'S GRANULOMA OF UTERUS 
C2188890|T047||CCS_10|FOLLICULAR LYMPHOMA OF UTERUS
C2188890|T047||CCS_10|FOLLICULAR LYMPHOMA OF UTERUS 
C2188901|T047||CCS_10|ANGIOIMMUNOBLASTIC T-CELL LYMPHOMA OF UTERUS 
C2188901|T047||CCS_10|ANGIOIMMUNOBLASTIC T-CELL LYMPHOMA OF UTERUS
C2188901|T047||CCS_10|ANGIOIMMUNOBLASTIC LYMPHADENOPATHY WITH DYSPROTEINEMIA (AILD) OF UTERUS
C2019461|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF UTERUS 
C2019461|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF UTERUS
C2217768|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGE IC
C2217768|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGE IC 
C2217768|T047||CCS_10|MALIGNANT TUMOR OF UTERUS STAGE IC
C2217768|T047||CCS_10|UTERINE CANCER STAGE IC
C2217774|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGE IVA 
C2217774|T047||CCS_10|MALIGNANT NEOPLASM OF UTERUS STAGE IVA
C2217774|T047||CCS_10|MALIGNANT TUMOR OF UTERUS STAGE IVA
C2217774|T047||CCS_10|UTERINE CANCER STAGE IVA
C2082473|T047||CCS_10|PLEOMORPHIC CARCINOMA OF UTERUS 
C2082473|T047||CCS_10|PLEOMORPHIC CARCINOMA OF UTERUS
C2011273|T047||CCS_10|GIANT CELL CARCINOMA OF UTERUS 
C2011273|T047||CCS_10|GIANT CELL CARCINOMA OF UTERUS
C2142943|T047||CCS_10|PSEUDOSARCOMATOUS CARCINOMA OF UTERUS
C2142943|T047||CCS_10|PSEUDOSARCOMATOUS CARCINOMA OF UTERUS 
C2200280|T047||CCS_10|LYMPHOEPITHELIAL SQUAMOUS CELL CARCINOMA OF UTERUS 
C2200280|T047||CCS_10|LYMPHOEPITHELIAL SQUAMOUS CELL CARCINOMA OF UTERUS
C2211959|T047||CCS_10|ADENOID CYSTIC CARCINOMA OF UTERUS 
C2211959|T047||CCS_10|ADENOID CYSTIC CARCINOMA OF UTERUS
C2188877|T047||CCS_10|LYMPHOCYTE-RICH HODGKIN'S LYMPHOMA OF UTERUS 
C2188877|T047||CCS_10|LYMPHOCYTE-RICH HODGKIN'S LYMPHOMA OF UTERUS
C2188876|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION, DIFFUSE FIBROSIS OF UTERUS
C2188876|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION, DIFFUSE FIBROSIS OF UTERUS 
C2188882|T047||CCS_10|NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF UTERUS 
C2188882|T047||CCS_10|NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF UTERUS
C2188893|T047||CCS_10|GRADE 3 FOLLICULAR LYMPHOMA OF UTERUS 
C2188893|T047||CCS_10|GRADE 3 FOLLICULAR LYMPHOMA OF UTERUS
C2188879|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION, RETICULAR OF UTERUS 
C2188879|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION, RETICULAR OF UTERUS
C0153595|T047||CCS_10|MALIGNANT NEOPLASM OF UNDESCENDED TESTIS
C0153595|T047||CCS_10|MALIGNANT TUMOR OF UNDESCENDED TESTIS
C0153595|T047||CCS_10|MALIGNANT NEOPLASM OF UNDESCENDED TESTIS 
C0153595|T047||CCS_10|MALIGNANT NEOPLASM OF RETAINED TESTIS
C0153595|T047||CCS_10|MALIGNANT NEOPLASM OF RETAINED TESTIS 
C0153595|T047||CCS_10|MALIGNANT TUMOR OF RETAINED TESTIS
C0153595|T047||CCS_10|MAL NEO UNDESCEND TESTIS
C0153595|T047||CCS_10|MALIGNANT TUMOR OF RETAINED TESTIS 
C0153595|T047||CCS_10|MALIGNANT TUMOUR OF RETAINED TESTIS
C0153595|T047||CCS_10|MALIGNANT NEOPLASM OF UNDESCENDED TESTIS NOS 
C0153595|T047||CCS_10|CANCER OF INTRA-ABDOMINAL TESTIS
C0153595|T047||CCS_10|MALIGNANT NEOPLASM OF UNDESCENDED TESTIS NOS
C0153595|T047||CCS_10|MALIGNANT NEOPLASM OF TESTIS, UNDESCENDED
C0153595|T047||CCS_10|CANCER OF UNDESCENDED TESTIS
C0153595|T047||CCS_10|MALIGNANT TUMOUR OF UNDESCENDED TESTIS
C0153595|T047||CCS_10|MALIGNANT TUMOR OF UNDESCENDED TESTIS 
C0348906|T047||CCS_10|MALIGNANT NEOPLASM OF DESCENDED TESTIS
C0348906|T047||CCS_10|TESTICULAR NEOPLASM MALIGNANT DESCENDED TESTIS
C0348906|T047||CCS_10|MALIGNANT NEOPLASM OF DESCENDED TESTIS 
C0348906|T047||CCS_10|MALIGNANT NEOPLASM OF DESCENDED TESTIS 
C0348906|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF DESCENDED TESTIS 
C0348906|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF DESCENDED TESTIS
C0348906|T047||CCS_10|TESTICULAR NEOPLASM MALIGNANT DESCENDED TESTIS PRIMARY
C0348906|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF DESCENDED TESTIS 
C0348906|T047||CCS_10|MALIGNANT NEOPLASM OF TESTIS, DESCENDED
C0153594|T047||CCS_10|MALIGNANT NEOPLASM OF TESTIS
C0153594|T047||CCS_10|TESTICULAR CANCER
C0153594|T047||CCS_10|MALIGNANT NEOPLASM OF TESTIS, UNSPECIFIED
C0153594|T047||CCS_10|TESTICULAR CANCER 
C0153594|T047||CCS_10|MALIGNANT NEOPLASM OF TESTIS 
C0153594|T047||CCS_10|CANCERS, TESTIS
C0153594|T047||CCS_10|TESTIS CANCERS
C0153594|T047||CCS_10|CANCER, TESTICULAR
C0153594|T047||CCS_10|CANCERS, TESTICULAR
C0153594|T047||CCS_10|TESTICULAR CANCERS
C0153594|T047||CCS_10|MALIGNANT TUMOR OF TESTIS
C0153594|T047||CCS_10|CANCER OF TESTIS
C0153594|T047||CCS_10|MALIGNANT NEOPLASM OF TESTIS NOS
C0153594|T047||CCS_10|MALIGNANT NEOPLASM OF TESTIS, UNSPECIFIED WHETHER DESCENDED OR UNDESCENDED
C0153594|T047||CCS_10|CANCER, TESTIS
C0153594|T047||CCS_10|MALIGNANT NEOPLASM OF TESTIS NOS 
C0153594|T047||CCS_10|TESTIS CANCER
C0153594|T047||CCS_10|TESTIS--CANCER
C0153594|T047||CCS_10|TESTIS NEOPLASM MALIGNANT
C0153594|T047||CCS_10|TESTICULAR NEOPLASMS MALIGNANT
C0153594|T047||CCS_10|CANCER OF THE TESTIS
C0153594|T047||CCS_10|CANCER OF THE TESTES
C0153594|T047||CCS_10|MALIGNANT TUMOUR OF TESTIS
C0153594|T047||CCS_10|MALIGNANT TUMOR OF TESTIS 
C0153594|T047||CCS_10|TESTICLE CANCER
C0153594|T047||CCS_10|MALIGNANT NEOPLASM OF TESTIS, NOS
C0153594|T047||CCS_10|MALIGNANT NEOPLASM OF THE TESTIS
C0153594|T047||CCS_10|MALIGNANT TESTICULAR NEOPLASM
C0153594|T047||CCS_10|MALIGNANT TESTICULAR TUMOR
C0153594|T047||CCS_10|MALIGNANT TUMOR OF THE TESTIS
C0153594|T047||CCS_10|NEOPLASM MALIG;TESTIS
C0153594|T047||CCS_10|MALIGNANT NEOSPLASM OF THE TESTIS
C0036631|T047||CCS_10|SEMINOMA
C0036631|T047||CCS_10|SEMINOMAS
C0036631|T047||CCS_10|TESTICULAR SEMINOMA
C0036631|T047||CCS_10|SEMINOMA OF TESTIS 
C0036631|T047||CCS_10|SEMINOMA OF TESTIS
C0036631|T047||CCS_10|SEMINOMA 
C0036631|T047||CCS_10|SEMINOMA (MORPHOLOGIC ABNORMALITY)
C0036631|T047||CCS_10|SEMINOMA, NO ICD-O SUBTYPE
C0036631|T047||CCS_10|SEMINOMA [DISEASE/FINDING]
C0036631|T047||CCS_10|[M]SEMINOMAS
C0036631|T047||CCS_10|SEMINOMA TESTIS
C0036631|T047||CCS_10|[M]SEMINOMAS (MORPHOLOGIC ABNORMALITY)
C0036631|T047||CCS_10|[M]SEMINOMA NOS
C0036631|T047||CCS_10|[M]SEMINOMA NOS (MORPHOLOGIC ABNORMALITY)
C0036631|T047||CCS_10|MALIGNANT NEOPLASM SEMINOMA
C0036631|T047||CCS_10|SEMINOMA 
C0036631|T047||CCS_10|SEMINOMA, NO ICD-O SUBTYPE (MORPHOLOGIC ABNORMALITY)
C0036631|T047||CCS_10|SEMINOMA, NO INTERNATIONAL CLASSIFICATION OF DISEASES FOR ONCOLOGY SUBTYPE
C0036631|T047||CCS_10|SEMINOMA, NO INTERNATIONAL CLASSIFICATION OF DISEASES FOR ONCOLOGY SUBTYPE (MORPHOLOGIC ABNORMALITY)
C0036631|T047||CCS_10|SEMINOMA, MALIGNANT
C0036631|T047||CCS_10|SEMINOMA, PURE
C0036631|T047||CCS_10|TESTICULAR SEMINOMA PURE NOS
C0036631|T047||CCS_10|TESTICULAR SEMINOMA (PURE)
C0036631|T047||CCS_10|SEMINOMA OF TESTIS 
C0036631|T047||CCS_10|SEMINOMA OF THE TESTIS
C0036631|T047||CCS_10|SEMINOMA, TESTICULAR
C0036631|T047||CCS_10|TESTICLE CANCER, SEMINOMA
C0036631|T047||CCS_10|TESTICULAR CANCER, SEMINOMA
C0036631|T047||CCS_10|TESTIS CANCER, SEMINOMA
C0036631|T047||CCS_10|SEMINOMA, NOS
C0036631|T047||CCS_10|TESTICULAR SEMINOMA PURE
C0855193|T047||CCS_10|TESTICULAR CHORIOCARCINOMA STAGE I
C0855193|T047||CCS_10|STAGE I TESTICULAR CHORIOCARCINOMA AJCC V7
C0855193|T047||CCS_10|STAGE I TESTICULAR CHORIOCARCINOMA AJCC V6
C0855193|T047||CCS_10|STAGE I TESTICULAR CHORIOCARCINOMA
C0853869|T047||CCS_10|TESTICULAR CHORIOCARCINOMA STAGE II
C0853869|T047||CCS_10|STAGE II TESTICULAR CHORIOCARCINOMA AJCC V6
C0853869|T047||CCS_10|STAGE II TESTICULAR CHORIOCARCINOMA AJCC V7
C0853869|T047||CCS_10|STAGE II TESTICULAR CHORIOCARCINOMA
C0855184|T047||CCS_10|TESTICULAR CHORIOCARCINOMA STAGE III
C0855184|T047||CCS_10|STAGE III TESTICULAR CHORIOCARCINOMA AJCC V6
C0855184|T047||CCS_10|STAGE III TESTICULAR CHORIOCARCINOMA AJCC V7
C0855184|T047||CCS_10|STAGE III TESTICULAR CHORIOCARCINOMA
C0855194|T047||CCS_10|TESTICULAR EMBRYONAL CARCINOMA STAGE I
C0855194|T047||CCS_10|STAGE I TESTICULAR EMBRYONAL CARCINOMA AJCC V6
C0855194|T047||CCS_10|STAGE I TESTICULAR EMBRYONAL CARCINOMA AJCC V7
C0855194|T047||CCS_10|STAGE I TESTICULAR EMBRYONAL CARCINOMA
C0855195|T047||CCS_10|TESTICULAR EMBRYONAL CARCINOMA STAGE II
C0855195|T047||CCS_10|STAGE II TESTICULAR EMBRYONAL CARCINOMA AJCC V6
C0855195|T047||CCS_10|STAGE II TESTICULAR EMBRYONAL CARCINOMA AJCC V7
C0855195|T047||CCS_10|STAGE II TESTICULAR EMBRYONAL CARCINOMA
C0855196|T047||CCS_10|TESTICULAR EMBRYONAL CARCINOMA STAGE III
C0855196|T047||CCS_10|STAGE III TESTICULAR EMBRYONAL CARCINOMA AJCC V7
C0855196|T047||CCS_10|STAGE III TESTICULAR EMBRYONAL CARCINOMA AJCC V6
C0855196|T047||CCS_10|STAGE III TESTICULAR EMBRYONAL CARCINOMA
C0855203|T047||CCS_10|TESTICULAR GERM CELL TUMOUR MIXED STAGE I
C0855203|T047||CCS_10|STAGE I TESTICULAR MIXED GERM CELL TUMOR AJCC V6
C0855203|T047||CCS_10|STAGE I TESTICULAR MIXED GERM CELL TUMOR AJCC V7
C0855203|T047||CCS_10|TESTICULAR GERM CELL TUMOR MIXED STAGE I
C0855203|T047||CCS_10|STAGE I TESTICULAR MIXED GERM CELL TUMOR
C0855199|T047||CCS_10|TESTICULAR GERM CELL TUMOUR MIXED STAGE II
C0855199|T047||CCS_10|STAGE II TESTICULAR MIXED GERM CELL TUMOR AJCC V7
C0855199|T047||CCS_10|STAGE II TESTICULAR MIXED GERM CELL TUMOR AJCC V6
C0855199|T047||CCS_10|TESTICULAR GERM CELL TUMOR MIXED STAGE II
C0855199|T047||CCS_10|STAGE II TESTICULAR MIXED GERM CELL TUMOR
C0855204|T047||CCS_10|TESTICULAR GERM CELL TUMOUR MIXED STAGE III
C0855204|T047||CCS_10|STAGE III TESTICULAR MIXED GERM CELL TUMOR AJCC V6
C0855204|T047||CCS_10|STAGE III TESTICULAR MIXED GERM CELL TUMOR AJCC V7
C0855204|T047||CCS_10|TESTICULAR GERM CELL TUMOR MIXED STAGE III
C0855204|T047||CCS_10|STAGE III TESTICULAR MIXED GERM CELL TUMOR
C0855205|T047||CCS_10|TESTICULAR MALIGNANT TERATOMA STAGE I
C0855206|T047||CCS_10|TESTICULAR MALIGNANT TERATOMA STAGE II
C0855207|T047||CCS_10|TESTICULAR MALIGNANT TERATOMA STAGE III
C0855208|T047||CCS_10|TESTICULAR SEMINOMA (PURE) STAGE I
C0855209|T047||CCS_10|TESTICULAR SEMINOMA (PURE) STAGE II
C0855210|T047||CCS_10|TESTICULAR SEMINOMA (PURE) STAGE III
C0855213|T047||CCS_10|TESTICULAR YOLK SAC TUMOUR STAGE I
C0855213|T047||CCS_10|STAGE I TESTICULAR YOLK SAC TUMOR AJCC V6
C0855213|T047||CCS_10|STAGE I TESTICULAR YOLK SAC TUMOR AJCC V7
C0855213|T047||CCS_10|TESTICULAR ENDODERMAL SINUS TUMOR STAGE I
C0855213|T047||CCS_10|TESTICULAR ENDODERMAL SINUS TUMOUR STAGE I
C0855213|T047||CCS_10|TESTICULAR YOLK SAC TUMOR STAGE I
C0855213|T047||CCS_10|STAGE I TESTICULAR YOLK SAC TUMOR
C0855214|T047||CCS_10|TESTICULAR YOLK SAC TUMOUR STAGE II
C0855214|T047||CCS_10|STAGE II TESTICULAR YOLK SAC TUMOR AJCC V6
C0855214|T047||CCS_10|STAGE II TESTICULAR YOLK SAC TUMOR AJCC V7
C0855214|T047||CCS_10|TESTICULAR ENDODERMAL SINUS TUMOUR STAGE II
C0855214|T047||CCS_10|TESTICULAR YOLK SAC TUMOR STAGE II
C0855214|T047||CCS_10|TESTICULAR ENDODERMAL SINUS TUMOR STAGE II
C0855214|T047||CCS_10|STAGE II TESTICULAR YOLK SAC TUMOR
C0855215|T047||CCS_10|TESTICULAR YOLK SAC TUMOUR STAGE III
C0855215|T047||CCS_10|STAGE III TESTICULAR YOLK SAC TUMOR AJCC V6
C0855215|T047||CCS_10|STAGE III TESTICULAR YOLK SAC TUMOR AJCC V7
C0855215|T047||CCS_10|TESTICULAR YOLK SAC TUMOR STAGE III
C0855215|T047||CCS_10|TESTICULAR ENDODERMAL SINUS TUMOR STAGE III
C0855215|T047||CCS_10|TESTICULAR ENDODERMAL SINUS TUMOUR STAGE III
C0855215|T047||CCS_10|STAGE III TESTICULAR YOLK SAC TUMOR
C0855197|T047||CCS_10|TESTICULAR CANCER (EXCLUDING GERM CELL OR TROPHOBLASTIC CANCER)
C0855197|T047||CCS_10|TESTICULAR CA. (NO GERM/TROPHO.)
C0855197|T047||CCS_10|TESTICULAR CANCER
C0855197|T047||CCS_10|TESTICULAR GERM CELL CANCER NOS
C0855197|T047||CCS_10|TESTICULAR MALIGNANT GERM CELL TUMOR NOS
C0855197|T047||CCS_10|TESTICULAR GERM CELL CANCER
C0855197|T047||CCS_10|MALIGNANT GERM CELL TUMOR OF TESTIS
C0855197|T047||CCS_10|MALIGNANT GERM CELL TUMOUR OF TESTIS
C0855197|T047||CCS_10|MALIGNANT GERM CELL TUMOR OF TESTIS 
C0855197|T047||CCS_10|TESTICULAR MALIGNANT GERM CELL TUMOR
C0855197|T047||CCS_10|MALIGNANT GERM CELL NEOPLASM OF TESTIS
C0855197|T047||CCS_10|MALIGNANT GERM CELL NEOPLASM OF THE TESTIS
C0855197|T047||CCS_10|MALIGNANT GERM CELL TUMOR OF THE TESTIS
C0855197|T047||CCS_10|MALIGNANT TESTICULAR GERM CELL NEOPLASM
C0855197|T047||CCS_10|MALIGNANT TESTICULAR GERM CELL TUMOR
C0238449|T047||CCS_10|CHORIOCARCINOMA OF TESTIS
C0238449|T047||CCS_10|CHORIOCARCINOMA OF TESTIS 
C0238449|T047||CCS_10|TESTICULAR CHORIOCARCINOMA
C0238449|T047||CCS_10|TESTICULAR CHORIOCARCINOMA NOS
C0238449|T047||CCS_10|CHORIOCARCINOMA OF TESTIS 
C0238449|T047||CCS_10|CHORIOCARCINOMA OF THE TESTIS
C0238449|T047||CCS_10|CHORIOCARCINOMA, TESTICULAR
C0238449|T047||CCS_10|TESTICLE CANCER, CHORIOCARCINOMA
C0238449|T047||CCS_10|TESTICULAR CANCER, CHORIOCARCINOMA
C0238449|T047||CCS_10|TESTIS CANCER, CHORIOCARCINOMA
C0238448|T047||CCS_10|EMBRYONAL CARCINOMA OF TESTIS 
C0238448|T047||CCS_10|EMBRYONAL CARCINOMA OF TESTIS
C0238448|T047||CCS_10|TESTICULAR EMBRYONAL CARCINOMA
C0238448|T047||CCS_10|TESTICULAR EMBRYONAL CARCINOMA NOS
C0238448|T047||CCS_10|EMBRYONAL CARCINOMA OF THE TESTIS
C0238448|T047||CCS_10|EMBRYONAL CARCINOMA, TESTICULAR
C0238448|T047||CCS_10|TESTICLE CANCER, EMBRYONAL
C0238448|T047||CCS_10|TESTICULAR CANCER, EMBRYONAL
C0238448|T047||CCS_10|TESTIS CANCER, EMBRYONAL
C2363951|T047||CCS_10|TESTICULAR GERM CELL CANCER METASTATIC
C1096715|T047||CCS_10|TESTICULAR CANCER METASTATIC
C1096715|T047||CCS_10|METASTATIC MALIGNANT TESTICULAR GERM CELL TUMOR
C1096715|T047||CCS_10|METASTATIC TESTICULAR CANCER
C2747856|T047||CCS_10|TESTICULAR CHORIOCARCINOMA RECURRENT
C0278841|T047||CCS_10|RECURRENT MALIGNANT TESTICULAR GERM CELL TUMOR
C0278841|T047||CCS_10|RECURRENT TESTICULAR CANCER
C0278841|T047||CCS_10|TESTIS CANCER RECURRENT
C0278841|T047||CCS_10|CANCER OF THE TESTIS, RECURRENT
C0278841|T047||CCS_10|CANCER OF THE TESTIS, RELAPSED
C0278841|T047||CCS_10|CARCINOMA OF THE TESTIS, RECURRENT
C0278841|T047||CCS_10|CARCINOMA OF THE TESTIS, RELAPSED
C0278841|T047||CCS_10|RECURRENT CANCER OF THE TESTIS
C0278841|T047||CCS_10|RECURRENT CARCINOMA OF THE TESTIS
C0278841|T047||CCS_10|RECURRENT OR REFRACTORY TESTICULAR CANCER
C0278841|T047||CCS_10|RECURRENT TESTIS CANCER
C0278841|T047||CCS_10|RELAPSED CANCER OF THE TESTIS
C0278841|T047||CCS_10|RELAPSED CARCINOMA OF THE TESTIS
C0278841|T047||CCS_10|RELAPSED TESTICULAR CANCER
C0278841|T047||CCS_10|RELAPSED TESTIS CANCER
C0278841|T047||CCS_10|TESTICLE CANCER, RECURRENT
C0278841|T047||CCS_10|TESTICLE CANCER, REFRACTORY
C0278841|T047||CCS_10|TESTICLE CANCER, RELAPSED
C0278841|T047||CCS_10|TESTICULAR CANCER, RECURRENT
C0278841|T047||CCS_10|TESTICULAR CANCER, RELAPSED
C0278841|T047||CCS_10|TESTIS CANCER, RECURRENT
C0278841|T047||CCS_10|TESTIS CANCER, RELAPSED
C0278841|T047||CCS_10|RECURRENT CANCER OF TESTIS
C0278841|T047||CCS_10|RELAPSED CANCER OF TESTIS
C2845878|T047||CCS_10|MALIGNANT NEOPLASM OF UNSPECIFIED TESTIS, UNSPECIFIED WHETHER DESCENDED OR UNDESCENDED
C2845878|T047||CCS_10|MALIG NEOPLASM OF UNSP TESTIS, UNSP DESCENDED OR UNDESCENDED
C2845879|T047||CCS_10|MALIGNANT NEOPLASM OF RIGHT TESTIS, UNSPECIFIED WHETHER DESCENDED OR UNDESCENDED
C2845879|T047||CCS_10|MALIG NEOPLM OF RIGHT TESTIS, UNSP DESCENDED OR UNDESCENDED
C2845880|T047||CCS_10|MALIGNANT NEOPLASM OF LEFT TESTIS, UNSPECIFIED WHETHER DESCENDED OR UNDESCENDED
C2845880|T047||CCS_10|MALIG NEOPLASM OF LEFT TESTIS, UNSP DESCENDED OR UNDESCENDED
C2212306|T047||CCS_10|TESTICULAR NEOPLASM MALIGNANT SMALL CELL TYPE
C2212306|T047||CCS_10|MALIGNANT SMALL CELL NEOPLASM OF TESTIS 
C2212306|T047||CCS_10|MALIGNANT SMALL CELL NEOPLASM OF TESTIS
C2011413|T047||CCS_10|GIANT CELL TYPE NEOPLASM OF TESTIS 
C2011413|T047||CCS_10|GIANT CELL TYPE NEOPLASM OF TESTIS
C2011413|T047||CCS_10|TESTICULAR NEOPLASM MALIGNANT GIANT CELL TYPE
C2018694|T047||CCS_10|TESTICULAR NEOPLASM MALIGNANT SPINDLE CELL TYPE
C2018694|T047||CCS_10|SPINDLE CELL TYPE NEOPLASM OF TESTIS 
C2018694|T047||CCS_10|SPINDLE CELL TYPE NEOPLASM OF TESTIS
C2075654|T047||CCS_10|TESTICULAR NEOPLASM MALIGNANT CLEAR CELL TYPE
C2075654|T047||CCS_10|CLEAR CELL TYPE NEOPLASM OF TESTIS
C2075654|T047||CCS_10|CLEAR CELL TYPE NEOPLASM OF TESTIS 
C0677483|T047||CCS_10|CARCINOMA OF TESTIS 
C0677483|T047||CCS_10|CARCINOMA OF TESTIS
C0677483|T047||CCS_10|TESTICULAR CARCINOMA
C0677483|T047||CCS_10|CARCINOMA;TESTIS
C0677483|T047||CCS_10|TESTICULAR CA
C0677483|T047||CCS_10|CARCINOMA TESTIS
C0677483|T047||CCS_10|CARCINOMA TESTES
C0677483|T047||CCS_10|CARCINOMA OF THE TESTIS
C2212309|T047||CCS_10|ADENOCARCINOMA OF TESTIS
C2212309|T047||CCS_10|ADENOCARCINOMA OF TESTIS 
C2212309|T047||CCS_10|TESTICULAR ADENOCARCINOMA
C2212312|T047||CCS_10|MALIGNANT GONADAL NEOPLASM OF TESTIS
C2212312|T047||CCS_10|MALIGNANT GONADAL NEOPLASM OF TESTIS 
C1336727|T047||CCS_10|SARCOMA OF TESTIS 
C1336727|T047||CCS_10|SARCOMA OF TESTIS
C1336727|T047||CCS_10|SARCOMA OF THE TESTIS
C1336727|T047||CCS_10|TESTICULAR SARCOMA
C1336726|T047||CCS_10|TESTICULAR MYOSARCOMA RHABDOMYOSARCOMA
C1336726|T047||CCS_10|RHABDOMYOSARCOMA OF TESTIS 
C1336726|T047||CCS_10|RHABDOMYOSARCOMA OF TESTIS
C1336726|T047||CCS_10|RHABDOMYOSARCOMA OF THE TESTIS
C1336726|T047||CCS_10|TESTICULAR RHABDOMYOSARCOMA
C2242809|T047||CCS_10|GERMINOMA OF TESTIS
C2242809|T047||CCS_10|GERMINOMA OF TESTIS 
C1334154|T047||CCS_10|MALIGNANT TERATOMA OF TESTIS
C1334154|T047||CCS_10|MALIGNANT TERATOMA OF TESTIS 
C1334154|T047||CCS_10|TESTICULAR MALIGNANT TERATOMA
C1334154|T047||CCS_10|IMMATURE TERATOMA OF TESTIS
C1334154|T047||CCS_10|IMMATURE TERATOMA OF THE TESTIS
C1334154|T047||CCS_10|IMMATURE TESTICULAR TERATOMA
C1334154|T047||CCS_10|MALIGNANT TERATOMA OF THE TESTIS
C1334154|T047||CCS_10|MALIGNANT TESTICULAR TERATOMA
C1334154|T047||CCS_10|TESTICULAR IMMATURE TERATOMA
C1334154|T047||CCS_10|MALIGNANT TERATOMA OF TESTIS 
C2057624|T047||CCS_10|MALIGNANT EPITHELIOID TROPHOBLASTIC TUMOR OF TESTIS
C2057624|T047||CCS_10|MALIGNANT EPITHELIOID TROPHOBLASTIC TUMOR OF TESTIS 
C0349644|T047||CCS_10|PRIMARY TESTICULAR LYMPHOMA
C0349644|T047||CCS_10|MALIGNANT LYMPHOMA OF TESTIS 
C0349644|T047||CCS_10|MALIGNANT LYMPHOMA OF TESTIS
C0349644|T047||CCS_10|MALIGNANT LYMPHOMA OF TESTIS 
C0349644|T047||CCS_10|LYMPHOMA OF TESTIS
C0349644|T047||CCS_10|LYMPHOMA OF THE TESTIS
C0349644|T047||CCS_10|TESTICULAR LYMPHOMA
C2212324|T047||CCS_10|MALIGNANT PLASMACYTOMA OF TESTIS 
C2212324|T047||CCS_10|MALIGNANT PLASMACYTOMA OF TESTIS
C2212326|T047||CCS_10|MALIGNANT MASTOCYTOSIS OF TESTIS
C2212326|T047||CCS_10|MALIGNANT MASTOCYTOSIS OF TESTIS 
C2217647|T047||CCS_10|MALIGNANT NEOPLASM OF TESTIS STAGING
C2217647|T047||CCS_10|MALIGNANT NEOPLASM OF TESTIS STAGING 
C2217647|T047||CCS_10|MALIGNANT TESTICULAR NEOPLASM STAGING
C2217647|T047||CCS_10|MALIGNANT TUMOR OF TESTIS STAGING
C2217647|T047||CCS_10|TESTICULAR CANCER STAGING
C2188087|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF TESTIS 
C2188087|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF TESTIS
C2057597|T047||CCS_10|CHORIOCARCINOMA OF TESTIS WITH OTHER GERM CELL ELEMENTS 
C2057597|T047||CCS_10|CHORIOCARCINOMA OF TESTIS WITH OTHER GERM CELL ELEMENTS
C2057597|T047||CCS_10|TESTICULAR CHORIOCARCINOMA COMBINED WITH OTHER GERM CELL ELEMENTS
C2057494|T047||CCS_10|TERATOCARCINOMA OF TESTIS 
C2057494|T047||CCS_10|TERATOCARCINOMA OF TESTIS
C2057494|T047||CCS_10|TESTICULAR TERATOCARCINOMA
C0334517|T047||CCS_10|SPERMATOCYTIC SEMINOMA
C0334517|T047||CCS_10|SPERMATOCYTOMA
C0334517|T047||CCS_10|SPERMATOCYTIC SEMINOMA (MORPHOLOGIC ABNORMALITY)
C0334517|T047||CCS_10|TESTICULAR SPERMATOCYTIC SEMINOMA
C0279708|T047||CCS_10|YOLK SAC TUMOR OF TESTIS 
C0279708|T047||CCS_10|YOLK SAC TUMOR OF TESTIS
C0279708|T047||CCS_10|TESTICULAR YOLK SAC TUMOUR
C0279708|T047||CCS_10|TESTICULAR YOLK SAC TUMOR
C0279708|T047||CCS_10|TESTICLE CANCER, YOLK SAC TUMOR
C0279708|T047||CCS_10|TESTICULAR CANCER, YOLK SAC TUMOR
C0279708|T047||CCS_10|TESTIS CANCER, YOLK SAC TUMOR
C0279708|T047||CCS_10|YOLK SAC TUMOR OF THE TESTIS
C0279708|T047||CCS_10|YOLK SAC TUMOR, TESTICULAR
C0279708|T047||CCS_10|ENDODERMAL SINUS NEOPLASM OF TESTIS
C0279708|T047||CCS_10|ENDODERMAL SINUS NEOPLASM OF THE TESTIS
C0279708|T047||CCS_10|ENDODERMAL SINUS TUMOR OF TESTIS
C0279708|T047||CCS_10|ENDODERMAL SINUS TUMOR OF THE TESTIS
C0279708|T047||CCS_10|TESTICULAR ENDODERMAL SINUS NEOPLASM
C0279708|T047||CCS_10|TESTICULAR ENDODERMAL SINUS TUMOR
C0279708|T047||CCS_10|TESTICULAR YOLK SAC NEOPLASM
C0279708|T047||CCS_10|YOLK SAC NEOPLASM OF TESTIS
C0279708|T047||CCS_10|YOLK SAC NEOPLASM OF THE TESTIS
C1336720|T047||CCS_10|MALIGNANT MIXED GERM CELL TUMOR OF TESTIS 
C1336720|T047||CCS_10|MALIGNANT MIXED GERM CELL TUMOR OF TESTIS
C1336720|T047||CCS_10|TESTICULAR GERM CELL TUMOUR MIXED
C1336720|T047||CCS_10|TESTICULAR GERM CELL TUMOR MIXED
C1336720|T047||CCS_10|MIXED GERM CELL NEOPLASM OF TESTIS
C1336720|T047||CCS_10|MIXED GERM CELL NEOPLASM OF THE TESTIS
C1336720|T047||CCS_10|MIXED GERM CELL TUMOR OF TESTIS
C1336720|T047||CCS_10|MIXED GERM CELL TUMOR OF THE TESTIS
C1336720|T047||CCS_10|TESTICULAR GERM CELL TUMOR (MIXED)
C1336720|T047||CCS_10|TESTICULAR MIXED GERM CELL NEOPLASM
C1336720|T047||CCS_10|TESTICULAR MIXED GERM CELL TUMOR
C3646009|T047||CCS_10|TESTICULAR MALIGNANT NEOPLASM SECONDARY
C3646009|T047||CCS_10|SECONDARY MALIGNANT TESTICULAR NEOPLASM 
C3646009|T047||CCS_10|SECONDARY MALIGNANT TESTICULAR NEOPLASM
C3646010|T047||CCS_10|PRIMARY MALIGNANT TESTICULAR NEOPLASM
C3646010|T047||CCS_10|TESTICULAR MALIGNANT NEOPLASM PRIMARY
C3646010|T047||CCS_10|PRIMARY MALIGNANT TESTICULAR NEOPLASM 
C2315963|T047||CCS_10|TESTICULAR NEOPLASM MALIGNANT NON-SEMINOMATOUS
C2315963|T047||CCS_10|NON-SEMINOMATOUS MALIGNANT NEOPLASM OF TESTIS 
C2315963|T047||CCS_10|NON-SEMINOMATOUS MALIGNANT NEOPLASM OF TESTIS
C2315963|T047||CCS_10|NON-SEMINOMATOUS MALIGNANT NEOPLASM OF TESTIS 
C0346236|T047||CCS_10|MALIGNANT NEOPLASM OF ECTOPIC TESTIS
C0346236|T047||CCS_10|MALIGNANT NEOPLASM OF ECTOPIC TESTIS 
C0346236|T047||CCS_10|MALIGNANT TUMOR OF ECTOPIC TESTIS
C0346236|T047||CCS_10|CANCER OF ECTOPIC TESTIS
C0346236|T047||CCS_10|MALIGNANT TUMOUR OF ECTOPIC TESTIS
C0346236|T047||CCS_10|MALIGNANT TUMOR OF ECTOPIC TESTIS 
C0346241|T047||CCS_10|MALIGNANT NEOPLASM OF TUNICA VAGINALIS 
C0346241|T047||CCS_10|MALIGNANT NEOPLASM OF TUNICA VAGINALIS
C0346241|T047||CCS_10|MALIGNANT TUMOR OF TUNICA VAGINALIS
C0346241|T047||CCS_10|MALIGNANT TUMOUR OF TUNICA VAGINALIS
C0346241|T047||CCS_10|MALIGNANT TUMOR OF TUNICA VAGINALIS 
C0347003|T047||CCS_10|METASTATIC NEOPLASM TO THE TESTIS
C0347003|T047||CCS_10|METASTASES TO TESTICLE
C0347003|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM IN THE TESTIS
C0347003|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO THE TESTIS
C0347003|T047||CCS_10|METASTASIS TO TESTIS
C0347003|T047||CCS_10|METASTATIC TUMOR TO TESTIS
C0347003|T047||CCS_10|METASTATIC TUMOUR TO TESTIS
C0347003|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF TESTIS
C0347003|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO TESTIS
C0347003|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF TESTIS 
C0347003|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO TESTIS, NOS
C0347003|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF TESTIS, NOS
C0347003|T047||CCS_10|METASTATIC TUMOR TO THE TESTIS
C1304869|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF TESTIS 
C1304869|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF TESTIS
C0153596|T047||CCS_10|MALIG NEO TESTIS NEC
C0153596|T047||CCS_10|MALIGNANT NEOPLASM OF OTHER AND UNSPECIFIED TESTIS
C0153596|T047||CCS_10|MALIGNANT NEOPLASM OF TESTIS, OTHER AND UNSPECIFIED
C0852641|T047||CCS_10|TESTIS CANCER (EXCL GERM CELL)
C0852641|T047||CCS_10|TESTIS CANCER (EXCLUDING GERM CELL)
C1387440|T047||CCS_10|SEMINOMA; ANAPLASTIC, UNSPECIFIED SITE
C1387440|T047||CCS_10|ANAPLASTIC; SEMINOMA, UNSPECIFIED SITE
C1388417|T047||CCS_10|MALIGNANT; ANDROBLASTOMA, UNSPECIFIED SITE, MALE
C1388417|T047||CCS_10|MALIGNANT; ARRHENOBLASTOMA, UNSPECIFIED SITE, MALE
C1388417|T047||CCS_10|ANDROBLASTOMA; MALIGNANT, UNSPECIFIED SITE, MALE
C1388417|T047||CCS_10|ARRHENOBLASTOMA; MALIGNANT, UNSPECIFIED SITE, MALE
C1391898|T047||CCS_10|CARCINOMA; CHORION, UNSPECIFIED SITE, MALE
C1391898|T047||CCS_10|CHORION; CARCINOMA, UNSPECIFIED SITE, MALE
C1391920|T047||CCS_10|CARCINOMA; LEYDIG CELL, UNSPECIFIED SITE, MALE
C1391920|T047||CCS_10|LEYDIG CELL; CARCINOMA, UNSPECIFIED SITE, MALE
C1391943|T047||CCS_10|CARCINOMA; SERTOLI CELL, UNSPECIFIED SITE
C1391943|T047||CCS_10|SERTOLI CELL; CARCINOMA, UNSPECIFIED SITE
C1391944|T047||CCS_10|CARCINOMA; SERTOLI CELL, UNSPECIFIED SITE, MALE
C1391944|T047||CCS_10|SERTOLI CELL; CARCINOMA, UNSPECIFIED SITE, MALE
C1392523|T047||CCS_10|CHORIOCARCINOMA; MALE
C1392523|T047||CCS_10|CHORIOCARCINOMA; UNSPECIFIED SITE, MALE
C1395770|T047||CCS_10|TUMOR; YOLK SAC, UNSPECIFIED SITE, MALE
C1395770|T047||CCS_10|YOLK SAC; TUMOR, UNSPECIFIED SITE, MALE
C1395936|T047||CCS_10|DYSGERMINOMA; UNSPECIFIED SITE, MALE
C1396368|T047||CCS_10|EMBRYOMA; MALIGNANT, TESTIS
C1396368|T047||CCS_10|MALIGNANT; EMBRYOMA, TESTIS
C1396371|T047||CCS_10|EMBRYOMA; TESTIS
C1396371|T047||CCS_10|TESTIS; EMBRYOMA
C1396615|T047||CCS_10|ENDODERMAL; SINUS, TUMOR, UNSPECIFIED SITE, MALE
C1396615|T047||CCS_10|TUMOR; ENDODERMAL SINUS, UNSPECIFIED SITE, MALE
C1402881|T047||CCS_10|LEYDIG CELL; TUMOR, MALIGNANT, UNSPECIFIED SITE, MALE
C1402881|T047||CCS_10|TUMOR; LEYDIG CELL, MALIGNANT, UNSPECIFIED SITE, MALE
C0334528|T047||CCS_10|MALIGNANT TROPHOBLASTIC TERATOMA
C0334528|T047||CCS_10|TROPHOBLASTIC MALIGNANT TERATOMA 
C0334528|T047||CCS_10|TROPHOBLASTIC MALIGNANT TERATOMA
C0334528|T047||CCS_10|MALIGNANT TERATOMA, TROPHOBLASTIC
C0334528|T047||CCS_10|MALIGNANT TERATOMA, TROPHOBLASTIC (MORPHOLOGIC ABNORMALITY)
C0334528|T047||CCS_10|MALIGNANT; TERATOMA, TROPHOBLASTIC, UNSPECIFIED SITE
C0334528|T047||CCS_10|TERATOMA; MALIGNANT, TROPHOBLASTIC, UNSPECIFIED SITE
C0014145|T047||CCS_10|ENDODERMAL SINUS TUMOR
C0014145|T047||CCS_10|ENDODERMAL SINUS TUMORS
C0014145|T047||CCS_10|TUMOR, ENDODERMAL SINUS
C0014145|T047||CCS_10|TUMOR, YOLK SAC
C0014145|T047||CCS_10|TUMORS, ENDODERMAL SINUS
C0014145|T047||CCS_10|TUMORS, YOLK SAC
C0014145|T047||CCS_10|YOLK SAC TUMORS
C0014145|T047||CCS_10|YOLK SAC TUMOR 
C0014145|T047||CCS_10|YOLK SAC TUMOR
C0014145|T047||CCS_10|YOLK SAC TUMOUR SITE UNSPECIFIED
C0014145|T047||CCS_10|ENDODERMAL SINUS TUMOR [DISEASE/FINDING]
C0014145|T047||CCS_10|YOLK SAC TUMOR, MALIGNANT
C0014145|T047||CCS_10|YOLK SAC NEOPLASM
C0014145|T047||CCS_10|ENDODERMAL SINUS NEOPLASM
C0014145|T047||CCS_10|YOLK SAC TUMOR SITE UNSPECIFIED
C0014145|T047||CCS_10|ENDODERMAL SINUS TUMOUR SITE UNSPECIFIED
C0014145|T047||CCS_10|ENDODERMAL SINUS TUMOR SITE UNSPECIFIED
C0014145|T047||CCS_10|POLYVESICULAR VITELLINE TUMOR
C0014145|T047||CCS_10|ORCHIOBLASTOMA
C0014145|T047||CCS_10|EMBRYONAL CARCINOMA, INFANTILE
C0014145|T047||CCS_10|ENDODERMAL SINUS TUMOUR
C0014145|T047||CCS_10|INFANTILE EMBRYONAL CARCINOMA
C0014145|T047||CCS_10|POLYVESICULAR VITELLINE TUMOUR
C0014145|T047||CCS_10|YOLK SAC TUMOUR
C0014145|T047||CCS_10|ENDODERMAL SINUS TUMOR (MORPHOLOGIC ABNORMALITY)
C0014145|T047||CCS_10|HEPATOID YOLK SAC TUMOR
C0014145|T047||CCS_10|HEPATOID YOLK SAC TUMOUR
C0014145|T047||CCS_10|YOLK SAC TUMOR 
C1405366|T047||CCS_10|POLYVESICULAR; TUMOR, UNSPECIFIED SITE, MALE
C1405366|T047||CCS_10|TUMOR; POLYVESICULAR, UNSPECIFIED SITE, MALE
C1409893|T047||CCS_10|SEMINOMA; UNSPECIFIED SITE
C1409893|T047||CCS_10|SPERMATOCYTOMA; UNSPECIFIED SITE
C1409698|T047||CCS_10|SEMINOMA; SPERMATOCYTIC, UNSPECIFIED SITE
C1409698|T047||CCS_10|SPERMATOCYTIC; SEMINOMA, UNSPECIFIED SITE
C0238451|T047||CCS_10|TERATOMA, TESTICULAR
C0238451|T047||CCS_10|TESTICULAR TERATOMA
C0238451|T047||CCS_10|TERATOMA OF TESTIS
C0238451|T047||CCS_10|TERATOMA OF TESTIS 
C0238451|T047||CCS_10|TERATOMA OF TESTES
C0238451|T047||CCS_10|TERATOMA OF THE TESTIS
C0238451|T047||CCS_10|TESTICLE CANCER, TERATOMA
C0238451|T047||CCS_10|TESTICULAR CANCER, TERATOMA
C0238451|T047||CCS_10|TESTIS CANCER, TERATOMA
C0238451|T047||CCS_10|TERATOMA; TESTIS
C0238451|T047||CCS_10|TESTIS; TERATOMA
C0280256|T047||CCS_10|STAGE, TESTICULAR CANCER
C0280256|T047||CCS_10|TESTICULAR CANCER STAGE
C0279869|T047||CCS_10|CELLULAR DIAGNOSIS, TESTICULAR CANCER
C0279869|T047||CCS_10|TESTICULAR CANCER CELLULAR DIAGNOSIS
C1336711|T047||CCS_10|TESTICULAR LEUKEMIA
C1515289|T047||CCS_10|MALIGNANT TESTICULAR SEX CORD-STROMAL TUMOR
C2212316|T047||CCS_10|MAST CELL SARCOMA OF TESTIS 
C2212316|T047||CCS_10|MAST CELL SARCOMA OF TESTIS
C2057633|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF TESTIS
C2057633|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF TESTIS 
C0153597|T047||CCS_10|MALIGNANT NEOPLASM OF PENIS AND OTHER MALE GENITAL ORGANS
C0153597|T047||CCS_10|MALIGNANT NEOPLASM OF PENIS AND OTHER MALE GENITAL ORGANS 
C0153597|T047||CCS_10|MALIGNANT NEOPLASM OF PENIS AND OTHER MALE GENITAL ORGAN NOS
C0153597|T047||CCS_10|MALIGNANT NEOPLASM OF PENIS AND OTHER MALE GENITAL ORGAN NOS 
C0376358|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE
C0376358|T047||CCS_10|PROSTATE CANCER
C0376358|T047||CCS_10|PROSTATIC CANCER
C0376358|T047||CCS_10|CANCER OF PROSTATE
C0376358|T047||CCS_10|CANCER, PROSTATE
C0376358|T047||CCS_10|CANCERS, PROSTATE
C0376358|T047||CCS_10|PROSTATE CANCERS
C0376358|T047||CCS_10|CANCER, PROSTATIC
C0376358|T047||CCS_10|CANCERS, PROSTATIC
C0376358|T047||CCS_10|PROSTATIC CANCERS
C0376358|T047||CCS_10|PROSTATE CANCER 
C0376358|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE GLAND 
C0376358|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE GLAND
C0376358|T047||CCS_10|CA PROSTATE
C0376358|T047||CCS_10|MALIGNANT TUMOR OF PROSTATE GLAND
C0376358|T047||CCS_10|MALIGN NEOPL PROSTATE
C0376358|T047||CCS_10|PROSTATIC NEOPLASMS MALIGNANT
C0376358|T047||CCS_10|MALIGNANT PROSTATIC TUMOR
C0376358|T047||CCS_10|MALIGNANT TUMOUR OF PROSTATE
C0376358|T047||CCS_10|CA - CANCER OF PROSTATE
C0376358|T047||CCS_10|MALIGNANT TUMOR OF PROSTATE
C0376358|T047||CCS_10|MALIGNANT PROSTATIC TUMOUR
C0376358|T047||CCS_10|MALIGNANT TUMOR OF PROSTATE 
C0376358|T047||CCS_10|PROSTATE--CANCER
C0376358|T047||CCS_10|-- PROSTATE CANCER
C0376358|T047||CCS_10|PROSTATE CANCER NOS
C0376358|T047||CCS_10|CANCER OF THE PROSTATE
C0376358|T047||CCS_10|MALIGNANT NEOPLASM OF THE PROSTATE
C0376358|T047||CCS_10|MALIGNANT PROSTATE NEOPLASM
C0376358|T047||CCS_10|MALIGNANT PROSTATE TUMOR
C0376358|T047||CCS_10|MALIGNANT TUMOR OF THE PROSTATE
C0376358|T047||CCS_10|NEOPLASM MALIG;PROSTATE
C0376358|T047||CCS_10|MALIGNANT NEOSPLASM OF THE PROSTATE
C0497581|T047|31|CCS_10|MALIGNANT NEOPLASM OF OTHER AND UNSPECIFIED MALE GENITAL ORGANS|CANCER OF OTHER MALE GENITAL ORGANS
C0497581|T047|31|CCS_10|OTHER MALE GENITAL MALIGNANT NEOPLASM|CANCER OF OTHER MALE GENITAL ORGANS
C0497581|T047|31|CCS_10|CANCER OF OTHER MALE GENITAL ORGANS|CANCER OF OTHER MALE GENITAL ORGANS
C0497581|T047|31|CCS_10|MALIGNANT NEOPLASM OF OTHER MALE GENITAL ORGAN|CANCER OF OTHER MALE GENITAL ORGANS
C0497581|T047|31|CCS_10|MALIGNANT NEOPLASM OF OTHER MALE GENITAL ORGAN NOS |CANCER OF OTHER MALE GENITAL ORGANS
C0497581|T047|31|CCS_10|MALIGNANT NEOPLASM OF OTHER MALE GENITAL ORGAN NOS|CANCER OF OTHER MALE GENITAL ORGANS
C0497581|T047|31|CCS_10|MALIGNANT NEOPLASM OF OTHER MALE GENITAL ORGAN |CANCER OF OTHER MALE GENITAL ORGANS
C0153601|T047||CCS_10|MALIGNANT NEOPLASM OF PENIS
C0153601|T047||CCS_10|MALIGNANT NEOPLASM OF PENIS, UNSPECIFIED
C0153601|T047||CCS_10|MALIGNANT NEOPLASM OF PENIS 
C0153601|T047||CCS_10|MALIGNANT PENILE NEOPLASM
C0153601|T047||CCS_10|CANCER, PENILE
C0153601|T047||CCS_10|CANCERS, PENILE
C0153601|T047||CCS_10|PENILE CANCERS
C0153601|T047||CCS_10|CANCERS, PENIS
C0153601|T047||CCS_10|PENIS CANCERS
C0153601|T047||CCS_10|MALIGNANT TUMOR OF PENIS
C0153601|T047||CCS_10|PENILE CANCER
C0153601|T047||CCS_10|MALIG NEO PENIS NOS
C0153601|T047||CCS_10|CANCER, PENIS
C0153601|T047||CCS_10|PENILE NEOPLASMS MALIGNANT
C0153601|T047||CCS_10|CA PENIS 
C0153601|T047||CCS_10|MALIGNANT NEOPLASM OF PENIS, PART UNSPECIFIED 
C0153601|T047||CCS_10|CA PENIS
C0153601|T047||CCS_10|MALIGNANT NEOPLASM OF PENIS, PART UNSPECIFIED
C0153601|T047||CCS_10|CANCER OF PENIS
C0153601|T047||CCS_10|PENILE CA
C0153601|T047||CCS_10|CA - CANCER OF PENIS
C0153601|T047||CCS_10|MALIGNANT TUMOUR OF PENIS
C0153601|T047||CCS_10|PENIS--CANCER
C0153601|T047||CCS_10|PENILE MALIGNANT NEOPLASM NOS
C0153601|T047||CCS_10|PENILE MALIGNANT NEOPLASM
C0153601|T047||CCS_10|PENIS CANCER
C0153601|T047||CCS_10|CANCER OF THE PENIS
C0153601|T047||CCS_10|MALIGNANT TUMOR OF PENIS 
C0153601|T047||CCS_10|MALIGNANT NEOPLASM OF PENIS, NOS
C0153601|T047||CCS_10|MALIGNANT NEOPLASM OF THE PENIS
C0153601|T047||CCS_10|MALIGNANT PENILE TUMOR
C0153601|T047||CCS_10|MALIGNANT TUMOR OF THE PENIS
C0153606|T047|2.8|CCS_10|MALIGNANT NEOPLASM OF MALE GENITAL ORGAN, UNSPECIFIED|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALIGNANT TUMOR OF MALE GENITAL ORGAN|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALIGNANT NEOPLASM OF MALE GENITAL ORGAN|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALE GENITAL CANCER|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALE GENITAL CANCER |CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALIGNANT NEOPLASMS OF MALE GENITAL ORGANS|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALIGNANT TUMOR OF MALE GENITALIA|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MAL NEO MALE GENITAL NOS|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|CANCER OF MALE GENITAL ORGANS|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALIGNANT NEOPLASMS OF MALE GENITAL ORGANS (C60-C63)|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALIGNANT NEOPLASM OF MALE GENITALIA|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALIGNANT NEOPLASM OF THE MALE GENITAL ORGANS |CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALIGNANT NEOPLASM OF THE MALE GENITAL ORGANS|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALIGNANT NEOPLASM OF MALE GENITAL ORGANS|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|GENITAL CANCER MALE|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|[X]MALIGNANT NEOPLASM OF MALE GENITAL ORGANS |CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|[X]MALIGNANT NEOPLASM OF MALE GENITAL ORGAN, UNSPECIFIED |CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|[X]MALIGNANT NEOPLASM OF MALE GENITAL ORGAN, UNSPECIFIED|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|[X]MALIGNANT NEOPLASM OF MALE GENITAL ORGANS|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALE REPROD. SYSTEM CANCER, NOS|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALE REPRODUCTIVE SYSTEM CANCER, NOS|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALIGNANT NEOPLASM OF MALE GENITAL ORGAN, SITE UNSPECIFIED|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALIGNANT TUMOUR OF MALE GENITAL ORGAN|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALIGNANT TUMOR OF MALE GENITAL ORGAN |CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALIGNANT NEOPLASM OF MALE GENITAL ORGAN, NOS|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALIGNANT MALE REPRODUCTIVE SYSTEM NEOPLASM|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALIGNANT MALE REPRODUCTIVE SYSTEM TUMOR|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALIGNANT NEOPLASM OF MALE REPRODUCTIVE SYSTEM|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALIGNANT NEOPLASM OF THE MALE REPRODUCTIVE SYSTEM|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALIGNANT TUMOR OF MALE REPRODUCTIVE SYSTEM|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALIGNANT TUMOR OF THE MALE REPRODUCTIVE SYSTEM|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALIGNANT NEOPLASM OF MALE GENITAL ORGAN OR TRACT NOS|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|NEOPLASM MALIG;GENITAL SYS;M|CANCER OF MALE GENITAL ORGANS
C0153606|T047|2.8|CCS_10|MALIGNANT NEOSPLASM OF THE MALE GENITAL SYSTEM|CANCER OF MALE GENITAL ORGANS
C2217869|T047||CCS_10|MALE GENITAL NEOPLASM MALIGNANT SMALL CELL TYPE
C2217869|T047||CCS_10|MALIGNANT SMALL CELL NEOPLASM OF MALE GENITALIA
C2217869|T047||CCS_10|MALIGNANT SMALL CELL NEOPLASM OF MALE GENITALIA 
C2011384|T047||CCS_10|GIANT CELL TYPE NEOPLASM OF MALE GENITALIA 
C2011384|T047||CCS_10|GIANT CELL TYPE NEOPLASM OF MALE GENITALIA
C2018667|T047||CCS_10|SPINDLE CELL TYPE NEOPLASM OF MALE GENITALIA
C2018667|T047||CCS_10|SPINDLE CELL TYPE NEOPLASM OF MALE GENITALIA 
C2075627|T047||CCS_10|CLEAR CELL TYPE NEOPLASM OF MALE GENITALIA
C2075627|T047||CCS_10|CLEAR CELL TYPE NEOPLASM OF MALE GENITALIA 
C2007032|T047||CCS_10|CARCINOMA OF MALE GENITALIA
C2007032|T047||CCS_10|CARCINOMA OF MALE GENITALIA 
C2215312|T047||CCS_10|ADENOCARCINOMA OF MALE GENITALIA
C2215312|T047||CCS_10|ADENOCARCINOMA OF MALE GENITALIA 
C2219527|T047||CCS_10|SARCOMA OF MALE GENITALIA 
C2219527|T047||CCS_10|SARCOMA OF MALE GENITALIA
C2230877|T047||CCS_10|FIBROSARCOMA OF MALE GENITALIA 
C2230877|T047||CCS_10|FIBROSARCOMA OF MALE GENITALIA
C2184067|T047||CCS_10|LIPOSARCOMA OF MALE GENITALIA 
C2184067|T047||CCS_10|LIPOSARCOMA OF MALE GENITALIA
C2230880|T047||CCS_10|MYOSARCOMA OF MALE GENITALIA
C2230880|T047||CCS_10|MYOSARCOMA OF MALE GENITALIA 
C2007077|T047||CCS_10|CARCINOSARCOMA OF MALE GENITALIA
C2007077|T047||CCS_10|CARCINOSARCOMA OF MALE GENITALIA 
C2216612|T047||CCS_10|MALIGNANT MESENCHYMOMA OF MALE GENITALIA
C2216612|T047||CCS_10|MALIGNANT MESENCHYMOMA OF MALE GENITALIA 
C2216469|T047||CCS_10|MARGINAL ZONE B-CELL LYMPHOMA OF MALE GENITALIA
C2216469|T047||CCS_10|MARGINAL ZONE B-CELL LYMPHOMA OF MALE GENITALIA 
C2216535|T047||CCS_10|MALIGNANT FIBROUS HISTIOCYTOMA OF MALE GENITALIA
C2216535|T047||CCS_10|MALIGNANT FIBROUS HISTIOCYTOMA OF MALE GENITALIA 
C2230882|T047||CCS_10|MULLERIAN MIXED TUMOR OF MALE GENITALIA 
C2230882|T047||CCS_10|MULLERIAN MIXED TUMOR OF MALE GENITALIA
C2216616|T047||CCS_10|MALIGNANT MESODERMAL MIXED TUMOR OF MALE GENITALIA 
C2216616|T047||CCS_10|MALIGNANT MESODERMAL MIXED TUMOR OF MALE GENITALIA
C2188071|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF MALE GENITALIA 
C2188071|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF MALE GENITALIA
C2230874|T047||CCS_10|BASALOID CARCINOMA OF MALE GENITALIA
C2230874|T047||CCS_10|BASALOID CARCINOMA OF MALE GENITALIA 
C2230874|T047||CCS_10|BASALOID CARCINOMA OF MALE GENITAL TRACT
C2216459|T047||CCS_10|FIBROBLASTIC LIPOSARCOMA OF MALE GENITALIA 
C2216459|T047||CCS_10|FIBROBLASTIC LIPOSARCOMA OF MALE GENITALIA
C1306367|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF MALE GENITAL ORGAN 
C1306367|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF MALE GENITAL ORGAN
C1306367|T047||CCS_10|MALE GENITAL MALIGNANT NEOPLASM PRIMARY
C1306367|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF MALE GENITAL ORGAN 
C0348369|T047||CCS_10|MALIGNANT NEOPLASM OVERLAPPING MALE GENITAL ORGAN SITE
C0348369|T047||CCS_10|OVERLAPPING LESION OF MALE GENITAL ORGANS
C0348369|T047||CCS_10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF MALE GENITAL ORGANS
C0348369|T047||CCS_10|MALIGNANT NEOPLASM OF OVRLP SITES OF MALE GENITAL ORGANS
C0348369|T047||CCS_10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF MALE GENITAL ORGANS 
C0348369|T047||CCS_10|MALE GENITAL NEOPLASM MALIGNANT OVERLAPPING SITES
C0348369|T047||CCS_10|MALIGNANT NEOPLASM, OVERLAPPING LESION OF MALE GENITAL ORGANS
C0348369|T047||CCS_10|[X]MALIGNANT NEOPLASM OF OVERLAPPING LESION OF MALE GENITAL ORGANS
C0348369|T047||CCS_10|[X]MALIGNANT NEOPLASM OF OVERLAPPING LESION OF MALE GENITAL ORGANS 
C0348369|T047||CCS_10|MALIGNANT NEOPLASM, OVERLAPPING LESION OF MALE GENITAL ORGANS 
C0348369|T047||CCS_10|OVERLAPPING MALIGNANT NEOPLASM OF MALE GENITAL ORGANS 
C0348369|T047||CCS_10|OVERLAPPING MALIGNANT NEOPLASM OF MALE GENITAL ORGANS
C0686232|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF VAS DEFERENS
C0686232|T047||CCS_10|SPERMATIC CORD NEOPLASM MALIGNANT VAS DEFERENS SECONDARY
C0686232|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF VAS DEFERENS 
C0686232|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO VAS DEFERENS
C0686232|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF VAS DEFERENS 
C0864963|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF SCROTUM
C0864963|T047||CCS_10|CANCER OF SCROTAL SKIN
C0864963|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF SCROTUM 
C0864963|T047||CCS_10|SCROTAL NEOPLASM MALIGNANT OF SKIN
C0864963|T047||CCS_10|MALIGNANT NEOPLASM OF SCROTAL SKIN
C0864963|T047||CCS_10|MALIGNANT NEOPLASM OF SCROTAL SKIN 
C0346225|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF PENIS NOS
C0346225|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF PENIS
C0346225|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF PENIS 
C0346225|T047||CCS_10|PENILE NEOPLASM MALIGNANT OF SKIN
C0346225|T047||CCS_10|CANCER OF PENILE SKIN
C0346225|T047||CCS_10|MALIGNANT TUMOR OF PENILE SKIN
C0346225|T047||CCS_10|MALIGNANT TUMOR OF SKIN OF PENIS
C0346225|T047||CCS_10|MALIGNANT TUMOUR OF PENILE SKIN
C0346225|T047||CCS_10|MALIGNANT TUMOUR OF SKIN OF PENIS
C0346225|T047||CCS_10|MALIGNANT TUMOR OF SKIN OF PENIS 
C0153602|T047||CCS_10|MALIGNANT NEOPLASM OF EPIDIDYMIS
C0153602|T047||CCS_10|MALIGNANT TUMOR OF EPIDIDYMIS
C0153602|T047||CCS_10|MALIGNANT NEOPLASM OF EPIDIDYMIS 
C0153602|T047||CCS_10|CANCER OF EPIDIDYMIS
C0153602|T047||CCS_10|MALIG NEO EPIDIDYMIS
C0153602|T047||CCS_10|EPIDIDYMAL CANCER
C0153602|T047||CCS_10|MALIGNANT EPIDIDYMAL NEOPLASM NOS
C0153602|T047||CCS_10|MALIGNANT TUMOUR OF EPIDIDYMIS
C0153602|T047||CCS_10|MALIGNANT TUMOR OF EPIDIDYMIS 
C0153602|T047||CCS_10|MALIGNANT EPIDIDYMAL NEOPLASM
C0153602|T047||CCS_10|MALIGNANT EPIDIDYMAL TUMOR
C0153602|T047||CCS_10|MALIGNANT NEOPLASM OF THE EPIDIDYMIS
C0153602|T047||CCS_10|MALIGNANT TUMOR OF THE EPIDIDYMIS
C0346216|T047||CCS_10|MALIGNANT NEOPLASM OF SEMINAL VESICLE 
C0346216|T047||CCS_10|MALIGNANT NEOPLASM OF SEMINAL VESICLE
C0346216|T047||CCS_10|MALIGNANT TUMOR OF SEMINAL VESICLE
C0346216|T047||CCS_10|MALIGNANT TUMOUR OF SEMINAL VESICLE
C0346216|T047||CCS_10|MALIGNANT TUMOR OF SEMINAL VESICLE 
C0153603|T047||CCS_10|MALIGNANT NEOPLASM OF SPERMATIC CORD
C0153603|T047||CCS_10|MALIGNANT NEOPLASM OF SPERMATIC CORD 
C0153603|T047||CCS_10|MALIGNANT TUMOR OF SPERMATIC CORD
C0153603|T047||CCS_10|MAL NEO SPERMATIC CORD
C0153603|T047||CCS_10|SPERMATIC CORD CA
C0153603|T047||CCS_10|MALIGNANT TUMOUR OF SPERMATIC CORD
C0153603|T047||CCS_10|MALIGNANT TUMOR OF SPERMATIC CORD 
C0153603|T047||CCS_10|MALIGNANT NEOPLASM OF THE SPERMATIC CORD
C0153603|T047||CCS_10|MALIGNANT SPERMATIC CORD NEOPLASM
C0153603|T047||CCS_10|MALIGNANT SPERMATIC CORD TUMOR
C0153603|T047||CCS_10|MALIGNANT TUMOR OF THE SPERMATIC CORD
C0347000|T047||CCS_10|MALE GENITAL MALIGNANT NEOPLASM SECONDARY
C0347000|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF MALE GENITAL ORGAN 
C0347000|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF MALE GENITAL ORGAN
C0347000|T047||CCS_10|CANCER METASTATIC TO MALE GENITAL ORGAN
C0347000|T047||CCS_10|CANCER METASTATIC TO MALE GENITALIA
C0347000|T047||CCS_10|METASTASIS TO MALE GENITAL ORGAN
C0347000|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO MALE GENITAL ORGAN
C0347000|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF MALE GENITAL ORGAN 
C0347000|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO MALE GENITAL ORGAN, NOS
C0347000|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF MALE GENITAL ORGAN, NOS
C0348368|T047||CCS_10|MALIGNANT NEOPLASM OF OTHER SPECIFIED MALE GENITAL ORGANS
C0348368|T047||CCS_10|OTHER SPECIFIED MALE GENITAL ORGANS
C0348368|T047||CCS_10|[X]MALIGNANT NEOPLASM OF OTHER SPECIFIED MALE GENITAL ORGANS
C0348368|T047||CCS_10|[X]MALIGNANT NEOPLASM OF OTHER SPECIFIED MALE GENITAL ORGANS 
C1398495|T047||CCS_10|GENITAL ORGANS; MELANOMA, MALE (EXTERNAL)
C1398495|T047||CCS_10|MELANOMA; GENITAL ORGANS, MALE (EXTERNAL)
C0863024|T047||CCS_10|ADENOCARCINOMA OF THE RETE TESTIS
C0863024|T047||CCS_10|ADENOCARCINOMA OF RETE TESTIS
C0863024|T047||CCS_10|RETE TESTIS ADENOCARCINOMA
C1519233|T047||CCS_10|SEMINAL VESICLE ADENOCARCINOMA
C1335705|T047||CCS_10|RECURRENT MALE REPRODUCTIVE SYSTEM CARCINOMA
C1335705|T047||CCS_10|RECURRENT MALE REPRODUCTIVE SYSTEM CANCER
C0746787|T047||CCS_10|MALIGNANT NEOPLASM OF NECK
C0746787|T047||CCS_10|NECK CANCER
C0746787|T047||CCS_10|MALIGNANT NEOPLASM OF NECK 
C0746787|T047||CCS_10|MALIGNANT NEOPLASM OF NECK NOS
C0746787|T047||CCS_10|MALIGNANT NEOPLASM OF NECK NOS 
C0746787|T047||CCS_10|NECK--CANCER
C0746787|T047||CCS_10|CANCER OF NECK
C0746787|T047||CCS_10|CANCER OF THE NECK
C0746787|T047||CCS_10|MALIGNANT TUMOR OF NECK
C0746787|T047||CCS_10|MALIGNANT TUMOUR OF NECK
C0746787|T047||CCS_10|MALIGNANT TUMOR OF NECK 
C0746787|T047||CCS_10|MALIGNANT NEOPLASM OF NECK, NOS
C0746787|T047||CCS_10|MALIGNANT NECK NEOPLASM
C0746787|T047||CCS_10|MALIGNANT NECK TUMOR
C0746787|T047||CCS_10|MALIGNANT NEOPLASM OF THE NECK
C0746787|T047||CCS_10|MALIGNANT TUMOR OF THE NECK
C2711842|T047||CCS_10|ADENOCARCINOMA OF HEAD AND NECK
C2711842|T047||CCS_10|ADENOCARCINOMA OF HEAD AND NECK 
C2711842|T047||CCS_10|ADENOCARCINOMA OF HEAD AND NECK 
C2711842|T047||CCS_10|MALIGNANT NEOPLASM OF ILL-DEFINED SITE HEAD AND NECK ADENOCARCINOMA
C1263914|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF FACE 
C1263914|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF FACE
C1263914|T047||CCS_10|NEOPLASM - PNS MALIGNANT FACE PRIMARY
C1263914|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF FACE 
C0153744|T047||CCS_10|HODGKIN'S SARCOMA OF LYMPH NODES OF HEAD, FACE, AND NECK
C0153744|T047||CCS_10|HODGKINS SARCOMA HEAD
C0153744|T047||CCS_10|HODGKIN SARCOMA OF LYMPH NODES OF HEAD, FACE AND NECK
C0153744|T047||CCS_10|HODGKIN SARCOMA OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0153744|T047||CCS_10|HODGKIN'S SARCOMA INVOLVING LYMPH NODES OF HEAD, FACE, AND NECK
C0153744|T047||CCS_10|HODGKIN'S SARCOMA, LYMPH NODES OF HEAD, FACE, AND NECK
C0153744|T047||CCS_10|HODGKIN SARCOMA OF LYMPH NODES OF HEAD, FACE, OR NECK
C0153744|T047||CCS_10|HODGKIN SARCOMA OF LYMPH NODES OF HEAD, FACE, OR NECK 
C0153744|T047||CCS_10|HODGKIN'S SARCOMA OF LYMPH NODES OF HEAD, FACE AND NECK
C0153744|T047||CCS_10|HODGKIN'S SARCOMA OF LYMPH NODES OF HEAD, FACE AND/OR NECK 
C0153744|T047||CCS_10|HODGKIN'S SARCOMA OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0153744|T047||CCS_10|HODGKIN'S SARCOMA OF LYMPH NODES OF HEAD, FACE AND NECK 
C0153744|T047||CCS_10|HODGKIN'S SARCOMA INVOLVING LYMPH NODES OF HEAD, FACE AND NECK
C0587226|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF TONGUE 
C0587226|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF TONGUE
C0587226|T047||CCS_10|TONGUE CANCER METASTATIC
C0587226|T047||CCS_10|TONGUE NEOPLASM MALIGNANT SECONDARY
C0587226|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF TONGUE 
C0587226|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO TONGUE
C0587226|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO TONGUE, NOS
C0587226|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF TONGUE, NOS
C0346931|T047||CCS_10|MALIGNANT NEOPLASM OF NASOLACRIMAL DUCT
C0346931|T047||CCS_10|MALIGNANT NEOPLASM OF NASOLACRIMAL DUCT 
C0346931|T047||CCS_10|MALIGNANT TUMOR OF NASOLACRIMAL DUCT
C0346931|T047||CCS_10|MALIGNANT NEOPLASM OF NASOLACRIMAL DUCT 
C0153379|T047||CCS_10|MALIGNANT NEOPLASM OF RETROMOLAR AREA
C0153379|T047||CCS_10|MALIGNANT NEOPLASM OF RETROMOLAR AREA 
C0153379|T047||CCS_10|MALIGNANT RETROMOLAR AREA NEOPLASM
C0153379|T047||CCS_10|MALIGNANT TUMOR OF RETROMOLAR AREA
C0153379|T047||CCS_10|MALIG NEO RETROMOLAR
C0153379|T047||CCS_10|MALIGNANT TUMOUR OF RETROMOLAR AREA
C0153379|T047||CCS_10|MALIGNANT TUMOR OF RETROMOLAR AREA 
C0349031|T047||CCS_10|MELANOMA IN SITU OF SCALP AND NECK
C0349031|T047||CCS_10|SKIN NEOPLASM MELANOMA IN SITU OF SCALP AND NECK
C0349031|T047||CCS_10|MELANOMA IN SITU OF SCALP AND NECK 
C0349031|T047||CCS_10|MELANOMA IN SITU OF SCALP AND NECK 
C0220636|T047||CCS_10|MALIGNANT NEOPLASM OF SALIVARY GLAND
C0220636|T047||CCS_10|MALIGNANT NEOPLASM OF SALIVARY GLAND DUCT
C0220636|T047||CCS_10|MALIGNANT NEOPLASM OF SALIVARY GLAND 
C0220636|T047||CCS_10|CANCERS, SALIVARY GLAND
C0220636|T047||CCS_10|SALIVARY GLAND CANCERS
C0220636|T047||CCS_10|MALIGNANT TUMOR OF SALIVARY GLAND
C0220636|T047||CCS_10|MAL NEO SALIVARY NOS
C0220636|T047||CCS_10|CANCER, SALIVARY GLAND
C0220636|T047||CCS_10|SALIVARY GLAND NEOPLASMS MALIGNANT
C0220636|T047||CCS_10|SALIVARY GLAND CANCER
C0220636|T047||CCS_10|SALIVARY GLANDS--CANCER
C0220636|T047||CCS_10|SALIVARY GLAND CANCER NOS
C0220636|T047||CCS_10|MALIGNANT SALIVARY GLAND CANCER
C0220636|T047||CCS_10|MALIGNANT SALIVARY GLAND NEOPLASM
C0220636|T047||CCS_10|MALIGNANT NEOPLASM OF SALIVARY GLAND, UNSPECIFIED
C0220636|T047||CCS_10|CANCER OF THE SALIVARY GLAND
C0220636|T047||CCS_10|CA - CANCER OF SALIVARY GLAND
C0220636|T047||CCS_10|CANCER OF SALIVARY GLAND
C0220636|T047||CCS_10|MALIGNANT TUMOUR OF SALIVARY GLAND
C0220636|T047||CCS_10|MALIGNANT TUMOR OF SALIVARY GLAND 
C0220636|T047||CCS_10|MALIGNANT NEOPLASM OF THE SALIVARY GLAND
C0220636|T047||CCS_10|MALIGNANT SALIVARY GLAND TUMOR
C0220636|T047||CCS_10|MALIGNANT TUMOR OF THE SALIVARY GLAND
C0220636|T047||CCS_10|MALIGNANT NEOPLASM OF SALIVARY GLAND NOS
C0684535|T047||CCS_10|BONE NEOPLASM, MALIGNANT - FACE SECONDARY
C0684535|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BONE OF FACE
C0684535|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BONE OF FACE 
C0684535|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO BONE OF FACE
C0684535|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BONE OF FACE 
C0684535|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO BONE OF FACE, NOS
C0684535|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BONE OF FACE, NOS
C0585362|T047||CCS_10|MALIGNANT SQUAMOUS CELL NEOPLASM OF ORAL CAVITY 
C0585362|T047||CCS_10|MALIGNANT SQUAMOUS CELL NEOPLASM OF ORAL CAVITY
C0585362|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE ORAL CAVITY
C0585362|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF MOUTH
C0585362|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF MOUTH 
C0585362|T047||CCS_10|MOUTH SCC
C0585362|T047||CCS_10|MOUTH SQUAMOUS CELL CARCINOMA
C0585362|T047||CCS_10|ORAL CAVITY SCC
C0585362|T047||CCS_10|ORAL CAVITY SQUAMOUS CELL CARCINOMA
C0585362|T047||CCS_10|SCC OF MOUTH
C0585362|T047||CCS_10|SCC OF ORAL CAVITY
C0585362|T047||CCS_10|SCC OF THE MOUTH
C0585362|T047||CCS_10|SCC OF THE ORAL CAVITY
C0585362|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF ORAL CAVITY
C0585362|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE MOUTH
C0686635|T047||CCS_10|SECONDARY AND UNSPECIFIED MALIGNANT NEOPLASM OF SUBMENTAL LYMPH NODES 
C0686635|T047||CCS_10|SECONDARY AND UNSPECIFIED MALIGNANT NEOPLASM OF SUBMENTAL LYMPH NODES
C0686635|T047||CCS_10|LYMPH NODE NEOPLASM MALIGNANT SECONDARY FACE SUBMENTAL
C0686635|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SUBMENTAL LYMPH NODES
C0686635|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SUBMENTAL LYMPH NODES 
C0686635|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO SUBMENTAL LYMPH NODES
C0686635|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SUBMENTAL LYMPH NODES 
C0153802|T047||CCS_10|MYCOSIS FUNGOIDES OF LYMPH NODES OF HEAD, FACE, AND NECK
C0153802|T047||CCS_10|MYCOSIS FUNGOIDES OF HEAD, FACE, AND NECK
C0153802|T047||CCS_10|MYCOSIS FUNGOIDES OF HEAD, FACE, AND NECK 
C0153802|T047||CCS_10|MYCOSIS FUNGOIDES HEAD
C0153802|T047||CCS_10|MYCOSIS FUNGOIDES, LYMPH NODES OF HEAD, FACE, AND NECK
C0153802|T047||CCS_10|MYCOSIS FUNGOIDES INVOLVING LYMPH NODES OF HEAD, FACE, AND NECK
C0153802|T047||CCS_10|MYCOSIS FUNGOIDES OF THE LYMPH NODES OF HEAD, FACE AND NECK 
C0153802|T047||CCS_10|MYCOSIS FUNGOIDES OF THE LYMPH NODES OF HEAD, FACE AND NECK
C0153802|T047||CCS_10|MYCOSIS FUNGOIDES OF LYMPH NODES OF HEAD, FACE AND/OR NECK 
C0153802|T047||CCS_10|MYCOSIS FUNGOIDES OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0153802|T047||CCS_10|MYCOSIS FUNGOIDES INVOLVING LYMPH NODES OF HEAD, FACE AND NECK
C0684747|T047||CCS_10|MALIGNANT NEOPLASM OF MUSCLE OF HEAD PRIMARY
C0684747|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF MUSCLE OF HEAD 
C0684747|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF MUSCLE OF HEAD
C0684747|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF MUSCLE OF HEAD 
C0339112|T047||CCS_10|BOWEN DISEASE OF EYELID
C0339112|T047||CCS_10|BOWEN'S DISEASE OF EYELID
C0339112|T047||CCS_10|BOWEN'S DISEASE OF EYELID 
C0339112|T047||CCS_10|BOWEN'S DISEASE OF EYELID 
C0686633|T047||CCS_10|SECONDARY AND UNSPECIFIED MALIGNANT NEOPLASM OF SUBMANDIBULAR LYMPH NODES 
C0686633|T047||CCS_10|SECONDARY AND UNSPECIFIED MALIGNANT NEOPLASM OF SUBMANDIBULAR LYMPH NODES
C0686633|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SUBMANDIBULAR LYMPH NODES
C0686633|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SUBMANDIBULAR LYMPH NODES 
C0686633|T047||CCS_10|LYMPH NODE NEOPLASM MALIGNANT SECONDARY NECK SUBMANDIBULAR
C0686633|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO SUBMANDIBULAR LYMPH NODES
C0686633|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SUBMANDIBULAR LYMPH NODES 
C0684530|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SPHENOID BONE
C0684530|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SPHENOID BONE 
C0684530|T047||CCS_10|BONE NEOPLASM, MALIGNANT - SKULL SPHENOID BONE SECONDARY
C0684530|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO SPHENOID BONE
C0684530|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SPHENOID BONE 
C0153712|T047||CCS_10|BURKITT'S LYMPHOMA OF LYMPH NODES OF HEAD, FACE, AND NECK 
C0153712|T047||CCS_10|BURKITT'S LYMPHOMA OF HEAD, FACE, AND NECK
C0153712|T047||CCS_10|BURKITT'S LYMPHOMA OF LYMPH NODES OF HEAD, FACE, AND NECK
C0153712|T047||CCS_10|BURKITT'S TUMOR HEAD
C0153712|T047||CCS_10|BURKITT LYMPHOMA OF LYMPH NODES OF HEAD, FACE AND NECK
C0153712|T047||CCS_10|BURKITT LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK
C0153712|T047||CCS_10|BURKITT'S TUMOR OR LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK
C0153712|T047||CCS_10|BURKITT'S TUMOR OR LYMPHOMA INVOLVING LYMPH NODES OF HEAD, FACE, AND NECK
C0153712|T047||CCS_10|BURKITT'S TUMOUR OR LYMPHOMA INVOLVING LYMPH NODES OF HEAD, FACE, AND NECK
C0153712|T047||CCS_10|BURKITT'S LYMPHOMA OF LYMPH NODES OF HEAD, FACE AND NECK
C0153712|T047||CCS_10|BURKITT'S LYMPHOMA OF LYMPH NODES OF HEAD, FACE AND NECK 
C0153712|T047||CCS_10|BURKITT'S TUMOR OR LYMPHOMA INVOLVING LYMPH NODES OF HEAD, FACE AND NECK
C0686010|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF ORAL CAVITY
C0686010|T047||CCS_10|ORAL CAVITY MALIGNANT NEOPLASM SECONDARY
C0686010|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF ORAL CAVITY 
C0686010|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO MOUTH
C0686010|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF MOUTH 
C0686010|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF MOUTH
C0686010|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO MOUTH, NOS
C0686010|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF MOUTH, NOS
C0563210|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF SKIN OF CHEEK
C0563210|T047||CCS_10|SKIN NEOPLASM FACE MALIGNANT SQUAMOUS CELL CARCINOMA CHEEK
C0563210|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF SKIN OF CHEEK 
C0563210|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF SKIN OF CHEEK 
C0684922|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF UPPER RESPIRATORY TRACT
C0684922|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF UPPER RESPIRATORY TRACT 
C0684922|T047||CCS_10|MALIGNANT NEOPLASM UPPER RESPIRATORY TRACT SECONDARY
C0684922|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO UPPER RESPIRATORY TRACT
C0684922|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF UPPER RESPIRATORY TRACT 
C0684922|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO UPPER RESPIRATORY TRACT, NOS
C0684922|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF UPPER RESPIRATORY TRACT, NOS
C1306049|T047||CCS_10|HYPOPHARYNGEAL NEOPLASM MALIGNANT POSTCRICOID REGION PRIMARY
C1306049|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF POSTCRICOID REGION
C1306049|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF POSTCRICOID REGION 
C1306049|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF POSTCRICOID REGION 
C0153728|T047||CCS_10|HODGKIN'S PARAGRANULOMA OF LYMPH NODES OF HEAD, FACE, AND NECK
C0153728|T047||CCS_10|HODGKINS PARAGRAN HEAD
C0153728|T047||CCS_10|HODGKIN PARAGRANULOMA OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0153728|T047||CCS_10|HODGKIN'S PARAGRANULOMA, LYMPH NODES OF HEAD, FACE, AND NECK
C0153728|T047||CCS_10|HODGKIN'S PARAGRANULOMA INVOLVING LYMPH NODES OF HEAD, FACE, AND NECK
C0153728|T047||CCS_10|HODGKIN'S PARAGRANULOMA OF LYMPH NODES OF HEAD, FACE, AND NECK 
C0153728|T047||CCS_10|HODGKIN DISEASE PARAGRANULOMA - HEAD, FACE, & NECK
C0153728|T047||CCS_10|HODGKIN PARAGRANULOMA OF LYMPH NODES OF HEAD, FACE, & NECK 
C0153728|T047||CCS_10|HODGKIN PARAGRANULOMA OF LYMPH NODES OF HEAD, FACE, & NECK
C0153728|T047||CCS_10|HODGKIN'S PARAGRANULOMA OF LYMPH NODES OF HEAD, FACE AND/OR NECK 
C0153728|T047||CCS_10|HODGKIN'S PARAGRANULOMA OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0153728|T047||CCS_10|HODGKIN'S PARAGRANULOMA INVOLVING LYMPH NODES OF HEAD, FACE AND NECK
C0686024|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF PALATE
C0686024|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF PALATE 
C0686024|T047||CCS_10|PALATE NEOPLASM MALIGNANT SECONDARY
C0686024|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO PALATE
C0686024|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF PALATE 
C0686024|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO PALATE, NOS
C0686024|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF PALATE, NOS
C0686492|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF MASTOID AIR CELLS 
C0686492|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF MASTOID AIR CELLS
C0686492|T047||CCS_10|BONE NEOPLASM, MALIGNANT - SKULL AND FACE, MASTOID AIR CELLS SECONDARY
C0686492|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO MASTOID AIR CELLS
C0686492|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF MASTOID AIR CELLS 
C1304846|T047||CCS_10|MALIGNANT NEOPLASM OF NECK PRIMARY
C1304846|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF NECK
C1304846|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF NECK 
C1304846|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF NECK 
C0346980|T047||CCS_10|SECONDARY MALIGNANT SKIN NEOPLASM OF HEAD 
C0346980|T047||CCS_10|SKIN NEOPLASM HEAD SECONDARY
C0346980|T047||CCS_10|SECONDARY MALIGNANT SKIN NEOPLASM OF HEAD
C0346980|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SKIN OF HEAD
C0346980|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SKIN OF HEAD 
C0496755|T047||CCS_10|MALIGNANT NEOPLASM OF TIP AND LATERAL BORDER OF TONGUE
C0496755|T047||CCS_10|MALIGNANT NEOPLASM OF BORDER OF TONGUE
C0496755|T047||CCS_10|MALIGNANT NEOPLASM OF TIP AND LATERAL BORDER OF TONGUE 
C0496755|T047||CCS_10|MALIGNANT TUMOR OF TIP AND LATERAL BORDER OF TONGUE
C0496755|T047||CCS_10|MAL NEO TIP/LAT TONGUE
C0496755|T047||CCS_10|MALIGNANT NEOPLASM OF TIP AND/OR LATERAL BORDER OF TONGUE
C0496755|T047||CCS_10|TONGUE NEOPLASM MALIGNANT BORDER
C0496755|T047||CCS_10|MALIGNANT NEOPLASM OF BORDER OF TONGUE 
C0496755|T047||CCS_10|MALIGNANT NEOPLASM OF TONGUE, TIP AND LATERAL BORDER
C0496755|T047||CCS_10|MALIGNANT NEOPLASM OF BORDER OF TONGUE 
C0496755|T047||CCS_10|MALIGNANT NEOPLASM OF TONGUE, TIP AND LATERAL BORDER 
C0685133|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BLOOD VESSEL OF FACE
C0685133|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BLOOD VESSEL OF FACE 
C0685133|T047||CCS_10|NEOPLASM - SOFT TISSUE TYPES BLOOD VESSEL MALIGNANT OF FACE SECONDARY
C0685133|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO BLOOD VESSEL OF FACE
C0685133|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BLOOD VESSEL OF FACE 
C0153644|T047||CCS_10|MALIGNANT CRANIAL NERVE NEOPL
C0153644|T047||CCS_10|CRANIAL NERVE NEOPL MALIGNANT
C0153644|T047||CCS_10|NEOPL CRANIAL NERVE MALIGNANT
C0153644|T047||CCS_10|MALIGNANT NEOPLASM OF CRANIAL NERVE
C0153644|T047||CCS_10|MALIGNANT NEOPLASM OF CRANIAL NERVE 
C0153644|T047||CCS_10|MALIGNANT TUMOR OF CRANIAL NERVE
C0153644|T047||CCS_10|MAL NEO CRANIAL NERVES
C0153644|T047||CCS_10|MALIGNANT NEOPLASM OF CRANIAL NERVE NOS
C0153644|T047||CCS_10|MALIGNANT NEOPLASM OF CRANIAL NERVES NOS
C0153644|T047||CCS_10|MALIGNANT NEOPLASM OF CRANIAL NERVES NOS 
C0153644|T047||CCS_10|MALIGNANT NEOPLASM OF CRANIAL NERVES
C0153644|T047||CCS_10|MALIGNANT CRANIAL NERVE NEOPLASM NOS
C0153644|T047||CCS_10|MALIGNANT CRANIAL NERVE NEOPLASM
C0153644|T047||CCS_10|TUMORS, CRANIAL NERVE, MALIGNANT
C0153644|T047||CCS_10|MALIGNANT CRANIAL NERVE TUMORS
C0153644|T047||CCS_10|MALIGNANT CRANIAL NERVE NEOPLASMS
C0153644|T047||CCS_10|NEOPLASMS, CRANIAL NERVE, MALIGNANT
C0153644|T047||CCS_10|CRANIAL NERVE TUMORS, MALIGNANT
C0153644|T047||CCS_10|CRANIAL NERVE NEOPLASMS, MALIGNANT
C0153644|T047||CCS_10|MALIGNANT TUMOUR OF CRANIAL NERVE
C0153644|T047||CCS_10|MALIGNANT TUMOR OF CRANIAL NERVE 
C0153644|T047||CCS_10|MALIGNANT NEOPLASM OF CRANIAL NERVE, NOS
C0153644|T047||CCS_10|CRANIAL NERVE NEOPLASM, MALIGNANT
C0153644|T047||CCS_10|MALIGNANT CRANIAL NERVE TUMOR
C0153644|T047||CCS_10|MALIGNANT NEOPLASM OF THE CRANIAL NERVE
C0153644|T047||CCS_10|MALIGNANT TUMOR OF THE CRANIAL NERVE
C0686408|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF CRANIAL NERVE
C0686408|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF CRANIAL NERVE 
C0686408|T047||CCS_10|CRANIAL NERVE NEOPLASM MALIGNANT SECONDARY
C0686408|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO CRANIAL NERVE
C0686408|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF CRANIAL NERVE 
C0686408|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO CRANIAL NERVE, NOS
C0686408|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF CRANIAL NERVE, NOS
C0153696|T047||CCS_10|RETICULOSARCOMA HEAD
C0153696|T047||CCS_10|RETICULOSARCOMA, LYMPH NODES OF HEAD, FACE, AND NECK
C0153696|T047||CCS_10|RETICULOSARCOMA INVOLVING LYMPH NODES OF HEAD, FACE, AND NECK
C0153696|T047||CCS_10|RETICULOSARCOMA OF LYMPH NODES OF HEAD, FACE, AND NECK 
C0153696|T047||CCS_10|RETICULOSARCOMA OF LYMPH NODES OF HEAD, FACE, AND NECK
C0153696|T047||CCS_10|RETICULOSARCOMA OF LYMPH NODES OF HEAD, FACE AND NECK
C0153696|T047||CCS_10|RETICULOSARCOMA OF LYMPH NODES OF HEAD, FACE AND NECK 
C0153696|T047||CCS_10|RETICULOSARCOMA INVOLVING LYMPH NODES OF HEAD, FACE AND NECK
C0684941|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF ACCESSORY SINUS 
C0684941|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF ACCESSORY SINUS
C0684941|T047||CCS_10|ACCESSORY SINUS NEOPLASM MALIGNANT SECONDARY
C0684941|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO ACCESSORY SINUS
C0684941|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF ACCESSORY SINUS 
C0684941|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO ACCESSORY SINUS, NOS
C0684941|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF ACCESSORY SINUS, NOS
C0686623|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF LYMPH NODES OF FACE
C0686623|T047||CCS_10|LYMPH NODE NEOPLASM MALIGNANT SECONDARY FACE
C0686623|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF LYMPH NODES OF FACE 
C0686623|T047||CCS_10|CANCER METASTATIC TO LYMPH NODES OF FACE
C0686623|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO LYMPH NODES OF FACE
C0686623|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF LYMPH NODES OF FACE 
C0686623|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO LYMPH NODES OF FACE, NOS
C0686623|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF LYMPH NODES OF FACE, NOS
C0685136|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BLOOD VESSEL OF NECK
C0685136|T047||CCS_10|NEOPLASM - SOFT TISSUE TYPES BLOOD VESSEL MALIGNANT OF NECK SECONDARY
C0685136|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BLOOD VESSEL OF NECK 
C0685136|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO BLOOD VESSEL OF NECK
C0685136|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BLOOD VESSEL OF NECK 
C0345614|T047||CCS_10|MALIGNANT NEOPLASM OF MINOR SALIVARY GLAND
C0345614|T047||CCS_10|MALIGNANT NEOPLASM OF MINOR SALIVARY GLAND 
C0345614|T047||CCS_10|MALIGNANT TUMOR OF MINOR SALIVARY GLAND
C0345614|T047||CCS_10|MALIGNANT SALIVARY GLAND NEOPLASM MINOR 
C0345614|T047||CCS_10|MALIGNANT SALIVARY GLAND NEOPLASM MINOR
C0345614|T047||CCS_10|MALIGNANT TUMOUR OF MINOR SALIVARY GLAND
C0345614|T047||CCS_10|MALIGNANT TUMOR OF MINOR SALIVARY GLAND 
C0345614|T047||CCS_10|MALIGNANT MINOR SALIVARY GLAND NEOPLASM
C0345614|T047||CCS_10|MALIGNANT MINOR SALIVARY GLAND TUMOR
C0345614|T047||CCS_10|MALIGNANT NEOPLASM OF THE MINOR SALIVARY GLAND
C0345614|T047||CCS_10|MALIGNANT TUMOR OF THE MINOR SALIVARY GLAND
C0686608|T047||CCS_10|OROPHARYNGEAL NEOPLASM TONSIL MALIGNANT SECONDARY
C0686608|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF OF TONSIL
C0686608|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF OF TONSIL 
C0686608|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO PALATINE TONSIL
C0686608|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO TONSIL
C0686608|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF PALATINE TONSIL
C0686608|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF TONSIL
C0686608|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF TONSIL 
C0346575|T047||CCS_10|MALIGNANT TUMOUR POSTERIOR MARGIN NASAL SEPTUM AND CHOANAE
C0346575|T047||CCS_10|MALIGNANT TUMOR POSTERIOR MARGIN NASAL SEPTUM AND CHOANAE 
C0346575|T047||CCS_10|MALIGNANT NEOPLASM OF POSTERIOR MARGIN OF NASAL SEPTUM AND CHOANAE
C0346575|T047||CCS_10|MALIGNANT TUMOR POSTERIOR MARGIN NASAL SEPTUM AND CHOANAE
C0346575|T047||CCS_10|NASAL CAVITY NEOPLASM MALIGNANT OF POSTERIOR MARGIN OF SEPTUM AND CHOANAE
C0346575|T047||CCS_10|MALIGNANT NEOPLASM OF POSTERIOR MARGIN OF NASAL SEPTUM AND CHOANAE 
C0346575|T047||CCS_10|MALIGNANT TUMOR OF POSTERIOR MARGIN OF NASAL SEPTUM AND CHOANAE
C0346575|T047||CCS_10|MALIGNANT TUMOUR OF POSTERIOR MARGIN OF NASAL SEPTUM AND CHOANAE
C0346575|T047||CCS_10|MALIGNANT TUMOR OF POSTERIOR MARGIN OF NASAL SEPTUM AND CHOANAE 
C0346726|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF EAR AND EXTERNAL AURICULAR CANAL
C0346726|T047||CCS_10|SKIN OF EAR AND EXTERNAL AURICULAR CANAL
C0346726|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF EAR AND EXTERNAL AUDITORY CANAL
C0346726|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF EAR AND EXTERNAL AUDITORY CANAL 
C0346726|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF EAR AND EXTERNAL AURICULAR CANAL 
C0346726|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF EAR AND EXTERNAL AURICULAR CANAL NOS 
C0346726|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF EAR AND EXTERNAL AURICULAR CANAL NOS
C0346726|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF EXTERNAL EAR AND AUDITORY CANAL 
C0346726|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF EXTERNAL EAR AND AUDITORY CANAL
C0346726|T047||CCS_10|SKIN NEOPLASM EXTERNAL EAR MALIGNANT AND AUDITORY CANAL
C0685135|T047||CCS_10|MALIGNANT NEOPLASM OF BLOOD VESSEL OF NECK
C0685135|T047||CCS_10|NEOPLASM - SOFT TISSUE TYPES BLOOD VESSEL MALIGNANT OF NECK PRIMARY
C0685135|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF BLOOD VESSEL OF NECK
C0685135|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF BLOOD VESSEL OF NECK 
C0685135|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF BLOOD VESSEL OF NECK 
C0346323|T047||CCS_10|OPTIC NERVE
C0346323|T047||CCS_10|MALIGNANT NEOPLASM OF OPTIC NERVE
C0346323|T047||CCS_10|MALIGNANT TUMOR OF OPTIC NERVE
C0346323|T047||CCS_10|MALIGNANT OPTIC NERVE NEOPL
C0346323|T047||CCS_10|MALIGNANT TUMOUR OF OPTIC NERVE
C0346323|T047||CCS_10|MALIGNANT TUMOUR OF OPTIC NERVE 
C0346323|T047||CCS_10|MALIGNANT OPTIC NERVE TUMOR
C0346323|T047||CCS_10|TUMOR, OPTIC NERVE, MALIGNANT
C0346323|T047||CCS_10|OPTIC NERVE TUMOR, MALIGNANT
C0346323|T047||CCS_10|TUMOR, MALIGNANT, OPTIC NERVE
C0346323|T047||CCS_10|MALIGNANT OPTIC NERVE NEOPLASM
C0346323|T047||CCS_10|MALIGNANT TUMOR OF OPTIC NERVE 
C0153654|T047||CCS_10|MALIGNANT NEOPLASM OF PITUITARY GLAND AND CRANIOPHARYNGEAL DUCT
C0153654|T047||CCS_10|MALIG NEO PITUITARY
C0153654|T047||CCS_10|MALIGNANT NEOPLASM OF PITUITARY GLAND OR CRANIOPHARYNGEAL DUCT NOS 
C0153654|T047||CCS_10|MALIGNANT NEOPLASM OF PITUITARY GLAND OR CRANIOPHARYNGEAL DUCT NOS
C0153654|T047||CCS_10|MALIGNANT NEOPLASM OF PITUITARY GLAND AND CRANIOPHARYNGEAL DUCT 
C0153654|T047||CCS_10|MALIGNANT NEOPLASM OF PITUITARY GLAND AND CRANIOPHARYNGEAL DUCT 
C0685130|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BLOOD VESSEL OF HEAD
C0685130|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BLOOD VESSEL OF HEAD 
C0685130|T047||CCS_10|NEOPLASM - SOFT TISSUE TYPES BLOOD VESSEL MALIGNANT OF HEAD SECONDARY
C0685130|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO BLOOD VESSEL OF HEAD
C0685130|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BLOOD VESSEL OF HEAD 
C0496788|T047||CCS_10|MIDDLE EAR
C0496788|T047||CCS_10|MALIGNANT NEOPLASM OF MIDDLE EAR
C0496788|T047||CCS_10|AUDITORY NEOPLASM MALIGNANT OF MIDDLE EAR
C0496788|T047||CCS_10|MALIGNANT NEOPLASM OF MIDDLE EAR 
C0496788|T047||CCS_10|MALIGNANT MIDDLE EAR NEOPLASM NOS
C0496788|T047||CCS_10|MALIGNANT MIDDLE EAR NEOPLASM
C0496788|T047||CCS_10|MALIGNANT TUMOR OF MIDDLE EAR
C0496788|T047||CCS_10|MALIGNANT TUMOUR OF MIDDLE EAR
C0496788|T047||CCS_10|MALIGNANT TUMOR OF MIDDLE EAR 
C0496788|T047||CCS_10|MALIGNANT MIDDLE EAR TUMOR
C0496788|T047||CCS_10|MALIGNANT NEOPLASM OF THE MIDDLE EAR
C0496788|T047||CCS_10|MALIGNANT TUMOR OF THE MIDDLE EAR
C0684689|T047||CCS_10|SOFT TISSUE NEOPLASM HEAD MALIGNANT SECONDARY
C0684689|T047||CCS_10|SECONDARY MALIGNANT SOFT TISSUE NEOPLASM OF HEAD
C0684689|T047||CCS_10|SECONDARY MALIGNANT SOFT TISSUE NEOPLASM OF HEAD 
C0684689|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO SOFT TISSUES OF HEAD
C0684689|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SOFT TISSUES OF HEAD
C0684689|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SOFT TISSUES OF HEAD 
C0153752|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC-HISTIOCYTIC PREDOMINANCE OF LYMPH NODES OF HEAD, FACE, AND NECK
C0153752|T047||CCS_10|HODG LYMPH-HISTIO HEAD
C0153752|T047||CCS_10|HODGKIN DISEASE, LYMPHOCYTIC-HISTIOCYTIC PREDOMINANCE OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0153752|T047||CCS_10|HODGKIN DISEASE, LYMPHOCYTIC-HISTIOCYTIC PREDOMINANCE OF LYMPH NODES OF HEAD, FACE AND NECK
C0153752|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC-HISTIOCYTIC PREDOMINANCE INVOLVING LYMPH NODES OF HEAD, FACE, AND NECK
C0153752|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC-HISTIOCYTIC PREDOMINANCE, LYMPH NODES OF HEAD, FACE, AND NECK
C0153752|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC-HISTIOCYTIC PREDOMINANCE OF LYMPH NODES OF HEAD, FACE, OR NECK
C0153752|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC-HISTIOCYTIC PREDOMINANCE OF LYMPH NODES OF HEAD, FACE, AND NECK 
C0153752|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC-HISTIOCYTIC PREDOMINANCE OF LYMPH NODES OF HEAD, FACE AND NECK
C0153752|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC-HISTIOCYTIC PREDOMINANCE OF LYMPH NODES OF HEAD, FACE AND/OR NECK 
C0153752|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC-HISTIOCYTIC PREDOMINANCE OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0153752|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC-HISTIOCYTIC PREDOMINANCE OF LYMPH NODES OF HEAD, FACE AND NECK 
C0153752|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC-HISTIOCYTIC PREDOMINANCE INVOLVING LYMPH NODES OF HEAD, FACE AND NECK
C0153688|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BRAIN AND SPINAL CORD
C0153688|T047||CCS_10|SEC MAL NEO BRAIN/SPINE
C0153688|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM BRAIN AND SPINAL CORD
C0153688|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM BRAIN AND SPINAL CORD 
C0153688|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BRAIN OR SPINAL CORD NOS 
C0153688|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BRAIN OR SPINAL CORD NOS
C0153688|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BRAIN AND SPINAL CORD 
C0685132|T047||CCS_10|MALIGNANT NEOPLASM OF BLOOD VESSEL OF FACE
C0685132|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF BLOOD VESSEL OF FACE
C0685132|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF BLOOD VESSEL OF FACE 
C0685132|T047||CCS_10|NEOPLASM - SOFT TISSUE TYPES BLOOD VESSEL MALIGNANT OF FACE PRIMARY
C0685132|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF BLOOD VESSEL OF FACE 
C0684756|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF MUSCLE OF NECK 
C0684756|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF MUSCLE OF NECK
C0684756|T047||CCS_10|MALIGNANT NEOPLASM OF MUSCLE OF NECK SECONDARY
C0684756|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO MUSCLE OF NECK
C0684756|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF MUSCLE OF NECK 
C0684692|T047||CCS_10|SECONDARY MALIGNANT SOFT TISSUE NEOPLASM OF FACE
C0684692|T047||CCS_10|SOFT TISSUE NEOPLASM FACE MALIGNANT SECONDARY
C0684692|T047||CCS_10|SECONDARY MALIGNANT SOFT TISSUE NEOPLASM OF FACE 
C0684692|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO SOFT TISSUES OF FACE
C0684692|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SOFT TISSUES OF FACE
C0684692|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SOFT TISSUES OF FACE 
C0346124|T047||CCS_10|MALIGNANT NEOPLASM OF SOFT TISSUES OF HEAD
C0346124|T047||CCS_10|MALIGNANT SOFT TISSUE NEOPLASM OF HEAD
C0346124|T047||CCS_10|MALIGNANT SOFT TISSUE NEOPLASM OF HEAD 
C0346124|T047||CCS_10|SOFT TISSUE NEOPLASM HEAD MALIGNANT
C0346124|T047||CCS_10|MALIGNANT TUMOR OF SOFT TISSUE OF HEAD
C0346124|T047||CCS_10|MALIGNANT TUMOUR OF SOFT TISSUE OF HEAD
C0346124|T047||CCS_10|MALIGNANT NEOPLASM OF SOFT TISSUE OF HEAD
C0346124|T047||CCS_10|MALIGNANT TUMOR OF SOFT TISSUE OF HEAD 
C0349038|T047||CCS_10|MALIGNANT NEOPLASM OVERLAPPING NASOPHARYNX SITE
C0349038|T047||CCS_10|OVERLAPPING LESION OF NASOPHARYNX
C0349038|T047||CCS_10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF NASOPHARYNX
C0349038|T047||CCS_10|MALIGNANT NEOPLASM, OVERLAPPING LESION OF NASOPHARYNX 
C0349038|T047||CCS_10|MALIGNANT NEOPLASM, OVERLAPPING LESION OF NASOPHARYNX
C0349038|T047||CCS_10|OVERLAPPING MALIGNANT NEOPLASM OF NASOPHARYNGEAL WALL
C0349038|T047||CCS_10|OVERLAPPING MALIGNANT NEOPLASM OF NASOPHARYNX 
C0349038|T047||CCS_10|OVERLAPPING MALIGNANT NEOPLASM OF NASOPHARYNX
C1263917|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF NECK
C1263917|T047||CCS_10|NEOPLASM - PNS MALIGNANT NECK PRIMARY
C1263917|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF NECK 
C1263917|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF NECK 
C0345628|T047||CCS_10|MALIGNANT NEOPLASM OF MASTOID AIR CELLS
C0345628|T047||CCS_10|BONE NEOPLASM, MALIGNANT - SKULL AND FACE, MASTOID AIR CELLS
C0345628|T047||CCS_10|MALIGNANT NEOPLASM OF MASTOID AIR CELLS 
C0345628|T047||CCS_10|MALIGNANT TUMOR OF MASTOID AIR CELLS
C0345628|T047||CCS_10|MALIGNANT TUMOUR OF MASTOID AIR CELLS
C0345628|T047||CCS_10|MALIGNANT TUMOR OF MASTOID AIR CELLS 
C0153704|T047||CCS_10|LYMPHOSARCOMA OF LYMPH NODES OF HEAD, FACE AND/OR NECK -RETIRED-
C0153704|T047||CCS_10|LYMPHOSARCOMA HEAD
C0153704|T047||CCS_10|LYMPHOSARCOMA INVOLVING LYMPH NODES OF HEAD, FACE, AND NECK
C0153704|T047||CCS_10|LYMPHOSARCOMA, LYMPH NODES OF HEAD, FACE, AND NECK
C0153704|T047||CCS_10|LYMPHOSARCOMA OF LYMPH NODES OF HEAD, FACE, AND NECK
C0153704|T047||CCS_10|LYMPHOSARCOMA OF LYMPH NODES OF HEAD, FACE AND/OR NECK 
C0153704|T047||CCS_10|LYMPHOSARCOMA OF HEAD, FACE, AND NECK LYMPH NODES
C0153704|T047||CCS_10|LYMPHOSARCOMA OF LYMPH NODES OF HEAD, FACE, AND NECK 
C0153704|T047||CCS_10|LYMPHOSARCOMA OF LYMPH NODES OF HEAD, FACE AND NECK
C0153704|T047||CCS_10|LYMPHOSARCOMA OF LYMPH NODES OF HEAD, FACE AND NECK 
C0153704|T047||CCS_10|LYMPHOSARCOMA INVOLVING LYMPH NODES OF HEAD, FACE AND NECK
C0345586|T047||CCS_10|ORAL CAVITY NEOPLASM MALIGNANT LABIAL SULCUS, LOWER
C0345586|T047||CCS_10|MALIGNANT NEOPLASM OF LOWER LABIAL SULCUS 
C0345586|T047||CCS_10|MALIGNANT NEOPLASM OF LOWER LABIAL SULCUS
C0345586|T047||CCS_10|MALIGNANT TUMOR OF LOWER LABIAL SULCUS
C0345586|T047||CCS_10|MALIGNANT TUMOUR OF LOWER LABIAL SULCUS
C0345586|T047||CCS_10|MALIGNANT TUMOR OF LOWER LABIAL SULCUS 
C0686641|T047||CCS_10|SECONDARY AND UNSPECIFIED MALIGNANT NEOPLASM OF INFRACLAVICULAR LYMPH NODES
C0686641|T047||CCS_10|SECONDARY AND UNSPECIFIED MALIGNANT NEOPLASM OF INFRACLAVICULAR LYMPH NODES 
C0686641|T047||CCS_10|LYMPH NODE NEOPLASM MALIGNANT SECONDARY NECK INFRACLAVICULAR
C0686641|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF INFRACLAVICULAR LYMPH NODES 
C0686641|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF INFRACLAVICULAR LYMPH NODES
C0686641|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO INFRACLAVICULAR LYMPH NODES
C0686641|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF INFRACLAVICULAR LYMPH NODES 
C0153354|T047||CCS_10|MALIGNANT NEOPLASM OF ANTERIOR TWO-THIRDS OF TONGUE, PART UNSPECIFIED
C0153354|T047||CCS_10|ANTERIOR TWO-THIRDS OF TONGUE, PART UNSPECIFIED
C0153354|T047||CCS_10|MALIGNANT NEOPLASM OF ANTERIOR TWO-THIRDS OF TONGUE
C0153354|T047||CCS_10|MALIGNANT NEOPLASM OF ANTERIOR TWO-THIRDS OF TONGUE 
C0153354|T047||CCS_10|MALIGNANT TUMOR OF ANTERIOR TWO-THIRDS OF TONGUE
C0153354|T047||CCS_10|MAL NEO ANT 2/3 TONGUE
C0153354|T047||CCS_10|MALIGNANT NEOPLASM OF MOBILE PART OF TONGUE NOS
C0153354|T047||CCS_10|MALIG NEOPLASM OF ANTERIOR TWO-THIRDS OF TONGUE, PART UNSP
C0153354|T047||CCS_10|MALIGNANT NEOPLASM OF ANTERIOR 2/3 OF TONGUE UNSPECIFIED
C0153354|T047||CCS_10|MALIGNANT TUMOUR OF MOBILE PART OF TONGUE
C0153354|T047||CCS_10|MALIGNANT TUMOR OF MOBILE PART OF TONGUE
C0153354|T047||CCS_10|MALIGNANT NEOPLASM OF ANTERIOR 2/3 OF TONGUE UNSPECIFIED 
C0153354|T047||CCS_10|MALIGNANT TUMOUR OF ANTERIOR TWO-THIRDS OF TONGUE
C0153354|T047||CCS_10|MALIGNANT TUMOR OF ANTERIOR TWO-THIRDS OF TONGUE 
C0153354|T047||CCS_10|MALIGNANT NEOPLASM OF ANTERIOR TWO-THIRDS OF TONGUE, NOS
C0153736|T047||CCS_10|HODGKIN'S GRANULOMA OF LYMPH NODES OF HEAD, FACE, AND NECK
C0153736|T047||CCS_10|HODGKINS GRANULOM HEAD
C0153736|T047||CCS_10|HODGKIN GRANULOMA OF LYMPH NODES OF HEAD, FACE AND NECK
C0153736|T047||CCS_10|HODGKIN GRANULOMA OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0153736|T047||CCS_10|HODGKIN'S GRANULOMA, LYMPH NODES OF HEAD, FACE, AND NECK
C0153736|T047||CCS_10|HODGKIN'S GRANULOMA INVOLVING LYMPH NODES OF HEAD, FACE, AND NECK
C0153736|T047||CCS_10|HODGKIN DISEASE GRANULOMA - HEAD, FACE, & NECK
C0153736|T047||CCS_10|HODGKIN GRANULOMA OF LYMPH NODES OF HEAD, FACE, & NECK 
C0153736|T047||CCS_10|HODGKIN GRANULOMA OF LYMPH NODES OF HEAD, FACE, & NECK
C0153736|T047||CCS_10|HODGKIN'S GRANULOMA OF LYMPH NODES OF HEAD, FACE AND NECK
C0153736|T047||CCS_10|HODGKIN'S GRANULOMA OF LYMPH NODES OF HEAD, FACE AND/OR NECK 
C0153736|T047||CCS_10|HODGKIN'S GRANULOMA OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0153736|T047||CCS_10|HODGKIN'S GRANULOMA OF LYMPH NODES OF HEAD, FACE AND NECK 
C0153736|T047||CCS_10|HODGKIN'S GRANULOMA INVOLVING LYMPH NODES OF HEAD, FACE AND NECK
C0684554|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF CERVICAL VERTEBRAL COLUMN 
C0684554|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF CERVICAL VERTEBRAL COLUMN
C0684554|T047||CCS_10|BONE NEOPLASM, MALIGNANT - VERTEBRAL COLUMN CERVICAL SECONDARY
C0684554|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO CERVICAL VERTEBRAL COLUMN
C0684554|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF CERVICAL VERTEBRAL COLUMN 
C0347957|T047||CCS_10|CONNECTIVE AND SOFT TISSUE OF HEAD, FACE AND NECK
C0347957|T047||CCS_10|MALIGNANT NEOPLASM OF CONNECTIVE AND SOFT TISSUE OF HEAD, FACE AND NECK
C0347957|T047||CCS_10|MALIG NEOPLM OF CONN AND SOFT TISSUE OF HEAD, FACE AND NECK
C0347957|T047||CCS_10|MALIGNANT NEOPLASM OF CONNECTIVE AND SOFT TISSUE OF HEAD, FACE, AND NECK 
C0347957|T047||CCS_10|MALIGNANT NEOPLASM OF CONNECTIVE AND SOFT TISSUE OF HEAD, FACE, AND NECK
C0347957|T047||CCS_10|MALIGNANT NEOPLASM OF CONNECTIVE AND SOFT TISSUE OF HEAD, FACE AND NECK 
C0153768|T047||CCS_10|HODGKIN'S DISEASE, MIXED CELLULARITY OF LYMPH NODES OF HEAD, FACE, AND NECK
C0153768|T047||CCS_10|HODGKIN'S DISEASE, MIXED CELLULARITY, INVOLVING LYMPH NODES OF HEAD, FACE, AND NECK.
C0153768|T047||CCS_10|HODGKINS MIX CELL HEAD
C0153768|T047||CCS_10|HODGKIN DISEASE, MIXED CELLULARITY OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0153768|T047||CCS_10|HODGKIN DISEASE, MIXED CELLULARITY OF LYMPH NODES OF HEAD, FACE AND NECK
C0153768|T047||CCS_10|HODGKIN'S DISEASE, MIXED CELLULARITY, LYMPH NODES OF HEAD, FACE, AND NECK
C0153768|T047||CCS_10|HODGKIN'S DISEASE, MIXED CELLULARITY, INVOLVING LYMPH NODES OF HEAD, FACE, AND NECK
C0153768|T047||CCS_10|MIXED CELLULARITY HODGKIN'S LYMPHOMA OF LYMPH NODES OF HEAD, FACE, AND NECK
C0153768|T047||CCS_10|HODGKIN'S LYMPHOMA MIXED CELLULARITY OF HEAD, FACE, AND NECK
C0153768|T047||CCS_10|MIXED CELLULARITY HODGKIN'S LYMPHOMA OF LYMPH NODES OF HEAD, FACE, AND NECK 
C0153768|T047||CCS_10|HODGKIN'S DISEASE, MIXED CELLULARITY OF LYMPH NODES OF HEAD, FACE AND NECK
C0153768|T047||CCS_10|HODGKIN'S DISEASE, MIXED CELLULARITY OF LYMPH NODES OF HEAD, FACE AND/OR NECK 
C0153768|T047||CCS_10|HODGKIN'S DISEASE, MIXED CELLULARITY OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0153768|T047||CCS_10|HODGKIN'S DISEASE, MIXED CELLULARITY OF LYMPH NODES OF HEAD, FACE AND NECK 
C0153768|T047||CCS_10|HODGKIN'S DISEASE, MIXED CELLULARITY, INVOLVING LYMPH NODES OF HEAD, FACE AND NECK
C1263911|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF HEAD
C1263911|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF HEAD 
C1263911|T047||CCS_10|NEOPLASM - PNS MALIGNANT HEAD PRIMARY
C1263911|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF HEAD 
C0346322|T047||CCS_10|MALIGNANT OPTIC NERVE SHEATH NEOPL
C0346322|T047||CCS_10|OPTIC NERVE SHEATH NEOPL MALIGNANT
C0346322|T047||CCS_10|MALIGNANT NEOPLASM OF OPTIC NERVE (II) AND SHEATH
C0346322|T047||CCS_10|MALIGNANT NEOPLASM OF OPTIC NERVE (II) AND SHEATH 
C0346322|T047||CCS_10|MALIGNANT NEOPLASM OF OPTIC NERVE SHEATH 
C0346322|T047||CCS_10|NEOPLASM - MALIGNANT OF OPTIC NERVE (II) AND SHEATH
C0346322|T047||CCS_10|MALIGNANT NEOPLASM OF OPTIC NERVE SHEATH
C0346322|T047||CCS_10|MALIGNANT OPTIC NERVE SHEATH TUMORS
C0346322|T047||CCS_10|OPTIC NERVE SHEATH NEOPLASMS, MALIGNANT
C0346322|T047||CCS_10|OPTIC NERVE SHEATH TUMORS, MALIGNANT
C0346322|T047||CCS_10|MALIGNANT OPTIC NERVE SHEATH NEOPLASMS
C0346322|T047||CCS_10|MALIGNANT TUMOR OF OPTIC NERVE AND SHEATH
C0346322|T047||CCS_10|MALIGNANT TUMOR OF OPTIC NERVE SHEATH
C0346322|T047||CCS_10|MALIGNANT TUMOUR OF OPTIC NERVE AND SHEATH
C0346322|T047||CCS_10|MALIGNANT TUMOUR OF OPTIC NERVE SHEATH
C0346322|T047||CCS_10|MALIGNANT TUMOR OF OPTIC NERVE AND SHEATH 
C0346322|T047||CCS_10|MALIGNANT TUMOR OF OPTIC NERVE SHEATH 
C0684520|T047||CCS_10|BONE NEOPLASM, MALIGNANT - SKULL SECONDARY
C0684520|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SKULL
C0684520|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SKULL 
C0684520|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO BONE OF SKULL
C0684520|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BONE OF SKULL 
C0684520|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BONE OF SKULL
C0684520|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO BONE OF SKULL, NOS
C0684520|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF BONE OF SKULL, NOS
C0206115|T047||CCS_10|WAGR SYNDROME
C0206115|T047||CCS_10|SYNDROME, WAGR
C0206115|T047||CCS_10|WAGR SYNDROMES
C0206115|T047||CCS_10|WAGR
C0206115|T047||CCS_10|WILMS TUMOR, ANIRIDIA, GENITOURINARY ANOMALIES, AND MENTAL RETARDATION SYNDROME
C0206115|T047||CCS_10|COMPLEX, WAGR
C0206115|T047||CCS_10|CONTIGUOUS GENE SYNDROME, WAGR
C0206115|T047||CCS_10|WAGR COMPLEX
C0206115|T047||CCS_10|WILMS TUMOR-ANIRIDIA-GENITOURINARY ANOMALIES-MR SYNDROME
C0206115|T047||CCS_10|WAGR CONTIGUOUS GENE SYNDROME
C0206115|T047||CCS_10|WAGR SYNDROME [DISEASE/FINDING]
C0206115|T047||CCS_10|WILMS TUMOR, ANIRIDIA, GENITOURINARY ANOMALIES, MENTAL RETARDATION SYNDROME
C0206115|T047||CCS_10|WILMS TUMOR-ANIRIDIA-GONADOBLASTOMA-MENTAL RETARDATION SYNDROME
C0206115|T047||CCS_10|WAGR COMPLICES
C0206115|T047||CCS_10|CHROMOSOME 11P13 DELETION SYNDROME
C0206115|T047||CCS_10|11P PARTIAL MONOSOMY SYNDROME
C0206115|T047||CCS_10|ANOMALY OF CHROMOSOME PAIR 11P PARTIAL MONOSOMY SYNDROME
C0206115|T047||CCS_10|11P PARTIAL MONOSOMY SYNDROME 
C0206115|T047||CCS_10|WILMS TUMOR-ANIRIDIA-GENITAL ANOMALIES-RETARDATION SYNDROME
C0206115|T047||CCS_10|WILMS TUMOR-ANIRIDIA-GENITOURINARY ANOMALIES-MENTAL RETARDATION SYNDROME
C0206115|T047||CCS_10|ANIRIDIA-WILMS TUMOR ASSOCIATION
C0206115|T047||CCS_10|ANIRIDIA-WILMS TUMOUR ASSOCIATION
C0206115|T047||CCS_10|11P PARTIAL MONOSOMY SYNDROME 
C0496763|T047||CCS_10|MALIGNANT NEOPLASM OF MAJOR SALIVARY GLANDS
C0496763|T047||CCS_10|MALIGNANT NEOPLASM OF MAJOR SALIVARY GLAND
C0496763|T047||CCS_10|MALIGNANT NEOPLASM OF MAJOR SALIVARY GLAND, UNSPECIFIED
C0496763|T047||CCS_10|MALIGNANT NEOPLASM OF SALIVARY GLAND (MAJOR) NOS
C0496763|T047||CCS_10|MALIGNANT NEOPLASM OF MAJOR SALIVARY GLAND NOS
C0496763|T047||CCS_10|MALIGNANT NEOPLASM OF MAJOR SALIVARY GLAND NOS 
C0496763|T047||CCS_10|MALIGNANT SALIVARY GLAND NEOPLASM MAJOR
C0496763|T047||CCS_10|MALIGNANT NEOPLASM OF MAJOR SALIVARY GLAND 
C0496763|T047||CCS_10|MALIGNANT TUMOR OF MAJOR SALIVARY GLAND
C0496763|T047||CCS_10|MALIGNANT TUMOUR OF MAJOR SALIVARY GLAND
C0496763|T047||CCS_10|MALIGNANT TUMOR OF MAJOR SALIVARY GLAND 
C0496763|T047||CCS_10|MALIGNANT NEOPLASM OF MAJOR SALIVARY GLAND, NOS
C0496763|T047||CCS_10|MALIGNANT MAJOR SALIVARY GLAND NEOPLASM
C0496763|T047||CCS_10|MALIGNANT MAJOR SALIVARY GLAND TUMOR
C0496763|T047||CCS_10|MALIGNANT NEOPLASM OF THE MAJOR SALIVARY GLAND
C0496763|T047||CCS_10|MALIGNANT TUMOR OF THE MAJOR SALIVARY GLAND
C0684967|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF POSTCRICOID REGION 
C0684967|T047||CCS_10|HYPOPHARYNGEAL NEOPLASM MALIGNANT POSTCRICOID REGION SECONDARY
C0684967|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF POSTCRICOID REGION
C0684967|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO POSTCRICOID REGION
C0684967|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF POSTCRICOID REGION 
C1305982|T047||CCS_10|CRANIAL NERVE NEOPLASM MALIGNANT PRIMARY
C1305982|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF CRANIAL NERVE 
C1305982|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF CRANIAL NERVE
C1305982|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF CRANIAL NERVE 
C1304838|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF UPPER RESPIRATORY TRACT
C1304838|T047||CCS_10|MALIGNANT NEOPLASM UPPER RESPIRATORY TRACT PRIMARY
C1304838|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF UPPER RESPIRATORY TRACT 
C1304838|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF UPPER RESPIRATORY TRACT 
C0346776|T047||CCS_10|MALIGNANT MELANOMA OF THE CHIN 
C0346776|T047||CCS_10|MALIGNANT MELANOMA OF THE CHIN
C0346776|T047||CCS_10|MALIGNANT MELANOMA OF CHIN
C0346776|T047||CCS_10|MALIGNANT MELANOMA OF SKIN OF CHIN
C0346776|T047||CCS_10|MALIGNANT MELANOMA OF CHIN 
C0346776|T047||CCS_10|MALIGNANT MELANOMA OF SKIN OF CHIN 
C0347013|T047||CCS_10|METASTASIS TO NERVOUS SYSTEM AND EYE 
C0347013|T047||CCS_10|MALIGNANT NEOPLASM METASTATIC CANCER TO NERVOUS SYSTEM AND EYE
C0347013|T047||CCS_10|METASTASIS TO NERVOUS SYSTEM AND EYE
C0347013|T047||CCS_10|METASTASIS TO NERVOUS SYSTEM AND EYE 
C0153810|T047||CCS_10|SÉZARY'S DISEASE OF LYMPH NODES OF HEAD, FACE AND NECK
C0153810|T047||CCS_10|SÉZARY'S DISEASE OF LYMPH NODES OF HEAD, FACE AND NECK 
C0153810|T047||CCS_10|SÉZARY'S DISEASE OF LYMPH NODES OF HEAD, FACE, AND NECK
C0153810|T047||CCS_10|SEZARY SYNDROME OF HEAD, FACE, AND NECK 
C0153810|T047||CCS_10|SEZARY SYNDROME OF HEAD, FACE, AND NECK
C0153810|T047||CCS_10|SEZARY'S DISEASE OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0153810|T047||CCS_10|SEZARY'S DISEASE HEAD
C0153810|T047||CCS_10|SÉZARY DISEASE OF LYMPH NODES OF HEAD, FACE AND NECK
C0153810|T047||CCS_10|SÉZARY DISEASE OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0153810|T047||CCS_10|SÉZARY DISEASE, LYMPH NODES OF HEAD, FACE, AND NECK
C0153810|T047||CCS_10|SEZARY'S DISEASE, LYMPH NODES OF HEAD, FACE, AND NECK
C0153810|T047||CCS_10|SEZARY'S DISEASE INVOLVING LYMPH NODES OF HEAD, FACE, AND NECK
C0153810|T047||CCS_10|SÉZARY'S DISEASE OF LYMPH NODES OF HEAD, FACE AND/OR NECK 
C0153810|T047||CCS_10|SEZARY'S DISEASE INVOLVING LYMPH NODES OF HEAD, FACE AND NECK
C0685010|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF LARYNGEAL ASPECT OF ARYEPIGLOTTIC FOLD
C0685010|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF LARYNGEAL ASPECT OF ARYEPIGLOTTIC FOLD 
C0685010|T047||CCS_10|MALIGNANT NEOPLASM SUPRAGLOTTIS LARYNGEAL ASPECT OF ARYEPIGLOTTIC FOLD SECONDARY
C0685010|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO LARYNGEAL ASPECT OF ARYEPIGLOTTIC FOLD
C0685010|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF LARYNGEAL ASPECT OF ARYEPIGLOTTIC FOLD 
C3647449|T047||CCS_10|MALIGNANT NEOPLASM OF ANTERIOR WALL OF NASOPHARYNX
C3647449|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF ANTERIOR WALL OF NASOPHARYNX 
C3647449|T047||CCS_10|PRIMARY MALIGNANT NASOPHARYNGEAL NEOPLASM OF ANTERIOR WALL
C3647449|T047||CCS_10|PRIMARY MALIGNANT NASOPHARYNGEAL NEOPLASM OF ANTERIOR WALL 
C3647449|T047||CCS_10|NASOPHARYNGEAL NEOPLASM ANTERIOR WALL, MALIGNANT PRIMARY
C3647449|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF ANTERIOR WALL OF NASOPHARYNX
C0686627|T047||CCS_10|SECONDARY AND UNSPECIFIED MALIGNANT NEOPLASM OF OCCIPITAL LYMPH NODES 
C0686627|T047||CCS_10|SECONDARY AND UNSPECIFIED MALIGNANT NEOPLASM OF OCCIPITAL LYMPH NODES
C0686627|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF OCCIPITAL LYMPH NODES
C0686627|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF OCCIPITAL LYMPH NODES 
C0686627|T047||CCS_10|LYMPH NODE NEOPLASM MALIGNANT SECONDARY HEAD OCCIPITAL
C0686627|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO OCCIPITAL LYMPH NODES
C0686627|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF OCCIPITAL LYMPH NODES 
C0018197|T047||CCS_10|GRANULOMA, LETHAL MIDLINE
C0018197|T047||CCS_10|GRANULOMAS, LETHAL MIDLINE
C0018197|T047||CCS_10|LETHAL MIDLINE GRANULOMAS
C0018197|T047||CCS_10|MIDLINE GRANULOMA, LETHAL
C0018197|T047||CCS_10|MIDLINE GRANULOMAS, LETHAL
C0018197|T047||CCS_10|LETHAL MIDLINE GRANULOMA
C0018197|T047||CCS_10|LETHAL MIDLINE GRANULOMA 
C0018197|T047||CCS_10|MIDLINE LETHAL GRANULOMA OF NASAL CAVITY AND PARANASAL SINUS
C0018197|T047||CCS_10|MIDLINE LETHAL GRANULOMA OF THE NASAL CAVITY AND PARANASAL SINUS
C0018197|T047||CCS_10|NASAL CAVITY AND PARANASAL SINUS LETHAL MIDLINE GRANULOMA
C0018197|T047||CCS_10|GRANULOMA, LETHAL MIDLINE [DISEASE/FINDING]
C0018197|T047||CCS_10|IDIOPATHIC MIDLINE GRANULOMA
C0018197|T047||CCS_10|LETHAL MIDLINE GRANULOMA OF FACE
C0018197|T047||CCS_10|MALIGNANT GRANULOMA OF FACE
C0018197|T047||CCS_10|LETHAL MIDLINE GRANULOMA 
C0018197|T047||CCS_10|PARANASAL SINUS AND NASAL CAVITY MIDLINE LETHAL GRANULOMA
C0018197|T047||CCS_10|LETHAL MIDLINE RETICULOSIS
C0018197|T047||CCS_10|MIDLINE LETHAL GRANULOMA, PARANASAL SINUS AND NASAL CAVITY
C0018197|T047||CCS_10|NASAL CAVITY AND PARANASAL SINUS MIDLINE LETHAL GRANULOMA
C0018197|T047||CCS_10|GRANULOMA; MIDLINE
C0018197|T047||CCS_10|MIDLINE; GRANULOMA
C0018197|T047||CCS_10|MIDFACIAL NECROTISING LESION
C0153381|T047||CCS_10|MALIGNANT NEOPLASM OF MOUTH
C0153381|T047||CCS_10|MALIGNANT NEOPLASM OF MOUTH, UNSPECIFIED
C0153381|T047||CCS_10|MALIGNANT NEOPLASM OF ORAL CAVITY 
C0153381|T047||CCS_10|MALIGNANT NEOPLASM OF ORAL CAVITY
C0153381|T047||CCS_10|MALIGNANT ORAL CAVITY NEOPLASMS
C0153381|T047||CCS_10|CANCERS, MOUTH
C0153381|T047||CCS_10|MOUTH CANCERS
C0153381|T047||CCS_10|CANCER, ORAL
C0153381|T047||CCS_10|CANCERS, ORAL
C0153381|T047||CCS_10|ORAL CANCERS
C0153381|T047||CCS_10|MALIGNANT TUMOR OF ORAL CAVITY
C0153381|T047||CCS_10|MALIG NEOPLASM MOUTH NOS
C0153381|T047||CCS_10|MALIGNANT NEOPLASM OF ORAL CAVITY NOS
C0153381|T047||CCS_10|CANCER, MOUTH
C0153381|T047||CCS_10|MOUTH CANCER
C0153381|T047||CCS_10|MALIGNANT TUMOUR OF MOUTH
C0153381|T047||CCS_10|CANCER OF ORAL CAVITY
C0153381|T047||CCS_10|CA - MOUTH CANCER
C0153381|T047||CCS_10|MALIGNANT NEOPLASM OF MOUTH NOS 
C0153381|T047||CCS_10|MALIGNANT TUMOR OF MOUTH
C0153381|T047||CCS_10|MALIGNANT NEOPLASM OF MOUTH NOS
C0153381|T047||CCS_10|MALIGNANT TUMOUR OF ORAL CAVITY
C0153381|T047||CCS_10|MOUTH--CANCER
C0153381|T047||CCS_10|ORAL NEOPLASM MALIGNANT
C0153381|T047||CCS_10|ORAL CANCER
C0153381|T047||CCS_10|CANCER OF THE MOUTH
C0153381|T047||CCS_10|MALIGNANT TUMOR OF ORAL CAVITY 
C0153381|T047||CCS_10|MALIGNANT NEOPLASM OF MOUTH, NOS
C0153381|T047||CCS_10|MALIGNANT MOUTH NEOPLASM
C0153381|T047||CCS_10|MALIGNANT MOUTH TUMOR
C0153381|T047||CCS_10|MALIGNANT NEOPLASM OF THE MOUTH
C0153381|T047||CCS_10|MALIGNANT ORAL CAVITY NEOPLASM
C0153381|T047||CCS_10|MALIGNANT ORAL CAVITY TUMOR
C0153381|T047||CCS_10|MALIGNANT ORAL NEOPLASM
C0153381|T047||CCS_10|MALIGNANT TUMOR OF THE MOUTH
C0153381|T047||CCS_10|CANCER OF MOUTH
C0684992|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF VOCAL CORD
C0684992|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF VOCAL CORD 
C0684992|T047||CCS_10|LARYNGEAL NEOPLASM VOCAL CORD MALIGNANT SECONDARY
C0684992|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO VOCAL CORD
C0684992|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF VOCAL CORD 
C0684748|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF MUSCLE OF HEAD
C0684748|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF MUSCLE OF HEAD 
C0684748|T047||CCS_10|MALIGNANT NEOPLASM OF MUSCLE OF HEAD SECONDARY
C0684748|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO MUSCLE OF HEAD
C0684748|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF MUSCLE OF HEAD 
C0240803|T047||CCS_10|PRIMARY CEREBRAL LYMPHOMA
C0240803|T047||CCS_10|PRIMARY LYMPHOMA OF CEREBRUM
C0240803|T047||CCS_10|PRIMARY LYMPHOMA OF THE CEREBRUM
C0240803|T047||CCS_10|PRIMARY LYMPHOMA, BRAIN
C0240803|T047||CCS_10|MALIGNANT LYMPHOMA OF BRAIN 
C0240803|T047||CCS_10|MALIGNANT LYMPHOMA OF BRAIN
C0240803|T047||CCS_10|NEOPLASM - BRAIN CEREBRUM, MALIGNANT PRIMARY LYMPHOMA
C0240803|T047||CCS_10|PRIMARY CEREBRAL LYMPHOMA 
C0240803|T047||CCS_10|PRIMARY MALIGNANT LYMPHOMA OF BRAIN 
C0240803|T047||CCS_10|PRIMARY MALIGNANT LYMPHOMA OF BRAIN
C0240803|T047||CCS_10|MALIGNANT NEOPLASM LYMPHOMA OF BRAIN PRIMARY
C0240803|T047||CCS_10|BRAIN LYMPHOMA
C0240803|T047||CCS_10|CEREBRAL LYMPHOMA
C0240803|T047||CCS_10|PRIMARY CEREBRAL LYMPHOMA 
C0686612|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF ADENOID 
C0686612|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF ADENOID
C0686612|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO ADENOID
C0686612|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF ADENOID 
C0686507|T047||CCS_10|METASTATIC NEOPLASM TO THE PARATHYROID
C0686507|T047||CCS_10|METASTATIC PARATHYROID NEOPLASM
C0686507|T047||CCS_10|METASTATIC MALIGNANT PARATHYROID GLAND NEOPLASM
C0686507|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF PARATHYROID GLAND 
C0686507|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF PARATHYROID GLAND
C0686507|T047||CCS_10|PARATHYROID NEOPLASM MALIGNANT SECONDARY
C0686507|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM IN THE PARATHYROID GLANDS
C0686507|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO THE PARATHYROID GLANDS
C0686507|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO PARATHYROID GLAND
C0686507|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF PARATHYROID GLAND 
C0686507|T047||CCS_10|METASTASIS TO THE PARATHYROID GLAND
C0686507|T047||CCS_10|METASTATIC NEOPLASM OF PARATHYROID GLAND
C0686507|T047||CCS_10|METASTATIC NEOPLASM OF PARATHYROID
C0686507|T047||CCS_10|METASTATIC NEOPLASM OF THE PARATHYROID GLAND
C0686507|T047||CCS_10|METASTATIC NEOPLASM OF THE PARATHYROID
C0686507|T047||CCS_10|METASTATIC NEOPLASM TO THE PARATHYROID GLAND
C0686507|T047||CCS_10|METASTATIC PARATHYROID GLAND NEOPLASM
C0686507|T047||CCS_10|METASTATIC PARATHYROID GLAND TUMOR
C0686507|T047||CCS_10|METASTATIC PARATHYROID TUMOR
C0686507|T047||CCS_10|METASTATIC TUMOR OF PARATHYROID GLAND
C0686507|T047||CCS_10|METASTATIC TUMOR OF PARATHYROID
C0686507|T047||CCS_10|METASTATIC TUMOR OF THE PARATHYROID GLAND
C0686507|T047||CCS_10|METASTATIC TUMOR OF THE PARATHYROID
C0686507|T047||CCS_10|METASTATIC TUMOR TO THE PARATHYROID GLAND
C0686507|T047||CCS_10|METASTATIC TUMOR TO THE PARATHYROID
C0153776|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION OF LYMPH NODES OF HEAD, FACE, AND NECK
C0153776|T047||CCS_10|LYMPHOCYTE DEPLETION HODGKIN'S DISEASE OF LYMPH NODES OF HEAD, FACE, OR NECK
C0153776|T047||CCS_10|LYMPHOCYTE DEPLETION HODGKIN'S DISEASE OF LYMPH NODES OF HEAD, FACE, OR NECK 
C0153776|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION, INVOLVING LYMPH NODES OF HEAD, FACE, AND NECK.
C0153776|T047||CCS_10|HODG LYMPH DEPLET HEAD
C0153776|T047||CCS_10|HODGKIN DISEASE, LYMPHOCYTIC DEPLETION OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0153776|T047||CCS_10|HODGKIN DISEASE, LYMPHOCYTIC DEPLETION OF LYMPH NODES OF HEAD, FACE AND NECK
C0153776|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION, LYMPH NODES OF HEAD, FACE, AND NECK
C0153776|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION, INVOLVING LYMPH NODES OF HEAD, FACE, AND NECK
C0153776|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION OF LYMPH NODES OF HEAD, FACE AND NECK
C0153776|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION OF LYMPH NODES OF HEAD, FACE AND/OR NECK 
C0153776|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0153776|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION OF LYMPH NODES OF HEAD, FACE AND NECK 
C0153776|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION, INVOLVING LYMPH NODES OF HEAD, FACE AND NECK
C0685991|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO SUBMAXILLARY GLAND
C0685991|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SUBMAXILLARY GLAND
C0685991|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF SUBMAXILLARY GLAND 
C1304847|T047||CCS_10|JAW NEOPLASM MALIGNANT PRIMARY
C1304847|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF JAW 
C1304847|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF JAW
C1304847|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF JAW 
C0153350|T047||CCS_10|MALIGNANT NEOPLASM OF BASE OF TONGUE
C0153350|T047||CCS_10|MALIGNANT NEOPLASM OF BASE OF TONGUE 
C0153350|T047||CCS_10|MALIGNANT TUMOR OF BASE OF TONGUE
C0153350|T047||CCS_10|MAL NEO TONGUE BASE
C0153350|T047||CCS_10|MALIGNANT NEOPLASM OF POSTERIOR THIRD OF TONGUE
C0153350|T047||CCS_10|MALIGNANT NEOPLASM OF FIXED PART OF TONGUE NOS
C0153350|T047||CCS_10|MALIGNANT NEOPLASM OF FIXED PART OF TONGUE NOS 
C0153350|T047||CCS_10|MALIGNANT TUMOR OF FIXED PART OF TONGUE
C0153350|T047||CCS_10|MALIGNANT TUMOR OF POSTERIOR THIRD OF TONGUE
C0153350|T047||CCS_10|MALIGNANT TUMOR OF TONGUE POSTERIOR TO VALLATE PAPILLAE
C0153350|T047||CCS_10|MALIGNANT TUMOUR OF BASE OF TONGUE
C0153350|T047||CCS_10|MALIGNANT TUMOUR OF FIXED PART OF TONGUE
C0153350|T047||CCS_10|MALIGNANT TUMOUR OF POSTERIOR THIRD OF TONGUE
C0153350|T047||CCS_10|MALIGNANT TUMOUR OF TONGUE POSTERIOR TO VALLATE PAPILLAE
C0153350|T047||CCS_10|MALIGNANT TUMOR OF BASE OF TONGUE 
C0153350|T047||CCS_10|MALIGNANT BASE OF TONGUE NEOPLASM
C0153350|T047||CCS_10|MALIGNANT BASE OF TONGUE TUMOR
C0153350|T047||CCS_10|MALIGNANT BASE OF THE TONGUE NEOPLASM
C0153350|T047||CCS_10|MALIGNANT BASE OF THE TONGUE TUMOR
C0153350|T047||CCS_10|MALIGNANT NEOPLASM OF POSTERIOR TONGUE
C0153350|T047||CCS_10|MALIGNANT NEOPLASM OF THE BASE OF THE TONGUE
C0153350|T047||CCS_10|MALIGNANT NEOPLASM OF THE POSTERIOR TONGUE
C0153350|T047||CCS_10|MALIGNANT POSTERIOR TONGUE NEOPLASM
C0153350|T047||CCS_10|MALIGNANT POSTERIOR TONGUE TUMOR
C0153350|T047||CCS_10|MALIGNANT TUMOR OF POSTERIOR TONGUE
C0153350|T047||CCS_10|MALIGNANT TUMOR OF THE BASE OF THE TONGUE
C0153350|T047||CCS_10|MALIGNANT TUMOR OF THE POSTERIOR TONGUE
C0345741|T047||CCS_10|MALIGNANT NEOPLASM OF FALSE VOCAL CORD
C0345741|T047||CCS_10|MALIGNANT NEOPLASM OF VENTRICULAR BANDS OF LARYNX
C0345741|T047||CCS_10|LARYNGEAL NEOPLASM FALSE VOCAL CORD MALIGNANT
C0345741|T047||CCS_10|MALIGNANT NEOPLASM OF FALSE VOCAL CORD 
C0345741|T047||CCS_10|MALIGNANT TUMOR OF FALSE CORD
C0345741|T047||CCS_10|MALIGNANT TUMOR OF VENTRICULAR BAND
C0345741|T047||CCS_10|MALIGNANT TUMOR OF VESTIBULAR FOLD
C0345741|T047||CCS_10|MALIGNANT TUMOUR OF FALSE CORD
C0345741|T047||CCS_10|MALIGNANT TUMOUR OF VENTRICULAR BAND
C0345741|T047||CCS_10|MALIGNANT TUMOUR OF VESTIBULAR FOLD
C0345741|T047||CCS_10|MALIGNANT TUMOR OF FALSE CORD 
C0345741|T047||CCS_10|MALIGNANT NEOPLASM OF FALSE VOCAL CORDS
C0686013|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF FLOOR OF MOUTH
C0686013|T047||CCS_10|FLOOR OF MOUTH MALIGNANT NEOPLASM SECONDARY
C0686013|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF FLOOR OF MOUTH 
C0686013|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF FLOOR OF MOUTH 
C0686013|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO FLOOR OF MOUTH
C0686013|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO FLOOR OF MOUTH, NOS
C0686013|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF FLOOR OF MOUTH, NOS
C0345756|T047||CCS_10|PHARYNGEAL NEOPLASM MALIGNANT PARAPHARYNEGAL SPACE
C0345756|T047||CCS_10|MALIGNANT NEOPLASM OF PARAPHARYNGEAL SPACE
C0345756|T047||CCS_10|MALIGNANT NEOPLASM OF PARAPHARYNGEAL SPACE 
C0345756|T047||CCS_10|MALIGNANT TUMOR OF PARAPHARYNGEAL SPACE
C0345756|T047||CCS_10|MALIGNANT TUMOUR OF PARAPHARYNGEAL SPACE
C0345756|T047||CCS_10|MALIGNANT TUMOR OF PARAPHARYNGEAL SPACE 
C0685129|T047||CCS_10|MALIGNANT NEOPLASM OF BLOOD VESSEL OF HEAD
C0685129|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF BLOOD VESSEL OF HEAD 
C0685129|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF BLOOD VESSEL OF HEAD
C0685129|T047||CCS_10|NEOPLASM - SOFT TISSUE TYPES BLOOD VESSEL MALIGNANT OF HEAD PRIMARY
C0685129|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF BLOOD VESSEL OF HEAD 
C0153405|T047||CCS_10|MALIGNANT NEOPLASM OF PHARYNX
C0153405|T047||CCS_10|MALIGNANT NEOPLASM OF PHARYNX, UNSPECIFIED
C0153405|T047||CCS_10|PHARYNX, UNSPECIFIED
C0153405|T047||CCS_10|MALIGNANT NEOPLASM OF PHARYNX 
C0153405|T047||CCS_10|MALIGNANT PHARYNGEAL NEOPLASM
C0153405|T047||CCS_10|CANCER, PHARNYX
C0153405|T047||CCS_10|CANCERS, PHARNYX
C0153405|T047||CCS_10|PHARNYX CANCERS
C0153405|T047||CCS_10|CANCER, PHARYNGEAL
C0153405|T047||CCS_10|CANCERS, PHARYNGEAL
C0153405|T047||CCS_10|PHARYNGEAL CANCERS
C0153405|T047||CCS_10|PHARYNX CANCER
C0153405|T047||CCS_10|PHARYNX CANCERS
C0153405|T047||CCS_10|PHARYNGEAL CANCER
C0153405|T047||CCS_10|MALIGNANT TUMOR OF PHARYNX
C0153405|T047||CCS_10|MAL NEO PHARYNX NOS
C0153405|T047||CCS_10|MALIGNANT NEOPLASM OF PHARYNX UNSPECIFIED 
C0153405|T047||CCS_10|MALIGNANT NEOPLASM OF PHARYNX UNSPECIFIED
C0153405|T047||CCS_10|PHARYNX--CANCER
C0153405|T047||CCS_10|PHARYNGEAL CANCER STAGE UNSPECIFIED
C0153405|T047||CCS_10|PHARYNX NEOPLASM MALIGNANT
C0153405|T047||CCS_10|CANCER OF THE PHARYNX
C0153405|T047||CCS_10|PHARNYX CANCER
C0153405|T047||CCS_10|MALIGNANT TUMOUR OF PHARYNX
C0153405|T047||CCS_10|CA - CANCER OF PHARYNX
C0153405|T047||CCS_10|CANCER OF PHARYNX
C0153405|T047||CCS_10|MALIGNANT TUMOR OF PHARYNX 
C0153405|T047||CCS_10|MALIGNANT NEOPLASM OF PHARYNX, NOS
C0153405|T047||CCS_10|MALIGNANT PHARYNGEAL TUMOR
C0153405|T047||CCS_10|MALIGNANT PHARYNX NEOPLASM
C0153405|T047||CCS_10|MALIGNANT PHARYNX TUMOR
C0153405|T047||CCS_10|MALIGNANT TUMOR OF THE PHARYNX
C0346825|T047||CCS_10|MALIGNANT TUMOR OF SOFT TISSUE OF HEAD, FACE AND NECK
C0346825|T047||CCS_10|MALIGNANT TUMOUR OF SOFT TISSUE OF HEAD, FACE AND NECK
C0346825|T047||CCS_10|MALIGNANT TUMOR OF SOFT TISSUE OF HEAD, FACE AND NECK 
C0153760|T047||CCS_10|HODGKIN'S DISEASE, NODULAR SCLEROSIS OF LYMPH NODES OF HEAD, FACE, AND NECK
C0153760|T047||CCS_10|HODGKIN'S DISEASE, NODULAR SCLEROSIS, INVOLVING LYMPH NODES OF HEAD, FACE, AND NECK.
C0153760|T047||CCS_10|HODG NODUL SCLERO HEAD
C0153760|T047||CCS_10|HODGKIN DISEASE, NODULAR SCLEROSIS OF LYMPH NODES OF HEAD, FACE AND NECK
C0153760|T047||CCS_10|HODGKIN DISEASE, NODULAR SCLEROSIS OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0153760|T047||CCS_10|HODGKIN'S DISEASE, NODULAR SCLEROSIS, LYMPH NODES OF HEAD, FACE, AND NECK
C0153760|T047||CCS_10|HODGKIN'S DISEASE, NODULAR SCLEROSIS, INVOLVING LYMPH NODES OF HEAD, FACE, AND NECK
C0153760|T047||CCS_10|NODULAR SCLEROSING HODGKIN'S DISEASE OF LYMPH NODES OF HEAD, FACE, AND NECK
C0153760|T047||CCS_10|NODULAR SCLEROSIS HODGKIN'S LYMPHOMA OF LYMPH NODES OF HEAD, FACE, AND NECK
C0153760|T047||CCS_10|NODULAR SCLEROSING HODGKIN'S DISEASE OF LYMPH NODES OF HEAD, FACE, AND NECK 
C0153760|T047||CCS_10|HODGKIN'S DISEASE, NODULAR SCLEROSIS OF LYMPH NODES OF HEAD, FACE AND NECK
C0153760|T047||CCS_10|HODGKIN'S DISEASE, NODULAR SCLEROSIS OF LYMPH NODES OF HEAD, FACE AND/OR NECK 
C0153760|T047||CCS_10|HODGKIN'S DISEASE, NODULAR SCLEROSIS OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0153760|T047||CCS_10|HODGKIN'S DISEASE, NODULAR SCLEROSIS OF LYMPH NODES OF HEAD, FACE AND NECK 
C0153760|T047||CCS_10|HODGKIN'S DISEASE, NODULAR SCLEROSIS, INVOLVING LYMPH NODES OF HEAD, FACE AND NECK
C0153794|T047||CCS_10|NODULAR LYMPHOMA HEAD
C0153794|T047||CCS_10|NODULAR LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK
C0153794|T047||CCS_10|NODULAR LYMPHOMA INVOLVING LYMPH NODES OF HEAD, FACE, AND NECK
C0153794|T047||CCS_10|NODULAR LYMPHOMA OF LYMPH NODES OF HEAD, FACE, AND NECK 
C0153794|T047||CCS_10|NODULAR LYMPHOMA OF LYMPH NODES OF HEAD, FACE, AND NECK
C0153794|T047||CCS_10|NODULAR LYMPHOMA OF LYMPH NODES OF HEAD, FACE, AND NECK 
C0153794|T047||CCS_10|NODULAR LYMPHOMA OF LYMPH NODES OF HEAD, FACE AND NECK
C0153794|T047||CCS_10|NODULAR LYMPHOMA OF LYMPH NODES OF HEAD, FACE AND NECK 
C0153794|T047||CCS_10|NODULAR LYMPHOMA INVOLVING LYMPH NODES OF HEAD, FACE AND NECK
C1290119|T047||CCS_10|MELANOMA IN SITU OF FACE 
C1290119|T047||CCS_10|MELANOMA IN SITU OF FACE
C1290119|T047||CCS_10|FACE; MELANOMA IN SITU
C1290119|T047||CCS_10|MELANOMA IN SITU; FACE
C0751255|T047||CCS_10|MALIGNANT NEOPLASM OF JAW
C0751255|T047||CCS_10|MALIGNANT NEOPLASM OF JAW 
C0751255|T047||CCS_10|CANCERS, JAW
C0751255|T047||CCS_10|JAW CANCERS
C0751255|T047||CCS_10|MALIGNANT TUMOR OF JAW
C0751255|T047||CCS_10|CANCER, JAW
C0751255|T047||CCS_10|MALIGNANT NEOPLASM OF JAW NOS
C0751255|T047||CCS_10|MALIGNANT NEOPLASM OF JAW NOS 
C0751255|T047||CCS_10|JAWS--CANCER
C0751255|T047||CCS_10|JAW CANCER
C0751255|T047||CCS_10|CANCER OF THE JAW
C0751255|T047||CCS_10|MALIGNANT NEOPLASM OF JAW, NOS
C0751255|T047||CCS_10|CANCER OF JAW
C0346944|T047||CCS_10|MALIGNANT NEOPLASM OF SUPRACLAVICULAR FOSSA NOS
C0346944|T047||CCS_10|MALIGNANT NEOPLASM OF SUPRACLAVICULAR FOSSA NOS 
C1299284|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF FALSE VOCAL CORD
C1299284|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF FALSE VOCAL CORD 
C1299284|T047||CCS_10|LARYNGEAL NEOPLASM FALSE VOCAL CORD MALIGNANT PRIMARY
C1299284|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF FALSE VOCAL CORD 
C0751177|T047||CCS_10|MALIGNANT NEOPLASM OF HEAD
C0751177|T047||CCS_10|HEAD CANCER
C0751177|T047||CCS_10|MALIGNANT NEOPLASM OF HEAD NOS
C0751177|T047||CCS_10|MALIGNANT NEOPLASM OF HEAD NOS 
C0751177|T047||CCS_10|MALIGNANT NEOPLASM OF ILL-DEFINED SITE HEAD
C0751177|T047||CCS_10|MALIGNANT NEOPLASM OF HEAD 
C0751177|T047||CCS_10|HEAD--CANCER
C0751177|T047||CCS_10|CANCER OF HEAD
C0751177|T047||CCS_10|CANCER OF THE HEAD
C0751177|T047||CCS_10|MALIGNANT NEOPLASM OF HEAD, NOS
C0349019|T047||CCS_10|MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF HEAD, FACE AND NECK
C0349019|T047||CCS_10|PERIPHERAL NERVES OF HEAD, FACE AND NECK
C0349019|T047||CCS_10|MALIGNANT NEOPLASM OF PRPH NERVES OF HEAD, FACE AND NECK
C0349019|T047||CCS_10|MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF HEAD, FACE, AND NECK 
C0349019|T047||CCS_10|MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF HEAD, FACE, AND NECK
C0349019|T047||CCS_10|NEOPLASM - PNS PERIPHERAL MALIGNANT HEAD FACE AND NECK
C0349019|T047||CCS_10|MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF HEAD, FACE AND NECK 
C0587060|T047||CCS_10|MALIGNANT MELANOMA OF HEAD AND NECK
C0587060|T047||CCS_10|MALIGNANT MELANOMA OF HEAD AND NECK 
C0587060|T047||CCS_10|MALIGNANT MELANOMA OF HEAD AND NECK 
C0587060|T047||CCS_10|MALIGNANT NEOPLASM OF ILL-DEFINED SITE HEAD AND NECK MELANOMA
C0346568|T047||CCS_10|MALIGNANT NEOPLASM OF EAR, NOSE, AND THROAT 
C0346568|T047||CCS_10|MALIGNANT NEOPLASM OF ILL-DEFINED SITE EAR, NOSE, AND THROAT
C0346568|T047||CCS_10|MALIGNANT NEOPLASM OF EAR, NOSE, AND THROAT
C0346568|T047||CCS_10|MALIGNANT TUMOR OF EAR, NOSE AND THROAT
C0346568|T047||CCS_10|MALIGNANT TUMOUR OF EAR, NOSE AND THROAT
C0346568|T047||CCS_10|MALIGNANT TUMOR OF EAR, NOSE AND THROAT 
C0496836|T047||CCS_10|MALIGNANT NEOPLASM OF EYE, UNSPECIFIED
C0496836|T047||CCS_10|MALIGNANT TUMOR OF EYE
C0496836|T047||CCS_10|MALIGNANT NEOPLASM OF EYE
C0496836|T047||CCS_10|MALIGNANT NEOPLASM OF EYE 
C0496836|T047||CCS_10|EYE CANCER 
C0496836|T047||CCS_10|EYE CANCER
C0496836|T047||CCS_10|MALIGNANT EYE NEOPLASM
C0496836|T047||CCS_10|CANCERS, EYE
C0496836|T047||CCS_10|EYE CANCERS
C0496836|T047||CCS_10|MALIGN NEOPL EYE NOS
C0496836|T047||CCS_10|MALIGNANT NEOPLASM OF UNSPECIFIED SITE OF EYE
C0496836|T047||CCS_10|CANCER, EYE
C0496836|T047||CCS_10|MALIGNANT TUMOUR OF EYE
C0496836|T047||CCS_10|MALIGNANT NEOPLASM OF EYE NOS
C0496836|T047||CCS_10|CA EYE
C0496836|T047||CCS_10|MALIGNANT NEOPLASM OF EYE NOS 
C0496836|T047||CCS_10|EYE--CANCER
C0496836|T047||CCS_10|MALIGNANT EYE CANCER, NOS
C0496836|T047||CCS_10|MALIGNANT NEOPLASM OF EYE, PART UNSPECIFIED
C0496836|T047||CCS_10|MALIGNANT EYE NEOPLASM NOS
C0496836|T047||CCS_10|CANCER OF THE EYE
C0496836|T047||CCS_10|MALIGNANT TUMOR OF EYE 
C0496836|T047||CCS_10|OCULAR CANCER
C0496836|T047||CCS_10|MALIGNANT NEOPLASM OF EYE, NOS
C0496836|T047||CCS_10|CANCER OF EYE
C0496836|T047||CCS_10|EYE NEOPLASM, MALIGNANT
C0496836|T047||CCS_10|MALIGNANT EYE TUMOR
C0496836|T047||CCS_10|MALIGNANT NEOPLASM OF THE EYE
C0496836|T047||CCS_10|MALIGNANT OCULAR NEOPLASM
C0496836|T047||CCS_10|MALIGNANT OCULAR TUMOR
C0496836|T047||CCS_10|MALIGNANT TUMOR OF THE EYE
C0496836|T047||CCS_10|NEOPLASM MALIG;EYE
C0496836|T047||CCS_10|MALIGNANT NEOSPLASM OF THE EYE
C0153645|T047||CCS_10|MALIGNANT NEOPLASM OF CEREBRAL MENINGES
C0153645|T047||CCS_10|MALIGNANT NEOPLASM OF CEREBRAL MENINGES 
C0153645|T047||CCS_10|MALIGNANT TUMOR OF CEREBRAL MENINGES
C0153645|T047||CCS_10|MAL NEO CEREBRAL MENING
C0153645|T047||CCS_10|MALIGNANT NEOPLASM OF CEREBRAL MENINGES NOS 
C0153645|T047||CCS_10|MALIGNANT NEOPLASM OF CEREBRAL MENINGES NOS
C0153645|T047||CCS_10|CANCER OF THE CEREBRAL MENINGES
C0153645|T047||CCS_10|MALIGNANT NEOPLASM OF CEREBRAL MENINGES 
C0346653|T047||CCS_10|MALIGNANT NEOPLASM OF BONES OF SKULL AND FACE
C0346653|T047||CCS_10|MALIGNANT NEOPLASM OF BONES OF SKULL AND FACE NOS 
C0346653|T047||CCS_10|MALIGNANT NEOPLASM OF BONES OF SKULL AND FACE NOS
C0346653|T047||CCS_10|BONE NEOPLASM, MALIGNANT - SKULL AND FACE
C0346653|T047||CCS_10|MALIGNANT NEOPLASM OF BONES OF SKULL AND FACE 
C0346653|T047||CCS_10|MALIGNANT NEOPLASM OF BONES OF SKULL AND FACE 
C0178247|T047||CCS_10|MALIGNANT NEOPLASM OF LIP, ORAL CAVITY AND PHARYNX 
C0178247|T047||CCS_10|MALIGNANT NEOPLASM OF LIP, ORAL CAVITY AND/OR PHARYNX 
C0178247|T047||CCS_10|MALIGNANT NEOPLASMS OF LIP, ORAL CAVITY AND PHARYNX
C0178247|T047||CCS_10|MALIGNANT NEOPLASMS OF LIP, ORAL CAVITY AND PHARYNX (C00-C14)
C0178247|T047||CCS_10|MALIGNANT NEOPLASM OF LIP, ORAL CAVITY AND PHARYNX
C0178247|T047||CCS_10|MALIGNANT NEOPLASM OF LIP, ORAL CAVITY AND PHARYNX NOS
C0178247|T047||CCS_10|CA LIP, ORAL, PHARYNX NOS
C0178247|T047||CCS_10|MALIGNANT NEOPLASM: [LIP] OR [ORAL CAVITY] OR [PHARYNX] 
C0178247|T047||CCS_10|CA LIP, ORAL, PHARYNX
C0178247|T047||CCS_10|MALIGNANT NEOPLASM: [LIP] OR [ORAL CAVITY] OR [PHARYNX]
C0178247|T047||CCS_10|CA LIP, ORAL, PHARYNX NOS 
C0178247|T047||CCS_10|MALIGNANT NEOPLASM OF LIP, ORAL CAVITY AND PHARYNX NOS 
C0178247|T047||CCS_10|MALIGNANT NEOPLASM OF LIP, ORAL CAVITY, AND/OR PHARYNX 
C0178247|T047||CCS_10|MALIGNANT NEOPLASM OF LIP, ORAL CAVITY, AND/OR PHARYNX
C0178247|T047||CCS_10|MALIGNANT NEOPLASM OF LIP, ORAL CAVITY, AND PHARYNX
C1828015|T047||CCS_10|MALIGNANT TUMOR OF EYELID 
C1828015|T047||CCS_10|MALIGNANT NEOPLASM OF EYELID 
C1828015|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF EYELID 
C1828015|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF EYELID
C1828015|T047||CCS_10|MALIGNANT NEOPLASM OF EYELID
C1828015|T047||CCS_10|SKIN NEOPLASM EYELID MALIGNANT
C1828015|T047||CCS_10|MALIGNANT NEOPLASM OF SKIN OF EYELID 
C1828015|T047||CCS_10|MALIGNANT NEOPLASM OF EYELID 
C1828015|T047||CCS_10|NEOPLASM OF OCULAR ADNEXA EYELID MALIGNANT
C1828015|T047||CCS_10|MALIGNANT TUMOR OF EYELID
C1828015|T047||CCS_10|MALIGNANT TUMOUR OF EYELID
C1828015|T047||CCS_10|MALIGNANT EYELID NEOPLASM
C1828015|T047||CCS_10|MALIGNANT EYELID TUMOR
C1828015|T047||CCS_10|MALIGNANT NEOPLASM OF THE EYELID
C1828015|T047||CCS_10|MALIGNANT TUMOR OF THE EYELID
C0684808|T047||CCS_10|MALIGNANT NEOPLASM OF FACE
C0684808|T047||CCS_10|MALIGNANT NEOPLASM OF FACE 
C0684808|T047||CCS_10|MALIGNANT TUMOR OF FACE
C0684808|T047||CCS_10|MALIGNANT TUMOUR OF FACE
C0684808|T047||CCS_10|MALIGNANT TUMOR OF FACE 
C0684808|T047||CCS_10|MALIGNANT NEOPLASM OF FACE, NOS
C0153627|T047||CCS_10|MALIGNANT NEOPLASM OF LACRIMAL GLAND
C0153627|T047||CCS_10|MALIGNANT NEOPLASM OF LACRIMAL GLAND 
C0153627|T047||CCS_10|LACRIMAL GLAND NEOPLASM MALIGNANT
C0153627|T047||CCS_10|MAL NEO LACRIMAL GLAND
C0153627|T047||CCS_10|MALIGNANT TUMOUR OF LACRIMAL GLAND
C0153627|T047||CCS_10|MALIGNANT TUMOUR OF LACRIMAL GLAND 
C0153627|T047||CCS_10|MALIGNANT TUMOR OF LACRIMAL GLAND
C0153627|T047||CCS_10|MALIGNANT TUMOR OF LACRIMAL GLAND 
C0153627|T047||CCS_10|MALIGNANT LACRIMAL GLAND NEOPLASM
C0153627|T047||CCS_10|MALIGNANT LACRIMAL GLAND TUMOR
C0153627|T047||CCS_10|MALIGNANT NEOPLASM OF THE LACRIMAL GLAND
C0153627|T047||CCS_10|MALIGNANT TUMOR OF THE LACRIMAL GLAND
C0153626|T047||CCS_10|MALIGNANT NEOPLASM OF ORBIT
C0153626|T047||CCS_10|MALIGNANT TUMOR OF ORBIT
C0153626|T047||CCS_10|MALIGNANT NEOPLASM OF ORBIT 
C0153626|T047||CCS_10|MALIGN NEOPL ORBIT
C0153626|T047||CCS_10|MALIGNANT NEOPLASM OF ORBIT NOS
C0153626|T047||CCS_10|MALIGNANT NEOPLASM OF ORBIT NOS 
C0153626|T047||CCS_10|MALIGNANT ORBITAL TUMOR
C0153626|T047||CCS_10|MALIGNANT ORBITAL TUMOUR
C0153626|T047||CCS_10|MALIGNANT TUMOUR OF ORBIT
C0153626|T047||CCS_10|MALIGNANT TUMOR OF ORBIT 
C0153626|T047||CCS_10|MALIGNANT NEOPLASM OF THE ORBIT
C0153626|T047||CCS_10|MALIGNANT ORBIT NEOPLASM
C0153626|T047||CCS_10|MALIGNANT ORBIT TUMOR
C0153626|T047||CCS_10|MALIGNANT ORBITAL NEOPLASM
C0153626|T047||CCS_10|MALIGNANT TUMOR OF THE ORBIT
C0686574|T047||CCS_10|MALIGNANT MAST CELL TUMORS INVOLVING LYMPH NODES OF HEAD, FACE, AND NECK
C0686574|T047||CCS_10|MALIGNANT MAST CELL TUMOR OF LYMPH NODES OF HEAD, FACE, AND NECK
C0686574|T047||CCS_10|MALIGNANT MASTOCYTOSIS OF HEAD, FACE, AND NECK 
C0686574|T047||CCS_10|MALIGNANT MASTOCYTOSIS OF HEAD, FACE, AND NECK
C0686574|T047||CCS_10|MAL MASTOCYTOSIS HEAD
C0686574|T047||CCS_10|MALIGNANT MAST CELL TUMORS, LYMPH NODES OF HEAD, FACE, AND NECK
C0686574|T047||CCS_10|MAST CELL MALIGNANCY OF LYMPH NODES OF HEAD, FACE, AND NECK
C0686574|T047||CCS_10|MAST CELL MALIGNANCY OF LYMPH NODES OF HEAD, FACE AND NECK
C0686574|T047||CCS_10|MAST CELL MALIGNANCY OF LYMPH NODES OF HEAD, FACE, AND NECK 
C0686574|T047||CCS_10|MALIGNANT MAST CELL TUMOR OF LYMPH NODES OF HEAD, FACE AND/OR NECK 
C0686574|T047||CCS_10|MALIGNANT MAST CELL TUMOR OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0686574|T047||CCS_10|MALIGNANT MAST CELL TUMOUR OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0686574|T047||CCS_10|MAST CELL MALIGNANCY OF LYMPH NODES OF HEAD, FACE AND NECK 
C0686574|T047||CCS_10|MALIGNANT MAST CELL TUMORS INVOLVING LYMPH NODES OF HEAD, FACE AND NECK
C0346903|T047||CCS_10|MALIGNANT NEOPLASM OF CEREBRUM
C0346903|T047||CCS_10|MALIGNANT NEOPLASM OF CEREBRUM 
C0346903|T047||CCS_10|MALIGNANT NEOPLASM OF CEREBRAL HEMISPHERE 
C0346903|T047||CCS_10|MALIGNANT NEOPLASM OF CEREBRAL HEMISPHERE
C0346903|T047||CCS_10|MALIGNANT TUMOR OF CEREBRAL HEMISPHERE
C0346903|T047||CCS_10|CEREBRAL TUMOR (MALIGNANT)
C0346903|T047||CCS_10|CEREBRAL TUMOR - MALIGNANT 
C0346903|T047||CCS_10|CEREBRUM CA 
C0346903|T047||CCS_10|MALIGNANT CEREBRAL TUMOR
C0346903|T047||CCS_10|MALIGNANT NEOPLASM OF CEREBRUM NOS
C0346903|T047||CCS_10|CEREBRUM CA
C0346903|T047||CCS_10|CEREBRAL TUMOUR (MALIGNANT)
C0346903|T047||CCS_10|CEREBRAL TUMOUR - MALIGNANT
C0346903|T047||CCS_10|MALIGNANT NEOPLASM OF CEREBRUM NOS 
C0346903|T047||CCS_10|CEREBRAL TUMOR - MALIGNANT
C0346903|T047||CCS_10|MALIGNANT CEREBRAL TUMOUR
C0346903|T047||CCS_10|MALIGNANT NEOPLASM OF CEREBRUM 
C0346903|T047||CCS_10|BRAIN TUMOR MALIGNANT OF CEREBRUM
C0346903|T047||CCS_10|MALIGNANT NEOPLASM OF CEREBRUM, NOS
C0346903|T047||CCS_10|MALIGNANT CEREBRAL HEMISPHERIC NEOPLASM
C0346903|T047||CCS_10|MALIGNANT CEREBRAL HEMISPHERIC TUMOR
C0346903|T047||CCS_10|MALIGNANT CEREBRAL NEOPLASM
C0346903|T047||CCS_10|MALIGNANT NEOPLASM OF CEREBRAL HEMISPHERES
C0346903|T047||CCS_10|MALIGNANT NEOPLASM OF THE CEREBRAL HEMISPHERES
C0346903|T047||CCS_10|MALIGNANT NEOPLASM OF THE CEREBRUM
C0346903|T047||CCS_10|MALIGNANT TUMOR OF CEREBRAL HEMISPHERES
C0346903|T047||CCS_10|MALIGNANT TUMOR OF CEREBRUM
C0346903|T047||CCS_10|MALIGNANT TUMOR OF THE CEREBRAL HEMISPHERES
C0346903|T047||CCS_10|MALIGNANT TUMOR OF THE CEREBRUM
C0346903|T047||CCS_10|CEREBRAL CANCER
C0580284|T047||CCS_10|METASTASIS TO HEAD AND NECK LYMPH NODE
C0580284|T047||CCS_10|METASTASIS TO HEAD AND NECK LYMPH NODE 
C0580284|T047||CCS_10|METASTASIS TO HEAD AND NECK LYMPH NODE 
C0580284|T047||CCS_10|METASTATIC CANCER TO HEAD AND NECK LYMPH NODE
C1306467|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF HEAD 
C1306467|T047||CCS_10|MALIGNANT NEOPLASM OF ILL-DEFINED SITE HEAD PRIMARY
C1306467|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF HEAD
C1306467|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF HEAD 
C0349750|T047||CCS_10|EYE NEOPLASM MALIGNANT LACRIMAL DRAINAGE STRUCTURE
C0349750|T047||CCS_10|MALIGNANT NEOPLASM OF LACRIMAL DRAINAGE STRUCTURE 
C0349750|T047||CCS_10|MALIGNANT NEOPLASM OF LACRIMAL DRAINAGE STRUCTURE
C0349750|T047||CCS_10|MALIGNANT TUMOR OF LACRIMAL DRAINAGE STRUCTURE
C0349750|T047||CCS_10|MALIGNANT TUMOUR OF LACRIMAL DRAINAGE STRUCTURE
C0349750|T047||CCS_10|MALIGNANT TUMOR OF LACRIMAL DRAINAGE STRUCTURE 
C0684805|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF HEAD
C0684805|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF HEAD 
C0684805|T047||CCS_10|MALIGNANT NEOPLASM OF ILL-DEFINED SITE HEAD SECONDARY
C0684805|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO HEAD
C0684805|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF HEAD 
C0684805|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO HEAD, NOS
C0684805|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF HEAD, NOS
C0432547|T047||CCS_10|LETTERER-SIWE DISEASE OF LYMPH NODES OF HEAD, FACE, AND NECK
C0432547|T047||CCS_10|LETTERER-SIWE DISEASE OF HEAD, FACE, OR NECK
C0432547|T047||CCS_10|LETTERER-SIWE DISEASE OF HEAD, FACE, OR NECK 
C0432547|T047||CCS_10|LETTERER-SIWE DIS HEAD
C0432547|T047||CCS_10|LETTERER-SIWE DISEASE, LYMPH NODES OF HEAD, FACE, AND NECK
C0432547|T047||CCS_10|LETTERER-SIWE DISEASE INVOLVING LYMPH NODES OF HEAD, FACE, AND NECK
C0432547|T047||CCS_10|LETTERER-SIWE DISEASE OF LYMPH NODES OF HEAD, FACE AND NECK
C0432547|T047||CCS_10|LETTERER-SIWE DISEASE OF LYMPH NODES OF HEAD, FACE AND NECK 
C0432547|T047||CCS_10|LETTERER-SIWE DISEASE OF LYMPH NODES OF HEAD, FACE AND/OR NECK 
C0432547|T047||CCS_10|LETTERER-SIWE DISEASE OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0432547|T047||CCS_10|LETTERER-SIWE DISEASE INVOLVING LYMPH NODES OF HEAD, FACE AND NECK
C0432538|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF LYMPH NODES OF HEAD, FACE, AND NECK
C0432538|T047||CCS_10|MAL HISTIOCYTOSIS HEAD
C0432538|T047||CCS_10|MALIGNANT HISTIOCYTOSIS, LYMPH NODES OF HEAD, FACE, AND NECK
C0432538|T047||CCS_10|MALIGNANT HISTIOCYTOSIS INVOLVING LYMPH NODES OF HEAD, FACE, AND NECK
C0432538|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF LYMPH NODES OF HEAD, FACE, AND NECK 
C0432538|T047||CCS_10|RETICULOENDOTHELIAL SYSTEM MALIGNANT HISTIOCYTOSIS LYMPH NODE HEAD, FACE, NECK
C0432538|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF LYMPH NODES OF HEAD, FACE AND NECK
C0432538|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF LYMPH NODES OF HEAD, FACE AND/OR NECK 
C0432538|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0432538|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF LYMPH NODES OF HEAD, FACE AND NECK 
C0432538|T047||CCS_10|MALIGNANT HISTIOCYTOSIS INVOLVING LYMPH NODES OF HEAD, FACE AND NECK
C0432556|T047||CCS_10|LYMPHOMA OF HEAD, FACE, AND NECK
C0432556|T047||CCS_10|LYMPHOMA OF HEAD, FACE, AND NECK 
C0432556|T047||CCS_10|MALIGNANT LYMPHOMA NOS OF LYMPH NODES OF HEAD, FACE AND NECK 
C0432556|T047||CCS_10|MALIGNANT LYMPHOMA NOS OF LYMPH NODES OF HEAD, FACE AND NECK
C0432556|T047||CCS_10|MALIGNANT LYMPHOMA OF LYMPH NODES OF HEAD, FACE AND/OR NECK 
C0432556|T047||CCS_10|MALIGNANT LYMPHOMA OF LYMPH NODES OF HEAD, FACE AND/OR NECK
C0432556|T047||CCS_10|MALIGNANT LYMPHOMA, NOS OF LYMPH NODES OF HEAD, FACE, AND NECK
C1719786|T047||CCS_10|MALIGNANT LYMPHOMA OF THE EYE REGION 
C1719786|T047||CCS_10|MALIGNANT LYMPHOMA OF THE EYE REGION
C1827431|T047||CCS_10|SARCOMA OF HEAD AND NECK 
C1827431|T047||CCS_10|SARCOMA OF HEAD AND NECK
C1827431|T047||CCS_10|MALIGNANT NEOPLASM SARCOMA OF HEAD AND NECK 
C1827431|T047||CCS_10|MALIGNANT NEOPLASM SARCOMA OF HEAD AND NECK
C0007107|T047||CCS_10|MALIGNANT NEOPLASM OF LARYNX
C0007107|T047||CCS_10|LARYNGEAL CANCER
C0007107|T047||CCS_10|MALIGNANT NEOPLASM OF LARYNX, UNSPECIFIED
C0007107|T047||CCS_10|MALIGNANT NEOPLASM OF LARYNX 
C0007107|T047||CCS_10|MALIGNANT LARYNGEAL NEOPLASM
C0007107|T047||CCS_10|CANCER, LARYNGEAL
C0007107|T047||CCS_10|CANCERS, LARYNGEAL
C0007107|T047||CCS_10|LARYNGEAL CANCERS
C0007107|T047||CCS_10|CANCERS, LARYNX
C0007107|T047||CCS_10|LARYNX CANCERS
C0007107|T047||CCS_10|MALIGNANT TUMOR OF LARYNX
C0007107|T047||CCS_10|CANCER OF LARYNX
C0007107|T047||CCS_10|MALIGNANT NEO LARYNX NOS
C0007107|T047||CCS_10|CANCER, LARYNX
C0007107|T047||CCS_10|LARYNGEAL NEOPLASMS MALIGNANT
C0007107|T047||CCS_10|LARYNGEAL CANCER 
C0007107|T047||CCS_10|MALIGNANT NEOPLASM OF LARYNX NOS 
C0007107|T047||CCS_10|CA LARYNX - NOS
C0007107|T047||CCS_10|MALIGNANT NEOPLASM OF LARYNX NOS
C0007107|T047||CCS_10|CA LARYNX - NOS 
C0007107|T047||CCS_10|MALIGNANT TUMOUR OF LARYNX
C0007107|T047||CCS_10|CA - CANCER OF LARYNX
C0007107|T047||CCS_10|LARYNX--CANCER
C0007107|T047||CCS_10|LARYNGEAL CANCER NOS
C0007107|T047||CCS_10|LARYNX CANCER
C0007107|T047||CCS_10|LARYNX NEOPLASM MALIGNANT
C0007107|T047||CCS_10|CANCER OF THE LARYNX
C0007107|T047||CCS_10|MALIGNANT TUMOR OF LARYNX 
C0007107|T047||CCS_10|MALIGNANT NEOPLASM OF LARYNX, NOS
C0007107|T047||CCS_10|MALIGNANT LARYNGEAL TUMOR
C0007107|T047||CCS_10|MALIGNANT LARYNX NEOPLASM
C0007107|T047||CCS_10|MALIGNANT LARYNX TUMOR
C0007107|T047||CCS_10|MALIGNANT NEOPLASM OF THE LARYNX
C0007107|T047||CCS_10|MALIGNANT TUMOR OF THE LARYNX
C0007107|T047||CCS_10|NEOPLASM MALIG;LARYNX
C0007107|T047||CCS_10|MALIGNANT NEOSPLASM OF THE LARYNX
C0220635|T047||CCS_10|SQUAMOUS CELL CARCINOMA METASTATIC IN THE NECK WITH OCCULT PRIMARY
C0220635|T047||CCS_10|SQUAMOUS CELL CARCINOMA METASTATIC TO THE NECK WITH OCCULT PRIMARY
C0220635|T047||CCS_10|EPIDERMOID CARCINOMA METASTATIC TO THE NECK WITH OCCULT PRIMARY
C0220635|T047||CCS_10|METASTATIC SQUAMOUS NECK CANCER WITH OCCULT PRIMARY
C0220635|T047||CCS_10|NECK CANCER, METASTATIC SQUAMOUS WITH OCCULT PRIMARY
C0220635|T047||CCS_10|OCCULT PRIMARY CANCER METASTATIC SQUAMOUS TO THE NECK
C0238301|T047||CCS_10|CANCER, NASOPHARYNGEAL
C0238301|T047||CCS_10|CANCERS, NASOPHARYNGEAL
C0238301|T047||CCS_10|NASOPHARYNGEAL CANCERS
C0238301|T047||CCS_10|CANCERS, NASOPHARYNX
C0238301|T047||CCS_10|NASOPHARYNX CANCERS
C0238301|T047||CCS_10|CANCER, NASOPHARYNX
C0238301|T047||CCS_10|CANCER OF NASOPHARYNX
C0238301|T047||CCS_10|NASOPHARYNGEAL CANCER
C0238301|T047||CCS_10|NASOPHARYNX--CANCER
C0238301|T047||CCS_10|CANCER OF THE NASOPHARYNX
C0238301|T047||CCS_10|NASOPHARYNX CANCER
C0238301|T047||CCS_10|CA - CANCER OF NASOPHARYNX
C1710095|T047||CCS_10|SINONASAL CARCINOMA
C1710095|T047||CCS_10|NASAL CAVITY AND PARANASAL SINUS CARCINOMA
C1710095|T047||CCS_10|PARANASAL SINUS AND NASAL CAVITY CANCER
C1710095|T047||CCS_10|NASAL CAVITY AND PARANASAL SINUS CANCER
C0153398|T047||CCS_10|MALIGNANT NEOPLASM OF HYPOPHARYNX
C0153398|T047||CCS_10|MALIGNANT NEOPLASM OF HYPOPHARYNX, UNSPECIFIED
C0153398|T047||CCS_10|MALIGNANT NEOPLASM OF HYPOPHARYNX 
C0153398|T047||CCS_10|MALIGNANT HYPOPHARYNGEAL NEOPLASM
C0153398|T047||CCS_10|CANCER, HYPOPHARYNGEAL
C0153398|T047||CCS_10|CANCERS, HYPOPHARYNGEAL
C0153398|T047||CCS_10|HYPOPHARYNGEAL CANCERS
C0153398|T047||CCS_10|MALIGNANT TUMOR OF HYPOPHARYNX
C0153398|T047||CCS_10|MAL NEO HYPOPHARYNX NOS
C0153398|T047||CCS_10|MALIGNANT NEOPLASM OF HYPOPHARYNX, UNSPECIFIED SITE
C0153398|T047||CCS_10|HYPOPHARYNGEAL CANCER
C0153398|T047||CCS_10|MALIGNANT NEOPLASM OF HYPOPHARYNX NOS 
C0153398|T047||CCS_10|MALIGNANT TUMOUR OF HYPOPHARYNX
C0153398|T047||CCS_10|MALIGNANT NEOPLASM OF HYPOPHARYNX NOS
C0153398|T047||CCS_10|MALIGNANT TUMOUR OF HYPOPHARYNX 
C0153398|T047||CCS_10|HYPOPHARYNX--CANCER
C0153398|T047||CCS_10|MALIGNANT NEOPLASM OF LARYNGOPHARYNX
C0153398|T047||CCS_10|MALIGNANT TUMOR OF LARYNGOPHARYNX
C0153398|T047||CCS_10|MALIGNANT TUMOUR OF LARYNGOPHARYNX
C0153398|T047||CCS_10|MALIGNANT TUMOR OF HYPOPHARYNX 
C0153398|T047||CCS_10|HYPOPHARYNX CANCER
C0153398|T047||CCS_10|MALIGNANT NEOPLASM OF HYPOPHARYNX, NOS
C0153398|T047||CCS_10|MALIGNANT HYPOPHARYNGEAL TUMOR
C0153398|T047||CCS_10|MALIGNANT NEOPLASM OF THE HYPOPHARYNX
C0153398|T047||CCS_10|MALIGNANT TUMOR OF THE HYPOPHARYNX
C0687150|T047||CCS_10|PARATHYROID CARCINOMA
C0687150|T047||CCS_10|PARATHYROID GLAND CARCINOMA
C0687150|T047||CCS_10|PARATHYROID CARCINOMAS
C0687150|T047||CCS_10|CARCINOMA OF PARATHYROID GLAND 
C0687150|T047||CCS_10|ADENOCARCINOMA OF PARATHYROID GLAND
C0687150|T047||CCS_10|ADENOCARCINOMA OF PARATHYROID GLAND 
C0687150|T047||CCS_10|CARCINOMA OF PARATHYROID GLAND
C0687150|T047||CCS_10|CANCERS, PARATHYROID
C0687150|T047||CCS_10|PARATHYROID CANCERS
C0687150|T047||CCS_10|PARATHYROID ADENOCARCINOMA
C0687150|T047||CCS_10|PARATHYROID GLAND CANCER
C0687150|T047||CCS_10|CANCER, PARATHYROID
C0687150|T047||CCS_10|PARATHYROID CANCER
C0687150|T047||CCS_10|PARATHYROID CANCER, NOS
C0687150|T047||CCS_10|PRTC
C0687150|T047||CCS_10|CANCER OF PARATHYROID
C0687150|T047||CCS_10|CANCER OF THE PARATHYROID
C0687150|T047||CCS_10|PARATHYROID CARCINOMA 
C0687150|T047||CCS_10|CARCINOMA OF THE PARATHYROID
C0687150|T047||CCS_10|PARATHYROID GLAND ADENOCARCINOMA
C0687150|T047||CCS_10|ADENOCARCINOMA OF PARATHYROID
C0687150|T047||CCS_10|ADENOCARCINOMA OF THE PARATHYROID GLAND
C0687150|T047||CCS_10|ADENOCARCINOMA OF THE PARATHYROID
C0687150|T047||CCS_10|CANCER OF PARATHYROID GLAND
C0687150|T047||CCS_10|CANCER OF THE PARATHYROID GLAND
C0687150|T047||CCS_10|CARCINOMA OF PARATHYROID
C0687150|T047||CCS_10|CARCINOMA OF THE PARATHYROID GLAND
C0687150|T047||CCS_10|CARCINOMA, PARATHYROID
C0687150|T047||CCS_10|CARCINOMAS, PARATHYROID
C2349952|T047||CCS_10|CARCINOMA OF OROPHARYNX 
C2349952|T047||CCS_10|CARCINOMA OF OROPHARYNX
C2349952|T047||CCS_10|OROPHARYNGEAL CARCINOMA
C2349952|T047||CCS_10|OROPHARNYX CANCER
C2349952|T047||CCS_10|OROPHARNYX CANCERS
C2349952|T047||CCS_10|CANCER, OROPHARYNGEAL
C2349952|T047||CCS_10|CANCERS, OROPHARYNGEAL
C2349952|T047||CCS_10|OROPHARYNGEAL CANCERS
C2349952|T047||CCS_10|CANCER, OROPHARYNX
C2349952|T047||CCS_10|CANCERS, OROPHARYNX
C2349952|T047||CCS_10|OROPHARYNX CANCERS
C2349952|T047||CCS_10|OROPHARYNGEAL CANCER
C2349952|T047||CCS_10|CANCER OF THE OROPHARYNX
C2349952|T047||CCS_10|OROPHARYNX CANCER
C2349952|T047||CCS_10|OROPHARYNX CARCINOMA
C2349952|T047||CCS_10|CANCER OF OROPHARYNX
C2349952|T047||CCS_10|CARCINOMA OF THE OROPHARYNX
C2349952|T047||CCS_10|CANCER OF OROPHARNYX
C0220641|T047||CCS_10|ORAL CANCER
C0220641|T047||CCS_10|ORAL CARCINOMA
C0220641|T047||CCS_10|LIP AND ORAL CAVITY CARCINOMA
C0220641|T047||CCS_10|LIP AND ORAL CAVITY CANCER
C0220641|T047||CCS_10|ORAL CAVITY AND LIP CANCER
C0496842|T047||CCS_10|MALIGNANT NEOPLASM OF PITUITARY GLAND
C0496842|T047||CCS_10|MALIGNANT NEOPLASM OF PITUITARY GLAND 
C0496842|T047||CCS_10|MALIGNANT PITUITARY NEOPLASM
C0496842|T047||CCS_10|MALIGNANT TUMOR OF PITUITARY GLAND
C0496842|T047||CCS_10|PITUITARY CANCER
C0496842|T047||CCS_10|MALIGNANT PITUITARY TUMOUR
C0496842|T047||CCS_10|PITUITARY TUMOR MALIGNANT
C0496842|T047||CCS_10|MALIGNANT PITUITARY TUMOR
C0496842|T047||CCS_10|PITUITARY TUMOUR MALIGNANT NOS
C0496842|T047||CCS_10|PITUITARY TUMOUR MALIGNANT
C0496842|T047||CCS_10|PITUITARY TUMOR MALIGNANT NOS
C0496842|T047||CCS_10|MALIGNANT TUMOUR OF PITUITARY GLAND
C0496842|T047||CCS_10|CA - CANCER OF PITUITARY GLAND
C0496842|T047||CCS_10|CANCER OF PITUITARY GLAND
C0496842|T047||CCS_10|MALIGNANT TUMOR OF PITUITARY GLAND 
C0496842|T047||CCS_10|MALIGNANT NEOPLASM OF PITUITARY
C0496842|T047||CCS_10|MALIGNANT NEOPLASM OF THE PITUITARY GLAND
C0496842|T047||CCS_10|MALIGNANT NEOPLASM OF THE PITUITARY
C0496842|T047||CCS_10|MALIGNANT PITUITARY GLAND NEOPLASM
C0496842|T047||CCS_10|MALIGNANT PITUITARY GLAND TUMOR
C0496842|T047||CCS_10|MALIGNANT TUMOR OF PITUITARY
C0496842|T047||CCS_10|MALIGNANT TUMOR OF THE PITUITARY GLAND
C0496842|T047||CCS_10|MALIGNANT TUMOR OF THE PITUITARY
C0496842|T047||CCS_10|PITUITARY NEOPLASMS, MALIGNANT
C0496842|T047||CCS_10|PITUITARY TUMOR, MALIGNANT
C0153656|T047||CCS_10|MALIGNANT NEOPLASM OF CAROTID BODY
C0153656|T047||CCS_10|CAROTID BODY TUMOR MALIGNANT
C0153656|T047||CCS_10|MALIGNANT NEOPLASM OF CAROTID BODY 
C0153656|T047||CCS_10|MAL NEO CAROTID BODY
C0153656|T047||CCS_10|MALIGNANT NEOPLASM OF CAROTID BODY 
C0153656|T047||CCS_10|CANCER OF CAROTID BODY
C0153656|T047||CCS_10|CHEMODECTOMA, MALIGNANT
C0153656|T047||CCS_10|MALIGNANT CAROTID BODY NEOPLASM
C0153656|T047||CCS_10|MALIGNANT TUMOR OF CAROTID BODY
C0153656|T047||CCS_10|MALIGNANT TUMOR OF THE CAROTID BODY
C0153656|T047||CCS_10|MALIGNANT CAROTID BODY TUMOR
C0153656|T047||CCS_10|MALIGNANT NEOPLASM OF THE CAROTID BODY
C0153656|T047||CCS_10|MALIGNANT CAROTID BODY TUMOUR
C0153656|T047||CCS_10|MALIGNANT CAROTID BODY TUMOR (MORPHOLOGIC ABNORMALITY)
C0153656|T047||CCS_10|MALIGNANT CAROTID BODY PARAGANGLIOMA
C0153474|T047||CCS_10|MALIGNANT NEOPLASM OF ACCESSORY SINUS, UNSPECIFIED
C0153474|T047||CCS_10|MALIGNANT TUMOR OF NASAL SINUSES
C0153474|T047||CCS_10|MALIGNANT NEOPLASM OF ACCESSORY SINUSES
C0153474|T047||CCS_10|MALIGNANT NEOPLASM OF ACCESSORY SINUS
C0153474|T047||CCS_10|MALIGNANT NEOPLASM OF ACCESSORY SINUS 
C0153474|T047||CCS_10|NASAL SINUS CANCER
C0153474|T047||CCS_10|MALIGNANT TUMOR OF ACCESSORY SINUS
C0153474|T047||CCS_10|MAL NEO ACCESS SINUS NOS
C0153474|T047||CCS_10|MALIGNANT NEOPLASM OF ACCESSORY SINUS NOS 
C0153474|T047||CCS_10|MALIGNANT NEOPLASM OF ACCESSORY SINUS NOS
C0153474|T047||CCS_10|MALIGNANT TUMOUR OF NASAL SINUSES
C0153474|T047||CCS_10|MALIGNANT TUMOR OF NASAL SINUSES 
C0153474|T047||CCS_10|MALIGNANT NEOPLASM OF ACCESSORY SINUS, NOS
C0153474|T047||CCS_10|MALIGNANT ACCESSORY SINUS NEOPLASM
C0153474|T047||CCS_10|MALIGNANT ACCESSORY SINUS TUMOR
C0153474|T047||CCS_10|MALIGNANT NEOPLASM OF PARANASAL SINUS
C0153474|T047||CCS_10|MALIGNANT NEOPLASM OF THE ACCESSORY SINUS
C0153474|T047||CCS_10|MALIGNANT NEOPLASM OF THE PARANASAL SINUS
C0153474|T047||CCS_10|MALIGNANT PARANASAL SINUS NEOPLASM
C0153474|T047||CCS_10|MALIGNANT PARANASAL SINUS TUMOR
C0153474|T047||CCS_10|MALIGNANT TUMOR OF PARANASAL SINUS
C0153474|T047||CCS_10|MALIGNANT TUMOR OF THE ACCESSORY SINUS
C0153474|T047||CCS_10|MALIGNANT TUMOR OF THE PARANASAL SINUS
C0728864|T047||CCS_10|MALIGNANT NEOPLASM OF NASAL CAVITY
C0728864|T047||CCS_10|MALIGNANT NEOPLASM OF NASAL CAVITY 
C0728864|T047||CCS_10|NASAL CAVITY CANCER 
C0728864|T047||CCS_10|NASAL CAVITY CANCER
C0728864|T047||CCS_10|MALIGNANT NASAL CAVITY NEOPLASM
C0728864|T047||CCS_10|MALIGNANT TUMOR OF NASAL CAVITY
C0728864|T047||CCS_10|MAL NEO NASAL CAVITIES
C0728864|T047||CCS_10|CANCER OF THE NASAL CAVITY
C0728864|T047||CCS_10|MALIGNANT NEOPLASM OF NASAL CAVITIES NOS 
C0728864|T047||CCS_10|MALIGNANT NEOPLASM OF NASAL CAVITIES NOS
C0728864|T047||CCS_10|MALIGNANT NEOPLASM OF NASAL CAVITIES
C0728864|T047||CCS_10|MALIGNANT TUMOUR OF NASAL CAVITY
C0728864|T047||CCS_10|MALIGNANT TUMOR OF NASAL CAVITY 
C0728864|T047||CCS_10|MALIGNANT NEOPLASM OF NASAL CAVITY, NOS
C0728864|T047||CCS_10|MALIGNANT NASAL CAVITY TUMOR
C0728864|T047||CCS_10|MALIGNANT NEOPLASM OF THE NASAL CAVITY
C0728864|T047||CCS_10|MALIGNANT TUMOR OF THE NASAL CAVITY
C3887461|T047||CCS_10|HEAD AND NECK CARCINOMA
C3887461|T047||CCS_10|CARCINOMA OF HEAD AND NECK
C3887461|T047||CCS_10|CARCINOMA OF THE HEAD AND NECK
C0347856|T047||CCS_10|MALIGNANT NEOPLASM OF GLOMUS JUGULARE
C0347856|T047||CCS_10|MALIGNANT NEOPLASM OF GLOMUS JUGULARE 
C0347856|T047||CCS_10|MALIGNANT TUMOR OF GLOMUS JUGULARE
C0347856|T047||CCS_10|MALIGNANT NEOPLASM OF GLOMUS JUGULARE 
C0347856|T047||CCS_10|GLOMUS JUGULARE NEOPLASM MALIGNANT PRIMARY
C0347856|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF GLOMUS JUGULARE 
C0347856|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF GLOMUS JUGULARE
C0347856|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF GLOMUS JUGULARE 
C0347856|T047||CCS_10|MALIGNANT GLOMUS JUGULARE NEOPLASM
C0347856|T047||CCS_10|MALIGNANT GLOMUS JUGULARE TUMOR
C0347856|T047||CCS_10|MALIGNANT JUGULOTYMPANIC PARAGANGLIOMA
C0347856|T047||CCS_10|MALIGNANT NEOPLASM OF THE GLOMUS JUGULARE
C0347856|T047||CCS_10|MALIGNANT TUMOR OF THE GLOMUS JUGULARE
C2350059|T047||CCS_10|CANCER OF EAR
C2350059|T047||CCS_10|MALIGNANT NEOPLASM OF EAR 
C2350059|T047||CCS_10|MALIGNANT NEOPLASM OF EAR
C2350059|T047||CCS_10|EAR NEOPLASM MALIGNANT
C2350059|T047||CCS_10|MALIGNANT NEOPLASM OF EAR 
C2350059|T047||CCS_10|NEOPLASM OF EAR MALIGNANT
C2350059|T047||CCS_10|EAR CANCER
C2350059|T047||CCS_10|CANCER OF THE EAR
C2350059|T047||CCS_10|MALIGNANT EAR NEOPLASM
C2350059|T047||CCS_10|MALIGNANT EAR TUMOR
C2350059|T047||CCS_10|MALIGNANT NEOPLASM OF THE EAR
C2350059|T047||CCS_10|MALIGNANT TUMOR OF EAR
C2350059|T047||CCS_10|MALIGNANT TUMOR OF THE EAR
C2350059|T047||CCS_10|NEOPLASM MALIG;EAR
C2350059|T047||CCS_10|MALIGNANT NEOSPLASM OF THE EAR
C1335975|T047||CCS_10|CHORDOMA OF SKULL BASE
C1335975|T047||CCS_10|CHORDOMA OF THE SKULL BASE
C1335975|T047||CCS_10|SKULL BASE CHORDOMA
C0153633|T047||CCS_10|MALIGNANT NEOPLASM OF BRAIN
C0153633|T047||CCS_10|MALIGNANT BRAIN NEOPLASM
C0153633|T047||CCS_10|MALIGNANT NEOPLASM OF BRAIN, UNSPECIFIED
C0153633|T047||CCS_10|BRAIN, UNSPECIFIED
C0153633|T047||CCS_10|MALIGNANT NEOPL BRAIN
C0153633|T047||CCS_10|NEOPL BRAIN MALIGNANT
C0153633|T047||CCS_10|BRAIN NEOPL MALIGNANT
C0153633|T047||CCS_10|MALIGNANT NEOPLASM OF BRAIN 
C0153633|T047||CCS_10|MALIGNANT NEOPLASM OF BRAIN 
C0153633|T047||CCS_10|BRAIN CANCER 
C0153633|T047||CCS_10|BRAIN CANCER
C0153633|T047||CCS_10|MALIGNANT BRAIN TUMOR
C0153633|T047||CCS_10|BRAIN CANCERS
C0153633|T047||CCS_10|CANCERS, BRAIN
C0153633|T047||CCS_10|BRAIN MALIGNANT NEOPLASM
C0153633|T047||CCS_10|BRAIN MALIGNANT NEOPLASMS
C0153633|T047||CCS_10|BRAIN NEOPLASM, MALIGNANT
C0153633|T047||CCS_10|MALIGNANT BRAIN NEOPLASMS
C0153633|T047||CCS_10|MALIGNANT NEOPLASM, BRAIN
C0153633|T047||CCS_10|CANCER OF BRAIN
C0153633|T047||CCS_10|MALIGNANT TUMOR OF BRAIN
C0153633|T047||CCS_10|MALIG NEO BRAIN NOS
C0153633|T047||CCS_10|CANCER, BRAIN
C0153633|T047||CCS_10|BRAIN CA
C0153633|T047||CCS_10|MALIGNANT NEOPLASM OF BRAIN NOS 
C0153633|T047||CCS_10|MALIGNANT BRAIN TUMOUR 
C0153633|T047||CCS_10|MALIGNANT BRAIN TUMOUR
C0153633|T047||CCS_10|MALIGNANT NEOPLASM OF BRAIN NOS
C0153633|T047||CCS_10|BRAIN--CANCER
C0153633|T047||CCS_10|MALIGNANT BRAIN NEOPLASM NOS
C0153633|T047||CCS_10|BRAIN NEOPLASM MALIGNANT
C0153633|T047||CCS_10|BRAIN NEOPLASMS, MALIGNANT
C0153633|T047||CCS_10|MALIGNANT NEOPLASMS, BRAIN
C0153633|T047||CCS_10|CANCER OF THE BRAIN
C0153633|T047||CCS_10|NEOPLASMS, BRAIN, MALIGNANT
C0153633|T047||CCS_10|MALIGNANT NEOPLASM OF BRAIN, NOS
C0153633|T047||CCS_10|MALIGNANT NEOPLASM OF THE BRAIN
C0153633|T047||CCS_10|MALIGNANT TUMOR OF THE BRAIN
C0153633|T047||CCS_10|NEOPLASM MALIG;BRAIN
C0153633|T047||CCS_10|MALIGNANT NEOSPLASM OF THE BRAIN
C0518967|T047||CCS_10|CARCINOMA OF HEAD OF PANCREAS
C0518967|T047||CCS_10|CARCINOMA OF HEAD OF PANCREAS 
C0518967|T047||CCS_10|PANCREATIC NEOPLASM MALIGNANT HEAD, CARCINOMA
C0518967|T047||CCS_10|CARCINOMA OF HEAD OF PANCREAS 
C0153459|T047||CCS_10|MALIGNANT NEOPLASM OF BODY OF PANCREAS
C0153459|T047||CCS_10|BODY OF PANCREAS
C0153459|T047||CCS_10|MAL NEO PANCREAS BODY
C0153459|T047||CCS_10|CA BODY OF PANCREAS
C0153459|T047||CCS_10|CA BODY OF PANCREAS 
C0153459|T047||CCS_10|PANCREATIC NEOPLASM MALIGNANT BODY
C0153459|T047||CCS_10|MALIGNANT NEOPLASM OF BODY OF PANCREAS 
C0153459|T047||CCS_10|MALIGNANT TUMOR OF BODY OF PANCREAS
C0153459|T047||CCS_10|MALIGNANT TUMOUR OF BODY OF PANCREAS
C0153459|T047||CCS_10|MALIGNANT TUMOR OF BODY OF PANCREAS 
C0153460|T047||CCS_10|MALIGNANT NEOPLASM OF TAIL OF PANCREAS
C0153460|T047||CCS_10|TAIL OF PANCREAS
C0153460|T047||CCS_10|MAL NEO PANCREAS TAIL
C0153460|T047||CCS_10|MALIGNANT NEOPLASM OF PANCREATIC TAIL
C0153460|T047||CCS_10|CA TAIL OF PANCREAS 
C0153460|T047||CCS_10|CA TAIL OF PANCREAS
C0153460|T047||CCS_10|MALIGNANT NEOPLASM OF TAIL OF PANCREAS 
C0153460|T047||CCS_10|PANCREATIC NEOPLASM MALIGNANT TAIL
C0153460|T047||CCS_10|MALIGNANT TUMOR OF TAIL OF PANCREAS
C0153460|T047||CCS_10|MALIGNANT TUMOUR OF TAIL OF PANCREAS
C0153460|T047||CCS_10|MALIGNANT TUMOR OF TAIL OF PANCREAS 
C0153458|T047||CCS_10|MALIGNANT NEOPLASM OF HEAD OF PANCREAS
C0153458|T047||CCS_10|HEAD OF PANCREAS
C0153458|T047||CCS_10|MAL NEO PANCREAS HEAD
C0153458|T047||CCS_10|MALIGNANT NEOPLASM OF HEAD OF PANCREAS 
C0153458|T047||CCS_10|PANCREATIC NEOPLASM MALIGNANT HEAD
C0153458|T047||CCS_10|CA HEAD OF PANCREAS 
C0153458|T047||CCS_10|MALIGNANT TUMOUR OF HEAD OF PANCREAS
C0153458|T047||CCS_10|CA HEAD OF PANCREAS
C0153458|T047||CCS_10|MALIGNANT TUMOR OF HEAD OF PANCREAS
C0153458|T047||CCS_10|CANCER OF HEAD OF PANCREAS
C0153458|T047||CCS_10|MALIGNANT TUMOR OF HEAD OF PANCREAS 
C1328479|T047||CCS_10|CARCINOMA, ISLET CELL
C1328479|T047||CCS_10|CARCINOMAS, ISLET CELL
C1328479|T047||CCS_10|ISLET CELL CARCINOMAS
C1328479|T047||CCS_10|ISLET CELL CARCINOMA
C1328479|T047||CCS_10|MALIGNANT NEOPLASM OF ISLETS OF LANGERHANS
C1328479|T047||CCS_10|ISLET CELL CARCINOMA OF PANCREAS
C1328479|T047||CCS_10|ISLET CELL CARCINOMA OF PANCREAS 
C1328479|T047||CCS_10|ISLET CELL CARCINOMA 
C1328479|T047||CCS_10|MAL NEO ISLET LANGERHANS
C1328479|T047||CCS_10|CARCINOMA, ISLET CELL [DISEASE/FINDING]
C1328479|T047||CCS_10|ISLET CELL TUMOR, MALIGNANT
C1328479|T047||CCS_10|HIGH GRADE PANCREATIC NEUROENDOCRINE CARCINOMA
C1328479|T047||CCS_10|POORLY DIFFERENTIATED PANCREATIC ENDOCRINE CARCINOMA
C1328479|T047||CCS_10|PANCREATIC NEC G3
C1328479|T047||CCS_10|HIGH-GRADE PANCREATIC NEUROENDOCRINE CARCINOMA
C1328479|T047||CCS_10|PANCREATIC ENDOCRINE CARCINOMA
C1328479|T047||CCS_10|PANCREATIC NEUROENDOCRINE CARCINOMA
C1328479|T047||CCS_10|PANCREATIC NEC
C1328479|T047||CCS_10|ISLET CELL CANCER
C1328479|T047||CCS_10|CARCINOMA, ISLET CELL, MALIGNANT
C1328479|T047||CCS_10|PANCREATIC ENDOCRINE CANCER
C1328479|T047||CCS_10|PANCREATIC NEOPLASM MALIGNANT CARCINOMA ENDOCRINE PANCREAS
C1328479|T047||CCS_10|CARCINOMA OF ENDOCRINE PANCREAS
C1328479|T047||CCS_10|CARCINOMA OF ENDOCRINE PANCREAS 
C1328479|T047||CCS_10|MALIGNANT NEOPLASM ENDOCRINE GLANDS ISLETS OF LANGERHANS
C1328479|T047||CCS_10|MALIGNANT NEOPLASM OF ISLETS OF LANGERHANS 
C1328479|T047||CCS_10|PANCREATIC ENDOCRINE TUMOR, MALIGNANT
C1328479|T047||CCS_10|PANCREATIC ENDOCRINE TUMOUR, MALIGNANT
C1328479|T047||CCS_10|MALIGNANT ISLET CELL TUMOR
C1328479|T047||CCS_10|MALIGNANT PANCREATIC ENDOCRINE TUMOR
C1328479|T047||CCS_10|PANCREATIC ISLET CELL NEOPLASM MALIGNANT NOS
C1328479|T047||CCS_10|MALIGNANT PANCREATIC ISLET NEOPLASM
C1328479|T047||CCS_10|PANCREATIC ISLET CELL CARCINOMA
C1328479|T047||CCS_10|ISLET CELL ADENOCARCINOMA
C1328479|T047||CCS_10|ENDOCRINE PANCREATIC CARCINOMA
C1328479|T047||CCS_10|MALIGNANT ISLET CELL TUMOUR
C1328479|T047||CCS_10|MALIGNANT TUMOR OF ISLETS OF LANGERHANS
C1328479|T047||CCS_10|MALIGNANT TUMOUR OF ISLETS OF LANGERHANS
C1328479|T047||CCS_10|CARCINOMA OF ENDOCRINE PANCREAS 
C1328479|T047||CCS_10|ISLET CELL CARCINOMA (MORPHOLOGIC ABNORMALITY)
C1328479|T047||CCS_10|MALIGNANT TUMOR OF ISLETS OF LANGERHANS 
C1328479|T047||CCS_10|CANCER OF THE ENDOCRINE PANCREAS
C1328479|T047||CCS_10|CARCINOMA OF THE ENDOCRINE PANCREAS
C1328479|T047||CCS_10|ENDOCRINE PANCREATIC CANCER
C1328479|T047||CCS_10|CARCINOMA; ISLET CELL, PANCREAS
C1328479|T047||CCS_10|CARCINOMA; ISLET CELL, UNSPECIFIED SITE
C1328479|T047||CCS_10|ISLET CELL; CARCINOMA, PANCREAS
C1328479|T047||CCS_10|ISLET CELL; CARCINOMA, UNSPECIFIED SITE
C1328479|T047||CCS_10|PANCREAS; CARCINOMA, ISLET CELL
C1328479|T047||CCS_10|PANCREAS; ISLET CELL CARCINOMA
C1328479|T047||CCS_10|MALIGNANT NEOPLASM OF ISLETS OF LANGERHANS, ANY PART OF PANCREAS
C0496785|T047||CCS_10|MALIGNANT NEOPLASM OF OTHER PARTS OF PANCREAS
C0496785|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF OTHER PARTS OF PANCREAS 
C0496785|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF OTHER PARTS OF PANCREAS
C0153463|T047||CCS_10|MALIGNANT NEOPLASM OF OTHER SPECIFIED SITES OF PANCREAS
C0153463|T047||CCS_10|MALIG NEO PANCREAS NEC
C0153463|T047||CCS_10|MALIGNANT NEOPLASM OF OTHER SPECIFIED SITES OF PANCREAS 
C0153461|T047||CCS_10|MALIGNANT NEOPLASM OF PANCREATIC DUCT
C0153461|T047||CCS_10|MAL NEO PANCREATIC DUCT
C0153461|T047||CCS_10|PANCREATIC NEOPLASM MALIGNANT PANCREATIC DUCT
C0153461|T047||CCS_10|MALIGNANT NEOPLASM OF PANCREATIC DUCT 
C0153461|T047||CCS_10|MALIGNANT TUMOR OF PANCREATIC DUCT
C0153461|T047||CCS_10|MALIGNANT TUMOUR OF PANCREATIC DUCT
C0153461|T047||CCS_10|MALIGNANT TUMOR OF PANCREATIC DUCT 
C0153461|T047||CCS_10|MALIGNANT NEOPLASM OF DUCT OF WIRSUNG
C0496784|T047||CCS_10|MALIGNANT NEOPLASM OF ENDOCRINE PANCREAS
C0496784|T047||CCS_10|MALIGNANT NEOPLASM OF ENDOCRINE PANCREAS 
C0496784|T047||CCS_10|PANCREATIC NEOPLASM MALIGNANT ENDOCRINE PANCREAS
C0496784|T047||CCS_10|MALIGNANT TUMOR OF ENDOCRINE PANCREAS
C0496784|T047||CCS_10|MALIGNANT TUMOUR OF ENDOCRINE PANCREAS
C0496784|T047||CCS_10|MALIGNANT TUMOR OF ENDOCRINE PANCREAS 
C0349053|T047||CCS_10|MALIGNANT NEOPLASM OVERLAPPING PANCREAS SITE
C0349053|T047||CCS_10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF PANCREAS
C0349053|T047||CCS_10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF PANCREAS 
C0349053|T047||CCS_10|PANCREATIC NEOPLASM MALIGNANT OVERLAPPING SITES
C0349053|T047||CCS_10|MALIGNANT NEOPLASM, OVERLAPPING LESION OF PANCREAS
C0349053|T047||CCS_10|MALIGNANT NEOPLASM, OVERLAPPING LESION OF PANCREAS 
C0349053|T047||CCS_10|CANCER OF THE PANCREAS, OVERLAPPING SITES
C0349053|T047||CCS_10|OVERLAPPING MALIGNANT NEOPLASM OF PANCREAS 
C0349053|T047||CCS_10|OVERLAPPING MALIGNANT NEOPLASM OF PANCREAS
C0346647|T047||CCS_10|MALIGNANT NEOPLASM OF PANCREAS
C0346647|T047||CCS_10|PANCREATIC CANCER
C0346647|T047||CCS_10|MALIGNANT NEOPLASM OF PANCREAS, UNSPECIFIED
C0346647|T047||CCS_10|PANCREAS, UNSPECIFIED
C0346647|T047||CCS_10|MALIGNANT NEOPLASM OF PANCREAS 
C0346647|T047||CCS_10|MALIGNANT PANCREATIC NEOPLASM
C0346647|T047||CCS_10|CANCERS, PANCREAS
C0346647|T047||CCS_10|PANCREAS CANCERS
C0346647|T047||CCS_10|CANCER, PANCREATIC
C0346647|T047||CCS_10|CANCERS, PANCREATIC
C0346647|T047||CCS_10|PANCREATIC CANCERS
C0346647|T047||CCS_10|MALIGNANT TUMOR OF PANCREAS
C0346647|T047||CCS_10|MALIG NEO PANCREAS NOS
C0346647|T047||CCS_10|CANCER OF PANCREAS
C0346647|T047||CCS_10|CANCER, PANCREAS
C0346647|T047||CCS_10|CA PANCREAS NOS 
C0346647|T047||CCS_10|CA PANCREAS NOS
C0346647|T047||CCS_10|CA - CANCER OF PANCREAS
C0346647|T047||CCS_10|CA - PANCREATIC CANCER
C0346647|T047||CCS_10|MALIGNANT TUMOUR OF PANCREAS
C0346647|T047||CCS_10|MALIGNANT NEOPLASM OF PANCREAS NOS
C0346647|T047||CCS_10|MALIGNANT NEOPLASM OF PANCREAS NOS 
C0346647|T047||CCS_10|PANCREAS--CANCER
C0346647|T047||CCS_10|PANCREAS CANCER
C0346647|T047||CCS_10|NEOPLASM OF THE PANCREAS
C0346647|T047||CCS_10|CANCER OF THE PANCREAS
C0346647|T047||CCS_10|NEOPLASIA OF THE PANCREAS
C0346647|T047||CCS_10|PANCREAS NEOPLASM MALIGNANT
C0346647|T047||CCS_10|MALIGNANT NEOPLASM OF PANCREAS, PART UNSPECIFIED
C0346647|T047||CCS_10|MALIGNANT TUMOR OF PANCREAS 
C0346647|T047||CCS_10|MALIGNANT NEOPLASM OF PANCREAS, NOS
C0346647|T047||CCS_10|MALIGNANT NEOPLASM OF THE PANCREAS
C0346647|T047||CCS_10|NEOPLASM MALIG;PANCREAS
C0346647|T047||CCS_10|MALIGNANT NEOSPLASM OF THE PANCREAS
C2007079|T047||CCS_10|CARCINOSARCOMA OF PANCREAS 
C2007079|T047||CCS_10|CARCINOSARCOMA OF PANCREAS
C0235974|T047||CCS_10|PANCREATIC CARCINOMA
C0235974|T047||CCS_10|CARCINOMA OF PANCREAS 
C0235974|T047||CCS_10|CARCINOMA OF PANCREAS
C0235974|T047||CCS_10|CARCINOMA;PANCREAS
C0235974|T047||CCS_10|PANCREATIC CANCER
C0235974|T047||CCS_10|PANCREATIC ACINAR CARCINOMA
C0235974|T047||CCS_10|CARCINOMA OF PANCREAS 
C0235974|T047||CCS_10|EXOCRINE CANCER
C0235974|T047||CCS_10|PANCREATIC CANCER (NOT ISLETS)
C0235974|T047||CCS_10|PANCREATIC CANCER (EXCLUDING ISLETS), NOS
C0235974|T047||CCS_10|PANCREATIC CARCINOMA NOS
C0235974|T047||CCS_10|PANCREAS CARCINOMA
C0235974|T047||CCS_10|CANCER OF PANCREAS
C0235974|T047||CCS_10|CANCER OF THE PANCREAS
C0235974|T047||CCS_10|PANCREAS CANCER
C0235974|T047||CCS_10|EXOCRINE PANCREAS CARCINOMA
C0235974|T047||CCS_10|CARCINOMA OF THE PANCREAS
C2205484|T047||CCS_10|MALIGNANT SMALL CELL NEOPLASM OF PANCREAS 
C2205484|T047||CCS_10|PANCREATIC NEOPLASM MALIGNANT SMALL CELL TYPE
C2205484|T047||CCS_10|MALIGNANT SMALL CELL NEOPLASM OF PANCREAS
C2011344|T047||CCS_10|GIANT CELL TYPE NEOPLASM OF PANCREAS
C2011344|T047||CCS_10|GIANT CELL TYPE NEOPLASM OF PANCREAS 
C2018676|T047||CCS_10|SPINDLE CELL TYPE NEOPLASM OF PANCREAS 
C2018676|T047||CCS_10|SPINDLE CELL TYPE NEOPLASM OF PANCREAS
C2018676|T047||CCS_10|PANCREATIC NEOPLASM MALIGNANT SPINDLE CELL TYPE
C2075636|T047||CCS_10|CLEAR CELL TYPE NEOPLASM OF PANCREAS
C2075636|T047||CCS_10|PANCREATIC NEOPLASM MALIGNANT CLEAR CELL TYPE
C2075636|T047||CCS_10|CLEAR CELL TYPE NEOPLASM OF PANCREAS 
C3536762|T047||CCS_10|MALIGNANT CARCINOID TUMOR OF PANCREAS
C3536762|T047||CCS_10|MALIGNANT CARCINOID TUMOR OF PANCREAS 
C3536762|T047||CCS_10|MALIGNANT CARCINOID TUMOR OF PANCREAS 
C3536762|T047||CCS_10|MALIGNANT CARCINOID TUMOUR OF PANCREAS
C1096346|T047||CCS_10|SARCOMA OF PANCREAS 
C1096346|T047||CCS_10|SARCOMA OF PANCREAS
C1096346|T047||CCS_10|PANCREATIC SARCOMA
C1096346|T047||CCS_10|SARCOMA OF THE PANCREAS
C2205511|T047||CCS_10|MYOSARCOMA OF PANCREAS 
C2205511|T047||CCS_10|MYOSARCOMA OF PANCREAS
C2205516|T047||CCS_10|MALIGNANT LYMPHOMA OF PANCREAS 
C2205516|T047||CCS_10|MALIGNANT LYMPHOMA OF PANCREAS
C2205519|T047||CCS_10|MALIGNANT PLASMACYTOMA OF PANCREAS
C2205519|T047||CCS_10|MALIGNANT PLASMACYTOMA OF PANCREAS 
C2205521|T047||CCS_10|MALIGNANT MASTOCYTOSIS OF PANCREAS 
C2205521|T047||CCS_10|MALIGNANT MASTOCYTOSIS OF PANCREAS
C0281361|T047||CCS_10|PANCREATIC ADENOCARCINOMA
C0281361|T047||CCS_10|ADENOCARCINOMA OF PANCREAS
C0281361|T047||CCS_10|ADENOCARCINOMA OF PANCREAS 
C0281361|T047||CCS_10|ADENOCARCINOMA PANCREAS
C0281361|T047||CCS_10|ADENOCARCINOMA OF PANCREAS 
C0281361|T047||CCS_10|ADENOCARCINOMA - PANCREAS
C0281361|T047||CCS_10|ADENOCARCINOMA OF THE PANCREAS
C0281361|T047||CCS_10|PANCREAS ADENOCARCINOMA
C2062546|T047||CCS_10|MICROADENOMATOSIS OF PANCREAS 
C2062546|T047||CCS_10|MICROADENOMATOSIS OF PANCREAS
C2062546|T047||CCS_10|PANCREATIC MICROADENOMATOSIS
C0086768|T047||CCS_10|CHOLERA, PANCREATIC
C0086768|T047||CCS_10|VERNER MORRISON SYNDROME
C0086768|T047||CCS_10|SYNDROME, VERNER-MORRISON
C0086768|T047||CCS_10|VERNER-MORRISON SYNDROME DUE TO PANCREATIC NEOPLASM
C0086768|T047||CCS_10|VERNER-MORRISON SYNDROME DUE TO PANCREATIC NEOPLASM 
C0086768|T047||CCS_10|PANCREATIC CHOLERA (WDHA SYNDROME)
C0086768|T047||CCS_10|WDHA SYNDROMES
C0086768|T047||CCS_10|EXCESSIVE VASOACTIVE INTESTINAL PEPTIDE SECRETION 
C0086768|T047||CCS_10|EXCESSIVE VASOACTIVE INTESTINAL PEPTIDE SECRETION
C0086768|T047||CCS_10|VERNER-MORRISON SYNDROME
C0086768|T047||CCS_10|VIPOMA SYNDROME
C0086768|T047||CCS_10|WATERY DIARRHEA SYNDROME
C0086768|T047||CCS_10|WDHH
C0086768|T047||CCS_10|WATERY DIARRHEA, HYPOKALEMIA, AND ACHLORHYDRIA SYNDROME
C0086768|T047||CCS_10|WATERY DIARRHEA WITH HYPOKALEMIC ALKALOSIS
C0086768|T047||CCS_10|WDHA
C0086768|T047||CCS_10|WDHA SYNDROME
C0086768|T047||CCS_10|SYNDROME, VIPOMA
C0086768|T047||CCS_10|PSEUDOPANCREATIC CHOLERA SYNDROME
C0086768|T047||CCS_10|PANCREATIC CHOLERA
C0086768|T047||CCS_10|WERNER MORRISON SYNDROME
C0086768|T047||CCS_10|PSEUDOPANCREATIC CHOLERA SYNDROME 
C0086768|T047||CCS_10|VERNER-MORRISON SYNDROME 
C0086768|T047||CCS_10|ISLET CELL WDHA SYNDROME
C0086768|T047||CCS_10|PANCREATIC WDHA SYNDROME
C0086768|T047||CCS_10|EXCESSIVE VASOACTIVE INTESTINAL PEPTIDE SECRETION [AMBIGUOUS]
C1389637|T047||CCS_10|MALIGNANT BETA CELL TUMOR OF PANCREAS 
C1389637|T047||CCS_10|MALIGNANT BETA CELL TUMOR OF PANCREAS
C1389637|T047||CCS_10|MALIGNANT INSULINOMA OF PANCREAS
C1389637|T047||CCS_10|MALIGNANT PANCREATIC BETA CELL TUMOR
C1389637|T047||CCS_10|MALIGNANT INSULINOMA OF PANCREAS 
C1389637|T047||CCS_10|BETA-CELL; TUMOR, MALIGNANT, PANCREAS
C1389637|T047||CCS_10|INSULINOMA; MALIGNANT, PANCREAS
C1389637|T047||CCS_10|MALIGNANT; INSULINOMA, PANCREAS
C1389637|T047||CCS_10|PANCREAS; BETA-CELL TUMOR, MALIGNANT
C1389637|T047||CCS_10|PANCREAS; INSULINOMA, MALIGNANT
C1389637|T047||CCS_10|PANCREAS; MALIGNANT INSULINOMA
C1389637|T047||CCS_10|PANCREAS; TUMOR, BETA-CELL, MALIGNANT
C1389637|T047||CCS_10|TUMOR; BETA-CELL, MALIGNANT, PANCREAS
C1335315|T047||CCS_10|SEROUS CYSTADENOCARCINOMA OF PANCREAS
C1335315|T047||CCS_10|SEROUS CYSTADENOCARCINOMA OF PANCREAS 
C1335315|T047||CCS_10|PANCREATIC SEROUS CYSTADENOCARCINOMA
C1335315|T047||CCS_10|SEROUS CYSTADENOCARCINOMA OF THE PANCREAS
C2063876|T047||CCS_10|INVASIVE MUCINOUS CYSTADENOCARCINOMA OF PANCREAS 
C2063876|T047||CCS_10|INVASIVE MUCINOUS CYSTADENOCARCINOMA OF PANCREAS
C1335304|T047||CCS_10|INTRADUCTAL PAPILLARY-MUCINOUS CARCINOMA OF PANCREAS 
C1335304|T047||CCS_10|INTRADUCTAL PAPILLARY-MUCINOUS CARCINOMA OF PANCREAS
C1335304|T047||CCS_10|PANCREATIC INTRADUCTAL PAPILLARY-COLLOID CARCINOMA
C1335304|T047||CCS_10|PANCREATIC INTRADUCTAL PAPILLARY-COLLOIDAL CARCINOMA
C1335304|T047||CCS_10|INTRADUCTAL PAPILLARY-COLLOIDAL CARCINOMA OF THE PANCREAS
C1335304|T047||CCS_10|INTRADUCTAL PAPILLARY-MUCINOUS CARCINOMA OF THE PANCREAS
C1335304|T047||CCS_10|INTRADUCTAL PAPILLARY-COLLOID CARCINOMA OF PANCREAS
C1335304|T047||CCS_10|INTRADUCTAL PAPILLARY-COLLOID CARCINOMA OF THE PANCREAS
C1335304|T047||CCS_10|INTRADUCTAL PAPILLARY-COLLOIDAL CARCINOMA OF PANCREAS
C1335304|T047||CCS_10|PANCREATIC INTRADUCTAL PAPILLARY-MUCINOUS CARCINOMA
C2063878|T047||CCS_10|MIXED ACINAR-ENDOCRINE CARCINOMA OF PANCREAS 
C2063878|T047||CCS_10|MIXED ACINAR-ENDOCRINE CARCINOMA OF PANCREAS
C2063878|T047||CCS_10|MUCINOUS CARCINOID TUMOR OF THE PANCREAS
C2063878|T047||CCS_10|MIXED CARCINOID-ADENOCARCINOMA OF THE PANCREAS
C2063878|T047||CCS_10|MIXED ACINAR-ENDOCRINE CARCINOMA OF THE PANCREAS
C2063878|T047||CCS_10|MIXED ACINAR-NEUROENDOCRINE CARCINOMA OF THE PANCREAS
C2063878|T047||CCS_10|ACINAR-ISLET CELL TUMOR, MALIGNANT
C0334489|T047||CCS_10|PANCREATOBLASTOMA 
C0334489|T047||CCS_10|PANCREATOBLASTOMA
C0334489|T047||CCS_10|PANCREATOBLASTOMA 
C0334489|T047||CCS_10|[M]PANCREATOBLASTOMA
C0334489|T047||CCS_10|[M] PANCREATOBLASTOMA
C0334489|T047||CCS_10|PANCREATOBLASTOMA (MORPHOLOGIC ABNORMALITY)
C2205494|T047||CCS_10|SCIRRHOUS ADENOCARCINOMA OF PANCREAS 
C2205494|T047||CCS_10|SCIRRHOUS ADENOCARCINOMA OF PANCREAS
C2205494|T047||CCS_10|PANCREATIC NEOPLASM ADENOCARCINOMA SCIRRHOUS
C2037343|T047||CCS_10|PANCREATIC NEOPLASM ADENOCARCINOMA SUPERFICIAL SPREADING
C2037343|T047||CCS_10|SUPERFICIAL SPREADING ADENOCARCINOMA OF PANCREAS 
C2037343|T047||CCS_10|SUPERFICIAL SPREADING ADENOCARCINOMA OF PANCREAS
C2205495|T047||CCS_10|BASAL CELL ADENOCARCINOMA OF PANCREAS 
C2205495|T047||CCS_10|BASAL CELL ADENOCARCINOMA OF PANCREAS
C2033127|T047||CCS_10|PAPILLARY ADENOCARCINOMA OF PANCREAS 
C2033127|T047||CCS_10|PAPILLARY ADENOCARCINOMA OF PANCREAS
C2189643|T047||CCS_10|VILLOUS ADENOCARCINOMA OF PANCREAS 
C2189643|T047||CCS_10|VILLOUS ADENOCARCINOMA OF PANCREAS
C2205497|T047||CCS_10|ADENOCARCINOMA IN TUBULOVILLOUS ADENOMA OF PANCREAS
C2205497|T047||CCS_10|ADENOCARCINOMA IN TUBULOVILLOUS ADENOMA OF PANCREAS 
C2205498|T047||CCS_10|ADENOCARCINOMA IN ADENOMATOUS POLYP OF PANCREAS 
C2205498|T047||CCS_10|ADENOCARCINOMA IN ADENOMATOUS POLYP OF PANCREAS
C2205499|T047||CCS_10|MUCIN-PRODUCING ADENOCARCINOMA OF PANCREAS 
C2205499|T047||CCS_10|MUCIN-PRODUCING ADENOCARCINOMA OF PANCREAS
C2033012|T047||CCS_10|INTRADUCTAL PAPILLARY ADENOCARCINOMA OF PANCREAS WITH INVASION
C2033012|T047||CCS_10|INTRADUCTAL PAPILLARY ADENOCARCINOMA OF PANCREAS WITH INVASION 
C2205500|T047||CCS_10|ADENOCARCINOMA OF PANCREAS WITH METAPLASIA 
C2205500|T047||CCS_10|PANCREATIC ADENOCARCINOMA WITH METAPLASIA
C2205500|T047||CCS_10|ADENOCARCINOMA OF PANCREAS WITH METAPLASIA
C2205501|T047||CCS_10|ADENOCARCINOMA OF PANCREAS WITH SQUAMOUS METAPLASIA 
C2205501|T047||CCS_10|ADENOCARCINOMA OF PANCREAS WITH SQUAMOUS METAPLASIA
C2205501|T047||CCS_10|PANCREATIC ADENOCARCINOMA WITH SQUAMOUS METAPLASIA
C2033013|T047||CCS_10|ADENOCARCINOMA WITH CARTILAGINOUS OR OSSEOUS METAPLASIA OF PANCREAS
C2033013|T047||CCS_10|ADENOCARCINOMA OF PANCREAS WITH CARTILAGINOUS AND OSSEOUS METAPLASIA
C2033013|T047||CCS_10|ADENOCARCINOMA OF PANCREAS WITH CARTILAGINOUS AND OSSEOUS METAPLASIA 
C2033013|T047||CCS_10|PANCREATIC ADENOCARCINOMA WITH CARTILAGINOUS OR OSSEOUS METAPLASIA
C2033013|T047||CCS_10|PANCREATIC ADENOCARCINOMA WITH CARTILAGINOUS AND OSSEOUS METAPLASIA
C2205502|T047||CCS_10|PANCREATIC ADENOCARCINOMA METAPLASTIC SPINDLE CELL
C2205502|T047||CCS_10|PANCREATIC ADENOCARCINOMA WITH SPINDLE CELL METAPLASIA
C2205502|T047||CCS_10|ADENOCARCINOMA OF PANCREAS WITH SPINDLE CELL METAPLASIA 
C2205502|T047||CCS_10|ADENOCARCINOMA OF PANCREAS WITH SPINDLE CELL METAPLASIA
C2205503|T047||CCS_10|PANCREATIC ADENOCARCINOMA WITH APOCRINE METAPLASIA
C2205503|T047||CCS_10|ADENOCARCINOMA OF PANCREAS WITH APOCRINE METAPLASIA 
C2205503|T047||CCS_10|ADENOCARCINOMA OF PANCREAS WITH APOCRINE METAPLASIA
C2033014|T047||CCS_10|ADENOCARCINOMA OF PANCREAS WITH NEUROENDOCRINE DIFFERENTIATION 
C2033014|T047||CCS_10|ADENOCARCINOMA OF PANCREAS WITH NEUROENDOCRINE DIFFERENTIATION
C2033014|T047||CCS_10|PANCREATIC ADENOCARCINOMA WITH NEUROENDOCRINE DIFFERENTIATION
C2030694|T047||CCS_10|HEPATOID ADENOCARCINOMA OF PANCREAS
C2030694|T047||CCS_10|HEPATOID ADENOCARCINOMA OF PANCREAS 
C2170821|T047||CCS_10|TUBULAR ADENOCARCINOMA OF PANCREAS 
C2170821|T047||CCS_10|TUBULAR ADENOCARCINOMA OF PANCREAS
C2075534|T047||CCS_10|CLEAR CELL ADENOCARCINOMA OF PANCREAS
C2075534|T047||CCS_10|CLEAR CELL ADENOCARCINOMA OF PANCREAS 
C2063871|T047||CCS_10|MUCINOUS ADENOCARCINOMA OF PANCREAS
C2063871|T047||CCS_10|MUCINOUS ADENOCARCINOMA OF PANCREAS 
C2033034|T047||CCS_10|NONINVASIVE INTRADUCTAL PAPILLARY-MUCINOUS CARCINOMA OF PANCREAS 
C2033034|T047||CCS_10|NONINVASIVE INTRADUCTAL PAPILLARY-MUCINOUS CARCINOMA OF PANCREAS
C1518871|T047||CCS_10|INTRADUCTAL PAPILLARY-MUCINOUS CARCINOMA OF THE PANCREAS INVASIVE
C1518871|T047||CCS_10|INVASIVE INTRADUCTAL PAPILLARY-MUCINOUS CARCINOMA OF PANCREAS
C1518871|T047||CCS_10|INTRADUCTAL PAPILLARY-MUCINOUS CARCINOMA OF THE PANCREAS INVASIVE 
C1518871|T047||CCS_10|PANCREATIC INTRADUCTAL PAPILLARY-MUCINOUS NEOPLASM WITH AN ASSOCIATED INVASIVE CARCINOMA
C1518871|T047||CCS_10|PANCREATIC INVASIVE INTRADUCTAL PAPILLARY-MUCINOUS CARCINOMA
C1518871|T047||CCS_10|PANCREATIC INTRADUCTAL PAPILLARY MUCINOUS NEOPLASM WITH AN ASSOCIATED INVASIVE CARCINOMA
C1336861|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF PANCREAS 
C1336861|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF PANCREAS
C1336861|T047||CCS_10|PANCREATIC CARCINOSARCOMA
C1336861|T047||CCS_10|PLEOMORPHIC LARGE CELL PANCREATIC CARCINOMA
C1336861|T047||CCS_10|SARCOMATOID PANCREATIC CARCINOMA
C1336861|T047||CCS_10|UNDIFFERENTIATED (ANAPLASTIC) PANCREATIC CARCINOMA
C1336861|T047||CCS_10|SPINDLE CELL PANCREATIC CARCINOMA
C1336861|T047||CCS_10|UNDIFFERENTIATED PANCREATIC CARCINOMA
C1336861|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF THE PANCREAS
C2033249|T047||CCS_10|PAPILLARY CYSTADENOCARCINOMA OF PANCREAS 
C2033249|T047||CCS_10|PAPILLARY CYSTADENOCARCINOMA OF PANCREAS
C2033261|T047||CCS_10|PAPILLARY MUCINOUS CYSTADENOCARCINOMA OF PANCREAS 
C2033261|T047||CCS_10|PAPILLARY MUCINOUS CYSTADENOCARCINOMA OF PANCREAS
C2106547|T047||CCS_10|COMEDOCARCINOMA OF PANCREAS
C2106547|T047||CCS_10|COMEDOCARCINOMA OF PANCREAS 
C2205496|T047||CCS_10|ADENOCARCINOMA IN VILLOUS ADENOMA OF PANCREAS
C2205496|T047||CCS_10|ADENOCARCINOMA IN VILLOUS ADENOMA OF PANCREAS 
C2018503|T047||CCS_10|SPINDLE CELL SARCOMA OF PANCREAS
C2018503|T047||CCS_10|SPINDLE CELL SARCOMA OF PANCREAS 
C2011317|T047||CCS_10|GIANT CELL SARCOMA OF PANCREAS
C2011317|T047||CCS_10|GIANT CELL SARCOMA OF PANCREAS 
C2205507|T047||CCS_10|SMALL CELL SARCOMA OF PANCREAS 
C2205507|T047||CCS_10|SMALL CELL SARCOMA OF PANCREAS
C2205508|T047||CCS_10|EPITHELIOID SARCOMA OF PANCREAS 
C2205508|T047||CCS_10|EPITHELIOID SARCOMA OF PANCREAS
C2188140|T047||CCS_10|UNDIFFERENTIATED SARCOMA OF PANCREAS
C2188140|T047||CCS_10|UNDIFFERENTIATED SARCOMA OF PANCREAS 
C2182952|T047||CCS_10|DESMOPLASTIC SMALL ROUND CELL SARCOMA OF PANCREAS
C2182952|T047||CCS_10|DESMOPLASTIC SMALL ROUND CELL SARCOMA OF PANCREAS 
C2046335|T047||CCS_10|HISTIOCYTIC SARCOMA OF PANCREAS
C2046335|T047||CCS_10|HISTIOCYTIC SARCOMA OF PANCREAS 
C2111172|T047||CCS_10|LANGERHANS CELL SARCOMA OF PANCREAS 
C2111172|T047||CCS_10|LANGERHANS CELL SARCOMA OF PANCREAS
C2077758|T047||CCS_10|INTERDIGITATING DENDRITIC CELL SARCOMA OF PANCREAS
C2077758|T047||CCS_10|INTERDIGITATING DENDRITIC CELL SARCOMA OF PANCREAS 
C2205510|T047||CCS_10|FOLLICULAR DENDRITIC CELL SARCOMA OF PANCREAS
C2205510|T047||CCS_10|FOLLICULAR DENDRITIC CELL SARCOMA OF PANCREAS 
C2205513|T047||CCS_10|ANGIOMYOSARCOMA OF PANCREAS 
C2205513|T047||CCS_10|ANGIOMYOSARCOMA OF PANCREAS
C1409081|T047||CCS_10|MIXED ISLET CELL AND EXOCRINE ADENOCARCINOMA OF PANCREAS 
C1409081|T047||CCS_10|MIXED ISLET CELL AND EXOCRINE ADENOCARCINOMA OF PANCREAS
C1409081|T047||CCS_10|PANCREAS; ADENOCARCINOMA ISLET CELL, WITH EXOCRINE MIXED
C2033018|T047||CCS_10|NONINFILTRATING INTRADUCTAL CARCINOMA OF PANCREAS 
C2033018|T047||CCS_10|NONINFILTRATING INTRADUCTAL CARCINOMA OF PANCREAS
C2033017|T047||CCS_10|NONINFILTRATING INTRACYSTIC CARCINOMA OF PANCREAS 
C2033017|T047||CCS_10|NONINFILTRATING INTRACYSTIC CARCINOMA OF PANCREAS
C2033016|T047||CCS_10|INTRADUCTAL MICROPAPILLARY CARCINOMA OF PANCREAS 
C2033016|T047||CCS_10|INTRADUCTAL MICROPAPILLARY CARCINOMA OF PANCREAS
C2205485|T047||CCS_10|MALIGNANT EPITHELIOMA OF PANCREAS 
C2205485|T047||CCS_10|MALIGNANT EPITHELIOMA OF PANCREAS
C2111650|T047||CCS_10|LARGE CELL CARCINOMA OF PANCREAS
C2111650|T047||CCS_10|LARGE CELL CARCINOMA OF PANCREAS 
C2111737|T047||CCS_10|LARGE CELL NEUROENDOCRINE CARCINOMA OF PANCREAS 
C2111737|T047||CCS_10|LARGE CELL NEUROENDOCRINE CARCINOMA OF PANCREAS
C2111651|T047||CCS_10|PANCREATIC NEOPLASM CARCINOMA LARGE CELL WITH RHABDOID PHENOTYPE
C2111651|T047||CCS_10|LARGE CELL CARCINOMA OF PANCREAS WITH RHABDOID PHENOTYPE 
C2111651|T047||CCS_10|LARGE CELL CARCINOMA OF PANCREAS WITH RHABDOID PHENOTYPE
C2012101|T047||CCS_10|GLASSY CELL CARCINOMA OF PANCREAS
C2012101|T047||CCS_10|GLASSY CELL CARCINOMA OF PANCREAS 
C2082450|T047||CCS_10|PLEOMORPHIC CARCINOMA OF PANCREAS 
C2082450|T047||CCS_10|PLEOMORPHIC CARCINOMA OF PANCREAS
C2011260|T047||CCS_10|GIANT CELL CARCINOMA OF PANCREAS
C2011260|T047||CCS_10|GIANT CELL CARCINOMA OF PANCREAS 
C2018400|T047||CCS_10|SPINDLE CELL CARCINOMA OF PANCREAS
C2018400|T047||CCS_10|SPINDLE CELL CARCINOMA OF PANCREAS 
C2011225|T047||CCS_10|GIANT CELL AND SPINDLE CELL CARCINOMA OF PANCREAS
C2011225|T047||CCS_10|GIANT CELL AND SPINDLE CELL CARCINOMA OF PANCREAS 
C2142930|T047||CCS_10|PSEUDOSARCOMATOUS CARCINOMA OF PANCREAS
C2142930|T047||CCS_10|PSEUDOSARCOMATOUS CARCINOMA OF PANCREAS 
C2111812|T047||CCS_10|POLYGONAL CELL CARCINOMA OF PANCREAS
C2111812|T047||CCS_10|POLYGONAL CELL CARCINOMA OF PANCREAS 
C2205486|T047||CCS_10|SMALL CELL CARCINOMA OF PANCREAS
C2205486|T047||CCS_10|SMALL CELL CARCINOMA OF PANCREAS 
C2009884|T047||CCS_10|FUSIFORM TYPE SMALL CELL CARCINOMA OF PANCREAS 
C2009884|T047||CCS_10|FUSIFORM TYPE SMALL CELL CARCINOMA OF PANCREAS
C2033227|T047||CCS_10|PAPILLARY CARCINOMA OF PANCREAS
C2033227|T047||CCS_10|PAPILLARY CARCINOMA OF PANCREAS 
C2033304|T047||CCS_10|PAPILLARY SQUAMOUS CELL CARCINOMA OF PANCREAS
C2033304|T047||CCS_10|PAPILLARY SQUAMOUS CELL CARCINOMA OF PANCREAS 
C2189356|T047||CCS_10|VERRUCOUS CARCINOMA OF PANCREAS
C2189356|T047||CCS_10|VERRUCOUS CARCINOMA OF PANCREAS 
C2675993|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF PANCREAS 
C2675993|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF PANCREAS
C2675993|T047||CCS_10|PANCREATIC SQUAMOUS CELL CARCINOMA
C2675993|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE PANCREAS
C2109314|T047||CCS_10|KERATINIZING SQUAMOUS CELL CARCINOMA OF PANCREAS
C2109314|T047||CCS_10|KERATINIZING SQUAMOUS CELL CARCINOMA OF PANCREAS 
C2205487|T047||CCS_10|PANCREATIC CARCINOMA SQUAMOUS CELL LARGE CELL NONKERATINIZING
C2205487|T047||CCS_10|NONKERATINIZING LARGE CELL SQUAMOUS CARCINOMA CELL OF PANCREAS
C2205487|T047||CCS_10|NONKERATINIZING LARGE CELL SQUAMOUS CARCINOMA CELL OF PANCREAS 
C2205488|T047||CCS_10|NONKERATINIZING SMALL CELL SQUAMOUS CELL CARCINOMA OF PANCREAS 
C2205488|T047||CCS_10|NONKERATINIZING SMALL CELL SQUAMOUS CELL CARCINOMA OF PANCREAS
C2018561|T047||CCS_10|SPINDLE CELL SQUAMOUS CELL CARCINOMA OF PANCREAS 
C2018561|T047||CCS_10|SPINDLE CELL SQUAMOUS CELL CARCINOMA OF PANCREAS
C2205489|T047||CCS_10|ADENOID SQUAMOUS CELL CARCINOMA OF PANCREAS 
C2205489|T047||CCS_10|ADENOID SQUAMOUS CELL CARCINOMA OF PANCREAS
C2205490|T047||CCS_10|MICROINVASIVE SQUAMOUS CELL CARCINOMA OF PANCREAS
C2205490|T047||CCS_10|MICROINVASIVE SQUAMOUS CELL CARCINOMA OF PANCREAS 
C2019489|T047||CCS_10|PANCREATIC NEOPLASM CARCINOMA SQUAMOUS CELL WITH HORN FORMATION
C2019489|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF PANCREAS WITH HORN FORMATION
C2019489|T047||CCS_10|SQUAMOUS CELL CARCINOMA WITH HORN FORMATION OF PANCREAS
C2019489|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF PANCREAS WITH HORN FORMATION 
C2017452|T047||CCS_10|SOLID CARCINOMA OF PANCREAS
C2017452|T047||CCS_10|SOLID CARCINOMA OF PANCREAS 
C2007049|T047||CCS_10|CARCINOMA SIMPLEX OF PANCREAS 
C2007049|T047||CCS_10|CARCINOMA SIMPLEX OF PANCREAS
C2205491|T047||CCS_10|MUCOEPIDERMOID CARCINOMA OF PANCREAS 
C2205491|T047||CCS_10|MUCOEPIDERMOID CARCINOMA OF PANCREAS
C2076527|T047||CCS_10|INFILTRATING DUCTAL CARCINOMA OF PANCREAS
C2076527|T047||CCS_10|INFILTRATING DUCTAL CARCINOMA OF PANCREAS 
C2078054|T047||CCS_10|INTRACYSTIC CARCINOMA OF PANCREAS
C2078054|T047||CCS_10|INTRACYSTIC CARCINOMA OF PANCREAS 
C2047536|T047||CCS_10|HYPERSECRETORY CYSTIC CARCINOMA OF PANCREAS
C2047536|T047||CCS_10|HYPERSECRETORY CYSTIC CARCINOMA OF PANCREAS 
C2205492|T047||CCS_10|MEDULLARY CARCINOMA OF PANCREAS 
C2205492|T047||CCS_10|MEDULLARY CARCINOMA OF PANCREAS
C2182972|T047||CCS_10|DUCT CARCINOMA, DESMOPLASTIC TYPE, OF PANCREAS
C2182972|T047||CCS_10|DUCT CARCINOMA, DESMOPLASTIC TYPE, OF PANCREAS 
C2076531|T047||CCS_10|INFILTRATING DUCTULAR CARCINOMA OF PANCREAS 
C2076531|T047||CCS_10|INFILTRATING DUCTULAR CARCINOMA OF PANCREAS
C2205493|T047||CCS_10|EPITHELIAL-MYOEPITHELIAL CARCINOMA OF PANCREAS 
C2205493|T047||CCS_10|EPITHELIAL-MYOEPITHELIAL CARCINOMA OF PANCREAS
C2205506|T047||CCS_10|NEUROENDOCRINE CARCINOMA OF PANCREAS
C2205506|T047||CCS_10|NEUROENDOCRINE CARCINOMA OF PANCREAS 
C2205514|T047||CCS_10|EMBRYONAL CARCINOSARCOMA OF PANCREAS 
C2205514|T047||CCS_10|EMBRYONAL CARCINOSARCOMA OF PANCREAS
C1335317|T047||CCS_10|SIGNET RING CELL CARCINOMA OF PANCREAS
C1335317|T047||CCS_10|SIGNET RING CELL CARCINOMA OF PANCREAS 
C1335317|T047||CCS_10|PANCREATIC SIGNET RING CELL CARCINOMA
C1335317|T047||CCS_10|SIGNET RING CELL CARCINOMA OF THE PANCREAS
C1335299|T047||CCS_10|ADENOSQUAMOUS CARCINOMA OF PANCREAS
C1335299|T047||CCS_10|ADENOSQUAMOUS CARCINOMA OF PANCREAS 
C1335299|T047||CCS_10|PANCREATIC ADENOACANTHOMA
C1335299|T047||CCS_10|PANCREATIC MUCOEPIDERMOID CARCINOMA
C1335299|T047||CCS_10|PANCREATIC MIXED SQUAMOUS AND ADENOCARCINOMA
C1335299|T047||CCS_10|ADENOSQUAMOUS CARCINOMA OF THE PANCREAS
C1335299|T047||CCS_10|PANCREATIC ADENOSQUAMOUS CARCINOMA
C2063872|T047||CCS_10|ANAPLASTIC CARCINOMA OF PANCREAS
C2063872|T047||CCS_10|ANAPLASTIC CARCINOMA OF PANCREAS 
C2007059|T047||CCS_10|CARCINOMA OF PANCREAS WITH OSTEOCLAST-LIKE GIANT CELLS
C2007059|T047||CCS_10|CARCINOMA OF PANCREAS WITH OSTEOCLAST-LIKE GIANT CELLS 
C2007059|T047||CCS_10|PANCREATIC CARCINOMA WITH OSTEOCLAST-LIKE GIANT CELLS
C2007059|T047||CCS_10|PANCREATIC OSTEOCLAST-LIKE GIANT CELL CARCINOMA
C2007059|T047||CCS_10|UNDIFFERENTIATED PANCREATIC CARCINOMA WITH OSTEOCLAST-LIKE GIANT CELLS
C2007059|T047||CCS_10|OSTEOCLAST-LIKE GIANT CELL NEOPLASM OF PANCREAS
C2007059|T047||CCS_10|OSTEOCLAST-LIKE GIANT CELL NEOPLASM OF THE PANCREAS
C0279661|T047||CCS_10|ACINAR CELL CARCINOMA OF PANCREAS
C0279661|T047||CCS_10|ACINAR CELL CARCINOMA OF PANCREAS 
C0279661|T047||CCS_10|ACINAR CELL ADENOCARCINOMA OF THE PANCREAS
C0279661|T047||CCS_10|ADENOCARCINOMA, ACINAR CELL, PANCREATIC
C0279661|T047||CCS_10|PANCREAS CANCER, ACINAR CELL ADENOCARCINOMA
C0279661|T047||CCS_10|PANCREATIC CANCER, ACINAR CELL ADENOCARCINOMA
C0279661|T047||CCS_10|ACINAR CELL ADENOCARCINOMA OF PANCREAS
C0279661|T047||CCS_10|ACINAR CELL CARCINOMA OF THE PANCREAS
C0279661|T047||CCS_10|PANCREAS ACINAR CELL ADENOCARCINOMA
C0279661|T047||CCS_10|PANCREATIC ACINAR CELL ADENOCARCINOMA
C0279661|T047||CCS_10|PANCREATIC ACINAR CELL CARCINOMA
C1336029|T047||CCS_10|SOLID PSEUDOPAPILLARY CARCINOMA OF PANCREAS 
C1336029|T047||CCS_10|SOLID PSEUDOPAPILLARY CARCINOMA OF PANCREAS
C1336029|T047||CCS_10|PANCREATIC SOLID PSEUDOPAPILLARY CARCINOMA
C1336029|T047||CCS_10|SOLID PSEUDOPAPILLARY CARCINOMA OF THE PANCREAS
C3472164|T047||CCS_10|PRIMARY ADENOCARCINOMA OF PANCREAS 
C3472164|T047||CCS_10|PRIMARY ADENOCARCINOMA OF PANCREAS
C3532881|T047||CCS_10|INTRADUCTAL PAPILLARY MUCINOUS CARCINOMA IN SITU OF PANCREAS 
C3532881|T047||CCS_10|INTRADUCTAL PAPILLARY MUCINOUS NEOPLASM WITH HIGH GRADE DYSPLASIA
C3532881|T047||CCS_10|INTRADUCTAL PAPILLARY MUCINOUS CARCINOMA IN SITU OF PANCREAS
C0153454|T047||CCS_10|MALIGNANT NEOPLASM OF AMPULLA OF VATER
C0153454|T047||CCS_10|MAL NEO AMPULLA OF VATER
C0153454|T047||CCS_10|MALIGNANT NEOPLASM AMPULLA OF VATER
C0153454|T047||CCS_10|MALIGNANT NEOPLASM AMPULLA OF VATER 
C0153454|T047||CCS_10|MALIGNANT TUMOUR OF AMPULLA OF VATER
C0153454|T047||CCS_10|MALIGNANT TUMOR OF AMPULLA OF VATER
C0153454|T047||CCS_10|MALIGNANT TUMOR OF AMPULLA OF VATER 
C0153454|T047||CCS_10|MALIGNANT AMPULLA OF VATER NEOPLASM
C0153454|T047||CCS_10|MALIGNANT AMPULLA OF VATER TUMOR
C0153454|T047||CCS_10|MALIGNANT NEOPLASM OF THE AMPULLA OF VATER
C0153454|T047||CCS_10|MALIGNANT TUMOR OF THE AMPULLA OF VATER
C1282477|T047||CCS_10|PANCREATIC MALIGNANT NEOPLASM, LOCAL RECURRENCE
C1282477|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT NEOPLASM OF PANCREAS
C1282477|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT NEOPLASM OF PANCREAS 
C1282477|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOR OF PANCREAS 
C1282477|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOR OF PANCREAS
C1282477|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOUR OF PANCREAS
C0346976|T047||CCS_10|METASTATIC NEOPLASM TO THE PANCREAS
C0346976|T047||CCS_10|METASTASES TO PANCREAS
C0346976|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF PANCREAS
C0346976|T047||CCS_10|PANCREATIC MALIGNANT NEOPLASM SECONDARY
C0346976|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF PANCREAS 
C0346976|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO THE PANCREAS
C0346976|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM IN THE PANCREAS
C0346976|T047||CCS_10|CANCER METASTATIC TO PANCREAS
C0346976|T047||CCS_10|MALIGNANT NEOPLASM OF PANCREAS METASTATIC
C0346976|T047||CCS_10|PANCREAS NEOPLASM MALIGNANT METASTATIC
C0346976|T047||CCS_10|PANCREATIC CANCER METASTATIC
C0346976|T047||CCS_10|METASTASIS TO PANCREAS
C0346976|T047||CCS_10|PANCREATIC METASTASIS
C0346976|T047||CCS_10|SECONDARY MALIGNANT DEPOSIT IN PANCREAS
C0346976|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO PANCREAS
C0346976|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF PANCREAS 
C0346976|T047||CCS_10|METASTATIC PANCREAS CANCER
C0346976|T047||CCS_10|METASTATIC PANCREATIC CANCER
C0346976|T047||CCS_10|PANCREAS CANCER, METASTATIC
C0346976|T047||CCS_10|PANCREATIC CANCER, METASTATIC
C0346976|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO PANCREAS, NOS
C0346976|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF PANCREAS, NOS
C0346976|T047||CCS_10|METASTATIC CANCER TO THE PANCREAS
C0346976|T047||CCS_10|METASTATIC TUMOR TO THE PANCREAS
C0346976|T047||CCS_10|SECONDARY CANCER TO THE PANCREAS
C0346976|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM TO THE PANCREAS
C0346976|T047||CCS_10|SECONDARY MALIGNANT TUMOR TO THE PANCREAS
C0346648|T047||CCS_10|MALIGNANT NEOPLASM OF EXOCRINE PANCREAS
C0346648|T047||CCS_10|MALIGNANT NEOPLASM OF EXOCRINE PANCREAS 
C0346648|T047||CCS_10|PANCREATIC NEOPLASM MALIGNANT EXOCRINE
C0346648|T047||CCS_10|MALIGNANT TUMOR OF EXOCRINE PANCREAS
C0346648|T047||CCS_10|MALIGNANT TUMOUR OF EXOCRINE PANCREAS
C0346648|T047||CCS_10|PANCREATIC EXOCRINE CANCER
C0346648|T047||CCS_10|MALIGNANT TUMOR OF EXOCRINE PANCREAS 
C0346648|T047||CCS_10|MALIGNANT EXOCRINE PANCREAS NEOPLASM
C0346648|T047||CCS_10|MALIGNANT EXOCRINE PANCREAS TUMOR
C0346648|T047||CCS_10|MALIGNANT NEOPLASM OF THE EXOCRINE PANCREAS
C0346648|T047||CCS_10|MALIGNANT TUMOR OF THE EXOCRINE PANCREAS
C0346650|T047||CCS_10|MALIGNANT NEOPLASM OF ECTOPIC TISSUE OF PANCREAS
C0346650|T047||CCS_10|PANCREATIC NEOPLASM MALIGNANT OF ECTOPIC TISSUE
C0346650|T047||CCS_10|MALIGNANT NEOPLASM OF ECTOPIC TISSUE OF PANCREAS 
C0346650|T047||CCS_10|MALIGNANT NEOPLASM OF ECTOPIC PANCREATIC TISSUE
C0346650|T047||CCS_10|MALIGNANT NEOPLASM OF ECTOPIC PANCREATIC TISSUE 
C0346651|T047||CCS_10|MALIGNANT NEOPLASM OF SPECIFIED SITE OF PANCREAS NOS 
C0346651|T047||CCS_10|MALIGNANT NEOPLASM OF SPECIFIED SITE OF PANCREAS NOS
C1299297|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF PANCREAS
C1299297|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF PANCREAS 
C1299297|T047||CCS_10|PANCREATIC MALIGNANT NEOPLASM PRIMARY
C1299297|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF PANCREAS 
C2205515|T047||CCS_10|MALIGNANT MYOEPITHELIOMA OF PANCREAS
C2205515|T047||CCS_10|MALIGNANT MYOEPITHELIOMA OF PANCREAS 
C2205515|T047||CCS_10|MYOEPITHELIOMA OF PANCREAS
C3836561|T047||CCS_10|PANCREATIC CANCER, SOMATIC
C3836561|T047||CCS_10|PANCREATIC CANCER, SOMATIC 
C1851697|T047||CCS_10|PANCREATIC ISLET CELL ADENOMA
C4030391|T047||CCS_10|BIOPSY OF PANCREAS SHOWED VILLOUS ADENOCARCINOMA 
C4030391|T047||CCS_10|BIOPSY OF PANCREAS SHOWED VILLOUS ADENOCARCINOMA
C4030391|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM ADENOCARCINOMA VILLOUS
C4030470|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT INSULINOMA 
C4030470|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA ISLET CELL INSULINOMA
C4030470|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT INSULINOMA
C4030411|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SMALL CELL SARCOMA 
C4030411|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SMALL CELL SARCOMA
C4030411|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM SARCOMA SMALL CELL
C4030557|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOID SQUAMOUS CELL CARCINOMA 
C4030557|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOID SQUAMOUS CELL CARCINOMA
C4030557|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA SQUAMOUS CELL ADENOID
C4030400|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SQUAMOUS CELL CARCINOMA 
C4030400|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SQUAMOUS CELL CARCINOMA
C4030400|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA SQUAMOUS CELL
C4030506|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM LYMPHOMA HODGKIN'S
C4030506|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HODGKIN'S LYMPHOMA
C4030506|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HODGKIN'S LYMPHOMA 
C4030416|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM ADENOCARCINOMA SCIRRHOUS
C4030416|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SCIRRHOUS ADENOCARCINOMA 
C4030416|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SCIRRHOUS ADENOCARCINOMA
C4030419|T047||CCS_10|BIOPSY PANCREAS MALIG LYMPHOMA PRECURSOR CELL LYMPHOBLASTIC T-CELL
C4030419|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PRECURSOR T-CELL LYMPHOBLASTIC LYMPHOMA 
C4030419|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PRECURSOR T-CELL LYMPHOBLASTIC LYMPHOMA
C4030510|T047||CCS_10|BIOPSY OF PANCREAS SHOWED GRADE 3 FOLLICULAR LYMPHOMA
C4030510|T047||CCS_10|BIOPSY OF PANCREAS SHOWED GRADE 3 FOLLICULAR LYMPHOMA 
C4030510|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM LYMPHOMA FOLLICULAR GRADE 3
C4030482|T047||CCS_10|BIOPSY OF PANCREAS SHOWED LEIOMYOSARCOMA 
C4030482|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM MYOSARCOMA LEIOMYOSARCOMA
C4030482|T047||CCS_10|BIOPSY OF PANCREAS SHOWED LEIOMYOSARCOMA
C4030533|T047||CCS_10|BIOPSY OF PANCREAS SHOWED CARCINOSARCOMA 
C4030533|T047||CCS_10|BIOPSY OF PANCREAS SHOWED CARCINOSARCOMA
C4030533|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOSARCOMA
C4030481|T047||CCS_10|BIOPSY OF PANCREAS SHOWED LYMPHOCYTE-RICH HODGKIN'S LYMPHOMA
C4030481|T047||CCS_10|BIOPSY PANCREAS MALIG NEOPLASM LYMPHOMA HODGKIN'S LYMPHOCYTE-RICH
C4030481|T047||CCS_10|BIOPSY OF PANCREAS SHOWED LYMPHOCYTE-RICH HODGKIN'S LYMPHOMA 
C4030452|T047||CCS_10|BIOPSY PANCREAS MALIG NEOPLASM LYMPHOMA HODGKIN'S MIXED CELLULARITY
C4030452|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MIXED CELLULARITY HODGKIN'S LYMPHOMA
C4030452|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MIXED CELLULARITY HODGKIN'S LYMPHOMA 
C4030505|T047||CCS_10|BIOPSY PANCREAS MALIG LYMPHOMA HODGKIN'S NODULAR SCLEROSIS GRADE 1
C4030505|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HODGKIN'S LYMPHOMA WITH GRADE 1 NODULAR SCLEROSIS 
C4030505|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HODGKIN'S LYMPHOMA WITH GRADE 1 NODULAR SCLEROSIS
C4030497|T047||CCS_10|BIOPSY OF PANCREAS SHOWED INFILTRATING DUCTULAR CARCINOMA
C4030497|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA INFILTRATING DUCTULAR
C4030497|T047||CCS_10|BIOPSY OF PANCREAS SHOWED INFILTRATING DUCTULAR CARCINOMA 
C4030565|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOCARCINOMA IN TUBULOVILLOUS ADENOMA 
C4030565|T047||CCS_10|BIOPSY PANCREAS MALIG NEOPLASM ADENOCARCINOMA IN TUBULOVILLOUS ADENOMA
C4030565|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOCARCINOMA IN TUBULOVILLOUS ADENOMA
C4030562|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOCARCINOMA WITH CARTILAGINOUS AND OSSEOUS METAPLASIA 
C4030562|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOCARCINOMA WITH CARTILAGINOUS AND OSSEOUS METAPLASIA
C4030562|T047||CCS_10|BIOPSY PANCREAS MALIG ADENOCARCINOMA METAPLASTIC CARTILAGINOUS & OSSEOUS
C4030479|T047||CCS_10|BIOPSY PANCREAS MALIG NEOPLASM SARCOMA DESMOPLASTIC SMALL ROUND CELL
C4030479|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT DESMOPLASTIC SMALL ROUND CELL TUMOR 
C4030479|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT DESMOPLASTIC SMALL ROUND CELL TUMOR
C4030516|T047||CCS_10|BIOPSY OF PANCREAS SHOWED GIANT CELL CARCINOMA
C4030516|T047||CCS_10|BIOPSY OF PANCREAS SHOWED GIANT CELL CARCINOMA 
C4030516|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA GIANT CELL
C4030473|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT GLUCAGONOMA
C4030473|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT GLUCAGONOMA 
C4030473|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA ISLET CELL GLUCAGONOMA
C4030504|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HODGKIN'S LYMPHOMA WITH GRADE 2 NODULAR SCLEROSIS
C4030504|T047||CCS_10|BIOPSY PANCREAS MALIG LYMPHOMA HODGKIN'S NODULAR SCLEROSIS GRADE 2
C4030504|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HODGKIN'S LYMPHOMA WITH GRADE 2 NODULAR SCLEROSIS 
C4030456|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM LYMPHOMA MATURE T-CELL
C4030456|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MATURE T-CELL LYMPHOMA 
C4030456|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MATURE T-CELL LYMPHOMA
C4030487|T047||CCS_10|BIOPSY OF PANCREAS SHOWED LANGERHANS CELL SARCOMA
C4030487|T047||CCS_10|BIOPSY OF PANCREAS SHOWED LANGERHANS CELL SARCOMA 
C4030487|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM SARCOMA LANGERHANS CELL
C4030498|T047||CCS_10|BIOPSY OF PANCREAS SHOWED INFILTRATING DUCT CARCINOMA 
C4030498|T047||CCS_10|BIOPSY OF PANCREAS SHOWED INFILTRATING DUCT CARCINOMA
C4030498|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA INFILTRATING DUCT
C4030488|T047||CCS_10|BIOPSY OF PANCREAS SHOWED KERATINIZING SQUAMOUS CELL CARCINOMA 
C4030488|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA SQUAMOUS CELL KERATINIZING
C4030488|T047||CCS_10|BIOPSY OF PANCREAS SHOWED KERATINIZING SQUAMOUS CELL CARCINOMA
C4030532|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM ADENOCARCINOMA CLEAR CELL
C4030532|T047||CCS_10|BIOPSY OF PANCREAS SHOWED CLEAR CELL ADENOCARCINOMA
C4030532|T047||CCS_10|BIOPSY OF PANCREAS SHOWED CLEAR CELL ADENOCARCINOMA 
C4030417|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SARCOMA 
C4030417|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM SARCOMA
C4030417|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SARCOMA
C4030484|T047||CCS_10|BIOPSY OF PANCREAS SHOWED LARGE CELL NEUROENDOCRINE CARCINOMA 
C4030484|T047||CCS_10|BIOPSY PANCREAS MALIG NEOPLASM CARCINOMA LARGE CELL NEUROENDOCRINE
C4030484|T047||CCS_10|BIOPSY OF PANCREAS SHOWED LARGE CELL NEUROENDOCRINE CARCINOMA
C4030392|T047||CCS_10|BIOPSY OF PANCREAS SHOWED VERRUCOUS CARCINOMA
C4030392|T047||CCS_10|BIOPSY OF PANCREAS SHOWED VERRUCOUS CARCINOMA 
C4030392|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA VERRUCOUS
C4030422|T047||CCS_10|BIOPSY OF PANCREAS SHOWED POLYGONAL CELL CARCINOMA
C4030422|T047||CCS_10|BIOPSY OF PANCREAS SHOWED POLYGONAL CELL CARCINOMA 
C4030422|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA POLYGONAL CELL
C4030527|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA CYSTIC HYPERSECRETORY
C4030527|T047||CCS_10|BIOPSY OF PANCREAS SHOWED CYSTIC HYPERSECRETORY CARCINOMA 
C4030527|T047||CCS_10|BIOPSY OF PANCREAS SHOWED CYSTIC HYPERSECRETORY CARCINOMA
C4030513|T047||CCS_10|BIOPSY OF PANCREAS SHOWED GOBLET CELL CARCINOID TUMOR 
C4030513|T047||CCS_10|BIOPSY OF PANCREAS SHOWED GOBLET CELL CARCINOID TUMOR
C4030513|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOID TUMOR GOBLET CELL
C4030409|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SOLID CARCINOMA 
C4030409|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SOLID CARCINOMA
C4030409|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA SOLID
C4030450|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM ADENOCARCINOMA MUCINOUS
C4030450|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MUCINOUS ADENOCARCINOMA
C4030450|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MUCINOUS ADENOCARCINOMA 
C4030521|T047||CCS_10|BIOPSY OF PANCREAS SHOWED EPITHELIOID SARCOMA
C4030521|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM SARCOMA EPITHELIOID
C4030521|T047||CCS_10|BIOPSY OF PANCREAS SHOWED EPITHELIOID SARCOMA 
C4030571|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOCARCINOMA
C4030571|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOCARCINOMA 
C4030571|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM ADENOCARCINOMA
C4030425|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PAPILLARY SQUAMOUS CELL CARCINOMA
C4030425|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PAPILLARY SQUAMOUS CELL CARCINOMA 
C4030425|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA PAPILLARY SQUAMOUS CELL
C4030480|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT CLEAR CELL TYPE NEOPLASM
C4030480|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT CLEAR CELL TYPE NEOPLASM 
C4030480|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CLEAR CELL TYPE
C4030426|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PAPILLARY MUCINOUS CYSTADENOCARCINOMA 
C4030426|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PAPILLARY MUCINOUS CYSTADENOCARCINOMA
C4030426|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CYSTADENOCARCINOMA PAPILLARY MUCINOUS
C4030460|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT SOMATOSTATINOMA 
C4030460|T047||CCS_10|BIOPSY PANCREAS MALIG NEOPLASM CARCINOMA ISLET CELL SOMATOSTATINOMA
C4030460|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT SOMATOSTATINOMA
C4030458|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM LYMPHOMA MARGINAL ZONE B-CELL
C4030458|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MARGINAL ZONE B-CELL LYMPHOMA
C4030458|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MARGINAL ZONE B-CELL LYMPHOMA 
C4030573|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ACINAR CELL CYSTADENOCARCINOMA
C4030573|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ACINAR CELL CYSTADENOCARCINOMA 
C4030573|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM ACINAR CELL CYSTADENOCARCINOMA
C4030441|T047||CCS_10|BIOPSY OF PANCREAS SHOWED NEUROENDOCRINE CARCINOMA
C4030441|T047||CCS_10|BIOPSY OF PANCREAS SHOWED NEUROENDOCRINE CARCINOMA 
C4030441|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA NEUROENDOCRINE
C4030396|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SUPERFICIAL SPREADING ADENOCARCINOMA 
C4030396|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SUPERFICIAL SPREADING ADENOCARCINOMA
C4030396|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM ADENOCARCINOMA SUPERFICIAL SPREADING
C4030563|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOCARCINOMA WITH APOCRINE METAPLASIA
C4030563|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM ADENOCARCINOMA METAPLASTIC APOCRINE
C4030563|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOCARCINOMA WITH APOCRINE METAPLASIA 
C4030453|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MICROINVASIVE SQUAMOUS CELL CARCINOMA
C4030453|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MICROINVASIVE SQUAMOUS CELL CARCINOMA 
C4030453|T047||CCS_10|BIOPSY PANCREAS MALIG NEOPLASM CARCINOMA SQUAMOUS CELL MICROINVASIVE
C4030390|T047||CCS_10|BIOPSY OF PANCREAS SHOWED VIPOMA
C4030390|T047||CCS_10|BIOPSY OF PANCREAS SHOWED VIPOMA 
C4030390|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA ISLET CELL VIPOMA
C4030486|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA LARGE CELL
C4030486|T047||CCS_10|BIOPSY OF PANCREAS SHOWED LARGE CELL CARCINOMA 
C4030486|T047||CCS_10|BIOPSY OF PANCREAS SHOWED LARGE CELL CARCINOMA
C4030499|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HODGKIN'S SARCOMA 
C4030499|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM LYMPHOMA HODGKIN'S SARCOMA
C4030499|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HODGKIN'S SARCOMA
C4030431|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM PANCREATOBLASTOMA
C4030431|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PANCREATOBLASTOMA
C4030431|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PANCREATOBLASTOMA 
C4030523|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA EPITHELIAL-MYOEPITHELIAL
C4030523|T047||CCS_10|BIOPSY OF PANCREAS SHOWED EPITHELIAL-MYOEPITHELIAL CARCINOMA
C4030523|T047||CCS_10|BIOPSY OF PANCREAS SHOWED EPITHELIAL-MYOEPITHELIAL CARCINOMA 
C4030402|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM SARCOMA SPINDLE CELL
C4030402|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SPINDLE CELL SARCOMA 
C4030402|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SPINDLE CELL SARCOMA
C4030412|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA SMALL CELL FUSIFORM CELL
C4030412|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SMALL CELL CARCINOMA, FUSIFORM CELL 
C4030412|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SMALL CELL CARCINOMA, FUSIFORM CELL
C4030507|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HODGKIN'S GRANULOMA
C4030507|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM LYMPHOMA HODGKIN'S GRANULOMA
C4030507|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HODGKIN'S GRANULOMA 
C4030467|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT LYMPHOPLASMACYTIC LYMPHOMA
C4030467|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT LYMPHOPLASMACYTIC LYMPHOMA 
C4030467|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM LYMPHOMA LYMPHOPLASMACYTIC
C4030405|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA SOMATIC
C4030405|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SOMATIC CARCINOMA
C4030405|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SOMATIC CARCINOMA 
C4030508|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HISTIOCYTIC SARCOMA
C4030508|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HISTIOCYTIC SARCOMA 
C4030508|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM SARCOMA HISTIOCYTIC
C4030468|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT LYMPHOMA
C4030468|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM LYMPHOMA
C4030468|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT LYMPHOMA 
C4030414|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SIGNET RING CELL CARCINOMA
C4030414|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA SIGNET RING CELL
C4030414|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SIGNET RING CELL CARCINOMA 
C4030509|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM ADENOCARCINOMA HEPATOID
C4030509|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HEPATOID ADENOCARCINOMA
C4030509|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HEPATOID ADENOCARCINOMA 
C4030570|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM ADENOCARCINOMA IN ADENOMATOUS POLYP
C4030570|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOCARCINOMA IN ADENOMATOUS POLYP
C4030570|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOCARCINOMA IN ADENOMATOUS POLYP 
C4030524|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ENTEROCHROMAFFIN CELL CARCINOID TUMOR 
C4030524|T047||CCS_10|BIOPSY PANCREAS MALIG NEOPLASM CARCINOID TUMOR ENTEROCHROMAFFIN CELL
C4030524|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ENTEROCHROMAFFIN CELL CARCINOID TUMOR
C4030530|T047||CCS_10|BIOPSY OF PANCREAS SHOWED COMPOSITE CARCINOID TUMOR
C4030530|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOID TUMOR COMPOSITE
C4030530|T047||CCS_10|BIOPSY OF PANCREAS SHOWED COMPOSITE CARCINOID TUMOR 
C4030534|T047||CCS_10|BIOPSY PANCREAS MALIG CARCINOMA WITH OSTEOCLAST-LIKE GIANT CELLS
C4030534|T047||CCS_10|BIOPSY OF PANCREAS SHOWED CARCINOMA WITH OSTEOCLAST-LIKE GIANT CELLS
C4030534|T047||CCS_10|BIOPSY OF PANCREAS SHOWED CARCINOMA WITH OSTEOCLAST-LIKE GIANT CELLS 
C4030514|T047||CCS_10|BIOPSY OF PANCREAS SHOWED GLASSY CELL CARCINOMA 
C4030514|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA GLASSY CELL
C4030514|T047||CCS_10|BIOPSY OF PANCREAS SHOWED GLASSY CELL CARCINOMA
C4030401|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SPINDLE CELL SQUAMOUS CELL CARCINOMA
C4030401|T047||CCS_10|BIOPSY PANCREAS MALIG NEOPLASM CARCINOMA SQUAMOUS CELL SPINDLE CELL
C4030401|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SPINDLE CELL SQUAMOUS CELL CARCINOMA 
C4030418|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA PSEUDOSARCOMATOUS
C4030418|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PSEUDOSARCOMATOUS CARCINOMA
C4030418|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PSEUDOSARCOMATOUS CARCINOMA 
C4030469|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT LARGE B-CELL DIFFUSE LYMPHOMA 
C4030469|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM LYMPHOMA LARGE B-CELL DIFFUSE
C4030469|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT LARGE B-CELL DIFFUSE LYMPHOMA
C4030518|T047||CCS_10|BIOPSY OF PANCREAS SHOWED FOLLICULAR LYMPHOMA 
C4030518|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM LYMPHOMA FOLLICULAR
C4030518|T047||CCS_10|BIOPSY OF PANCREAS SHOWED FOLLICULAR LYMPHOMA
C4030465|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM MASTOCYTOSIS
C4030465|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT MASTOCYTOSIS
C4030465|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT MASTOCYTOSIS 
C4030555|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA ADENOSQUAMOUS
C4030555|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOSQUAMOUS CARCINOMA
C4030555|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOSQUAMOUS CARCINOMA 
C4030393|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM SARCOMA UNDIFFERENTIATED
C4030393|T047||CCS_10|BIOPSY OF PANCREAS SHOWED UNDIFFERENTIATED SARCOMA
C4030393|T047||CCS_10|BIOPSY OF PANCREAS SHOWED UNDIFFERENTIATED SARCOMA 
C4030449|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MUCINOUS CYSTADENOCARCINOMA 
C4030449|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CYSTADENOCARCINOMA MUCINOUS
C4030449|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MUCINOUS CYSTADENOCARCINOMA
C4030477|T047||CCS_10|BIOPSY PANCREAS MALIG NEOPLASM CARCINOMA ISLET CELL ENTEROGLUCAGONOMA
C4030477|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT ENTEROGLUCAGONOMA
C4030477|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT ENTEROGLUCAGONOMA 
C4030520|T047||CCS_10|BIOPSY OF PANCREAS SHOWED EXTRAMEDULLARY PLASMACYTOMA
C4030520|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM PLASMACYTOMA EXTRAMEDULLARY
C4030520|T047||CCS_10|BIOPSY OF PANCREAS SHOWED EXTRAMEDULLARY PLASMACYTOMA 
C4030413|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SMALL CELL CARCINOMA
C4030413|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SMALL CELL CARCINOMA 
C4030413|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA SMALL CELL
C4030525|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOSARCOMA EMBRYONAL
C4030525|T047||CCS_10|BIOPSY OF PANCREAS SHOWED EMBRYONAL CARCINOSARCOMA 
C4030525|T047||CCS_10|BIOPSY OF PANCREAS SHOWED EMBRYONAL CARCINOSARCOMA
C4030457|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MAST CELL SARCOMA
C4030457|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM SARCOMA MAST CELL
C4030457|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MAST CELL SARCOMA 
C4030519|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM SARCOMA FOLLICULAR DENDRITIC CELL
C4030519|T047||CCS_10|BIOPSY OF PANCREAS SHOWED FOLLICULAR DENDRITIC CELL SARCOMA
C4030519|T047||CCS_10|BIOPSY OF PANCREAS SHOWED FOLLICULAR DENDRITIC CELL SARCOMA 
C4030443|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM MYOSARCOMA LEIOMYOSARCOMA MYXOID
C4030443|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MYXOID LEIOMYOSARCOMA 
C4030443|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MYXOID LEIOMYOSARCOMA
C4030564|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM ADENOCARCINOMA IN VILLOUS ADENOMA
C4030564|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOCARCINOMA IN VILLOUS ADENOMA
C4030564|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOCARCINOMA IN VILLOUS ADENOMA 
C4030464|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOSARCOMA MYOEPITHELIOMA
C4030464|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT MYOEPITHELIOMA
C4030464|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT MYOEPITHELIOMA 
C4030502|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HODGKIN'S LYMPHOMA WITH LYMPHOCYTIC DEPLETION WITH DIFFUSE FIBROSIS
C4030502|T047||CCS_10|BIOPSY PANCREAS MALIG LYMPHOMA HODGKIN'S LYMPHOCYT DEPLET DIFFUSE FIBROSIS
C4030502|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HODGKIN'S LYMPHOMA WITH LYMPHOCYTIC DEPLETION WITH DIFFUSE FIBROSIS 
C4030500|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HODGKIN'S LYMPHOMA WITH NODULAR SCLEROSIS CELLULAR PHASE 
C4030500|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HODGKIN'S LYMPHOMA WITH NODULAR SCLEROSIS CELLULAR PHASE
C4030500|T047||CCS_10|BIOPSY PANCREAS MALIG LYMPHOMA HODGKIN'S NODULAR SCLEROSIS CELLULAR PHASE
C4030408|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SOLID PSEUDOPAPILLARY CARCINOMA
C4030408|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA SOLID PSEUDOPAPILLARY
C4030408|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SOLID PSEUDOPAPILLARY CARCINOMA 
C4030495|T047||CCS_10|BIOPSY OF PANCREAS SHOWED INTRACYSTIC CARCINOMA
C4030495|T047||CCS_10|BIOPSY OF PANCREAS SHOWED INTRACYSTIC CARCINOMA 
C4030495|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA INTRACYSTIC
C4030558|T047||CCS_10|BIOPSY PANCREAS MALIG NEOPLASM ADENOCARCINOMA METAPLASTIC SQUAMOUS
C4030558|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOCARCINOMA WITH SQUAMOUS METAPLASIA 
C4030558|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOCARCINOMA WITH SQUAMOUS METAPLASIA
C4030560|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOCARCINOMA WITH NEUROENDOCRINE DIFFERENTIATION
C4030560|T047||CCS_10|BIOPSY PANCREAS MALIG ADENOCARC METAPLASTIC NEUROENDOCRINE DIFFERENTIATION
C4030560|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOCARCINOMA WITH NEUROENDOCRINE DIFFERENTIATION 
C4030539|T047||CCS_10|BIOPSY OF PANCREAS SHOWED CARCINOMA 
C4030539|T047||CCS_10|BIOPSY OF PANCREAS SHOWED CARCINOMA
C4030539|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA
C4030403|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SPINDLE CELL CARCINOMA 
C4030403|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA SPINDLE CELL
C4030403|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SPINDLE CELL CARCINOMA
C4030517|T047||CCS_10|BIOPSY OF PANCREAS SHOWED GIANT CELL AND SPINDLE CELL CARCINOMA
C4030517|T047||CCS_10|BIOPSY OF PANCREAS SHOWED GIANT CELL AND SPINDLE CELL CARCINOMA 
C4030517|T047||CCS_10|BIOPSY PANCREAS MALIG NEOPLASM CARCINOMA GIANT CELL AND SPINDLE CELL
C4030483|T047||CCS_10|BIOPSY OF PANCREAS SHOWED LARGE CELL, NONKERATINIZING SQUAMOUS CELL CARCINOMA
C4030483|T047||CCS_10|BIOPSY OF PANCREAS SHOWED LARGE CELL, NONKERATINIZING SQUAMOUS CELL CARCINOMA 
C4030483|T047||CCS_10|BIOPSY PANCREAS MALIG CARCINOMA SQUAMOUS CELL LARGE CELL NONKERATINIZING
C4030410|T047||CCS_10|BIOPSY PANCREAS MALIG CARCINOMA SQUAMOUS CELL SMALL CELL NONKERATINIZING
C4030410|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SMALL CELL, NONKERATINIZING SQUAMOUS CELL CARCINOMA 
C4030410|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SMALL CELL, NONKERATINIZING SQUAMOUS CELL CARCINOMA
C4030475|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT GASTRINOMA 
C4030475|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT GASTRINOMA
C4030475|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA ISLET CELL GASTRINOMA
C4030472|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT HISTIOCYTOSIS 
C4030472|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT HISTIOCYTOSIS
C4030472|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM LYMPHOMA HISTIOCYTOSIS
C4030541|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM LYMPHOMA BURKITT'S
C4030541|T047||CCS_10|BIOPSY OF PANCREAS SHOWED BURKITT'S LYMPHOMA
C4030541|T047||CCS_10|BIOPSY OF PANCREAS SHOWED BURKITT'S LYMPHOMA 
C4030421|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PRECURSOR B-CELL LYMPHOBLASTIC LYMPHOMA
C4030421|T047||CCS_10|BIOPSY PANCREAS MALIG LYMPHOMA PRECURSOR CELL LYMPHOBLASTIC B-CELL
C4030421|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PRECURSOR B-CELL LYMPHOBLASTIC LYMPHOMA 
C4030444|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM MYOSARCOMA
C4030444|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MYOSARCOMA 
C4030444|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MYOSARCOMA
C4030446|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM ADENOCARCINOMA MUCIN-PRODUCING
C4030446|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MUCIN-PRODUCING ADENOCARCINOMA
C4030446|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MUCIN-PRODUCING ADENOCARCINOMA 
C4030526|T047||CCS_10|BIOPSY OF PANCREAS SHOWED DESMOPLASTIC TYPE DUCT CARCINOMA 
C4030526|T047||CCS_10|BIOPSY OF PANCREAS SHOWED DESMOPLASTIC TYPE DUCT CARCINOMA
C4030526|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA DUCT, DESMOPLASTIC TYPE
C4030429|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA PAPILLARY
C4030429|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PAPILLARY CARCINOMA 
C4030429|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PAPILLARY CARCINOMA
C4030548|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOID TUMOR ATYPICAL
C4030548|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ATYPICAL CARCINOID TUMOR
C4030548|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ATYPICAL CARCINOID TUMOR 
C4030461|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT SMALL CELL TYPE NEOPLASM
C4030461|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM SMALL CELL TYPE
C4030461|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT SMALL CELL TYPE NEOPLASM 
C4030394|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA UNDIFFERENTIATED
C4030394|T047||CCS_10|BIOPSY OF PANCREAS SHOWED UNDIFFERENTIATED CARCINOMA
C4030394|T047||CCS_10|BIOPSY OF PANCREAS SHOWED UNDIFFERENTIATED CARCINOMA 
C4030485|T047||CCS_10|BIOPSY OF PANCREAS SHOWED LARGE CELL CARCINOMA WITH RHABDOID PHENOTYPE
C4030485|T047||CCS_10|BIOPSY OF PANCREAS SHOWED LARGE CELL CARCINOMA WITH RHABDOID PHENOTYPE 
C4030485|T047||CCS_10|BIOPSY PANCREAS MALIG CARCINOMA LARGE CELL WITH RHABDOID PHENOTYPE
C4030529|T047||CCS_10|BIOPSY OF PANCREAS SHOWED COMPOSITE HODGKIN'S AND NON-HODGKIN'S LYMPHOMA 
C4030529|T047||CCS_10|BIOPSY OF PANCREAS SHOWED COMPOSITE HODGKIN'S AND NON-HODGKIN'S LYMPHOMA
C4030529|T047||CCS_10|BIOPSY PANCREAS MALIG LYMPHOMA COMPOSITE HODGKIN'S & NON-HODGKIN'S
C4030511|T047||CCS_10|BIOPSY OF PANCREAS SHOWED GRADE 2 FOLLICULAR LYMPHOMA
C4030511|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM LYMPHOMA FOLLICULAR GRADE 2
C4030511|T047||CCS_10|BIOPSY OF PANCREAS SHOWED GRADE 2 FOLLICULAR LYMPHOMA 
C4030420|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PRECURSOR CELL LYMPHOBLASTIC LYMPHOMA
C4030420|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PRECURSOR CELL LYMPHOBLASTIC LYMPHOMA 
C4030420|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM LYMPHOMA PRECURSOR CELL LYMPHOBLASTIC
C4030424|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PLASMACYTOMA 
C4030424|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM PLASMACYTOMA
C4030424|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PLASMACYTOMA
C4030574|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ACINAR CELL CARCINOMA
C4030574|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ACINAR CELL CARCINOMA 
C4030574|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA ACINAR CELL
C4030430|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PAPILLARY ADENOCARCINOMA 
C4030430|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM ADENOCARCINOMA PAPILLARY
C4030430|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PAPILLARY ADENOCARCINOMA
C4030478|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT ENTEROCHROMAFFIN-LIKE CELL CARCINOID TUMOR
C4030478|T047||CCS_10|BIOPSY PANCREAS MALIG CARCINOID TUMOR ENTEROCHROMAFFIN-LIKE CELL
C4030478|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT ENTEROCHROMAFFIN-LIKE CELL CARCINOID TUMOR 
C4030459|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT SPINDLE CELL TYPE NEOPLASM 
C4030459|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM SPINDLE CELL TYPE
C4030459|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT SPINDLE CELL TYPE NEOPLASM
C4030423|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PLEOMORPHIC CARCINOMA 
C4030423|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA PLEOMORPHIC
C4030423|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PLEOMORPHIC CARCINOMA
C4030528|T047||CCS_10|BIOPSY OF PANCREAS SHOWED CYSTADENOCARCINOMA
C4030528|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA CYSTADENOCARCINOMA
C4030528|T047||CCS_10|BIOPSY OF PANCREAS SHOWED CYSTADENOCARCINOMA 
C4030496|T047||CCS_10|BIOPSY OF PANCREAS SHOWED INTERDIGITATING DENDRITIC CELL SARCOMA
C4030496|T047||CCS_10|BIOPSY PANCREAS MALIG NEOPLASM SARCOMA INTERDIGITATING DENDRITIC CELL
C4030496|T047||CCS_10|BIOPSY OF PANCREAS SHOWED INTERDIGITATING DENDRITIC CELL SARCOMA 
C4030439|T047||CCS_10|BIOPSY OF PANCREAS SHOWED NON-HODGKIN'S LYMPHOMA
C4030439|T047||CCS_10|BIOPSY OF PANCREAS SHOWED NON-HODGKIN'S LYMPHOMA 
C4030439|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM LYMPHOMA NON-HODGKIN'S
C4030503|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HODGKIN'S LYMPHOMA WITH LYMPHOCYTIC DEPLETION
C4030503|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HODGKIN'S LYMPHOMA WITH LYMPHOCYTIC DEPLETION 
C4030503|T047||CCS_10|BIOPSY PANCREAS MALIG LYMPHOMA HODGKIN'S LYMPHOCYTIC DEPLETION
C4030531|T047||CCS_10|BIOPSY OF PANCREAS SHOWED COMEDOCARCINOMA 
C4030531|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA COMEDOCARCINOMA
C4030531|T047||CCS_10|BIOPSY OF PANCREAS SHOWED COMEDOCARCINOMA
C4030427|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PAPILLARY CYSTADENOCARCINOMA 
C4030427|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CYSTADENOCARCINOMA PAPILLARY
C4030427|T047||CCS_10|BIOPSY OF PANCREAS SHOWED PAPILLARY CYSTADENOCARCINOMA
C4030559|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOCARCINOMA WITH SPINDLE CELL METAPLASIA 
C4030559|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOCARCINOMA WITH SPINDLE CELL METAPLASIA
C4030559|T047||CCS_10|BIOPSY PANCREAS MALIG NEOPLASM ADENOCARCINOMA METAPLASTIC SPINDLE CELL
C4030572|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOID TUMOR ADENOCARCINOID
C4030572|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOCARCINOID TUMOR 
C4030572|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ADENOCARCINOID TUMOR
C4030466|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT MANTLE CELL LYMPHOMA
C4030466|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT MANTLE CELL LYMPHOMA 
C4030466|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM LYMPHOMA MANTLE CELL
C4030471|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT IMMUNOBLASTIC LARGE B-CELL DIFFUSE LYMPHOMA
C4030471|T047||CCS_10|BIOPSY PANCREAS MALIG LYMPHOMA LARGE B-CELL DIFFUSE IMMUNOBLASTIC
C4030471|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT IMMUNOBLASTIC LARGE B-CELL DIFFUSE LYMPHOMA 
C4030522|T047||CCS_10|BIOPSY OF PANCREAS SHOWED EPITHELIOID LEIOMYOSARCOMA
C4030522|T047||CCS_10|BIOPSY OF PANCREAS SHOWED EPITHELIOID LEIOMYOSARCOMA 
C4030522|T047||CCS_10|BIOPSY PANCREAS MALIG NEOPLASM MYOSARCOMA LEIOMYOSARCOMA EPITHELIOID
C4030454|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MEDULLARY CARCINOMA 
C4030454|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MEDULLARY CARCINOMA
C4030454|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA MEDULLARY
C4030547|T047||CCS_10|BIOPSY OF PANCREAS SHOWED BASAL CELL ADENOCARCINOMA 
C4030547|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM ADENOCARCINOMA BASAL CELL
C4030547|T047||CCS_10|BIOPSY OF PANCREAS SHOWED BASAL CELL ADENOCARCINOMA
C4030451|T047||CCS_10|BIOPSY PANCREAS MALIG MIXED ISLET CELL & EXOCRINE ADENOCARCINOMA
C4030451|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MIXED ISLET CELL AND EXOCRINE ADENOCARCINOMA 
C4030451|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MIXED ISLET CELL AND EXOCRINE ADENOCARCINOMA
C4030476|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT EPITHELIOMA 
C4030476|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA EPITHELIOMA
C4030476|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT EPITHELIOMA
C4030462|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT SMALL B-CELL LYMPHOCYTIC LYMPHOMA 
C4030462|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM LYMPHOMA SMALL B-CELL LYMPHOCYTIC
C4030462|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT SMALL B-CELL LYMPHOCYTIC LYMPHOMA
C4030501|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM LYMPHOMA HODGKIN'S NODULAR SCLEROSIS
C4030501|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HODGKIN'S LYMPHOMA WITH NODULAR SCLEROSIS 
C4030501|T047||CCS_10|BIOPSY OF PANCREAS SHOWED HODGKIN'S LYMPHOMA WITH NODULAR SCLEROSIS
C4030493|T047||CCS_10|BIOPSY PANCREAS MALIG ADENOCARCINOMA INTRADUCTAL PAPILLARY W/ INVASION
C4030493|T047||CCS_10|BIOPSY OF PANCREAS SHOWED INTRADUCTAL PAPILLARY ADENOCARCINOMA WITH INVASION 
C4030493|T047||CCS_10|BIOPSY OF PANCREAS SHOWED INTRADUCTAL PAPILLARY ADENOCARCINOMA WITH INVASION
C4030463|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT NEOPLASM
C4030463|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM
C4030463|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT NEOPLASM 
C4030490|T047||CCS_10|BIOPSY PANCREAS MALIG CARCINOMA INTRADUCTAL PAPILLARY-MUCINOUS INVASIVE
C4030490|T047||CCS_10|BIOPSY OF PANCREAS SHOWED INVASIVE INTRADUCTAL PAPILLARY-MUCINOUS CARCINOMA
C4030490|T047||CCS_10|BIOPSY OF PANCREAS SHOWED INVASIVE INTRADUCTAL PAPILLARY-MUCINOUS CARCINOMA 
C4030395|T047||CCS_10|BIOPSY OF PANCREAS SHOWED TUBULAR ADENOCARCINOMA
C4030395|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM ADENOCARCINOMA TUBULAR
C4030395|T047||CCS_10|BIOPSY OF PANCREAS SHOWED TUBULAR ADENOCARCINOMA 
C4030515|T047||CCS_10|BIOPSY OF PANCREAS SHOWED GIANT CELL SARCOMA 
C4030515|T047||CCS_10|BIOPSY OF PANCREAS SHOWED GIANT CELL SARCOMA
C4030515|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM SARCOMA GIANT CELL
C4030474|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM GIANT CELL TYPE
C4030474|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT GIANT CELL TYPE NEOPLASM 
C4030474|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MALIGNANT GIANT CELL TYPE NEOPLASM
C4030554|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ANAPLASTIC CARCINOMA 
C4030554|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ANAPLASTIC CARCINOMA
C4030554|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA ANAPLASTIC
C4030397|T047||CCS_10|BIOPSY PANCREAS MALIG CARCINOMA SQUAMOUS CELL WITH HORN FORMATION
C4030397|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SQUAMOUS CELL CARCINOMA WITH HORN FORMATION
C4030397|T047||CCS_10|BIOPSY OF PANCREAS SHOWED SQUAMOUS CELL CARCINOMA WITH HORN FORMATION 
C4030535|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA SIMPLEX
C4030535|T047||CCS_10|BIOPSY OF PANCREAS SHOWED CARCINOMA SIMPLEX 
C4030535|T047||CCS_10|BIOPSY OF PANCREAS SHOWED CARCINOMA SIMPLEX
C4030445|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MUCOEPIDERMOID CARCINOMA 
C4030445|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOMA MUCOEPIDERMOID
C4030445|T047||CCS_10|BIOPSY OF PANCREAS SHOWED MUCOEPIDERMOID CARCINOMA
C4030512|T047||CCS_10|BIOPSY OF PANCREAS SHOWED GRADE 1 FOLLICULAR LYMPHOMA
C4030512|T047||CCS_10|BIOPSY OF PANCREAS SHOWED GRADE 1 FOLLICULAR LYMPHOMA 
C4030512|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM LYMPHOMA FOLLICULAR GRADE 1
C4030550|T047||CCS_10|BIOPSY PANCREAS MALIG NEOPLASM LYMPHOMA MATURE T-CELL ANGIOIMMUNOBLASTIC
C4030550|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ANGIOIMMUNOBLASTIC T-CELL LYMPHOMA 
C4030550|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ANGIOIMMUNOBLASTIC T-CELL LYMPHOMA
C4030549|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ANGIOMYOSARCOMA 
C4030549|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM MYOSARCOMA ANGIOMYOSARCOMA
C4030549|T047||CCS_10|BIOPSY OF PANCREAS SHOWED ANGIOMYOSARCOMA
C4030540|T047||CCS_10|BIOPSY OF PANCREAS SHOWED CARCINOID TUMOR 
C4030540|T047||CCS_10|BIOPSY PANCREAS MALIGNANT NEOPLASM CARCINOID TUMOR
C4030540|T047||CCS_10|BIOPSY OF PANCREAS SHOWED CARCINOID TUMOR
C1409082|T047||CCS_10|PANCREAS; ISLET CELL ADENOCARCINOMA WITH EXOCRINE
C1386256|T047||CCS_10|ADENOCARCINOMA; ISLET CELL WITH EXOCRINE, UNSPECIFIED SITE
C1391905|T047||CCS_10|CARCINOMA; ISLET CELL, MET EXOCRINE, UNSPECIFIED SITE
C1396226|T047||CCS_10|ISLET CELL; ADENOCARCINOMA, MET EXOCRINE, UNSPECIFIED SITE
C1396227|T047||CCS_10|ISLET CELL; CARCINOMA WITH EXOCRINE, UNSPECIFIED SITE
C0279884|T047||CCS_10|CELLULAR DIAGNOSIS, PANCREATIC CANCER
C0279884|T047||CCS_10|PANCREAS CANCER CELLULAR DIAGNOSIS
C0279884|T047||CCS_10|PANCREATIC CANCER CELLULAR DIAGNOSIS
C0280222|T047||CCS_10|STAGE, PANCREATIC CANCER
C0280222|T047||CCS_10|PANCREATIC CANCER STAGE
C1335307|T047||CCS_10|MALIGNANT LYMPHOMA OF PANCREATIC LYMPH NODES 
C1335307|T047||CCS_10|MALIGNANT LYMPHOMA OF PANCREATIC LYMPH NODES
C1335307|T047||CCS_10|PANCREATIC LYMPHOMA
C1335307|T047||CCS_10|LYMPHOMA OF PANCREAS
C1335307|T047||CCS_10|LYMPHOMA OF THE PANCREAS
C1276580|T047||CCS_10|T2: TUMOR LIMITED TO PANCREAS AND > 2 CM IN GREATEST DIMENSION 
C1276580|T047||CCS_10|T2: TUMOR LIMITED TO PANCREAS AND > 2 CM IN GREATEST DIMENSION
C1276580|T047||CCS_10|T2: TUMOUR LIMITED TO PANCREAS AND > 2 CM IN GREATEST DIMENSION
C1276580|T047||CCS_10|T2: TUMOR LIMITED TO PANCREAS AND > 2 CM IN GREATEST DIMENSION (TUMOR STAGING)
C0341485|T047||CCS_10|MALIGNANT CYSTIC NEOPLASM OF EXOCRINE PANCREAS
C0341485|T047||CCS_10|PANCREATIC NEOPLASM MALIGNANT EXOCRINE CYSTIC
C0341485|T047||CCS_10|MALIGNANT CYSTIC NEOPLASM OF EXOCRINE PANCREAS 
C0341485|T047||CCS_10|MALIGNANT CYSTIC TUMOR OF EXOCRINE PANCREAS
C0341485|T047||CCS_10|MALIGNANT CYSTIC TUMOUR OF EXOCRINE PANCREAS
C0341485|T047||CCS_10|MALIGNANT CYSTIC TUMOR OF EXOCRINE PANCREAS 
C0238337|T047||CCS_10|CYSTADENOCARCINOMA OF PANCREAS 
C0238337|T047||CCS_10|CYSTADENOCARCINOMA OF PANCREAS
C0238337|T047||CCS_10|CYSTADENOCARCINOMA - PANCREAS
C0238337|T047||CCS_10|CYSTADENOCARCINOMA OF THE PANCREAS
C0238337|T047||CCS_10|CYSTADENOCARCINOMA PANCREAS
C0238337|T047||CCS_10|CYSTADENOCARCINOMA OF PANCREAS 
C0238337|T047||CCS_10|PANCREATIC CYSTADENOCARCINOMA
C0345933|T047||CCS_10|PANCREATIC CARCINOID TUMOR
C0345933|T047||CCS_10|CARCINOID NEOPLASM OF PANCREAS
C0345933|T047||CCS_10|CARCINOID NEOPLASM OF THE PANCREAS
C0345933|T047||CCS_10|CARCINOID TUMOR OF PANCREAS
C0345933|T047||CCS_10|CARCINOID TUMOR OF THE PANCREAS
C0345933|T047||CCS_10|PANCREATIC SEROTONIN PRODUCING NEOPLASM
C0345933|T047||CCS_10|EC CELL, SEROTONIN PRODUCING PANCREATIC NET
C0345933|T047||CCS_10|PANCREATIC SEROTONIN PRODUCING TUMOR
C0345933|T047||CCS_10|ENTEROCHROMAFFIN CELL SEROTONIN-PRODUCING PANCREATIC NEUROENDOCRINE TUMOR
C0345933|T047||CCS_10|EC CELL, SEROTONIN PRODUCING PANCREATIC NEUROENDOCRINE TUMOR
C0345933|T047||CCS_10|CARCINOID TUMOUR OF THE PANCREAS
C0345933|T047||CCS_10|CARCINOID TUMOUR OF PANCREAS
C0345933|T047||CCS_10|CARCINOID TUMOR OF PANCREAS 
C0345933|T047||CCS_10|SEROTONIN-PRODUCING TUMOR OF PANCREAS
C0345933|T047||CCS_10|SEROTONIN-PRODUCING TUMOR OF THE PANCREAS
C2033026|T047||CCS_10|LYMPHOCYTE-RICH HODGKIN'S LYMPHOMA OF PANCREAS 
C2033026|T047||CCS_10|LYMPHOCYTE-RICH HODGKIN'S LYMPHOMA OF PANCREAS
C2033030|T047||CCS_10|NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF PANCREAS 
C2033030|T047||CCS_10|NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF PANCREAS
C2033048|T047||CCS_10|GRADE 3 FOLLICULAR LYMPHOMA OF PANCREAS 
C2033048|T047||CCS_10|GRADE 3 FOLLICULAR LYMPHOMA OF PANCREAS
C2033055|T047||CCS_10|MATURE T-CELL LYMPHOMA OF PANCREAS 
C2033055|T047||CCS_10|MATURE T-CELL LYMPHOMA OF PANCREAS
C2046512|T047||CCS_10|PANCREATIC MALIGNANT LYMPHOMA HODGKIN'S AND NON-HODGKIN'S
C2046512|T047||CCS_10|COMPOSITE HODGKIN'S AND NON-HODGKIN'S LYMPHOMA OF PANCREAS 
C2046512|T047||CCS_10|COMPOSITE HODGKIN'S AND NON-HODGKIN'S LYMPHOMA OF PANCREAS
C2033052|T047||CCS_10|LYMPHOPLASMACYTIC LYMPHOMA OF PANCREAS
C2033052|T047||CCS_10|LYMPHOPLASMACYTIC LYMPHOMA OF PANCREAS 
C2033045|T047||CCS_10|FOLLICULAR LYMPHOMA OF PANCREAS
C2033045|T047||CCS_10|FOLLICULAR LYMPHOMA OF PANCREAS 
C2033046|T047||CCS_10|GRADE 1 FOLLICULAR LYMPHOMA OF PANCREAS 
C2033046|T047||CCS_10|GRADE 1 FOLLICULAR LYMPHOMA OF PANCREAS
C2046585|T047||CCS_10|HODGKIN'S GRANULOMA OF PANCREAS
C2046585|T047||CCS_10|HODGKIN'S GRANULOMA OF PANCREAS 
C2033058|T047||CCS_10|SMALL B-CELL LYMPHOCYTIC LYMPHOMA OF PANCREAS
C2033058|T047||CCS_10|SMALL B-CELL LYMPHOCYTIC LYMPHOMA OF PANCREAS 
C2033053|T047||CCS_10|MANTLE CELL LYMPHOMA OF PANCREAS
C2033053|T047||CCS_10|MANTLE CELL LYMPHOMA OF PANCREAS 
C2033051|T047||CCS_10|IMMUNOBLASTIC LARGE B-CELL DIFFUSE LYMPHOMA OF PANCREAS 
C2033051|T047||CCS_10|IMMUNOBLASTIC LARGE B-CELL DIFFUSE LYMPHOMA OF PANCREAS
C2113717|T047||CCS_10|PRECURSOR CELL LYMPHOBLASTIC LYMPHOMA OF PANCREAS 
C2113717|T047||CCS_10|PRECURSOR CELL LYMPHOBLASTIC LYMPHOMA OF PANCREAS
C2205509|T047||CCS_10|MAST CELL SARCOMA OF PANCREAS
C2205509|T047||CCS_10|MAST CELL SARCOMA OF PANCREAS 
C2033050|T047||CCS_10|LARGE B-CELL DIFFUSE LYMPHOMA OF PANCREAS 
C2033050|T047||CCS_10|LARGE B-CELL DIFFUSE LYMPHOMA OF PANCREAS
C2033047|T047||CCS_10|GRADE 2 FOLLICULAR LYMPHOMA OF PANCREAS
C2033047|T047||CCS_10|GRADE 2 FOLLICULAR LYMPHOMA OF PANCREAS 
C2113646|T047||CCS_10|PRECURSOR B-CELL LYMPHOBLASTIC LYMPHOMA OF PANCREAS 
C2113646|T047||CCS_10|PRECURSOR B-CELL LYMPHOBLASTIC LYMPHOMA OF PANCREAS
C2113786|T047||CCS_10|PRECURSOR T-CELL LYMPHOBLASTIC LYMPHOMA OF PANCREAS
C2113786|T047||CCS_10|PRECURSOR T-CELL LYMPHOBLASTIC LYMPHOMA OF PANCREAS 
C2033029|T047||CCS_10|MIXED CELLULARITY HODGKIN'S LYMPHOMA OF PANCREAS
C2033029|T047||CCS_10|MIXED CELLULARITY HODGKIN'S LYMPHOMA OF PANCREAS 
C2033033|T047||CCS_10|GRADE 2 NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF PANCREAS 
C2033033|T047||CCS_10|GRADE 2 NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF PANCREAS
C2033054|T047||CCS_10|MARGINAL ZONE B-CELL LYMPHOMA OF PANCREAS 
C2033054|T047||CCS_10|MARGINAL ZONE B-CELL LYMPHOMA OF PANCREAS
C2033056|T047||CCS_10|ANGIOIMMUNOBLASTIC T-CELL LYMPHOMA OF PANCREAS
C2033056|T047||CCS_10|ANGIOIMMUNOBLASTIC T-CELL LYMPHOMA OF PANCREAS 
C2033056|T047||CCS_10|ANGIOIMMUNOBLASTIC LYMPHADENOPATHY WITH DYSPROTEINEMIA (AILD) OF PANCREAS
C2033032|T047||CCS_10|GRADE 1 NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF PANCREAS
C2033032|T047||CCS_10|GRADE 1 NODULAR SCLEROSING HODGKIN'S LYMPHOMA OF PANCREAS 
C2033057|T047||CCS_10|NK/T-CELL LYMPHOMA OF PANCREAS 
C2033057|T047||CCS_10|NK/T-CELL LYMPHOMA OF PANCREAS
C2033027|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION OF PANCREAS 
C2033027|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION OF PANCREAS
C2033028|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION, DIFFUSE FIBROSIS OF PANCREAS
C2033028|T047||CCS_10|HODGKIN'S DISEASE, LYMPHOCYTIC DEPLETION, DIFFUSE FIBROSIS OF PANCREAS 
C2033031|T047||CCS_10|NODULAR SCLEROSING HODGKIN'S LYMPHOMA IN CELLULAR PHASE OF PANCREAS
C2033031|T047||CCS_10|NODULAR SCLEROSING HODGKIN'S LYMPHOMA IN CELLULAR PHASE OF PANCREAS 
C2046725|T047||CCS_10|HODGKIN'S SARCOMA OF PANCREAS 
C2046725|T047||CCS_10|HODGKIN'S SARCOMA OF PANCREAS
C2033049|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF PANCREAS
C2033049|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF PANCREAS 
C2205522|T047||CCS_10|SEZARY SYNDROME OF PANCREAS 
C2205522|T047||CCS_10|SEZARY SYNDROME OF PANCREAS
C0153620|T047||CCS_10|MALIGNANT NEOPLASM OF URETHRA
C0153620|T047||CCS_10|MALIGNANT NEOPLASM OF URETHRA 
C0153620|T047||CCS_10|MALIGNANT TUMOR OF URETHRA
C0153620|T047||CCS_10|MALIGN NEOPL URETHRA
C0153620|T047||CCS_10|MALIGNANT TUMOUR OF URETHRA
C0153620|T047||CCS_10|MALIGNANT TUMOUR OF URETHRA 
C0153620|T047||CCS_10|MALIGNANT URETHRAL TUMOR
C0153620|T047||CCS_10|MALIGNANT URETHRAL TUMOUR
C0153620|T047||CCS_10|MALIGNANT TUMOR OF URETHRA 
C0153620|T047||CCS_10|MALIGNANT NEOPLASM OF THE URETHRA
C0153620|T047||CCS_10|MALIGNANT TUMOR OF THE URETHRA
C0153620|T047||CCS_10|MALIGNANT URETHRA NEOPLASM
C0153620|T047||CCS_10|MALIGNANT URETHRA TUMOR
C0153620|T047||CCS_10|MALIGNANT URETHRAL NEOPLASM
C0153620|T047||CCS_10|NEOPLASM MALIG;URETHRA
C0153620|T047||CCS_10|MALIGNANT NEOSPLASM OF THE URETHRA
C0153621|T047||CCS_10|MALIGNANT NEOPLASM OF PARAURETHRAL GLANDS
C0153621|T047||CCS_10|PARAURETHRAL GLAND
C0153621|T047||CCS_10|MALIGNANT NEOPLASM OF PARAURETHRAL GLAND
C0153621|T047||CCS_10|MALIGNANT NEOPLASM OF PARAURETHRAL GLAND 
C0153621|T047||CCS_10|MALIGNANT TUMOR OF PARAURETHRAL GLAND
C0153621|T047||CCS_10|MAL NEO PARAURETHRAL
C0153621|T047||CCS_10|MALIGNANT TUMOUR OF PARAURETHRAL GLAND
C0153621|T047||CCS_10|MALIGNANT TUMOR OF PARAURETHRAL GLAND 
C0349055|T047||CCS_10|MALIGNANT NEOPLASM OVERLAPPING URINARY ORGAN SITE
C0349055|T047||CCS_10|OVERLAPPING LESION OF URINARY ORGANS
C0349055|T047||CCS_10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF URINARY ORGANS
C0349055|T047||CCS_10|MALIGNANT NEOPLASM OF URINARY ORGANS OVERLAPPING SITES
C0349055|T047||CCS_10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF URINARY ORGANS 
C0349055|T047||CCS_10|MALIGNANT NEOPLASM OF OVERLAPPING LESION OF URINARY ORGANS
C0349055|T047||CCS_10|MALIGNANT NEOPLASM OF OVERLAPPING LESION OF URINARY ORGANS 
C0348371|T047||CCS_10|MALIGNANT NEOPLASM OF URINARY ORGAN, UNSPECIFIED
C0348371|T047||CCS_10|URINARY ORGAN, UNSPECIFIED
C0348371|T047||CCS_10|MAL NEO URINARY NOS
C0348371|T047||CCS_10|CANCER OF URINARY ORGANS
C0348371|T047||CCS_10|MALIGNANT NEOPLASM OF URINARY ORGAN 
C0348371|T047||CCS_10|CANCER OF URINARY ORGAN
C0348371|T047||CCS_10|MALIGNANT NEOPLASM OF URINARY ORGAN
C0348371|T047||CCS_10|[X]MALIGNANT NEOPLASM OF URINARY ORGAN, UNSPECIFIED
C0348371|T047||CCS_10|[X]MALIGNANT NEOPLASM OF URINARY ORGAN, UNSPECIFIED 
C0348371|T047||CCS_10|URINARY ORGANS--CANCER
C0348371|T047||CCS_10|MALIGNANT NEOPLASM OF URINARY ORGAN, SITE UNSPECIFIED
C0346890|T047|34|CCS_10|MALIGNANT NEOPLASM OF OTHER AND UNSPECIFIED URINARY ORGANS|CANCER OF OTHER URINARY ORGANS
C0346890|T047|34|CCS_10|CANCER OF OTHER URINARY ORGANS|CANCER OF OTHER URINARY ORGANS
C0346890|T047|34|CCS_10|MALIGNANT NEOPLASM OF OTHER URINARY ORGANS |CANCER OF OTHER URINARY ORGANS
C0346890|T047|34|CCS_10|MALIGNANT NEOPLASM OF OTHER URINARY ORGANS|CANCER OF OTHER URINARY ORGANS
C0700101|T047||CCS_10|URETHRAL CARCINOMA
C0700101|T047||CCS_10|CARCINOMA OF URETHRA 
C0700101|T047||CCS_10|URETHRAL CARCINOMA 
C0700101|T047||CCS_10|CARCINOMA OF URETHRA
C0700101|T047||CCS_10|CANCERS, URETHRA
C0700101|T047||CCS_10|URETHRA CANCERS
C0700101|T047||CCS_10|CANCER, URETHRAL
C0700101|T047||CCS_10|CANCERS, URETHRAL
C0700101|T047||CCS_10|URETHRAL CANCERS
C0700101|T047||CCS_10|CARCINOMA;URETHRA
C0700101|T047||CCS_10|CANCER, URETHRA
C0700101|T047||CCS_10|URETHRAL CANCER
C0700101|T047||CCS_10|URETHRA CANCER
C0700101|T047||CCS_10|URETHRAL CANCER NOS
C0700101|T047||CCS_10|CANCER OF THE URETHRA
C0700101|T047||CCS_10|CA - CANCER OF URETHRA
C0700101|T047||CCS_10|URETHRAL CA
C0700101|T047||CCS_10|URETHRA CARCINOMA
C0700101|T047||CCS_10|CARCINOMA OF THE URETHRA
C0700101|T047||CCS_10|CANCER OF URETHRA
C0153619|T047||CCS_10|MALIGNANT NEOPLASM OF URETER
C0153619|T047||CCS_10|URETER, CANCER OF
C0153619|T047||CCS_10|MALIGNANT NEOPLASM OF URETER 
C0153619|T047||CCS_10|URETER CANCERS
C0153619|T047||CCS_10|CANCER, URETERAL
C0153619|T047||CCS_10|CANCERS, URETERAL
C0153619|T047||CCS_10|URETERAL CANCERS
C0153619|T047||CCS_10|MALIGNANT TUMOR OF URETER
C0153619|T047||CCS_10|URETERAL CANCER
C0153619|T047||CCS_10|MALIGN NEOPL URETER
C0153619|T047||CCS_10|MALIGNANT TUMOUR OF URETER 
C0153619|T047||CCS_10|MALIGNANT TUMOUR OF URETER
C0153619|T047||CCS_10|URETERS--CANCER
C0153619|T047||CCS_10|URETER CANCER
C0153619|T047||CCS_10|URETERIC CANCER
C0153619|T047||CCS_10|URETERIC CANCER NOS
C0153619|T047||CCS_10|CANCER OF THE URETER
C0153619|T047||CCS_10|URETER CA
C0153619|T047||CCS_10|CANCER OF URETER
C0153619|T047||CCS_10|MALIGNANT TUMOR OF URETER 
C0153619|T047||CCS_10|MALIGNANT NEOPLASM OF THE URETER
C0153619|T047||CCS_10|MALIGNANT TUMOR OF THE URETER
C0153619|T047||CCS_10|MALIGNANT URETER NEOPLASM
C0153619|T047||CCS_10|MALIGNANT URETER TUMOR
C0153619|T047||CCS_10|MALIGNANT URETERAL NEOPLASM
C0153619|T047||CCS_10|MALIGNANT URETERAL TUMOR
C0153619|T047||CCS_10|NEOPLASM MALIG;URETER
C0153619|T047||CCS_10|MALIGNANT NEOSPLASM OF THE URETER
C0153618|T047||CCS_10|MALIGNANT NEOPLASM OF RENAL PELVIS
C0153618|T047||CCS_10|MALIGNANT NEOPLASM OF RENAL PELVIS 
C0153618|T047||CCS_10|MALIGNANT TUMOR OF RENAL PELVIS
C0153618|T047||CCS_10|MALIG NEO RENAL PELVIS
C0153618|T047||CCS_10|MALIGNANT NEOPLASM OF RENAL PELVIS NOS
C0153618|T047||CCS_10|MALIGNANT NEOPLASM OF RENAL PELVIS NOS 
C0153618|T047||CCS_10|RENAL PELVIS CANCER NOS
C0153618|T047||CCS_10|MALIGNANT TUMOUR OF RENAL PELVIS
C0153618|T047||CCS_10|MALIGNANT TUMOR OF RENAL PELVIS 
C0153618|T047||CCS_10|MALIGNANT NEOPLASM OF THE RENAL PELVIS
C0153618|T047||CCS_10|MALIGNANT RENAL PELVIS NEOPLASM
C0153618|T047||CCS_10|MALIGNANT RENAL PELVIS TUMOR
C0153618|T047||CCS_10|MALIGNANT TUMOR OF THE RENAL PELVIS
C0153622|T047||CCS_10|MALIGNANT NEOPLASM OF OTHER SPECIFIED SITES OF URINARY ORGANS
C0153622|T047||CCS_10|MAL NEO URINARY NEC
C0494158|T047||CCS_10|MALIGNANT NEOPLASM OF KIDNEY, EXCEPT RENAL PELVIS
C0494158|T047||CCS_10|MALIG NEOPL KIDNEY
C0494158|T047||CCS_10|MALIGNANT NEOPLASM OF KIDNEY, EXCEPT PELVIS
C0494158|T047||CCS_10|MALIGNANT NEOPLASM OF KIDNEY, EXCL PELVIS
C0494158|T047||CCS_10|MALIGNANT NEOPLASM OF KIDNEY, EXCLUDING PELVIS
C0494158|T047||CCS_10|MALIGNANT NEOPLASM OF KIDNEY EXCEPT PELVIS
C0494158|T047||CCS_10|MALIGNANT KIDNEY NEOPLASM EXCEPT PELVIS
C0600079|T047||CCS_10|CARCINOMA OF URETER
C0600079|T047||CCS_10|CARCINOMA OF URETER 
C0600079|T047||CCS_10|URETER CARCINOMA
C0600079|T047||CCS_10|CARCINOMA;URETER
C0600079|T047||CCS_10|URETERAL CARCINOMA
C0600079|T047||CCS_10|CARCINOMA OF THE URETER
C0751571|T047||CCS_10|MALIGNANT URINARY SYSTEM NEOPLASM
C0751571|T047||CCS_10|MALIGNANT URINARY TRACT NEOPLASM
C0751571|T047||CCS_10|MALIGNANT NEOPLASM OF URINARY SYSTEM
C0751571|T047||CCS_10|MALIGNANT NEOPLASM OF URINARY ORGANS 
C0751571|T047||CCS_10|MALIGNANT NEOPLASM OF URINARY ORGANS
C0751571|T047||CCS_10|MALIGNANT NEOPLASMS OF URINARY TRACT
C0751571|T047||CCS_10|MALIGNANT TUMOR OF URINARY TRACT PROPER 
C0751571|T047||CCS_10|MALIGNANT TUMOR OF URINARY TRACT
C0751571|T047||CCS_10|MALIGNANT TUMOUR OF URINARY TRACT
C0751571|T047||CCS_10|MALIGNANT TUMOR OF URINARY TRACT PROPER
C0751571|T047||CCS_10|MALIGNANT TUMOR OF URINARY TRACT 
C0751571|T047||CCS_10|MALIGNANT TUMOUR OF URINARY TRACT PROPER
C0751571|T047||CCS_10|CANCERS, URINARY TRACT
C0751571|T047||CCS_10|URINARY TRACT CANCERS
C0751571|T047||CCS_10|CANCER, UROLOGIC
C0751571|T047||CCS_10|CANCERS, UROLOGIC
C0751571|T047||CCS_10|UROLOGIC CANCERS
C0751571|T047||CCS_10|CANCER, UROLOGICAL
C0751571|T047||CCS_10|CANCERS, UROLOGICAL
C0751571|T047||CCS_10|UROLOGICAL CANCERS
C0751571|T047||CCS_10|MALIGNANT NEOPLASM OF URINARY SYSTEM NOS
C0751571|T047||CCS_10|CANCER, URINARY TRACT
C0751571|T047||CCS_10|MALIGNANT NEOPLASMS OF URINARY TRACT (C64-C68)
C0751571|T047||CCS_10|[X]MALIGNANT NEOPLASM OF URINARY TRACT 
C0751571|T047||CCS_10|[X]MALIGNANT NEOPLASM OF URINARY TRACT
C0751571|T047||CCS_10|MALIGNANT NEOPLASM OF URINARY TRACT PROPER 
C0751571|T047||CCS_10|MALIGNANT NEOPLASM OF URINARY TRACT PROPER
C0751571|T047||CCS_10|MALIGNANT NEOPLASM URINARY SYSTEM
C0751571|T047||CCS_10|URINARY NEOPLASM MALIGNANT OF TRACT PROPER
C0751571|T047||CCS_10|MALIGNANT NEOPLASM OF URINARY SYSTEM 
C0751571|T047||CCS_10|UROTHELIAL/BLADDER CANCER, NOS
C0751571|T047||CCS_10|UROTHELIAL TRACT/BLADDER CANCER, NOS
C0751571|T047||CCS_10|MALIGNANT URINARY TRACT NEOPLASM NOS
C0751571|T047||CCS_10|CANCER OF THE URINARY TRACT
C0751571|T047||CCS_10|UROLOGICAL CANCER
C0751571|T047||CCS_10|UROLOGIC CANCER
C0751571|T047||CCS_10|URINARY TRACT CANCER
C0751571|T047||CCS_10|MALIGNANT NEOPLASM OF URINARY SYSTEM, NOS
C0751571|T047||CCS_10|CANCER OF URINARY TRACT
C0751571|T047||CCS_10|NEOPLASM MALIG;UROLOGICAL
C0751571|T047||CCS_10|MALIGNANT NEOSPLASM OF THE UROLOGICAL SYSTEM
C1276598|T047||CCS_10|TA: NONINVASIVE PAPILLARY CARCINOMA (URINARY TRACT) 
C1276598|T047||CCS_10|TA: NONINVASIVE PAPILLARY CARCINOMA (URINARY TRACT)
C1276598|T047||CCS_10|TA: NONINVASIVE PAPILLARY CARCINOMA (URINARY TRACT) (TUMOR STAGING)
C0023418|T047||CCS_10|LEUKEMIAS
C0023418|T047||CCS_10|LEUKEMIA
C0023418|T047||CCS_10|LEUKEMIA OF UNSPECIFIED CELL TYPE
C0023418|T047||CCS_10|LEUKAEMIA
C0023418|T047||CCS_10|LEUKAEMIA OF UNSPECIFIED CELL TYPE
C0023418|T047||CCS_10|LEUKAEMIA, UNSPECIFIED
C0023418|T047||CCS_10|LEUKEMIA, UNSPECIFIED
C0023418|T047||CCS_10|LEUKEMIA, DISEASE
C0023418|T047||CCS_10|LEUKAEMIA, DISEASE
C0023418|T047||CCS_10|LEUKEMIA 
C0023418|T047||CCS_10|LEUKAEMIA, NO ICD-O SUBTYPE
C0023418|T047||CCS_10|LEUKEMIA, NO ICD-O SUBTYPE
C0023418|T047||CCS_10|LEUKAEMIAS
C0023418|T047||CCS_10|LEUKEMIA NOS
C0023418|T047||CCS_10|LEUKEMIA [DISEASE/FINDING]
C0023418|T047||CCS_10|LEUKAEMIA OF UNSPECIFIED CELL TYPE 
C0023418|T047||CCS_10|[M]LEUKEMIA NOS
C0023418|T047||CCS_10|LEUKEMIA 
C0023418|T047||CCS_10|[M]LEUKAEMIA NOS
C0023418|T047||CCS_10|LEUKEMIA OF UNSPECIFIED CELL TYPE 
C0023418|T047||CCS_10|[M]LEUKEMIA UNSPECIFIED, NOS
C0023418|T047||CCS_10|[M]LEUKEMIA UNSPECIFIED, NOS (MORPHOLOGIC ABNORMALITY)
C0023418|T047||CCS_10|[M]LEUKAEMIA NOS 
C0023418|T047||CCS_10|LEUKEMIA NOS 
C0023418|T047||CCS_10|[M]LEUKEMIA NOS (MORPHOLOGIC ABNORMALITY)
C0023418|T047||CCS_10|[M]LEUKAEMIA UNSPECIFIED, NOS
C0023418|T047||CCS_10|LEUKAEMIA NOS
C0023418|T047||CCS_10|[M]LEUKAEMIAS UNSPECIFIED
C0023418|T047||CCS_10|[M]LEUKEMIAS UNSPECIFIED (MORPHOLOGIC ABNORMALITY)
C0023418|T047||CCS_10|[M]LEUKEMIAS UNSPECIFIED
C0023418|T047||CCS_10|LEUKEMIA, NO ICD-O SUBTYPE (MORPHOLOGIC ABNORMALITY)
C0023418|T047||CCS_10|LEUKEMIA, NO INTERNATIONAL CLASSIFICATION OF DISEASES FOR ONCOLOGY SUBTYPE (MORPHOLOGIC ABNORMALITY)
C0023418|T047||CCS_10|LEUKEMIA, NO INTERNATIONAL CLASSIFICATION OF DISEASES FOR ONCOLOGY SUBTYPE
C0023418|T047||CCS_10|LEUKEMIA, NOS
C0023418|T047||CCS_10|LEUKEMIA, MALIGNANT
C0023418|T047||CCS_10|-- LEUKEMIA
C0023418|T047||CCS_10|BLOOD (LEUKEMIA)
C0023418|T047||CCS_10|LEUKEMIAS, GENERAL
C0023418|T047||CCS_10|LEUKEMIA UNSPECIFIED
C0023418|T047||CCS_10|UNSPECIFIED LEUKEMIA WITHOUT MENTION OF REMISSION
C0023418|T047||CCS_10|UNSPECIFIED LEUKAEMIA WITHOUT MENTION OF REMISSION
C0023418|T047||CCS_10|LEUKAEMIA UNSPECIFIED
C0023418|T047||CCS_10|UNSPECIFIED LEUKAEMIA
C0023418|T047||CCS_10|UNSPECIFIED LEUKEMIA
C0023418|T047||CCS_10|LEUKAEMIA MORPHOLOGY
C0023418|T047||CCS_10|LEUKEMIA MORPHOLOGY
C0023418|T047||CCS_10|CHRONIC LEUKAEMIA [OBS]
C0023418|T047||CCS_10|CHRONIC LEUKEMIA [OBS]
C0023418|T047||CCS_10|LEUKEMIA, DISEASE 
C0023418|T047||CCS_10|ALEUKAEMIC LEUKAEMIA [OBS]
C0023418|T047||CCS_10|ALEUKEMIC LEUKEMIA [OBS]
C0023418|T047||CCS_10|SUBACUTE LEUKAEMIA [OBS]
C0023418|T047||CCS_10|SUBACUTE LEUKEMIA [OBS]
C0023418|T047||CCS_10|LEUKAEMIA, NOS
C0023418|T047||CCS_10|LEUKAEMIA, NOS, WITHOUT MENTION OF REMISSION
C0023418|T047||CCS_10|LEUKEMIA, NOS, WITHOUT MENTION OF REMISSION
C0023418|T047||CCS_10|LEUKEMIA, MORPHOLOGY (MORPHOLOGIC ABNORMALITY)
C0026764|T047||CCS_10|MULTIPLE MYELOMA
C0026764|T047||CCS_10|MULTIPLE MYELOMAS
C0026764|T047||CCS_10|MYELOMA, PLASMA CELL
C0026764|T047||CCS_10|MYELOMAS, MULTIPLE
C0026764|T047||CCS_10|PLASMA CELL MYELOMA
C0026764|T047||CCS_10|MYELOMATOSIS
C0026764|T047||CCS_10|MYELOMAS, PLASMA-CELL
C0026764|T047||CCS_10|PLASMA-CELL MYELOMA
C0026764|T047||CCS_10|PLASMA-CELL MYELOMAS
C0026764|T047||CCS_10|MULTIPLE MYELOMA / PLASMA CELL NEOPLASM
C0026764|T047||CCS_10|MYELOMA, MULTIPLE
C0026764|T047||CCS_10|MYELOMA
C0026764|T047||CCS_10|MULTIPLE MYELOMA 
C0026764|T047||CCS_10|MULTIPLE MYELOMA, NO ICD-O SUBTYPE
C0026764|T047||CCS_10|CELL MYELOMA, PLASMA
C0026764|T047||CCS_10|CELL MYELOMAS, PLASMA
C0026764|T047||CCS_10|PLASMA CELL MYELOMAS
C0026764|T047||CCS_10|MYELOMAS, PLASMA CELL
C0026764|T047||CCS_10|KAHLER'S DISEASE
C0026764|T047||CCS_10|MULTIPLE MYELOMA NOS
C0026764|T047||CCS_10|MULTIPLE MYELOMA [DISEASE/FINDING]
C0026764|T047||CCS_10|MYELOMA, PLASMA-CELL
C0026764|T047||CCS_10|MYELOMATOSES
C0026764|T047||CCS_10|DISEASE, KAHLER
C0026764|T047||CCS_10|MYELOMA-MULTIPLES
C0026764|T047||CCS_10|MYELOMA MULTIPLE
C0026764|T047||CCS_10|MYELOMA;MULTIPLE
C0026764|T047||CCS_10|MYELOMA-MULTIPLE
C0026764|T047||CCS_10|KAHLER DISEASE
C0026764|T047||CCS_10|MULTIPLE MYELOMA MYELOMATOSIS
C0026764|T047||CCS_10|MYELOMA 
C0026764|T047||CCS_10|MULTIPLE MYELOMA 
C0026764|T047||CCS_10|MULTIPLE MYELOMA, NO INTERNATIONAL CLASSIFICATION OF DISEASES FOR ONCOLOGY SUBTYPE (MORPHOLOGIC ABNORMALITY)
C0026764|T047||CCS_10|MULTIPLE MYELOMA, NO ICD-O SUBTYPE (MORPHOLOGIC ABNORMALITY)
C0026764|T047||CCS_10|MULTIPLE MYELOMA, NO INTERNATIONAL CLASSIFICATION OF DISEASES FOR ONCOLOGY SUBTYPE
C0026764|T047||CCS_10|MYELOMA, PLASMA CELL, MALIGNANT
C0026764|T047||CCS_10|MYELOMA, NOS
C0026764|T047||CCS_10|[M]PLASMA CELL MYELOMA
C0026764|T047||CCS_10|PERIPHERAL PLASMA CELL MYELOMA
C0026764|T047||CCS_10|MYELOMATOSIS MULTIPLE
C0026764|T047||CCS_10|PLASMACYTIC MYELOMA
C0026764|T047||CCS_10|PLASMA CELL NEOPLASM
C0026764|T047||CCS_10|NEOPLASM, PLASMA CELL
C0026764|T047||CCS_10|MULTIPLE MYELOMA AND OTHER PLASMA CELL NEOPLASMS
C0026764|T047||CCS_10|PLASMA CELL NEOPLASMS
C0026764|T047||CCS_10|MYELOMATA; MULTIPLE
C0026764|T047||CCS_10|MULTIPLE MYELOMA (CLINICAL)
C0026764|T047||CCS_10|MULTIPLE MYELOMA, MORPHOLOGY (MORPHOLOGIC ABNORMALITY)
C0019829|T047|37|CCS_10|DISEASE, HODGKIN|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN DISEASE|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S DISEASE|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|LYMPHOGRANULOMAS, MALIGNANT|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|MALIGNANT LYMPHOGRANULOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|MALIGNANT LYMPHOGRANULOMAS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|DISEASE, HODGKIN'S|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|DISEASE, HODGKINS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S DISEASE, UNSPECIFIED|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN LYMPHOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN DIS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKINS DIS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S LYMPHOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|LYMPHOMA, HODGKIN'S|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|LYMPHOMA, HODGKIN|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKINS LYMPHOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S GRANULOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S SARCOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|LYMPHOGRANULOMATOSIS (MALIGNANT)|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S PARAGRANULOMA, NOS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S DISEASE, NOS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN LYMPHOMA, NO ICD-O SUBTYPE|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S PARAGRANULOMA -RETIRED-|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|LYMPHOMAS HODGKIN'S DISEASE|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGINS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN SARCOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN GRANULOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN LYMPHOMA, UNSPECIFIED|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN DISEASE [DISEASE/FINDING]|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|GRANULOMA, HODGKINS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|GRANULOMA, HODGKIN|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKINS DISEASE|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|LYMPHOGRANULOMA, MALIGNANT|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|GRANULOMA, HODGKIN'S|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|GRANULOMA, MALIGNANT|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|DISEASE;HODGKINS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|LYMPHOMA;HODGKINS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|SARCOMA;HODGKINS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKINS GRANULOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|MALIGNANT GRANULOMAS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|MALIGNANT GRANULOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|LYMPHOGRANULOMATOSIS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S PARAGRANULOMA (MORPHOLOGIC ABNORMALITY)|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|[M]HODGKIN'S DISEASE NOS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S DISEASE NOS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S SARCOMA OF UNSPECIFIED SITE|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S PARAGRANULOMA OF UNSPECIFIED SITE|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S SARCOMA NOS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S GRANULOMA NOS |HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|[M]HODGKIN'S PARAGRANULOMA (MORPHOLOGIC ABNORMALITY)|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|[M]HODGKIN'S DISEASE NOS (MORPHOLOGIC ABNORMALITY)|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|[M]HODGKIN'S PARAGRANULOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|[M]LYMPHOGRANULOMA, MALIGNANT (MORPHOLOGIC ABNORMALITY)|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S PARAGRANULOMA |HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|[M]HODGKIN'S DISEASE NOS (& [LYMPHOGRANULOMA MALIGNANT])|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S DISEASE NOS, UNSPECIFIED SITE |HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S PARAGRANULOMA NOS |HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S GRANULOMA OF UNSPECIFIED SITE|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S SARCOMA NOS |HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S DISEASE NOS, UNSPECIFIED SITE|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S DISEASE NOS |HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S PARAGRANULOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|[M]LYMPHOGRANULOMA, MALIGNANT|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S PARAGRANULOMA OF UNSPECIFIED SITE |HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|[M]HODGKIN'S DISEASE NOS (& [LYMPHOGRANULOMA MALIGNANT]) |HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S PARAGRANULOMA NOS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S GRANULOMA NOS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S SARCOMA OF UNSPECIFIED SITE |HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|[M]HODGKIN'S DISEASE NOS |HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S DISEASE |HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S GRANULOMA OF UNSPECIFIED SITE |HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN LYMPHOMA, NO ICD-O SUBTYPE (MORPHOLOGIC ABNORMALITY)|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN LYMPHOMA, NO INTERNATIONAL CLASSIFICATION OF DISEASES FOR ONCOLOGY SUBTYPE|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN LYMPHOMA, NO INTERNATIONAL CLASSIFICATION OF DISEASES FOR ONCOLOGY SUBTYPE (MORPHOLOGIC ABNORMALITY)|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN LYMPHOMA, NOS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN DISEASE |HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN DISEASE SARCOMA |HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN DISEASE SARCOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN DISEASE GRANULOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN DISEASE GRANULOMA |HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN DISEASE PARAGRANULOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN DISEASE PARAGRANULOMA |HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|[M]HODGKIN'S DISEASE|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|[M]HODGKIN'S GRANULOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|[M]HODGKIN'S SARCOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|CHL|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|LYMPHOMA, HODGKIN, CLASSIC|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|LYMPHOMA, HODGKINS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S DISEASE, UNSPECIFIED TYPE|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN`S DISEASE|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|MALIGNANT HODGKIN'S LYMPHOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|MALIGNANT LYMPHOMA, HODGKIN'S|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HD - HODGKIN'S DISEASE|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN GRANULOMA [OBS] (MORPHOLOGIC ABNORMALITY)|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN GRANULOMA [OBS]|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN PARAGRANULOMA [OBS]|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN PARAGRANULOMA, NODULAR [OBS]|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN SARCOMA [OBS] (MORPHOLOGIC ABNORMALITY)|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN SARCOMA [OBS]|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S DISEASE (CLINICAL)|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S GRANULOMA (CLINICAL)|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S GRANULOMA |HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S PARAGRANULOMA (CLINICAL)|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S SARCOMA (CLINICAL)|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S SARCOMA |HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN; GRANULOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN; LYMPHOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN; PARAGRANULOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN; SARCOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|DISEASE; HODGKIN|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|GRANULOMA; HODGKIN|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|GRANULOMA; MALIGNANT|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|LYMPHOMA; HODGKIN|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|MALIGNANT; GRANULOMA|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|PARAGRANULOMA; HODGKIN|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|SARCOMA; HODGKIN|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S PARAGRANULOMA, NODULAR|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKIN'S LYMPHOMA NOS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|MALIGNANT LYMPHOGRANULOMATOSIS|HODGKIN`S DISEASE
C0019829|T047|37|CCS_10|HODGKINS SARCOMA|HODGKIN`S DISEASE
C0023448|T047||CCS_10|LYMPHOID LEUKEMIAS
C0023448|T047||CCS_10|LEUKEMIAS, LYMPHOCYTIC
C0023448|T047||CCS_10|LEUKEMIAS, LYMPHOID
C0023448|T047||CCS_10|LYMPHOCYTIC LEUKEMIAS
C0023448|T047||CCS_10|LEUKEMIA LYMPHATIC
C0023448|T047||CCS_10|LEUKEMIA LYMPHOCYTIC
C0023448|T047||CCS_10|LEUKEMIA LYMPHOID
C0023448|T047||CCS_10|LYMPHOID LEUKEMIA
C0023448|T047||CCS_10|LYMPHOCYTIC LEUKEMIA
C0023448|T047||CCS_10|LYMPHOID LEUKAEMIA
C0023448|T047||CCS_10|LYMPHOID LEUKAEMIA, UNSPECIFIED
C0023448|T047||CCS_10|LYMPHOID LEUKEMIA, UNSPECIFIED
C0023448|T047||CCS_10|LEUKEMIA, LYMPHOID
C0023448|T047||CCS_10|LYMPHATIC LEUKEMIA
C0023448|T047||CCS_10|LYMPHOBLASTIC LEUKEMIA
C0023448|T047||CCS_10|LYMPHOGENOUS LEUKEMIA
C0023448|T047||CCS_10|LYMPHOCYTIC LEUKEMIA 
C0023448|T047||CCS_10|LYMPHOID LEUKAEMIA, NO ICD-O SUBTYPE
C0023448|T047||CCS_10|LYMPHOID LEUKEMIA, NO ICD-O SUBTYPE
C0023448|T047||CCS_10|LYMPHOCYTIC LEUKAEMIA
C0023448|T047||CCS_10|LYMPHOID LEUKEMIA NOS
C0023448|T047||CCS_10|LEUKEMIA, LYMPHOCYTIC
C0023448|T047||CCS_10|LEUKEMIA, LYMPHOID [DISEASE/FINDING]
C0023448|T047||CCS_10|[M]LYMPHOID LEUKAEMIAS
C0023448|T047||CCS_10|[M]LYMPHOID LEUKEMIAS
C0023448|T047||CCS_10|LYMPHOID LEUKEMIA, DISEASE 
C0023448|T047||CCS_10|LYMPHOID LEUKAEMIA NOS
C0023448|T047||CCS_10|LYMPHOID LEUKEMIA NOS 
C0023448|T047||CCS_10|[M]LYMPHOID LEUKEMIAS (MORPHOLOGIC ABNORMALITY)
C0023448|T047||CCS_10|LYMPHOID LEUKEMIA, NO ICD-O SUBTYPE (MORPHOLOGIC ABNORMALITY)
C0023448|T047||CCS_10|LYMPHOID LEUKEMIA, NO INTERNATIONAL CLASSIFICATION OF DISEASES FOR ONCOLOGY SUBTYPE (MORPHOLOGIC ABNORMALITY)
C0023448|T047||CCS_10|LYMPHOID LEUKEMIA, NO INTERNATIONAL CLASSIFICATION OF DISEASES FOR ONCOLOGY SUBTYPE
C0023448|T047||CCS_10|LEUKEMIA, LYMPHOCYTIC, MALIGNANT
C0023448|T047||CCS_10|[M]LYMPHOID LEUKEMIA NOS
C0023448|T047||CCS_10|[M]LYMPHOID LEUKAEMIA NOS
C0023448|T047||CCS_10|LEUKAEMIA LYMPHOCYTIC
C0023448|T047||CCS_10|LEUKAEMIA LYMPHOID
C0023448|T047||CCS_10|UNSPECIFIED LYMPHOID LEUKEMIA
C0023448|T047||CCS_10|LYMPHOBLASTIC LEUKEMIA NOS
C0023448|T047||CCS_10|LYMPHATIC LEUKAEMIA
C0023448|T047||CCS_10|LEUKAEMIA LYMPHATIC
C0023448|T047||CCS_10|LYMPHOBLASTIC LEUKAEMIA NOS
C0023448|T047||CCS_10|UNSPECIFIED LYMPHOID LEUKAEMIA
C0023448|T047||CCS_10|ALEUKAEMIC LYMPHATIC LEUKAEMIA [OBS]
C0023448|T047||CCS_10|ALEUKAEMIC LYMPHOCYTIC LEUKAEMIA [OBS]
C0023448|T047||CCS_10|ALEUKAEMIC LYMPHOID LEUKAEMIA [OBS]
C0023448|T047||CCS_10|ALEUKEMIC LYMPHATIC LEUKEMIA [OBS]
C0023448|T047||CCS_10|ALEUKEMIC LYMPHOCYTIC LEUKEMIA [OBS]
C0023448|T047||CCS_10|ALEUKEMIC LYMPHOID LEUKEMIA [OBS]
C0023448|T047||CCS_10|LYMPHOID LEUKEMIA 
C0023448|T047||CCS_10|LYMPHOSARCOMA CELL LEUKAEMIA [OBS]
C0023448|T047||CCS_10|LYMPHOSARCOMA CELL LEUKEMIA [OBS]
C0023448|T047||CCS_10|LEUKEMIA; LYMPHATIC
C0023448|T047||CCS_10|LEUKEMIA; LYMPHOBLASTIC
C0023448|T047||CCS_10|LYMPHATIC; LEUKEMIA
C0023448|T047||CCS_10|LYMPHOBLASTIC; LEUKEMIA
C0023448|T047||CCS_10|LYMPHATIC LEUKEMIA, NOS
C0023448|T047||CCS_10|LYMPHOCYTIC LEUKEMIA, NOS
C0023448|T047||CCS_10|LYMPHOID LEUKEMIA, NOS
C0023448|T047||CCS_10|LYMPHOID LEUKEMIA, DISEASE [AMBIGUOUS]
C0598894|T047||CCS_10|MONOCYTIC LEUKEMIA
C0598894|T047||CCS_10|LEUKEMIA MONOCYTIC
C0598894|T047||CCS_10|MONOCYTIC LEUKAEMIA
C0598894|T047||CCS_10|MONOCYTIC LEUKAEMIA, UNSPECIFIED
C0598894|T047||CCS_10|MONOCYTIC LEUKEMIA, UNSPECIFIED
C0598894|T047||CCS_10|SCHILLING'S LEUKEMIA
C0598894|T047||CCS_10|MONOCYTIC LEUKEMIA 
C0598894|T047||CCS_10|MONOCYTIC LEUKAEMIA -RETIRED-
C0598894|T047||CCS_10|MONOCYTIC LEUKEMIA -RETIRED-
C0598894|T047||CCS_10|MONOCYTOID LEUKEMIA
C0598894|T047||CCS_10|MONOCYTIC LEUKEMIA, UNSPECIFIED NOS
C0598894|T047||CCS_10|MONOCYTIC LEUKEMIA (MORPHOLOGIC ABNORMALITY)
C0598894|T047||CCS_10|MONOCYTIC LEUKEMIA NOS
C0598894|T047||CCS_10|[M]MONOCYTIC LEUKAEMIAS
C0598894|T047||CCS_10|MONOCYTIC LEUKEMIA 
C0598894|T047||CCS_10|[M]MONOCYTIC LEUKEMIAS
C0598894|T047||CCS_10|[M]MONOCYTIC LEUKAEMIA NOS
C0598894|T047||CCS_10|[M]MONOCYTIC LEUKEMIAS (MORPHOLOGIC ABNORMALITY)
C0598894|T047||CCS_10|MONOCYTIC LEUKEMIA NOS 
C0598894|T047||CCS_10|[M]MONOCYTIC LEUKAEMIA NOS 
C0598894|T047||CCS_10|MONOCYTIC LEUKAEMIA NOS
C0598894|T047||CCS_10|[M]MONOCYTIC LEUKEMIA NOS
C0598894|T047||CCS_10|LEUKAEMIA MONOCYTIC NOS
C0598894|T047||CCS_10|UNSPECIFIED MONOCYTIC LEUKEMIA
C0598894|T047||CCS_10|LEUKEMIA MONOCYTIC NOS
C0598894|T047||CCS_10|UNSPECIFIED MONOCYTIC LEUKAEMIA
C0598894|T047||CCS_10|LEUKAEMIA MONOCYTIC
C0598894|T047||CCS_10|SCHILLING-TYPE MONOCYTIC LEUKEMIA
C0598894|T047||CCS_10|SCHILLING-TYPE MONOCYTIC LEUKAEMIA
C0598894|T047||CCS_10|LEUKEMIA; MONOCYTIC
C0598894|T047||CCS_10|MONOCYTIC; LEUKEMIA
C0598894|T047||CCS_10|MONOCYTIC LEUKEMIA, NOS
C0023470|T047||CCS_10|MYELOID LEUKEMIAS
C0023470|T047||CCS_10|GRANULOCYTIC LEUKEMIAS
C0023470|T047||CCS_10|LEUKEMIA, MYELOID
C0023470|T047||CCS_10|LEUKEMIAS, GRANULOCYTIC
C0023470|T047||CCS_10|LEUKEMIAS, MYELOCYTIC
C0023470|T047||CCS_10|LEUKEMIAS, MYELOGENOUS
C0023470|T047||CCS_10|LEUKEMIAS, MYELOID
C0023470|T047||CCS_10|MYELOCYTIC LEUKEMIAS
C0023470|T047||CCS_10|MYELOGENOUS LEUKEMIAS
C0023470|T047||CCS_10|MYELOID LEUKEMIA
C0023470|T047||CCS_10|LEUKEMIA GRANULOCYTIC
C0023470|T047||CCS_10|LEUKEMIA MYELOGENOUS
C0023470|T047||CCS_10|LEUKEMIA MYELOID
C0023470|T047||CCS_10|MYELOGENOUS LEUKEMIA
C0023470|T047||CCS_10|MYELOID LEUKAEMIA
C0023470|T047||CCS_10|MYELOID LEUKAEMIA, UNSPECIFIED
C0023470|T047||CCS_10|MYELOID LEUKEMIA, UNSPECIFIED
C0023470|T047||CCS_10|MYELOCYTIC LEUKEMIA
C0023470|T047||CCS_10|MYELOSIS
C0023470|T047||CCS_10|GRANULOCYTIC LEUKEMIA
C0023470|T047||CCS_10|MYELOID GRANULOCYTIC LEUKEMIA
C0023470|T047||CCS_10|MYELOGENOUS LEUKEMIA 
C0023470|T047||CCS_10|MYELOID LEUKEMIA - CATEGORY
C0023470|T047||CCS_10|MYELOID LEUKAEMIA - CATEGORY
C0023470|T047||CCS_10|LEUKEMIC GRANULOCYTIC
C0023470|T047||CCS_10|MYELOID LEUKEMIA, UNSPECIFIED NOS
C0023470|T047||CCS_10|LEUKEMIA, GRANULOCYTIC
C0023470|T047||CCS_10|LEUKEMIA, MYELOCYTIC
C0023470|T047||CCS_10|LEUKEMIA, MYELOGENOUS
C0023470|T047||CCS_10|LEUKEMIA, MYELOID [DISEASE/FINDING]
C0023470|T047||CCS_10|MYELOID LEUKEMIA NOS 
C0023470|T047||CCS_10|MYELOID LEUKAEMIA NOS
C0023470|T047||CCS_10|MYELOID LEUKEMIA NOS
C0023470|T047||CCS_10|[M]MYELOID LEUKEMIAS (MORPHOLOGIC ABNORMALITY)
C0023470|T047||CCS_10|[M]MYELOID LEUKAEMIAS
C0023470|T047||CCS_10|MYELOID LEUKEMIA, DISEASE 
C0023470|T047||CCS_10|[M]MYELOID LEUKEMIAS
C0023470|T047||CCS_10|GRANULOCYTIC LEUKEMIA 
C0023470|T047||CCS_10|MYELOID LEUKEMIA, NO ICD-O SUBTYPE (MORPHOLOGIC ABNORMALITY)
C0023470|T047||CCS_10|MYELOID LEUKEMIA, NO INTERNATIONAL CLASSIFICATION OF DISEASES FOR ONCOLOGY SUBTYPE
C0023470|T047||CCS_10|MYELOID LEUKEMIA, NO INTERNATIONAL CLASSIFICATION OF DISEASES FOR ONCOLOGY SUBTYPE (MORPHOLOGIC ABNORMALITY)
C0023470|T047||CCS_10|LEUKEMIA, GRANULOCYTIC, MALIGNANT
C0023470|T047||CCS_10|[M]MYELOID LEUKAEMIA NOS
C0023470|T047||CCS_10|[M]MYELOID LEUKEMIA NOS
C0023470|T047||CCS_10|NON-LYMPHOBLASTIC LEUKEMIA
C0023470|T047||CCS_10|NON-LYMPHOCYTIC LEUKEMIA
C0023470|T047||CCS_10|LEUKEMIA GRANULOCYTIC NOS
C0023470|T047||CCS_10|NON-LYMPHOBLASTIC LEUKEMIA NOS
C0023470|T047||CCS_10|UNSPECIFIED MYELOID LEUKEMIA
C0023470|T047||CCS_10|LEUKAEMIA GRANULOCYTIC
C0023470|T047||CCS_10|MYELOCYTIC LEUKAEMIA
C0023470|T047||CCS_10|UNSPECIFIED MYELOID LEUKAEMIA
C0023470|T047||CCS_10|LEUKAEMIA MYELOGENOUS
C0023470|T047||CCS_10|LEUKAEMIA MYELOID
C0023470|T047||CCS_10|NON-LYMPHOBLASTIC LEUKAEMIA NOS
C0023470|T047||CCS_10|LEUKAEMIA GRANULOCYTIC NOS
C0023470|T047||CCS_10|GRANULOCYTIC LEUKAEMIA
C0023470|T047||CCS_10|ALEUKAEMIC MONOCYTIC LEUKAEMIA [OBS]
C0023470|T047||CCS_10|ALEUKEMIC MONOCYTIC LEUKEMIA [OBS]
C0023470|T047||CCS_10|MYELOGENOUS LEUKAEMIA
C0023470|T047||CCS_10|MYELOID LEUKAEMIA 
C0023470|T047||CCS_10|MYELOID LEUKEMIA 
C0023470|T047||CCS_10|MYELOID LEUKEMIA 
C0023470|T047||CCS_10|MYELOID LEUKEMIA - CATEGORY (MORPHOLOGIC ABNORMALITY)
C0023470|T047||CCS_10|NON-LYMPHOCYTIC LEUKAEMIA
C0023470|T047||CCS_10|GRANULOCYTIC; LEUKEMIA
C0023470|T047||CCS_10|LEUKEMIA; GRANULOCYTIC
C0023470|T047||CCS_10|LEUKEMIA; MYELOCYTIC
C0023470|T047||CCS_10|LEUKEMIA; MYELOID
C0023470|T047||CCS_10|MYELOCYTIC; LEUKEMIA
C0023470|T047||CCS_10|MYELOID; LEUKEMIA
C0023470|T047||CCS_10|GRANULOCYTIC LEUKEMIA, NOS
C0023470|T047||CCS_10|MYELOCYTIC LEUKEMIA, NOS
C0023470|T047||CCS_10|MYELOGENOUS LEUKEMIA, NOS
C0023470|T047||CCS_10|MYELOID LEUKEMIA, NOS
C0023470|T047||CCS_10|MYELOID LEUKAEMIA, NOS
C0023470|T047||CCS_10|MYELOID LEUKEMIA, DISEASE [AMBIGUOUS]
C0023470|T047||CCS_10|MYELOID LEUKEMIA, MORPHOLOGY (MORPHOLOGIC ABNORMALITY)
C0348394|T047||CCS_10|DIFFUSE NON-HODGKIN'S LYMPHOMA, UNSPECIFIED
C0348394|T047||CCS_10|DIFFUSE NON-HODGKIN'S LYMPHOMA
C0348394|T047||CCS_10|DIFFUSE NON-HODGKIN LYMPHOMA
C0348394|T047||CCS_10|NONFOLLICULAR LYMPHOMA
C0348394|T047||CCS_10|[X]DIFFUSE NON-HODGKIN'S LYMPHOMA, UNSPECIFIED 
C0348394|T047||CCS_10|[X]DIFFUSE NON-HODGKIN'S LYMPHOMA, UNSPECIFIED
C0348394|T047||CCS_10|DIFFUSE NON-HODGKIN'S LYMPHOMA 
C0024301|T047||CCS_10|BRILL SYMMERS DISEASE
C0024301|T047||CCS_10|FOLLICULAR LYMPHOMAS
C0024301|T047||CCS_10|FOLLICULAR LYMPHOMAS, GIANT
C0024301|T047||CCS_10|GIANT FOLLICULAR LYMPHOMAS
C0024301|T047||CCS_10|LYMPHOMA, FOLLICULAR
C0024301|T047||CCS_10|LYMPHOMAS, FOLLICULAR
C0024301|T047||CCS_10|LYMPHOMAS, GIANT FOLLICULAR
C0024301|T047||CCS_10|LYMPHOMAS, NODULAR
C0024301|T047||CCS_10|NODULAR LYMPHOMAS
C0024301|T047||CCS_10|DISEASE, BRILL-SYMMERS
C0024301|T047||CCS_10|NODULAR LYMPHOMA
C0024301|T047||CCS_10|FOLLICULAR [NODULAR] NON-HODGKIN'S LYMPHOMA
C0024301|T047||CCS_10|FOLLICULAR NON-HODGKIN'S LYMPHOMA, UNSPECIFIED
C0024301|T047||CCS_10|FOLLICULAR NON-HODGKIN LYMPHOMA
C0024301|T047||CCS_10|GIANT FOLLIC LYMPHOMA
C0024301|T047||CCS_10|FOLLIC LYMPHOMA
C0024301|T047||CCS_10|FOLLIC LYMPHOMA GIANT
C0024301|T047||CCS_10|LYMPHOMA FOLLIC
C0024301|T047||CCS_10|LYMPHOMA GIANT FOLLIC
C0024301|T047||CCS_10|BRILL SYMMERS DIS
C0024301|T047||CCS_10|FOLLICULAR LYMPHOMA
C0024301|T047||CCS_10|NODULAR MALIGNANT LYMPHOMA 
C0024301|T047||CCS_10|NODULAR MALIGNANT LYMPHOMA
C0024301|T047||CCS_10|MALIGNANT LYMPHOMA, CENTROBLASTIC-CENTROCYTIC, FOLLICULAR -RETIRED-
C0024301|T047||CCS_10|GIANT FOLLICULAR LYMPHOSARCOMA 
C0024301|T047||CCS_10|NODULAR LYMPHOSARCOMA
C0024301|T047||CCS_10|GIANT FOLLICULAR LYMPHOSARCOMA
C0024301|T047||CCS_10|NODULAR LYMPHOSARCOMA 
C0024301|T047||CCS_10|FOLLICULAR LYMPHOMA, UNSPECIFIED
C0024301|T047||CCS_10|LYMPHOMA, NODULAR
C0024301|T047||CCS_10|BRILL-SYMMERS DISEASE
C0024301|T047||CCS_10|LYMPHOMA, GIANT FOLLICULAR
C0024301|T047||CCS_10|LYMPHOMA, FOLLICULAR [DISEASE/FINDING]
C0024301|T047||CCS_10|FOLLICULAR LYMPHOMA, GIANT
C0024301|T047||CCS_10|GIANT FOLLICULAR LYMPHOMA
C0024301|T047||CCS_10|FOLLICULAR LYMPHOMA 
C0024301|T047||CCS_10|MALIGNANT NEOPLASM NODULAR LYMPHOMA FOLLICULAR
C0024301|T047||CCS_10|(NODULAR LYMPHOMA: BRILL-SYMMERS DISEASE) OR (RETICULOSARCOMA - FOLLICULAR OR NODULAR) 
C0024301|T047||CCS_10|NODULAR LYMPHOMA NOS 
C0024301|T047||CCS_10|FOLLICULAR LYMPHOMA NOS
C0024301|T047||CCS_10|FOLLICULAR LYMPHOMA: [NON-HODGKIN'S] OR [NOS] 
C0024301|T047||CCS_10|NODULAR LYMPHOMA (BRILL - SYMMERS DISEASE)
C0024301|T047||CCS_10|[M]MALIGNANT LYMPHOMA, CENTROBLASTIC-CENTROCYTIC, FOLLICULAR
C0024301|T047||CCS_10|(NODULAR LYMPHOMA: BRILL-SYMMERS DISEASE) OR (RETICULOSARCOMA - FOLLICULAR OR NODULAR)
C0024301|T047||CCS_10|NODULAR LYMPHOMA OF UNSPECIFIED SITE
C0024301|T047||CCS_10|[M]MALIGNANT LYMPHOMA, CENTROBLASTIC-CENTROCYTIC, FOLLICULAR (MORPHOLOGIC ABNORMALITY)
C0024301|T047||CCS_10|[M]MALIGNANT LYMPHOMA, NODULAR NOS (& [BRILL - SYMMERS' DISEASE])
C0024301|T047||CCS_10|[M]MALIGNANT LYMPHOMA, NODULAR NOS
C0024301|T047||CCS_10|[M]FOLLICULAR LYMPHOSARCOMA NOS
C0024301|T047||CCS_10|[M]MALIGNANT LYMPHOMA, NODULAR NOS (& [BRILL - SYMMERS' DISEASE]) 
C0024301|T047||CCS_10|[M]GIANT FOLLICULAR LYMPHOMA
C0024301|T047||CCS_10|NODULAR LYMPHOMA NOS
C0024301|T047||CCS_10|FOLLICULAR NON-HODGKIN'S LYMPHOMA
C0024301|T047||CCS_10|[M]BRILL - SYMMERS' DISEASE
C0024301|T047||CCS_10|FOLLICULAR LYMPHOMA: [NON-HODGKIN'S] OR [NOS]
C0024301|T047||CCS_10|MALIGNANT LYMPHOMA, CENTROBLASTIC-CENTROCYTIC, FOLLICULAR (MORPHOLOGIC ABNORMALITY)
C0024301|T047||CCS_10|NODULAR LYMPHOMA OF UNSPECIFIED SITE 
C0024301|T047||CCS_10|RETICULOSARCOMA - FOLLICULAR OR NODULAR
C0024301|T047||CCS_10|MALIGNANT LYMPHOMA, CENTROBLASTIC-CENTROCYTIC, FOLLICULAR
C0024301|T047||CCS_10|[M]MALIGNANT LYMPHOMA, NODULAR NOS (MORPHOLOGIC ABNORMALITY)
C0024301|T047||CCS_10|[M]NODULAR LYMPHOSARCOMA NOS
C0024301|T047||CCS_10|FOLLICULAR MALIGNANT LYMPHOMA - CENTROBLASTIC-CENTROCYTIC
C0024301|T047||CCS_10|MALIGNANT NEOPLASM LYMPHOMA FOLLICULAR - CENTROBLASTIC-CENTROCYTIC
C0024301|T047||CCS_10|MALIGNANT NEOPLASM LYMPHOMA B-CELL LOW GRADE FOLLICULAR
C0024301|T047||CCS_10|FOLLICULAR MALIGNANT LYMPHOMA - CENTROBLASTIC-CENTROCYTIC 
C0024301|T047||CCS_10|FOLLICULAR LOW GRADE B-CELL LYMPHOMA 
C0024301|T047||CCS_10|FOLLICULAR LOW GRADE B-CELL LYMPHOMA
C0024301|T047||CCS_10|LYMPHOMA, FOLLICULAR, MALIGNANT
C0024301|T047||CCS_10|LYMPHOMA, FOLLICULAR CENTRE CELL
C0024301|T047||CCS_10|FOLLICULAR CENTRE CELL LYMPHOMA
C0024301|T047||CCS_10|FOLLICLE CENTER LYMPHOMA
C0024301|T047||CCS_10|NODULAR (FOLLICULAR) LYMPHOMA
C0024301|T047||CCS_10|MALIGNANT LYMPHOMA, NODULAR
C0024301|T047||CCS_10|MALIGNANT LYMPHOMA, FOLLICULAR
C0024301|T047||CCS_10|FOLLICULAR LYMPHOSARCOMA
C0024301|T047||CCS_10|BRILL - SYMMERS' DISEASE
C0024301|T047||CCS_10|GERMINOBLASTOMA, FOLLICULAR
C0024301|T047||CCS_10|FOLLICULAR LOW GRADE B-CELL LYMPHOMA 
C0024301|T047||CCS_10|FOLLICULAR LYMPHOMA (MORPHOLOGIC ABNORMALITY)
C0024301|T047||CCS_10|FOLLICULAR NON-HODGKIN'S LYMPHOMA 
C0024301|T047||CCS_10|MALIGNANT LYMPHOMA, CENTROBLASTIC-CENTROCYTIC, FOLLICULAR 
C0024301|T047||CCS_10|MALIGNANT LYMPHOMA, FOLLICLE CENTER, FOLLICULAR
C0024301|T047||CCS_10|MALIGNANT LYMPHOMA, FOLLICLE CENTER
C0024301|T047||CCS_10|MALIGNANT LYMPHOMA, FOLLICLE CENTRE, FOLLICULAR
C0024301|T047||CCS_10|MALIGNANT LYMPHOMA, FOLLICLE CENTRE
C0024301|T047||CCS_10|MALIGNANT LYMPHOMA, LYMPHOCYTIC, NODULAR
C0024301|T047||CCS_10|NODULAR LYMPHOMA 
C0024301|T047||CCS_10|FOLLICULAR; GERMINOBLASTOMA
C0024301|T047||CCS_10|FOLLICULAR; LYMPHOSARCOMA
C0024301|T047||CCS_10|GERMINOBLASTOMA; FOLLICULAR
C0024301|T047||CCS_10|BRILL-SYMMERS
C0024301|T047||CCS_10|LYMPHOCYTIC; LYMPHOMA, NODULAR
C0024301|T047||CCS_10|LYMPHOMA; FOLLICULAR
C0024301|T047||CCS_10|LYMPHOMA; LYMPHOCYTIC, NODULAR
C0024301|T047||CCS_10|LYMPHOMA; NODULAR, LYMPHOCYTIC
C0024301|T047||CCS_10|LYMPHOMA; NODULAR
C0024301|T047||CCS_10|LYMPHOSARCOMA; FOLLICULAR
C0024301|T047||CCS_10|NODULAR; LYMPHOMA, LYMPHOCYTIC
C0024301|T047||CCS_10|NODULAR; LYMPHOMA
C0024301|T047||CCS_10|MALIGNANT LYMPHOMA, FOLLICULAR, NOS
C0024301|T047||CCS_10|MALIGNANT LYMPHOMA, LYMPHOCYTIC, NODULAR, NOS
C0024301|T047||CCS_10|MALIGNANT LYMPHOMA, NODULAR, NOS
C0024301|T047||CCS_10|NODULAR LYMPHOCYTIC LYMPHOMA
C1264191|T047||CCS_10|MALIGNANT IMMUNOPROLIFERATIVE DISEASE, UNSPECIFIED
C1264191|T047||CCS_10|MALIGNANT IMMUNOPROLIFERATIVE DISEASES
C1264191|T047||CCS_10|MALIGNANT IMMUNOPROLIFERATIVE DISEASE
C1264191|T047||CCS_10|MALIGNANT IMMUNOPROLIFERATIVE DISEASE 
C1264191|T047||CCS_10|MALIGNANT IMMUNOPROLIFERATIVE DISEASE (CLINICAL)
C1264191|T047||CCS_10|MALIGNANT IMMUNOPROLIFERATIVE DISEASE 
C0494174|T047||CCS_10|MULTIPLE MYELOMA AND MALIGNANT PLASMA CELL NEOPLASMS
C0494176|T047||CCS_10|OTHER AND UNSPECIFIED MALIGNANT NEOPLASMS OF LYMPHOID, HAEMATOPOIETIC AND RELATED TISSUE
C0494176|T047||CCS_10|OTHER AND UNSPECIFIED MALIGNANT NEOPLASMS OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE
C0494172|T047||CCS_10|OTHER AND UNSPECIFIED TYPES OF NON-HODGKIN'S LYMPHOMA
C0494172|T047||CCS_10|OTHER SPECIFIED AND UNSPECIFIED TYPES OF NON-HODGKIN LYMPHOMA
C0494175|T047||CCS_10|OTHER LEUKAEMIAS OF SPECIFIED CELL TYPE
C0494175|T047||CCS_10|OTHER LEUKEMIAS OF SPECIFIED CELL TYPE
C0456860|T047||CCS_10|PERIPHERAL AND CUTANEOUS T-CELL LYMPHOMAS
C0456860|T047||CCS_10|MALIGNANT NEOPLASM LYMPHOMA CUTANEOUS / PERIPHERAL T-CELL
C0456860|T047||CCS_10|CUTANEOUS / PERIPHERAL T-CELL LYMPHOMA
C0456860|T047||CCS_10|CUTANEOUS / PERIPHERAL T-CELL LYMPHOMA 
C0456860|T047||CCS_10|CUTANEOUS/PERIPHERAL T-CELL LYMPHOMA
C0456860|T047||CCS_10|CUTANEOUS/PERIPHERAL T-CELL LYMPHOMA 
C2853945|T047||CCS_10|NON-FOLLICULAR LYMPHOMA
C0079774|T047||CCS_10|LYMPHOMA, PERIPHERAL T-CELL
C0079774|T047||CCS_10|LYMPHOMA, T-CELL, PERIPHERAL
C0079774|T047||CCS_10|LYMPHOMAS, PERIPHERAL T-CELL
C0079774|T047||CCS_10|PERIPHERAL T CELL LYMPHOMA
C0079774|T047||CCS_10|PERIPHERAL T-CELL LYMPHOMAS
C0079774|T047||CCS_10|T CELL LYMPHOMA, PERIPHERAL
C0079774|T047||CCS_10|T-CELL LYMPHOMAS, PERIPHERAL
C0079774|T047||CCS_10|PERIPHERAL T-CELL LYMPHOMA
C0079774|T047||CCS_10|MATURE T-CELL AND NK-CELL NON-HODGKIN'S LYMPHOMA
C0079774|T047||CCS_10|MATURE T-CELL AND NK-CELL NON-HODGKIN LYMPHOMA
C0079774|T047||CCS_10|MATURE T-CELL LYMPHOMA
C0079774|T047||CCS_10|MATURE T-CELL LYMPHOMA 
C0079774|T047||CCS_10|PERIPHERAL T-CELL LYMPHOMA, NO ICD-O SUBTYPE
C0079774|T047||CCS_10|PERIPHERAL T-CELL LYMPHOMA, NOT OTHERWISE SPECIFIED
C0079774|T047||CCS_10|PERIPHERAL T-CELL LYMPHOMA, NOS
C0079774|T047||CCS_10|MATURE T/NK-CELL LYMPHOMAS, UNSPECIFIED
C0079774|T047||CCS_10|MATURE T/NK-CELL LYMPHOMAS
C0079774|T047||CCS_10|LYMPHOMA, T-CELL, PERIPHERAL [DISEASE/FINDING]
C0079774|T047||CCS_10|T-CELL LYMPHOMA, PERIPHERAL
C0079774|T047||CCS_10|LYMPHOMA, T CELL, PERIPHERAL
C0079774|T047||CCS_10|[M] PERIPHERAL T-CELL LYMPHOMA NOS (MORPHOLOGIC ABNORMALITY)
C0079774|T047||CCS_10|PERIPHERAL T-CELL LYMPHOMA 
C0079774|T047||CCS_10|[M] PERIPHERAL T-CELL LYMPHOMA NOS
C0079774|T047||CCS_10|MATURE NK/T-CELL LYMPHOMA 
C0079774|T047||CCS_10|MATURE NK/T-CELL LYMPHOMA
C0079774|T047||CCS_10|MALIGNANT NEOPLASM LYMPHOMA MATURE NK/T-CELL
C0079774|T047||CCS_10|PERIPHERAL T-CELL LYMPHOMA, NO INTERNATIONAL CLASSIFICATION OF DISEASES FOR ONCOLOGY SUBTYPE (MORPHOLOGIC ABNORMALITY)
C0079774|T047||CCS_10|PERIPHERAL T-CELL LYMPHOMA, NO ICD-O SUBTYPE (MORPHOLOGIC ABNORMALITY)
C0079774|T047||CCS_10|PERIPHERAL T-CELL LYMPHOMA, NO INTERNATIONAL CLASSIFICATION OF DISEASES FOR ONCOLOGY SUBTYPE
C0079774|T047||CCS_10|PERIPHERAL T-CELL LYMPHOMA UNSPECIFIED
C0079774|T047||CCS_10|PERIPHERAL T-CELL LYMPHOMA UNSPECIFIED NOS
C0079774|T047||CCS_10|PERIPHERAL T-CELL LYMPHOMA (CLINICAL)
C0079774|T047||CCS_10|T-CELL; LYMPHOMA, PERIPHERAL
C0079774|T047||CCS_10|LYMPHOMA; T-CELL, PERIPHERAL
C0079774|T047||CCS_10|LYMPHOMA; PERIPHERAL T-CELL
C0079774|T047||CCS_10|PERIPHERAL; T-CELL LYMPHOMA
C0079774|T047||CCS_10|MATURE T-CELL NON-HODGKIN'S LYMPHOMA
C0079774|T047||CCS_10|MATURE T-CELL AND NK-CELL LYMPHOMA
C0079774|T047||CCS_10|MATURE T-AND NK-CELL LYMPHOMA
C0079774|T047||CCS_10|PTCL
C0079774|T047||CCS_10|PERIPHERAL T-CELL LYMPHOMA (MORPHOLOGIC ABNORMALITY)
C2854064|T047||CCS_10|OTHER SPECIFIED TYPES OF T/NK-CELL LYMPHOMA
C2854069|T047||CCS_10|MALIGNANT IMMUNOPROLIFERATIVE DISEASES AND CERTAIN OTHER B-CELL LYMPHOMAS
C0152276|T047||CCS_10|MYELOID SARCOMA
C0152276|T047||CCS_10|CHLOROMA
C0152276|T047||CCS_10|SARCOMAS, MYELOID
C0152276|T047||CCS_10|MYELOID SARCOMAS
C0152276|T047||CCS_10|SARCOMA, MYELOID
C0152276|T047||CCS_10|MYELOID SARCOMA, MORPHOLOGY
C0152276|T047||CCS_10|MYELOID SARCOMA, DISEASE
C0152276|T047||CCS_10|CHLOROMA 
C0152276|T047||CCS_10|GRANULOCYTIC SARCOMA 
C0152276|T047||CCS_10|LEUKEMIA MYELOID SARCOMA
C0152276|T047||CCS_10|LEUKEMIA MYELOID SARCOMA GRANULOCYTIC SARCOMA
C0152276|T047||CCS_10|GRANULOCYTIC SARCOMA
C0152276|T047||CCS_10|MYELOID SARCOMA 
C0152276|T047||CCS_10|LEUKEMIA MYELOID SARCOMA CHLOROMA
C0152276|T047||CCS_10|MYELOID SARCOMA NOS
C0152276|T047||CCS_10|MYELOID CELL TUMOR, EXTRAMEDULLARY
C0152276|T047||CCS_10|EXTRAMEDULLARY MYELOID CELL TUMOR
C0152276|T047||CCS_10|SARCOMA, GRANULOCYTIC
C0152276|T047||CCS_10|SARCOMA, MYELOID [DISEASE/FINDING]
C0152276|T047||CCS_10|CHLOROMAS
C0152276|T047||CCS_10|GRANULOCYTIC SARCOMAS
C0152276|T047||CCS_10|SARCOMAS, GRANULOCYTIC
C0152276|T047||CCS_10|MYELOID SARCOMA NOS 
C0152276|T047||CCS_10|SARCOMA, GRANULOCYTIC, MALIGNANT
C0152276|T047||CCS_10|SARCOMA, MYELOID, MALIGNANT
C0152276|T047||CCS_10|[M]MYELOID SARCOMA
C0152276|T047||CCS_10|[M]CHLOROMA
C0152276|T047||CCS_10|[M]GRANULOCYTIC SARCOMA
C0152276|T047||CCS_10|EXTRAMEDULLARY MYELOID TUMOR
C0152276|T047||CCS_10|CHLOROMA 
C0152276|T047||CCS_10|GRANULOCYTIC SARCOMA 
C0152276|T047||CCS_10|MYELOID SARCOMA, DISEASE 
C0152276|T047||CCS_10|MYELOID SARCOMA, MORPHOLOGY (MORPHOLOGIC ABNORMALITY)
C0152276|T047||CCS_10|MYELOSARCOMA
C0152276|T047||CCS_10|GRANULOCYTIC; SARCOMA
C0152276|T047||CCS_10|MYELOID; SARCOMA
C0152276|T047||CCS_10|SARCOMA; GRANULOCYTIC
C0152276|T047||CCS_10|SARCOMA; MYELOID
C0348393|T047|2.10|CCS_10|MALIGNANT NEOPLASM OF LYMPHOID, HAEMATOPOIETIC AND RELATED TISSUE, UNSPECIFIED|CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|MALIGNANT NEOPLASM OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE, UNSPECIFIED|CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|MALIGNANT NEOPLASMS OF LYMPHOID, HAEMATOPOIETIC AND RELATED TISSUE|CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|MALIGNANT NEOPLASMS OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE|CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE|CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|MALIGNANT NEOPLASMS OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE (C81-C96)|CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|MALIGNANT TUMOR OF LYMPHOID HEMOPOIETIC AND RELATED TISSUE|CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|MALIG NEOPLM OF LYMPHOID, HEMATPOETC AND REL TISSUE, UNSP|CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|[X]MALIGNANT NEOPLASM OF LYMPHOID, HAEMATOPOIETIC AND RELATED TISSUE, UNSPECIFIED|CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|MALIGNANT NEOPLASM OF LYMPHATIC AND HEMOPOIETIC TISSUE|CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|[X]MALIGNANT NEOPLASMS OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE |CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|[X]MALIGNANT NEOPLASMS OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE|CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|[X]MALIGNANT NEOPLASM OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE, UNSPECIFIED|CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|[X]MALIGNANT NEOPLASM OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE, UNSPECIFIED |CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|[X]MALIGNANT NEOPLASMS OF LYMPHOID, HAEMATOPOIETIC AND RELATED TISSUE|CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|MALIGNANT NEOPLASM OF LYMPHATIC AND HAEMOPOIETIC TISSUE|CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|MALIGNANT NEOPLASM OF LYMPHOID, HEMOPOIETIC AND/OR RELATED TISSUE |CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|MALIGNANT NEOPLASM OF LYMPHOID, HEMOPOIETIC AND/OR RELATED TISSUE|CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|MALIGNANT TUMOR OF LYMPHOID, HEMOPOIETIC AND/OR RELATED TISSUE|CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|MALIGNANT TUMOUR OF LYMPHOID HAEMOPOIETIC AND RELATED TISSUE|CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|HEMATOPOIETIC/LYMPHOID CANCER|CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|MALIGNANT TUMOR OF LYMPHOID, HEMOPOIETIC AND/OR RELATED TISSUE |CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|MALIGNANT TUMOR OF LYMPHOID HEMOPOIETIC AND RELATED TISSUE |CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348393|T047|2.10|CCS_10|MALIGNANT NEOPLASM OF LYMPHATIC AND HEMATOPOIETIC TISSUE|CANCER OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0021071|T047||CCS_10|ALPHA CHAIN DISEASE
C0021071|T047||CCS_10|IMMUNOPROLIFERATIVE SMALL INTESTINAL DISEASE
C0021071|T047||CCS_10|DISEASE, ALPHA-CHAIN
C0021071|T047||CCS_10|DISEASES, ALPHA-CHAIN
C0021071|T047||CCS_10|ALPHA-CHAIN DISEASES
C0021071|T047||CCS_10|ALPHA HEAVY CHAIN DISEASE
C0021071|T047||CCS_10|ALPHA CHAIN DIS
C0021071|T047||CCS_10|HEAVY CHAIN DIS IGA TYPE
C0021071|T047||CCS_10|IMMUNOPROLIFERATIVE SMALL INTESTINAL DIS
C0021071|T047||CCS_10|MEDITERRANEANL LYMPHOMA
C0021071|T047||CCS_10|ALPHA HEAVY CHAIN DISEASE, NOS
C0021071|T047||CCS_10|IMMUNOPROLIFERATIVE SMALL INTESTINAL DISEASE 
C0021071|T047||CCS_10|ALPHA HEAVY CHAIN DISEASE -RETIRED-
C0021071|T047||CCS_10|IMMUNOPROLIFERATIVE INTESTINAL DISEASE
C0021071|T047||CCS_10|MEDITERRANEAN LYMPHOMA
C0021071|T047||CCS_10|IMMUNOPROLIFERATIVE SMALL INTESTINAL DISEASE [DISEASE/FINDING]
C0021071|T047||CCS_10|LYMPHOMA, MEDITERRANEAN
C0021071|T047||CCS_10|HEAVY CHAIN DISEASE, IGA TYPE
C0021071|T047||CCS_10|ALPHA-CHAIN DISEASE
C0021071|T047||CCS_10|IPSID
C0021071|T047||CCS_10|[M] IMMUNOPROLIFERATIVE SMALL INTESTINAL DISEASE
C0021071|T047||CCS_10|[M] ALPHA HEAVY CHAIN DISEASE
C0021071|T047||CCS_10|ALPHA HEAVY CHAIN DISEASE 
C0021071|T047||CCS_10|[M] ALPHA HEAVY CHAIN DISEASE (MORPHOLOGIC ABNORMALITY)
C0021071|T047||CCS_10|[M] IMMUNOPROLIFERATIVE SMALL INTESTINAL DISEASE (MORPHOLOGIC ABNORMALITY)
C0021071|T047||CCS_10|ALPHA HEAVY CHAIN DISEASE 
C0021071|T047||CCS_10|ALPHA HEAVY CHAIN DISEASE, ENTERIC FORM 
C0021071|T047||CCS_10|HEAVY CHAIN DISEASE ALPHA, ENTERIC FORM
C0021071|T047||CCS_10|ALPHA HEAVY CHAIN DISEASE, ENTERIC FORM
C0021071|T047||CCS_10|HEAVY CHAIN DISEASE ALPHA
C0021071|T047||CCS_10|IMMUNOPROLIFERATIVE SMALL INTESTINAL DISEASE (CLINICAL)
C0021071|T047||CCS_10|IMMUNOPROLIFERATIVE SMALL INTESTINAL DISEASE 
C0021071|T047||CCS_10|IMMUNOPROLIFERATIVE SMALL INTESTINAL DISEASE (MORPHOLOGIC ABNORMALITY)
C0021071|T047||CCS_10|ALPHA HEAVY CHAIN DISEASE (CLINICAL)
C0021071|T047||CCS_10|ALPHA HEAVY CHAIN DISEASE, ENTERIC FORM 
C0021071|T047||CCS_10|MEDITERRANEAN LYMPHOMA (CLINICAL)
C0021071|T047||CCS_10|IGA HEAVY CHAIN DISEASE
C0021071|T047||CCS_10|DISEASE (OR DISORDER); ALPHA HEAVY CHAIN
C0021071|T047||CCS_10|DISEASE (OR DISORDER); HEAVY CHAIN, ALPHA
C0021071|T047||CCS_10|DISEASE (OR DISORDER); IMMUNOPROLIFERATIVE, SMALL INTESTINE
C0021071|T047||CCS_10|DISEASE; ALPHA HEAVY CHAIN
C0021071|T047||CCS_10|HEAVY CHAIN ALPHA
C0021071|T047||CCS_10|LYMPHOMA; MEDITERRANEAN
C0021071|T047||CCS_10|MEDITERRANEAN; LYMPHOMA
C0021071|T047||CCS_10|ALPHA HEAVY CHAIN; DISEASE
C0021071|T047||CCS_10|ALPHA; ALPHA HEAVY CHAIN DISEASE
C0021071|T047||CCS_10|IGA HEAVY CHAIN DISEASE, NOS
C0021071|T047||CCS_10|ALPHA HEAVY CHAIN DISEASE [DUP] 
C0021071|T047||CCS_10|MEDITERRANEAN ABDOMINAL LYMPHOMA
C0021071|T047||CCS_10|IMMUNOPROLIFERATIVE; DISEASE, SMALL INTESTINE
C0376545|T047||CCS_10|HEMATOLOGIC NEOPLASM
C0376545|T047||CCS_10|HEMATOLOGIC NEOPLASMS
C0376545|T047||CCS_10|HEMATOLOGICAL MALIGNANCY
C0376545|T047||CCS_10|HEMATOLOGICAL NEOPLASM
C0376545|T047||CCS_10|MALIGNANCIES, HEMATOLOGICAL
C0376545|T047||CCS_10|MALIGNANCY, HEMATOLOGICAL
C0376545|T047||CCS_10|NEOPLASM, HEMATOLOGIC
C0376545|T047||CCS_10|NEOPLASM, HEMATOLOGICAL
C0376545|T047||CCS_10|NEOPLASMS, HEMATOLOGICAL
C0376545|T047||CCS_10|HAEMATOLOGICAL MALIGNANCY
C0376545|T047||CCS_10|NEOPL HEMATOL
C0376545|T047||CCS_10|MALIGNANCY HEMATOL
C0376545|T047||CCS_10|HEMATOL NEOPL
C0376545|T047||CCS_10|HEMATOL MALIGNANCY
C0376545|T047||CCS_10|MALIGNANCIES HEMATOL
C0376545|T047||CCS_10|HEMATOL MALIGNANCIES
C0376545|T047||CCS_10|HEMATOLOGIC MALIGNANCY
C0376545|T047||CCS_10|MALIGNANCY, HEMATOLOGIC
C0376545|T047||CCS_10|HEMATOLOGIC MALIGNANCIES
C0376545|T047||CCS_10|HEMATOLOGICAL NEOPLASMS
C0376545|T047||CCS_10|HEMATOLOGICAL MALIGNANCIES
C0376545|T047||CCS_10|HEMATOLOGIC NEOPLASMS [DISEASE/FINDING]
C0376545|T047||CCS_10|MALIGNANCIES, HEMATOLOGIC
C0376545|T047||CCS_10|NEOPLASMS, HEMATOLOGIC
C0376545|T047||CCS_10|CARCINOMA;BLOOD
C0376545|T047||CCS_10|CARCINOMA;BONE;MARROW
C0376545|T047||CCS_10|BLOOD CANCER
C0376545|T047||CCS_10|HEMATOLOGIC MALIGNANCY 
C0376545|T047||CCS_10|HAEMATOLOGIC MALIGNANCY
C0376545|T047||CCS_10|HEMATOLOGIC CANCER
C0376545|T047||CCS_10|HAEMATOLOGIC NEOPLASM
C0376545|T047||CCS_10|HEMATOLOGIC NEOPLASM 
C0376545|T047||CCS_10|HEMATOLOGICAL TUMOR
C0376545|T047||CCS_10|MALIGNANT HEMATOLOGIC NEOPLASM
C0018854|T047||CCS_10|FRANKLINS DISEASE
C0018854|T047||CCS_10|FRANKLIN'S DISEASE
C0018854|T047||CCS_10|GAMMA CHAIN DISEASE
C0018854|T047||CCS_10|GAMMA-CHAIN DISEASES
C0018854|T047||CCS_10|GAMMA HEAVY CHAIN DISEASE
C0018854|T047||CCS_10|FRANKLINS DIS
C0018854|T047||CCS_10|FRANKLIN DIS
C0018854|T047||CCS_10|GAMMA HEAVY CHAIN DISEASE -RETIRED-
C0018854|T047||CCS_10|FRANKLIN DISEASE
C0018854|T047||CCS_10|GAMMA HEAVY CHAIN DISEASE 
C0018854|T047||CCS_10|[M] GAMMA HEAVY CHAIN DISEASE
C0018854|T047||CCS_10|GAMMA HEAVY CHAIN DISEASE (MORPHOLOGIC ABNORMALITY)
C0018854|T047||CCS_10|[M] GAMMA HEAVY CHAIN DISEASE (MORPHOLOGIC ABNORMALITY)
C0018854|T047||CCS_10|:: GAMMA HEAVY CHAIN DISEASE
C0018854|T047||CCS_10|HEAVY CHAIN DISEASE GAMMA
C0018854|T047||CCS_10|GAMMA HEAVY CHAIN DISEASE 
C0018854|T047||CCS_10|GAMMA HEAVY CHAIN DISEASE (CLINICAL)
C0018854|T047||CCS_10|DISEASE; GAMMA HEAVY CHAIN
C0018854|T047||CCS_10|GAMMA HEAVY CHAIN; DISEASE
C0018854|T047||CCS_10|HEAVY CHAIN GAMMA
C0018854|T047||CCS_10|IGG HEAVY CHAIN DISEASE
C0018854|T047||CCS_10|GAMMA HEAVY CHAIN DISEASE [DUP] 
C0018854|T047||CCS_10|GAMMA-CHAIN DISEASE
C0543670|T047||CCS_10|MALIGNANT WHITE BLOOD CELL DISORDER
C0543670|T047||CCS_10|MALIGNANT WHITE BLOOD CELL DISORDER 
C0543670|T047||CCS_10|MALIGNANT NEOPLASM WHITE BLOOD CELL DISORDER
C0543670|T047||CCS_10|MALIGNANT WHITE BLOOD CELL DISORDER 
C0474969|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHATIC OR HEMATOPOIETIC TISSUE OTHERWISE SPECIFIED 
C0474969|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHATIC OR HEMATOPOIETIC TISSUE OTHERWISE SPECIFIED
C0474969|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHATIC OR HAEMATOPOIETIC TISSUE OTHERWISE SPECIFIED
C0474970|T047||CCS_10|LYMPHATIC/HEMATOPOIETIC NEOPLASM
C0474970|T047||CCS_10|NEOPLASM OF LYMPHATIC OR HEMATOPOIETIC TISSUE
C0474970|T047||CCS_10|MALIGNANT NEOPLASM LYMPHATIC OR HAEMATOPOIETIC TISSUE NOS
C0474970|T047||CCS_10|MALIGNANT NEOPLASM LYMPHATIC OR HEMATOPOIETIC TISSUE NOS 
C0474970|T047||CCS_10|MALIGNANT NEOPLASM LYMPHATIC OR HEMATOPOIETIC TISSUE NOS
C0474970|T047||CCS_10|MALIGNANT LYMPHATIC/HEMATOPOIETIC NEOPLASM 
C0474970|T047||CCS_10|MALIGNANT LYMPHATIC/HEMATOPOIETIC NEOPLASM
C0348391|T047||CCS_10|OTHER MALIGNANT IMMUNOPROLIFERATIVE DISEASES
C0348391|T047||CCS_10|[X]OTHER MALIGNANT IMMUNOPROLIFERATIVE DISEASES
C0348391|T047||CCS_10|[X]OTHER MALIGNANT IMMUNOPROLIFERATIVE DISEASES 
C0348392|T047||CCS_10|OTHER SPECIFIED MALIGNANT NEOPLASMS OF LYMPHOID, HAEMATOPOIETIC AND RELATED TISSUE
C0348392|T047||CCS_10|OTHER SPECIFIED MALIGNANT NEOPLASMS OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE
C0348392|T047||CCS_10|OTH MALIG NEOPLM OF LYMPHOID, HEMATPOETC AND RELATED TISSUE
C0348392|T047||CCS_10|[X]OTHER SPECIFIED MALIGNANT NEOPLASMS OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE 
C0348392|T047||CCS_10|[X]OTHER SPECIFIED MALIGNANT NEOPLASMS OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE
C0348392|T047||CCS_10|[X]OTHER SPECIFIED MALIGNANT NEOPLASMS OF LYMPHOID, HAEMATOPOIETIC AND RELATED TISSUE
C0024299|T047||CCS_10|LYMPHOMAS
C0024299|T047||CCS_10|GERMINOBLASTIC SARCOMAS
C0024299|T047||CCS_10|GERMINOBLASTOMAS
C0024299|T047||CCS_10|LYMPHOMA
C0024299|T047||CCS_10|RETICULOLYMPHOSARCOMAS
C0024299|T047||CCS_10|SARCOMAS, GERMINOBLASTIC
C0024299|T047||CCS_10|LYMPHOMAS, MALIGNANT
C0024299|T047||CCS_10|MALIGNANT LYMPHOMAS
C0024299|T047||CCS_10|GERMINOBLASTIC SARCOMA
C0024299|T047||CCS_10|MALIGNANT LYMPHOMA
C0024299|T047||CCS_10|LYMPHOMA (HODGKIN AND NON-HODGKIN)
C0024299|T047||CCS_10|MALIGNANT LYMPHOMA - CATEGORY
C0024299|T047||CCS_10|MALIGNANT LYMPHOMA 
C0024299|T047||CCS_10|MALIGNANT LYMPHOMA 
C0024299|T047||CCS_10|MALIGNANT LYMPHOMA, NO ICD-O SUBTYPE
C0024299|T047||CCS_10|LYMPHOMA NOS
C0024299|T047||CCS_10|MALIGNANT LYMPHOMA NOS
C0024299|T047||CCS_10|GERMINOBLASTOMA
C0024299|T047||CCS_10|RETICULOLYMPHOSARCOMA
C0024299|T047||CCS_10|SARCOMA, GERMINOBLASTIC
C0024299|T047||CCS_10|LYMPHOMA, MALIGNANT
C0024299|T047||CCS_10|LYMPHOMA [DISEASE/FINDING]
C0024299|T047||CCS_10|LYMPHOMATOUS
C0024299|T047||CCS_10|MALIGNANT LYMPHOMA NOS OF UNSPECIFIED SITE
C0024299|T047||CCS_10|MALIGNANT LYMPHOMA NOS 
C0024299|T047||CCS_10|[M]RETICULOLYMPHOSARCOMA NOS
C0024299|T047||CCS_10|[M]MALIGNANT LYMPHOMA NOS 
C0024299|T047||CCS_10|MALIGNANT LYMPHOMA NOS OF UNSPECIFIED SITE 
C0024299|T047||CCS_10|LYMPHOMA MORPHOLOGY
C0024299|T047||CCS_10|[M]MALIGNANT LYMPHOMA NOS
C0024299|T047||CCS_10|LYMPHOMA MORPHOLOGY (MORPHOLOGIC ABNORMALITY)
C0024299|T047||CCS_10|LYMPHOSARCOMA
C0024299|T047||CCS_10|MALIGNANT LYMPHOMA, NO ICD-O SUBTYPE (MORPHOLOGIC ABNORMALITY)
C0024299|T047||CCS_10|MALIGNANT LYMPHOMA, NO INTERNATIONAL CLASSIFICATION OF DISEASES FOR ONCOLOGY SUBTYPE (MORPHOLOGIC ABNORMALITY)
C0024299|T047||CCS_10|MALIGNANT LYMPHOMA, NO INTERNATIONAL CLASSIFICATION OF DISEASES FOR ONCOLOGY SUBTYPE
C0024299|T047||CCS_10|LYMPHOMA, NOS
C0024299|T047||CCS_10|LYMPHOMA (HODGKIN'S AND NON-HODGKIN'S)
C0024299|T047||CCS_10|LYMPHOMA MALIGNANT
C0024299|T047||CCS_10|LYMPHOMA (CLINICAL)
C0024299|T047||CCS_10|MALIGNANT LYMPHOMA (CLINICAL)
C0024299|T047||CCS_10|MALIGNANT LYMPHOMA 
C0024299|T047||CCS_10|MALIGNANT LYMPHOMA - CATEGORY (MORPHOLOGIC ABNORMALITY)
C0024299|T047||CCS_10|MALIGNANT LYMPHOMA, NOS
C1306621|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF SPLEEN
C1306621|T047||CCS_10|SPLENIC NEOPLASM MALIGNANT PRIMARY
C1306621|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF SPLEEN 
C1306621|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF SPLEEN 
C0040028|T047||CCS_10|ESSENTIAL THROMBOCYTHEMIAS
C0040028|T047||CCS_10|HEMORRHAGIC THROMBOCYTHEMIAS
C0040028|T047||CCS_10|IDIOPATHIC THROMBOCYTHEMIAS
C0040028|T047||CCS_10|PRIMARY THROMBOCYTHEMIAS
C0040028|T047||CCS_10|THROMBOCYTHEMIAS, ESSENTIAL
C0040028|T047||CCS_10|THROMBOCYTHEMIAS, HEMORRHAGIC
C0040028|T047||CCS_10|THROMBOCYTHEMIAS, IDIOPATHIC
C0040028|T047||CCS_10|THROMBOCYTHEMIAS, PRIMARY
C0040028|T047||CCS_10|ESSENTIAL THROMBOCYTHEMIA
C0040028|T047||CCS_10|IDIOPATHIC THROMBOCYTHEMIA
C0040028|T047||CCS_10|HEMORRHAGIC THROMBOCYTHEMIA
C0040028|T047||CCS_10|ESSENTIAL (HAEMORRHAGIC) THROMBOCYTHAEMIA
C0040028|T047||CCS_10|ESSENTIAL (HEMORRHAGIC) THROMBOCYTHEMIA
C0040028|T047||CCS_10|ESSENTIAL THROMBOCYTHAEMIA
C0040028|T047||CCS_10|ESSENTIAL THROMBOCYTOSIS
C0040028|T047||CCS_10|ESSENTIAL HEMORRHAGIC THROMBOCYTHEMIA
C0040028|T047||CCS_10|IDIOPATHIC (HEMORRHAGIC) THROMBOCYTHEMIA
C0040028|T047||CCS_10|PRIMARY THROMBOCYTOSIS
C0040028|T047||CCS_10|PRIMARY THROMBOCYTHEMIA
C0040028|T047||CCS_10|ESSENTIAL THROMBOCYTHAEMIA 
C0040028|T047||CCS_10|ESSENTIAL THROMBOCYTHEMIA (CLINICAL)
C0040028|T047||CCS_10|ESSENTIAL THROMBOCYTOSIS 
C0040028|T047||CCS_10|ESSENTIAL THROMBOCYTHEMIA 
C0040028|T047||CCS_10|PRIMARY THROMBOCYTOSIS 
C0040028|T047||CCS_10|IDIOPATHIC THROMBOCYTHEMIA 
C0040028|T047||CCS_10|IDIOPATHIC THROMBOCYTHAEMIA -RETIRED-
C0040028|T047||CCS_10|IDIOPATHIC THROMBOCYTHEMIA -RETIRED-
C0040028|T047||CCS_10|ESSENTIAL HEMORRHAGIC THROMBOCYTHEMIA 
C0040028|T047||CCS_10|THROMBOCYTHEMIA, ESSENTIAL
C0040028|T047||CCS_10|IDEOPATHIC THROMBOCYTOSIS
C0040028|T047||CCS_10|ESSNTIAL THROMBOCYTHEMIA
C0040028|T047||CCS_10|IDIOPATHIC HEMORRHAGIC THROMBOCYTHEMIA
C0040028|T047||CCS_10|THROMBOCYTHEMIA, PRIMARY
C0040028|T047||CCS_10|THROMBOCYTHEMIA, IDIOPATHIC
C0040028|T047||CCS_10|THROMBOCYTHEMIA, ESSENTIAL [DISEASE/FINDING]
C0040028|T047||CCS_10|THROMBOCYTHEMIA, HEMORRHAGIC
C0040028|T047||CCS_10|THROMBOCYTOSIS;ESSENTIAL
C0040028|T047||CCS_10|THROMBOCYTOSES, PRIMARY
C0040028|T047||CCS_10|PRIMARY THROMBOCYTOSES
C0040028|T047||CCS_10|THROMBOCYTOSIS, PRIMARY
C0040028|T047||CCS_10|IDIOPATHIC THROMBOCYTHAEMIA
C0040028|T047||CCS_10|ESSENTIAL THROMBOCYTOSIS 
C0040028|T047||CCS_10|ET - ESSENTIAL THROMBOCYTHAEMIA
C0040028|T047||CCS_10|ESSENTIAL THROMBOCYTHAEMIA 
C0040028|T047||CCS_10|IDIOPATHIC THROMBOCYTHEMIA 
C0040028|T047||CCS_10|ET - ESSENTIAL THROMBOCYTHEMIA
C0040028|T047||CCS_10|IDIOPATHIC THROMBOCYTHAEMIA 
C0040028|T047||CCS_10|IDIOPATHIC THROMBOCYTHEMIA (MORPHOLOGIC ABNORMALITY)
C0040028|T047||CCS_10|[M]IDIOPATHIC THROMBOCYTHAEMIA
C0040028|T047||CCS_10|[M]IDIOPATHIC THROMBOCYTHEMIA
C0040028|T047||CCS_10|PRIMARY THROMBOCYTHAEMIA
C0040028|T047||CCS_10|IDIOPATHIC THROMBOCYTOSIS
C0040028|T047||CCS_10|ESSENTIAL HAEMORRHAGIC THROMBOCYTHAEMIA
C0040028|T047||CCS_10|IDIOPATHIC HAEMORRHAGIC THROMBOCYTHAEMIA
C0040028|T047||CCS_10|ESSENTIAL THROMBOCYTHEMIA 
C0040028|T047||CCS_10|ESSENTIAL THROMBOCYTHEMIA (MORPHOLOGIC ABNORMALITY)
C0040028|T047||CCS_10|THROMBOCYTOSIS; ESSENTIAL
C0040028|T047||CCS_10|ESSENTIAL THROMBOCYTHAEMIA (CLINICAL)
C0040028|T047||CCS_10|ESSENTIAL THROMBOCYTEMIA
C0040028|T047||CCS_10|ESSENTIAL THROMBOCYTHEMIA 
C3463824|T047||CCS_10|DYSMYELOPOIETIC SYNDROME
C3463824|T047||CCS_10|MYELODYSPLASTIC SYNDROMES
C3463824|T047||CCS_10|SYNDROME, DYSMYELOPOIETIC
C3463824|T047||CCS_10|SYNDROMES, DYSMYELOPOIETIC
C3463824|T047||CCS_10|SYNDROMES, MYELODYSPLASTIC
C3463824|T047||CCS_10|MYELODYSPLASTIC SYNDROME
C3463824|T047||CCS_10|SYNDROME, MYELODYSPLASTIC
C3463824|T047||CCS_10|MYELODYSPLASTIC SYNDROME, UNSPECIFIED
C3463824|T047||CCS_10|OLIGOBLASTIC LEUKEMIA
C3463824|T047||CCS_10|MYELODYSPLASIA
C3463824|T047||CCS_10|MYELODYSPLASTIC SYNDROME (MORPHOLOGY) -RETIRED-
C3463824|T047||CCS_10|MYELODYSPLASTIC SYNDROME (MORPHOLOGY)
C3463824|T047||CCS_10|MYELODYSPLASIA 
C3463824|T047||CCS_10|MYELODYSPLASTIC SYND NOS
C3463824|T047||CCS_10|MYELODYSPLASTIC SYNDROME/NEOPLASM
C3463824|T047||CCS_10|MYELODYSPLASTIC NEOPLASM
C3463824|T047||CCS_10|HEMATOPOEITIC - MYELODYSPLASTIC SYNDROME (MDS)
C3463824|T047||CCS_10|MYELODYSPLASTIC SYNDROMES [DISEASE/FINDING]
C3463824|T047||CCS_10|DYSMYELOPOIETIC SYNDROMES
C3463824|T047||CCS_10|MDS
C3463824|T047||CCS_10|PRELEUKEMIA
C3463824|T047||CCS_10|SMOLDERING LEUKEMIA
C3463824|T047||CCS_10|[X]MYELODYSPLASTIC SYNDROME, UNSPECIFIED
C3463824|T047||CCS_10|SMOULDERING LEUKAEMIA
C3463824|T047||CCS_10|MYELODYSPLASTIC SYNDROME 
C3463824|T047||CCS_10|PRELEUKAEMIA
C3463824|T047||CCS_10|MYELODYSPLASTIC SYNDROME (MORPHOLOGIC ABNORMALITY)
C3463824|T047||CCS_10|PRELEUKEMIC SYNDROME
C3463824|T047||CCS_10|MYELODYSPLASIA 
C3463824|T047||CCS_10|PRELEUKAEMIC SYNDROME
C3463824|T047||CCS_10|[X]MYELODYSPLASTIC SYNDROME, UNSPECIFIED 
C3463824|T047||CCS_10|[M]MYELODYSPLASTIC SYNDROME
C3463824|T047||CCS_10|MYELODYSPLASTIC SYNDROME 
C3463824|T047||CCS_10|MYELODYSPLASTIC SYNDROME, NOS
C3463824|T047||CCS_10|MYELODYSPLASTIC SYNDROME, SUSCEPTIBILITY TO
C3463824|T047||CCS_10|MYELOID DYSPLASIA
C3463824|T047||CCS_10|MYELODYSPLASTIC SYNDROME NOS
C3463824|T047||CCS_10|MDS - MYELODYSPLASTIC SYNDROME
C3463824|T047||CCS_10|MYELODYSPLASTIC SYNDROME (CLINICAL)
C3463824|T047||CCS_10|DYSMYELOPOIESIS
C3463824|T047||CCS_10|MYELODYSPLASTIC; SYNDROME
C3463824|T047||CCS_10|PRELEUKEMIC; SYNDROME
C3463824|T047||CCS_10|SYNDROME; MYELODYSPLASTIC
C3463824|T047||CCS_10|SYNDROME; PRELEUKEMIC
C0019613|T047||CCS_10|DISORDER, MALIGNANT HISTIOCYTIC
C0019613|T047||CCS_10|DISORDERS, MALIGNANT HISTIOCYTIC
C0019613|T047||CCS_10|HISTIOCYTIC DISORDER, MALIGNANT
C0019613|T047||CCS_10|HISTIOCYTIC DISORDERS, MALIGNANT
C0019613|T047||CCS_10|MALIGNANT HISTIOCYTIC DISORDER
C0019613|T047||CCS_10|MALIGNANT HISTIOCYTIC DISORDERS
C0019613|T047||CCS_10|HISTIOCYTIC DISORDERS, MALIGNANT [DISEASE/FINDING]
C0019613|T047||CCS_10|MALIG NEOPLASM HISTIOCYTIC DISORDER
C0019613|T047||CCS_10|MALIGNANT HISTIOCYTIC DISORDER 
C0019613|T047||CCS_10|MALIGNANT HISTIOCYTIC DISORDER 
C0341713|T047||CCS_10|LEUKEMIC INFILTRATE OF KIDNEY 
C0341713|T047||CCS_10|LEUKEMIC INFILTRATE OF KIDNEY
C0341713|T047||CCS_10|RENAL NEOPLASM MALIGNANT LEUKEMIC INFILTRATE
C0341713|T047||CCS_10|LEUKAEMIC INFILTRATE OF KIDNEY
C0341713|T047||CCS_10|LEUKEMIC INFILTRATE OF KIDNEY 
C1301145|T047||CCS_10|MAST CELL MALIGNANCY 
C1301145|T047||CCS_10|MAST CELL MALIGNANCY
C1301145|T047||CCS_10|MAST CELL MALIGNANCY 
C0024305|T047||CCS_10|LYMPHOMA, NON HODGKIN'S
C0024305|T047||CCS_10|LYMPHOMA, NON-HODGKIN
C0024305|T047||CCS_10|LYMPHOMA, NONHODGKIN
C0024305|T047||CCS_10|NON HODGKIN'S LYMPHOMA
C0024305|T047||CCS_10|NON-HODGKINS LYMPHOMA
C0024305|T047||CCS_10|NONHODGKIN'S LYMPHOMA
C0024305|T047||CCS_10|NON-HODGKIN'S LYMPHOMA, UNSPECIFIED TYPE
C0024305|T047||CCS_10|LYMPHOMA, NON HODGKIN
C0024305|T047||CCS_10|LYMPHOMA, NON HODGKINS
C0024305|T047||CCS_10|NON HODGKIN LYMPHOMA
C0024305|T047||CCS_10|NONHODGKINS LYMPHOMA
C0024305|T047||CCS_10|SMALL CLEAVED CELL (DIFFUSE) NON-HODGKIN'S LYMPHOMA
C0024305|T047||CCS_10|LYMPHOMA, NON-HODGKIN, FAMILIAL
C0024305|T047||CCS_10|NON-HODGKIN LYMPHOMA
C0024305|T047||CCS_10|THIS IS AN OK ABBREV.
C0024305|T047||CCS_10|NONHODGKIN LYMPHOMA
C0024305|T047||CCS_10|NON-HODGKIN'S LYMPHOMA
C0024305|T047||CCS_10|DIFFUSE SMALL CLEAVED CELL LYMPHOMA
C0024305|T047||CCS_10|LYMPHOMA SMALL CLEAVED DIFFUSE
C0024305|T047||CCS_10|SMALL CLEAVED CELL LYMPHOMA, DIFFUSE
C0024305|T047||CCS_10|DIFFUSE SMALL CLEAVED LYMPHOMA
C0024305|T047||CCS_10|SMALL CLEAVED LYMPHOMA DIFFUSE
C0024305|T047||CCS_10|MALIGNANT LYMPHOMA, NON-HODGKIN'S, NOS
C0024305|T047||CCS_10|NON-HODGKIN'S LYMPHOMA 
C0024305|T047||CCS_10|NON-HODGKIN LYMPHOMA - CATEGORY
C0024305|T047||CCS_10|MALIGNANT LYMPHOMA, SMALL CLEAVED CELL, DIFFUSE -RETIRED-
C0024305|T047||CCS_10|NON-HODGKIN LYMPHOMA, NO ICD-O SUBTYPE
C0024305|T047||CCS_10|NON-HODGKIN'S LYMPHOMA (NHL)
C0024305|T047||CCS_10|NON-HODGKIN LYMPHOMA NOS
C0024305|T047||CCS_10|LYMPHOMA, NONHODGKINS
C0024305|T047||CCS_10|LYMPHOMA, NON-HODGKIN'S
C0024305|T047||CCS_10|LYMPHOMA, NONHODGKIN'S
C0024305|T047||CCS_10|LYMPHOMA, NON-HODGKIN [DISEASE/FINDING]
C0024305|T047||CCS_10|LYMPHOMA, NON-HODGKINS
C0024305|T047||CCS_10|SMALL CLEAVED-CELL LYMPHOMA, DIFFUSE
C0024305|T047||CCS_10|LYMPHOMA, ATYPICAL DIFFUSE SMALL LYMPHOID
C0024305|T047||CCS_10|DIFFUSE SMALL CLEAVED-CELL LYMPHOMA
C0024305|T047||CCS_10|LYMPHOMA, SMALL CLEAVED CELL, DIFFUSE
C0024305|T047||CCS_10|LYMPHOMA, SMALL CLEAVED-CELL, DIFFUSE
C0024305|T047||CCS_10|LYMPHOMA;NON HODGKINS
C0024305|T047||CCS_10|[X]NON-HODGKIN'S LYMPHOMA, UNSPECIFIED TYPE 
C0024305|T047||CCS_10|[X]NON-HODGKIN'S LYMPHOMA, UNSPECIFIED TYPE
C0024305|T047||CCS_10|NON-HODGKIN'S LYMPHOMA NOS
C0024305|T047||CCS_10|[M]MALIGNANT LYMPHOMA, SMALL CLEAVED CELL, DIFFUSE (MORPHOLOGIC ABNORMALITY)
C0024305|T047||CCS_10|[M]MALIGNANT LYMPHOMA, SMALL CLEAVED CELL, DIFFUSE
C0024305|T047||CCS_10|NON-HODGKIN LYMPHOMA, NO INTERNATIONAL CLASSIFICATION OF DISEASES FOR ONCOLOGY SUBTYPE (MORPHOLOGIC ABNORMALITY)
C0024305|T047||CCS_10|NON-HODGKIN LYMPHOMA, NO ICD-O SUBTYPE (MORPHOLOGIC ABNORMALITY)
C0024305|T047||CCS_10|NON-HODGKIN LYMPHOMA, NO INTERNATIONAL CLASSIFICATION OF DISEASES FOR ONCOLOGY SUBTYPE
C0024305|T047||CCS_10|NHL, NOS
C0024305|T047||CCS_10|NON-HODGKIN LYMPHOMA, NOS
C0024305|T047||CCS_10|[M]NON-HODGKIN'S LYMPHOMA
C0024305|T047||CCS_10|[M]MALIGNANT LYMPHOMA, NON-HODGKIN'S TYPE
C0024305|T047||CCS_10|LYMPHOMA (NON-HODGKIN'S)
C0024305|T047||CCS_10|NON-HODGKIN`S LYMPHOMA
C0024305|T047||CCS_10|DIFFUSE NON-HODGKIN'S SMALL CLEAVED CELL (DIFFUSE) LYMPHOMA
C0024305|T047||CCS_10|MALIGNANT LYMPHOMA, NON-HODGKIN'S TYPE
C0024305|T047||CCS_10|NHL - NON-HODGKIN'S LYMPHOMA
C0024305|T047||CCS_10|MALIGNANT LYMPHOMA, CLEAVED CELL [OBS]
C0024305|T047||CCS_10|MALIGNANT LYMPHOMA, NON-HODGKIN'S
C0024305|T047||CCS_10|MALIGNANT LYMPHOMA, NON-HODGKIN
C0024305|T047||CCS_10|MALIGNANT LYMPHOMA, SMALL CELL, NONCLEAVED, DIFFUSE [OBS]
C0024305|T047||CCS_10|MALIGNANT LYMPHOMA, SMALL CLEAVED CELL [OBS]
C0024305|T047||CCS_10|MALIGNANT LYMPHOMA, SMALL CLEAVED CELL, DIFFUSE [OBS]
C0024305|T047||CCS_10|MALIGNANT LYMPHOMA, UNDIFFERENTIATED CELL TYPE [OBS]
C0024305|T047||CCS_10|MALIGNANT LYMPHOMA, UNDIFFERENTIATED CELL, NON-BURKITT [OBS]
C0024305|T047||CCS_10|NON-HODGKIN LYMPHOMA 
C0024305|T047||CCS_10|NON-HODGKIN LYMPHOMA - CATEGORY (MORPHOLOGIC ABNORMALITY)
C0024305|T047||CCS_10|NON-HODGKIN'S LYMPHOMA (CLINICAL)
C0024305|T047||CCS_10|NON-HODGKIN'S LYMPHOMA 
C0024305|T047||CCS_10|NON-HODGKIN'S LYMPHOMA - DISORDER
C0024305|T047||CCS_10|DIFFUSE; LYMPHOMA, SMALL CELL, CLEAVED
C0024305|T047||CCS_10|LYMPHOMA; DIFFUSE, SMALL CELL, CLEAVED
C0024305|T047||CCS_10|LYMPHOMA; NON-HODGKIN'S
C0024305|T047||CCS_10|LYMPHOMA; SMALL CELL, CLEAVED (DIFFUSE)
C0024305|T047||CCS_10|NON-HODGKIN'S; LYMPHOMA
C0024305|T047||CCS_10|SMALL CELL; LYMPHOMA, CLEAVED (DIFFUSE)
C0024305|T047||CCS_10|NON-HODGKIN'S LYMPHOMA, NOS
C0024305|T047||CCS_10|NON HODGKINS LYMPHOMA
C1292778|T047||CCS_10|CHRONIC MYELOPROLIFERATIVE DISEASE
C1292778|T047||CCS_10|MYELOPROLIFERATIVE DISEASE (CHRONIC) NOS
C1292778|T047||CCS_10|CHRONIC MYELOPROLIFERATIVE DISORDER
C1292778|T047||CCS_10|CHRONIC MYELOPROLIFERATIVE DISEASE -RETIRED-
C1292778|T047||CCS_10|CHRONIC MYELOPROLIFERATIVE DISEASE, NO ICD-O SUBTYPE
C1292778|T047||CCS_10|MYELOPROLIFERATIVE DISORDER
C1292778|T047||CCS_10|MYELOPROLIFERATIVE NEOPLASM
C1292778|T047||CCS_10|CHRONIC MYELOPROLIFERATIVE NEOPLASM
C1292778|T047||CCS_10|MYELOPROLIFERATIVE TUMOR
C1292778|T047||CCS_10|CHRONIC MYELOPROLIFERATIVE SYNDROME 
C1292778|T047||CCS_10|CHRONIC MYELOPROLIFERATIVE SYNDROME
C1292778|T047||CCS_10|MYELOPROLIFERATIVE SYNDROME CHRONIC
C1292778|T047||CCS_10|CHRONIC MYELOPROLIFERATIVE DISEASE, NO INTERNATIONAL CLASSIFICATION OF DISEASES FOR ONCOLOGY SUBTYPE
C1292778|T047||CCS_10|CHRONIC MYELOPROLIFERATIVE DISEASE, NO INTERNATIONAL CLASSIFICATION OF DISEASES FOR ONCOLOGY SUBTYPE (MORPHOLOGIC ABNORMALITY)
C1292778|T047||CCS_10|CHRONIC MYELOPROLIFERATIVE DISEASE, NO ICD-O SUBTYPE (MORPHOLOGIC ABNORMALITY)
C1292778|T047||CCS_10|MYELOPROLIFERATIVE NEOPLASM, NO ICD-O SUBTYPE
C1292778|T047||CCS_10|CHRONIC MYELOPROLIFERATIVE DISORDER (MORPHOLOGY)
C1292778|T047||CCS_10|PROBABLY OK
C1292778|T047||CCS_10|CHRONIC MYELOPROLIFERATIVE DISORDER (CLINICAL) 
C1292778|T047||CCS_10|CHRONIC MYELOPROLIFERATIVE DISORDER (CLINICAL)
C1292778|T047||CCS_10|CHRONIC MYELOPROLIFERATIVE DISORDER (MORPHOLOGIC ABNORMALITY)
C1292778|T047||CCS_10|CHRONIC MYELOPROLIFERATIVE DISORDERS
C1292778|T047||CCS_10|DISEASE (OR DISORDER); MYELOPROLIFERATIVE (CHRONIC)
C1292778|T047||CCS_10|MYELOPROLIFERATIVE; DISEASE (CHRONIC)
C1292778|T047||CCS_10|CMPD
C1292778|T047||CCS_10|CHRONIC MYELOPROLIFERATIVE DISEASE (MORPHOLOGIC ABNORMALITY)
C1292778|T047||CCS_10|CHRONIC MYELOPROLIFERATIVE DISEASE NOS
C1301355|T047||CCS_10|DISEASE, MYELOPROLIFERATIVE-MYELODISPLASTIC
C1301355|T047||CCS_10|DISEASES, MYELOPROLIFERATIVE-MYELODISPLASTIC
C1301355|T047||CCS_10|MYELODYSPLASTIC-MYELOPROLIFERATIVE DISEASES
C1301355|T047||CCS_10|MYELODYSPLASTIC-MYELOPROLIFERATIVE DISEASE
C1301355|T047||CCS_10|DISEASE, MYELODYSPLASTIC-MYELOPROLIFERATIVE
C1301355|T047||CCS_10|MYELODYSPLASTIC MYELOPROLIFERATIVE DISEASES
C1301355|T047||CCS_10|MYELOPROLIFERATIVE-MYELODISPLASTIC DISEASE
C1301355|T047||CCS_10|DISEASES, MYELODYSPLASTIC-MYELOPROLIFERATIVE
C1301355|T047||CCS_10|MYELOPROLIFERATIVE MYELODISPLASTIC DISEASES
C1301355|T047||CCS_10|MYELODYSPLASTIC/MYELOPROLIFERATIVE NEOPLASM
C1301355|T047||CCS_10|MYELODYSPLASTIC/MYELOPROLIFERATIVE DISEASE
C1301355|T047||CCS_10|MDS/MPN
C1301355|T047||CCS_10|MYELOPROLIFERATIVE-MYELODISPLASTIC DISEASES
C1301355|T047||CCS_10|MYELODYSPLASTIC-MYELOPROLIFERATIVE DISEASES [DISEASE/FINDING]
C1301355|T047||CCS_10|MYELODYSPLASTIC/MYELOPROLIFERATIVE DISEASE 
C1301355|T047||CCS_10|MYELODYSPLASTIC / MYELOPROLIFERATIVE DISEASE
C1301355|T047||CCS_10|MYELODYSPLASTIC / MYELOPROLIFERATIVE DISEASE 
C1301355|T047||CCS_10|BONE MARROW NEOPLASM MYELODYSPLASTIC / MYELOPROLIFERATIVE DISEASE
C1301355|T047||CCS_10|MYELODYSPLASTIC/MYELOPROLIFERATIVE DISEASE (MORPHOLOGIC ABNORMALITY)
C1301355|T047||CCS_10|MDS/MPD
C1301355|T047||CCS_10|MYELODYSPLASTIC/MYELOPROLIFERATIVE DISEASES
C1301355|T047||CCS_10|MDS-MPD
C1301355|T047||CCS_10|MPD-MDS
C1301355|T047||CCS_10|MPD/MDS
C1301355|T047||CCS_10|MYELODYSPLASTIC/MYELOPROLIFERATIVE DISORDERS
C1301355|T047||CCS_10|MYELODYSPLASTIC/MYELOPROLIFERATIVE DISORDER
C1301355|T047||CCS_10|MYELOPROLIFERATIVE/MYELODYSPLASTIC DISORDERS
C1301355|T047||CCS_10|MYELOPROLIFERATIVE/MYELODYSPLASTIC SYNDROMES
C0029812|T047||CCS_10|OTHER SPECIFIED LEUKAEMIAS
C0029812|T047||CCS_10|OTHER SPECIFIED LEUKEMIAS
C0029812|T047||CCS_10|OTHER SPECIFIED LEUKEMIA 
C0029812|T047||CCS_10|OTHER SPECIFIED LEUKEMIAS NOS
C0029812|T047||CCS_10|OTHER SPECIFIED LEUKEMIA NOS 
C0029812|T047||CCS_10|[X]OTHER SPECIFIED LEUKAEMIAS
C0029812|T047||CCS_10|OTHER SPECIFIED LEUKEMIA
C0029812|T047||CCS_10|OTHER SPECIFIED LEUKAEMIA
C0029812|T047||CCS_10|OTHER SPECIFIED LEUKEMIA NOS
C0029812|T047||CCS_10|[X]OTHER SPECIFIED LEUKEMIAS
C0029812|T047||CCS_10|[X]OTHER SPECIFIED LEUKEMIAS 
C0029812|T047||CCS_10|OTHER SPECIFIED LEUKAEMIA NOS
C1955727|T047||CCS_10|LYMPHOSARCOMA AND RETICULOSARCOMA AND OTHER SPECIFIED MALIGNANT TUMORS OF LYMPHATIC TISSUE
C0153867|T047||CCS_10|MULTIPLE MYELOMA AND IMMUNOPROLIFERATIVE NEOPLASMS
C0153867|T047||CCS_10|MULTIPLE MYELOMA AND IMMUNOPROLIFERATIVE DISEASE
C0153867|T047||CCS_10|MULTIPLE MYELOMA AND IMMUNOPROLIFERATIVE DISEASE 
C0153793|T047||CCS_10|OTHER MALIGNANT NEOPLASMS OF LYMPHOID AND HISTIOCYTIC TISSUE
C0153793|T047||CCS_10|OTHER MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE 
C0153793|T047||CCS_10|OTHER MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE
C0432564|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE
C0432564|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE 
C0432564|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND/OR HISTIOCYTIC TISSUE -RETIRED-
C0432564|T047||CCS_10|MALIGNANT TUMOR OF LYMPHOID AND HISTIOCYTIC TISSUE
C0432564|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND/OR HISTIOCYTIC TISSUE
C0432564|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND/OR HISTIOCYTIC TISSUE 
C0432564|T047||CCS_10|UNSPECIFIED MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE OF UNSPECIFIED SITE 
C0432564|T047||CCS_10|UNSPECIFIED MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE OF UNSPECIFIED SITE
C0432564|T047||CCS_10|MALIGNANT NEOPLASMS OF LYMPHOID AND HISTIOCYTIC TISSUE NOS 
C0432564|T047||CCS_10|MALIGNANT NEOPLASMS OF LYMPHOID AND HISTIOCYTIC TISSUE NOS
C0432564|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE, NOS
C2217148|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE OF HEAD, FACE, OR NECK 
C2217148|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE OF HEAD, FACE, OR NECK
C2217148|T047||CCS_10|MALIGNANT TUMOR OF LYMPHOID AND HISTIOCYTIC TISSUE OF HEAD, FACE, OR NECK
C2217152|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE OF INTRATHORACIC REGION 
C2217152|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE OF INTRATHORACIC REGION
C2217152|T047||CCS_10|MALIGNANT NEOPLASM OF INTRATHORACIC LYMPHOID AND HISTIOCYTIC TISSUE
C2217152|T047||CCS_10|MALIGNANT TUMOR OF LYMPHOID AND HISTIOCYTIC TISSUE OF INTRATHORACIC REGION
C2217150|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE OF INTRA-ABDOMINAL REGION 
C2217150|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE OF INTRA-ABDOMINAL REGION
C2217150|T047||CCS_10|MALIGNANT NEOPLASM OF INTRA-ABDOMINAL LYMPHOID AND HISTIOCYTIC TISSUE
C2217150|T047||CCS_10|MALIGNANT TUMOR OF LYMPHOID AND HISTIOCYTIC TISSUE OF INTRA-ABDOMINAL REGION
C2217147|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE OF AXILLA OR UPPER LIMB
C2217147|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE OF AXILLA OR UPPER LIMB 
C2217147|T047||CCS_10|MALIGNANT TUMOR OF LYMPHOID AND HISTIOCYTIC TISSUE OF AXILLA OR UPPER LIMB
C2217149|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE OF INGUINAL REGION OR LOWER LIMB 
C2217149|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE OF INGUINAL REGION OR LOWER LIMB
C2217149|T047||CCS_10|MALIGNANT TUMOR OF LYMPHOID AND HISTIOCYTIC TISSUE OF INGUINAL REGION OR LOWER LIMB
C2217151|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE OF INTRAPELVIC REGION 
C2217151|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE OF INTRAPELVIC REGION
C2217151|T047||CCS_10|MALIGNANT NEOPLASM OF INTRAPELVIC LYMPHOID AND HISTIOCYTIC TISSUE
C2217151|T047||CCS_10|MALIGNANT TUMOR OF LYMPHOID AND HISTIOCYTIC TISSUE OF INTRAPELVIC REGION
C2217154|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE OF SPLEEN
C2217154|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE OF SPLEEN 
C2217154|T047||CCS_10|MALIGNANT NEOPLASM OF SPLENIC LYMPHOID AND HISTIOCYTIC TISSUE
C2217154|T047||CCS_10|MALIGNANT TUMOR OF LYMPHOID AND HISTIOCYTIC TISSUE OF SPLEEN
C2217153|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE OF MULTIPLE SITES 
C2217153|T047||CCS_10|MALIGNANT NEOPLASM OF LYMPHOID AND HISTIOCYTIC TISSUE OF MULTIPLE SITES
C2217153|T047||CCS_10|MALIGNANT TUMOR OF LYMPHOID AND HISTIOCYTIC TISSUE OF MULTIPLE SITES
C0936223|T047||CCS_10|PROSTATE CANCER METASTATIC
C0936223|T047||CCS_10|METASTATIC PROSTATE CARCINOMA
C0936223|T047||CCS_10|METASTATIC PROSTATE CANCER
C0936223|T047||CCS_10|CARCINOMA OF THE PROSTATE METASTATIC
C0936223|T047||CCS_10|PROSTATIC CANCER METASTATIC
C0936223|T047||CCS_10|PROSTATE CARCINOMA METASTATIC
C0278838|T047||CCS_10|PROSTATE CANCER RECURRENT
C0278838|T047||CCS_10|RECURRENT PROSTATE CANCER
C0278838|T047||CCS_10|RECURRENT PROSTATE CARCINOMA
C0278838|T047||CCS_10|CARCINOMA OF THE PROSTATE RECURRENT
C0278838|T047||CCS_10|PROSTATIC CANCER RECURRENT
C0278838|T047||CCS_10|PROSTATE CANCER, RECURRENT
C0278838|T047||CCS_10|RECURRENT CANCER OF PROSTATE
C0278838|T047||CCS_10|RECURRENT CANCER OF THE PROSTATE
C0854969|T047||CCS_10|PROSTATE CANCER STAGE 0
C0854969|T047||CCS_10|PROSTATIC CANCER STAGE 0
C0278834|T047||CCS_10|PROSTATE CANCER STAGE I
C0278834|T047||CCS_10|STAGE I PROSTATE CARCINOMA
C0278834|T047||CCS_10|STAGE I PROSTATE CANCER AJCC V6
C0278834|T047||CCS_10|STAGE I PROSTATIC CANCER AJCC V6
C0278834|T047||CCS_10|PROSTATE CARCINOMA STAGE I AJCC V6
C0278834|T047||CCS_10|PROSTATE CANCER STAGE I AJCC V6
C0278834|T047||CCS_10|STAGE I PROSTATE CARCINOMA AJCC V6
C0278834|T047||CCS_10|CANCER OF PROSTATE STAGE I AJCC V6
C0278834|T047||CCS_10|CANCER OF THE PROSTATE STAGE I AJCC V6
C0278834|T047||CCS_10|STAGE I CANCER OF THE PROSTATE AJCC V6
C0278834|T047||CCS_10|STAGE I CANCER OF PROSTATE AJCC V6
C0278834|T047||CCS_10|STAGE I PROSTATIC CARCINOMA AJCC V6
C0278834|T047||CCS_10|STAGE I PROSTATE CANCER
C0278834|T047||CCS_10|PROSTATIC CANCER STAGE I
C0278834|T047||CCS_10|CARCINOMA OF THE PROSTATE STAGE I
C0278834|T047||CCS_10|CANCER OF THE PROSTATE, STAGE I
C0278834|T047||CCS_10|CARCINOMA OF THE PROSTATE, STAGE I
C0278834|T047||CCS_10|PROSTATE CANCER, STAGE I
C0278834|T047||CCS_10|STAGE I CANCER OF THE PROSTATE
C0278834|T047||CCS_10|STAGE I CARCINOMA OF THE PROSTATE
C0278835|T047||CCS_10|PROSTATE CANCER STAGE II
C0278835|T047||CCS_10|STAGE II PROSTATE CARCINOMA
C0278835|T047||CCS_10|CANCER OF THE PROSTATE STAGE II AJCC V6
C0278835|T047||CCS_10|PROSTATE CANCER STAGE II AJCC V6
C0278835|T047||CCS_10|STAGE II CANCER OF PROSTATE AJCC V6
C0278835|T047||CCS_10|STAGE II CANCER OF THE PROSTATE AJCC V6
C0278835|T047||CCS_10|STAGE II PROSTATE CARCINOMA AJCC V6
C0278835|T047||CCS_10|PROSTATE CARCINOMA STAGE II AJCC V6
C0278835|T047||CCS_10|STAGE II PROSTATE CANCER AJCC V6
C0278835|T047||CCS_10|STAGE II PROSTATIC CARCINOMA AJCC V6
C0278835|T047||CCS_10|STAGE II PROSTATIC CANCER AJCC V6
C0278835|T047||CCS_10|CANCER OF PROSTATE STAGE II AJCC V6
C0278835|T047||CCS_10|STAGE II PROSTATE CANCER
C0278835|T047||CCS_10|PROSTATIC CANCER STAGE II
C0278835|T047||CCS_10|CARCINOMA OF THE PROSTATE STAGE II
C0278835|T047||CCS_10|CANCER OF THE PROSTATE, STAGE II
C0278835|T047||CCS_10|CARCINOMA OF THE PROSTATE, STAGE II
C0278835|T047||CCS_10|PROSTATE CANCER, STAGE II
C0278835|T047||CCS_10|STAGE II CANCER OF THE PROSTATE
C0278835|T047||CCS_10|STAGE II CARCINOMA OF THE PROSTATE
C0278836|T047||CCS_10|PROSTATE CANCER STAGE III
C0278836|T047||CCS_10|STAGE III PROSTATE CARCINOMA
C0278836|T047||CCS_10|STAGE III PROSTATE CARCINOMA AJCC V6
C0278836|T047||CCS_10|STAGE III CANCER OF PROSTATE AJCC V6
C0278836|T047||CCS_10|CANCER OF PROSTATE STAGE III AJCC V6
C0278836|T047||CCS_10|PROSTATE CANCER STAGE III AJCC V6
C0278836|T047||CCS_10|STAGE III CANCER OF THE PROSTATE AJCC V6
C0278836|T047||CCS_10|PROSTATE CARCINOMA STAGE III AJCC V6
C0278836|T047||CCS_10|STAGE III PROSTATE CANCER AJCC V6
C0278836|T047||CCS_10|CANCER OF THE PROSTATE STAGE III AJCC V6
C0278836|T047||CCS_10|STAGE III PROSTATIC CANCER AJCC V6
C0278836|T047||CCS_10|STAGE III PROSTATIC CARCINOMA AJCC V6
C0278836|T047||CCS_10|STAGE III PROSTATE CANCER
C0278836|T047||CCS_10|CARCINOMA OF THE PROSTATE STAGE III
C0278836|T047||CCS_10|PROSTATIC CANCER STAGE III
C0278836|T047||CCS_10|CANCER OF THE PROSTATE, STAGE III
C0278836|T047||CCS_10|CARCINOMA OF THE PROSTATE, STAGE III
C0278836|T047||CCS_10|PROSTATE CANCER, STAGE III
C0278836|T047||CCS_10|STAGE III CANCER OF THE PROSTATE
C0278836|T047||CCS_10|STAGE III CARCINOMA OF THE PROSTATE
C0278837|T047||CCS_10|PROSTATE CANCER STAGE IV
C0278837|T047||CCS_10|STAGE IV PROSTATE CARCINOMA
C0278837|T047||CCS_10|STAGE IV PROSTATE CANCER AJCC V6
C0278837|T047||CCS_10|PROSTATE CANCER STAGE IV AJCC V6
C0278837|T047||CCS_10|STAGE IV CANCER OF PROSTATE AJCC V6
C0278837|T047||CCS_10|STAGE IV CANCER OF THE PROSTATE AJCC V6
C0278837|T047||CCS_10|PROSTATE CARCINOMA STAGE IV AJCC V6
C0278837|T047||CCS_10|STAGE IV PROSTATIC CANCER AJCC V6
C0278837|T047||CCS_10|CANCER OF PROSTATE STAGE IV AJCC V6
C0278837|T047||CCS_10|CANCER OF THE PROSTATE STAGE IV AJCC V6
C0278837|T047||CCS_10|STAGE IV PROSTATE CARCINOMA AJCC V6
C0278837|T047||CCS_10|STAGE IV PROSTATIC CARCINOMA AJCC V6
C0278837|T047||CCS_10|STAGE IV PROSTATE CANCER
C0278837|T047||CCS_10|CARCINOMA OF THE PROSTATE STAGE IV
C0278837|T047||CCS_10|PROSTATIC CANCER STAGE IV
C0278837|T047||CCS_10|CANCER OF THE PROSTATE, STAGE IV
C0278837|T047||CCS_10|CARCINOMA OF THE PROSTATE, STAGE IV
C0278837|T047||CCS_10|PROSTATE CANCER, STAGE IV
C0278837|T047||CCS_10|STAGE IV CANCER OF THE PROSTATE
C0278837|T047||CCS_10|STAGE IV CARCINOMA OF THE PROSTATE
C1297952|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING PROSTATE BY DIRECT EXTENSION FROM BLADDER 
C1297952|T047||CCS_10|PROSTATE GLAND MALIGNANT BY DIRECT EXTENSION FROM BLADDER
C1297952|T047||CCS_10|MALIGNANT NEOPLASM INVOLVING PROSTATE BY DIRECT EXTENSION FROM BLADDER
C1297952|T047||CCS_10|MALIGNANT TUMOR INVOLVING PROSTATE BY DIRECT EXTENSION FROM BLADDER 
C1297952|T047||CCS_10|MALIGNANT TUMOR INVOLVING PROSTATE BY DIRECT EXTENSION FROM BLADDER
C1297952|T047||CCS_10|MALIGNANT TUMOUR INVOLVING PROSTATE BY DIRECT EXTENSION FROM BLADDER
C2007082|T047||CCS_10|CARCINOSARCOMA OF PROSTATE GLAND 
C2007082|T047||CCS_10|CARCINOSARCOMA OF PROSTATE GLAND
C2212269|T047||CCS_10|MALIGNANT SMALL CELL NEOPLASM OF PROSTATE GLAND
C2212269|T047||CCS_10|PROSTATE GLAND NEOPLASM MALIGNANT SMALL CELL TYPE
C2212269|T047||CCS_10|MALIGNANT SMALL CELL NEOPLASM OF PROSTATE GLAND 
C2011401|T047||CCS_10|GIANT CELL TYPE NEOPLASM OF PROSTATE GLAND 
C2011401|T047||CCS_10|PROSTATE GLAND NEOPLASM MALIGNANT GIANT CELL TYPE
C2011401|T047||CCS_10|GIANT CELL TYPE NEOPLASM OF PROSTATE GLAND
C2018684|T047||CCS_10|SPINDLE CELL TYPE NEOPLASM OF PROSTATE GLAND
C2018684|T047||CCS_10|SPINDLE CELL TYPE NEOPLASM OF PROSTATE GLAND 
C2018684|T047||CCS_10|PROSTATE GLAND NEOPLASM MALIGNANT SPINDLE CELL TYPE
C2075644|T047||CCS_10|PROSTATE GLAND NEOPLASM MALIGNANT CLEAR CELL TYPE
C2075644|T047||CCS_10|CLEAR CELL TYPE NEOPLASM OF PROSTATE GLAND
C2075644|T047||CCS_10|CLEAR CELL TYPE NEOPLASM OF PROSTATE GLAND 
C0600139|T047||CCS_10|CARCINOMA OF PROSTATE
C0600139|T047||CCS_10|CARCINOMA OF PROSTATE GLAND
C0600139|T047||CCS_10|CARCINOMA OF PROSTATE GLAND 
C0600139|T047||CCS_10|PROSTATIC CARCINOMA
C0600139|T047||CCS_10|CARCINOMA;PROSTATE
C0600139|T047||CCS_10|CANCER OF PROSTATE
C0600139|T047||CCS_10|CARCINOMA OF PROSTATE 
C0600139|T047||CCS_10|PROSTATE CANCER, NOS
C0600139|T047||CCS_10|PROSTATE CANCER
C0600139|T047||CCS_10|PROSTATE CARCINOMA
C0600139|T047||CCS_10|CARCINOMA PROSTATE
C0600139|T047||CCS_10|CARCINOMA PROSTATIC
C0600139|T047||CCS_10|CA - CARCINOMA OF PROSTATE
C0600139|T047||CCS_10|CARCINOMA, PROSTATIC
C0600139|T047||CCS_10|CANCER OF THE PROSTATE
C0600139|T047||CCS_10|CARCINOMA OF THE PROSTATE
C2212291|T047||CCS_10|SARCOMA OF PROSTATE GLAND 
C2212291|T047||CCS_10|SARCOMA OF PROSTATE GLAND
C2212294|T047||CCS_10|FIBROSARCOMA OF PROSTATE GLAND
C2212294|T047||CCS_10|FIBROSARCOMA OF PROSTATE GLAND 
C2212297|T047||CCS_10|MYOSARCOMA OF PROSTATE GLAND
C2212297|T047||CCS_10|MYOSARCOMA OF PROSTATE GLAND 
C2142688|T047||CCS_10|MARGINAL ZONE B-CELL LYMPHOMA OF PROSTATE GLAND
C2142688|T047||CCS_10|MARGINAL ZONE B-CELL LYMPHOMA OF PROSTATE GLAND 
C2217386|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE GLAND STAGING
C2217386|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE GLAND STAGING 
C2217386|T047||CCS_10|MALIGNANT PROSTATIC NEOPLASM STAGING
C2217386|T047||CCS_10|PROSTATIC CANCER STAGING
C2217386|T047||CCS_10|MALIGNANT TUMOR OF PROSTATE GLAND STAGING
C0007112|T047||CCS_10|ADENOCARCINOMA OF PROSTATE GLAND
C0007112|T047||CCS_10|ADENOCARCINOMA OF PROSTATE GLAND 
C0007112|T047||CCS_10|PROSTATIC ADENOCARCINOMA
C0007112|T047||CCS_10|PROSTATE ADENOCARCINOMA
C0007112|T047||CCS_10|ADENOCARCINOMA OF PROSTATE
C0007112|T047||CCS_10|ADENOCARCINOMA OF PROSTATE 
C0007112|T047||CCS_10|ADENOCARCINOMA OF THE PROSTATE
C0007112|T047||CCS_10|ADENOCARCINOMA, PROSTATIC
C0007112|T047||CCS_10|PROSTATE CANCER, ADENOCARCINOMA
C2146665|T047||CCS_10|ACINAR CELL CARCINOMA OF PROSTATE GLAND 
C2146665|T047||CCS_10|ACINAR CELL CARCINOMA OF PROSTATE GLAND
C2146677|T047||CCS_10|ACINAR CELL CYSTADENOCARCINOMA OF PROSTATE GLAND
C2146677|T047||CCS_10|PROSTATE MALIGNANT CARCINOMA ACINAR CELL CYSTADENOCARCINOMA
C2146677|T047||CCS_10|ACINAR CELL CYSTADENOCARCINOMA OF PROSTATE GLAND 
C2033179|T047||CCS_10|PAPILLARY CARCINOMA IN SITU OF PROSTATE GLAND
C2033179|T047||CCS_10|PAPILLARY CARCINOMA IN SITU OF PROSTATE GLAND 
C2142680|T047||CCS_10|NONINVASIVE PAPILLARY SQUAMOUS CELL CARCINOMA IN SITU OF PROSTATE GLAND
C2142680|T047||CCS_10|PROSTATE GLAND CIS PAPILLARY SQUAMOUS CELL NONINVASIVE
C2142680|T047||CCS_10|NONINVASIVE PAPILLARY SQUAMOUS CELL CARCINOMA IN SITU OF PROSTATE GLAND 
C2019399|T047||CCS_10|SQUAMOUS CELL CARCINOMA IN SITU OF PROSTATE GLAND
C2019399|T047||CCS_10|SQUAMOUS CELL CARCINOMA IN SITU OF PROSTATE GLAND 
C2019400|T047||CCS_10|SQUAMOUS CELL CARCINOMA IN SITU OF PROSTATE GLAND WITH QUESTIONABLE STROMAL INVASION 
C2019400|T047||CCS_10|PROSTATE CARCINOMA IN SITU SQUAMOUS CELL WITH QUESTIONABLE STROMAL INVASION
C2019400|T047||CCS_10|SQUAMOUS CELL CARCINOMA IN SITU OF PROSTATE GLAND WITH QUESTIONABLE STROMAL INVASION
C2145436|T047||CCS_10|TRANSITIONAL CELL CARCINOMA IN SITU OF PROSTATE GLAND
C2145436|T047||CCS_10|TRANSITIONAL CELL CARCINOMA IN SITU OF PROSTATE GLAND 
C2142681|T047||CCS_10|NONINVASIVE PAPILLARY TRANSITIONAL CELL CARCINOMA IN SITU OF PROSTATE GLAND
C2142681|T047||CCS_10|PROSTATE GLAND CIS PAPILLARY TRANSITIONAL CELL NONINVASIVE
C2142681|T047||CCS_10|NONINVASIVE PAPILLARY TRANSITIONAL CELL CARCINOMA IN SITU OF PROSTATE GLAND 
C2142714|T047||CCS_10|NONINFILTRATING INTRADUCTAL PAPILLARY ADENOCARCINOMA IN SITU OF PROSTATE GLAND
C2142714|T047||CCS_10|NONINFILTRATING INTRADUCTAL PAPILLARY ADENOCARCINOMA IN SITU OF PROSTATE GLAND 
C2142714|T047||CCS_10|PROSTATE NONINFILTRATING INTRADUCTAL PAPILLARY ADENOCARCINOMA IN SITU
C2142679|T047||CCS_10|PROSTATE GLAND CIS NONINFILTRATING INTRACYSTIC CARCINOMA
C2142679|T047||CCS_10|NONINFILTRATING INTRACYSTIC CARCINOMA IN SITU OF PROSTATE GLAND
C2142679|T047||CCS_10|NONINFILTRATING INTRACYSTIC CARCINOMA IN SITU OF PROSTATE GLAND 
C2142677|T047||CCS_10|PROSTATE GLAND CARCINOMA IN SITU INTRADUCTAL MICROPAPILLARY
C2142677|T047||CCS_10|INTRADUCTAL MICROPAPILLARY CARCINOMA IN SITU OF PROSTATE GLAND 
C2142677|T047||CCS_10|INTRADUCTAL MICROPAPILLARY CARCINOMA IN SITU OF PROSTATE GLAND
C2212270|T047||CCS_10|MALIGNANT EPITHELIOMA OF PROSTATE GLAND 
C2212270|T047||CCS_10|MALIGNANT EPITHELIOMA OF PROSTATE GLAND
C2111662|T047||CCS_10|LARGE CELL CARCINOMA OF PROSTATE GLAND
C2111662|T047||CCS_10|LARGE CELL CARCINOMA OF PROSTATE GLAND 
C2111743|T047||CCS_10|LARGE CELL NEUROENDOCRINE CARCINOMA OF PROSTATE GLAND 
C2111743|T047||CCS_10|LARGE CELL NEUROENDOCRINE CARCINOMA OF PROSTATE GLAND
C2111663|T047||CCS_10|LARGE CELL CARCINOMA OF PROSTATE GLAND WITH RHABDOID PHENOTYPE
C2111663|T047||CCS_10|LARGE CELL CARCINOMA OF PROSTATE GLAND WITH RHABDOID PHENOTYPE 
C2111663|T047||CCS_10|PROSTATE MALIGNANT CARCINOMA LARGE CELL WITH RHABDOID PHENOTYPE
C2012107|T047||CCS_10|GLASSY CELL CARCINOMA OF PROSTATE GLAND
C2012107|T047||CCS_10|GLASSY CELL CARCINOMA OF PROSTATE GLAND 
C2188081|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF PROSTATE GLAND
C2188081|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF PROSTATE GLAND 
C2212271|T047||CCS_10|ANAPLASTIC CARCINOMA OF PROSTATE GLAND
C2212271|T047||CCS_10|ANAPLASTIC CARCINOMA OF PROSTATE GLAND 
C2082456|T047||CCS_10|PLEOMORPHIC CARCINOMA OF PROSTATE GLAND 
C2082456|T047||CCS_10|PLEOMORPHIC CARCINOMA OF PROSTATE GLAND
C2011261|T047||CCS_10|GIANT CELL CARCINOMA OF PROSTATE GLAND 
C2011261|T047||CCS_10|GIANT CELL CARCINOMA OF PROSTATE GLAND
C2018401|T047||CCS_10|SPINDLE CELL CARCINOMA OF PROSTATE GLAND 
C2018401|T047||CCS_10|SPINDLE CELL CARCINOMA OF PROSTATE GLAND
C2011226|T047||CCS_10|GIANT CELL AND SPINDLE CELL CARCINOMA OF PROSTATE GLAND 
C2011226|T047||CCS_10|GIANT CELL AND SPINDLE CELL CARCINOMA OF PROSTATE GLAND
C2011226|T047||CCS_10|PROSTATE MALIGNANT CARCINOMA GIANT CELL AND SPINDLE CELL
C2142931|T047||CCS_10|PSEUDOSARCOMATOUS CARCINOMA OF PROSTATE GLAND 
C2142931|T047||CCS_10|PSEUDOSARCOMATOUS CARCINOMA OF PROSTATE GLAND
C2111813|T047||CCS_10|POLYGONAL CELL CARCINOMA OF PROSTATE GLAND
C2111813|T047||CCS_10|POLYGONAL CELL CARCINOMA OF PROSTATE GLAND 
C2142712|T047||CCS_10|CARCINOMA OF PROSTATE GLAND WITH OSTEOCLAST-LIKE GIANT CELLS 
C2142712|T047||CCS_10|CARCINOMA OF PROSTATE GLAND WITH OSTEOCLAST-LIKE GIANT CELLS
C2142712|T047||CCS_10|PROSTATIC CARCINOMA WITH OSTEOCLAST-LIKE GIANT CELLS
C2033229|T047||CCS_10|PAPILLARY CARCINOMA OF PROSTATE GLAND
C2033229|T047||CCS_10|PAPILLARY CARCINOMA OF PROSTATE GLAND 
C2033307|T047||CCS_10|PAPILLARY SQUAMOUS CELL CARCINOMA OF PROSTATE GLAND 
C2033307|T047||CCS_10|PAPILLARY SQUAMOUS CELL CARCINOMA OF PROSTATE GLAND
C2189358|T047||CCS_10|VERRUCOUS CARCINOMA OF PROSTATE GLAND 
C2189358|T047||CCS_10|VERRUCOUS CARCINOMA OF PROSTATE GLAND
C2109317|T047||CCS_10|PROSTATE MALIGNANT CARCINOMA SQUAMOUS CELL KERATINIZING
C2109317|T047||CCS_10|KERATINIZING SQUAMOUS CELL CARCINOMA OF PROSTATE GLAND 
C2109317|T047||CCS_10|KERATINIZING SQUAMOUS CELL CARCINOMA OF PROSTATE GLAND
C2212272|T047||CCS_10|NONKERATINIZING LARGE CELL SQUAMOUS CARCINOMA CELL OF PROSTATE GLAND
C2212272|T047||CCS_10|PROSTATE MALIGNANT CARCINOMA SQUAMOUS CELL LARGE CELL NONKERATINIZING
C2212272|T047||CCS_10|NONKERATINIZING LARGE CELL SQUAMOUS CARCINOMA CELL OF PROSTATE GLAND 
C2212273|T047||CCS_10|NONKERATINIZING SMALL CELL SQUAMOUS CELL CARCINOMA OF PROSTATE GLAND 
C2212273|T047||CCS_10|PROSTATE MALIGNANT CARCINOMA SQUAMOUS CELL SMALL CELL NONKERATINIZING
C2212273|T047||CCS_10|NONKERATINIZING SMALL CELL SQUAMOUS CELL CARCINOMA OF PROSTATE GLAND
C2018564|T047||CCS_10|SPINDLE CELL SQUAMOUS CELL CARCINOMA OF PROSTATE GLAND 
C2018564|T047||CCS_10|SPINDLE CELL SQUAMOUS CELL CARCINOMA OF PROSTATE GLAND
C2018564|T047||CCS_10|PROSTATE MALIGNANT CARCINOMA SQUAMOUS CELL SPINDLE CELL
C2212275|T047||CCS_10|MICROINVASIVE SQUAMOUS CELL CARCINOMA OF PROSTATE GLAND 
C2212275|T047||CCS_10|PROSTATE MALIGNANT CARCINOMA SQUAMOUS CELL MICROINVASIVE
C2212275|T047||CCS_10|MICROINVASIVE SQUAMOUS CELL CARCINOMA OF PROSTATE GLAND
C2019492|T047||CCS_10|PROSTATE MALIGNANT CARCINOMA SQUAMOUS CELL WITH HORN FORMATION
C2019492|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF PROSTATE GLAND WITH HORN FORMATION
C2019492|T047||CCS_10|SQUAMOUS CELL CARCINOMA WITH HORN FORMATION OF PROSTATE GLAND
C2019492|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF PROSTATE GLAND WITH HORN FORMATION 
C2009885|T047||CCS_10|FUSIFORM TYPE SMALL CELL CARCINOMA OF PROSTATE GLAND
C2009885|T047||CCS_10|FUSIFORM TYPE SMALL CELL CARCINOMA OF PROSTATE GLAND 
C2182974|T047||CCS_10|DUCT CARCINOMA, DESMOPLASTIC TYPE, OF PROSTATE GLAND 
C2182974|T047||CCS_10|DUCT CARCINOMA, DESMOPLASTIC TYPE, OF PROSTATE GLAND
C2145466|T047||CCS_10|TRANSITIONAL CELL CARCINOMA OF PROSTATE GLAND 
C2145466|T047||CCS_10|TRANSITIONAL CELL CARCINOMA OF PROSTATE GLAND
C2018609|T047||CCS_10|SPINDLE CELL TRANSITIONAL CELL CARCINOMA OF PROSTATE GLAND 
C2018609|T047||CCS_10|PROSTATE MALIGNANT CARCINOMA TRANSITIONAL CELL SPINDLE CELL
C2018609|T047||CCS_10|SPINDLE CELL TRANSITIONAL CELL CARCINOMA OF PROSTATE GLAND
C2212276|T047||CCS_10|PROSTATE GLAND MALIGNANT CARCINOMA SCHNEIDERIAN
C2212276|T047||CCS_10|SCHNEIDERIAN CARCINOMA OF PROSTATE GLAND
C2212276|T047||CCS_10|SCHNEIDERIAN CARCINOMA OF PROSTATE GLAND 
C2212277|T047||CCS_10|BASALOID CARCINOMA OF PROSTATE GLAND
C2212277|T047||CCS_10|BASALOID CARCINOMA OF PROSTATE GLAND 
C2075845|T047||CCS_10|CLOACOGENIC CARCINOMA OF PROSTATE GLAND 
C2075845|T047||CCS_10|CLOACOGENIC CARCINOMA OF PROSTATE GLAND
C2033335|T047||CCS_10|PROSTATE MALIGNANT CARCINOMA TRANSITIONAL CELL PAPILLARY
C2033335|T047||CCS_10|PAPILLARY TRANSITIONAL CELL CARCINOMA OF PROSTATE GLAND
C2033335|T047||CCS_10|PAPILLARY TRANSITIONAL CELL CARCINOMA OF PROSTATE GLAND 
C2212278|T047||CCS_10|MICROPAPILLARY TRANSITIONAL CELL CARCINOMA OF PROSTATE GLAND 
C2212278|T047||CCS_10|MICROPAPILLARY TRANSITIONAL CELL CARCINOMA OF PROSTATE GLAND
C2212279|T047||CCS_10|ADENOID CYSTIC CARCINOMA OF PROSTATE GLAND
C2212279|T047||CCS_10|ADENOID CYSTIC CARCINOMA OF PROSTATE GLAND 
C2138458|T047||CCS_10|CRIBRIFORM CARCINOMA OF PROSTATE GLAND 
C2138458|T047||CCS_10|CRIBRIFORM CARCINOMA OF PROSTATE GLAND
C2142686|T047||CCS_10|PROSTATE GLAND MALIGNANT CARCINOMA INTRACYSTIC
C2142686|T047||CCS_10|PROSTATE GLAND MALIGNANT CARCINOMA INTRACYSTIC 
C2212280|T047||CCS_10|ADENOSQUAMOUS CARCINOMA OF PROSTATE GLAND
C2212280|T047||CCS_10|ADENOSQUAMOUS CARCINOMA OF PROSTATE GLAND 
C2212281|T047||CCS_10|EPITHELIAL-MYOEPITHELIAL CARCINOMA OF PROSTATE GLAND
C2212281|T047||CCS_10|EPITHELIAL-MYOEPITHELIAL CARCINOMA OF PROSTATE GLAND 
C2212282|T047||CCS_10|MEDULLARY CARCINOMA OF PROSTATE GLAND
C2212282|T047||CCS_10|MEDULLARY CARCINOMA OF PROSTATE GLAND 
C2212283|T047||CCS_10|SCIRRHOUS ADENOCARCINOMA OF PROSTATE GLAND
C2212283|T047||CCS_10|SCIRRHOUS ADENOCARCINOMA OF PROSTATE GLAND 
C2212283|T047||CCS_10|PROSTATE GLAND MALIGNANT ADENOCARCINOMA SCIRRHOUS
C2037349|T047||CCS_10|SUPERFICIAL SPREADING ADENOCARCINOMA OF PROSTATE 
C2037349|T047||CCS_10|SUPERFICIAL SPREADING ADENOCARCINOMA OF PROSTATE
C2033129|T047||CCS_10|PAPILLARY ADENOCARCINOMA OF PROSTATE GLAND
C2033129|T047||CCS_10|PAPILLARY ADENOCARCINOMA OF PROSTATE GLAND 
C2189645|T047||CCS_10|VILLOUS ADENOCARCINOMA OF PROSTATE GLAND
C2189645|T047||CCS_10|VILLOUS ADENOCARCINOMA OF PROSTATE GLAND 
C2212285|T047||CCS_10|MUCINOUS ADENOCARCINOMA OF PROSTATE GLAND
C2212285|T047||CCS_10|MUCINOUS ADENOCARCINOMA OF PROSTATE GLAND 
C2212286|T047||CCS_10|MUCIN-PRODUCING ADENOCARCINOMA OF PROSTATE GLAND
C2212286|T047||CCS_10|MUCIN-PRODUCING ADENOCARCINOMA OF PROSTATE GLAND 
C2018507|T047||CCS_10|SPINDLE CELL SARCOMA OF PROSTATE GLAND 
C2018507|T047||CCS_10|SPINDLE CELL SARCOMA OF PROSTATE GLAND
C2011321|T047||CCS_10|GIANT CELL SARCOMA OF PROSTATE GLAND
C2011321|T047||CCS_10|GIANT CELL SARCOMA OF PROSTATE GLAND 
C2212292|T047||CCS_10|SMALL CELL SARCOMA OF PROSTATE GLAND 
C2212292|T047||CCS_10|SMALL CELL SARCOMA OF PROSTATE GLAND
C2212293|T047||CCS_10|EPITHELIOID SARCOMA OF PROSTATE GLAND 
C2212293|T047||CCS_10|EPITHELIOID SARCOMA OF PROSTATE GLAND
C2188144|T047||CCS_10|UNDIFFERENTIATED SARCOMA OF PROSTATE GLAND 
C2188144|T047||CCS_10|UNDIFFERENTIATED SARCOMA OF PROSTATE GLAND
C2142687|T047||CCS_10|DESMOPLASTIC SMALL ROUND CELL TUMOR OF PROSTATE GLAND
C2142687|T047||CCS_10|DESMOPLASTIC SMALL ROUND CELL TUMOR OF PROSTATE GLAND 
C2170822|T047||CCS_10|TUBULAR ADENOCARCINOMA OF PROSTATE GLAND
C2170822|T047||CCS_10|TUBULAR ADENOCARCINOMA OF PROSTATE GLAND 
C2212295|T047||CCS_10|FIBROMYXOSARCOMA OF PROSTATE GLAND
C2212295|T047||CCS_10|FIBROMYXOSARCOMA OF PROSTATE GLAND 
C2212296|T047||CCS_10|FASCIAL FIBROSARCOMA OF PROSTATE GLAND 
C2212296|T047||CCS_10|FASCIAL FIBROSARCOMA OF PROSTATE GLAND
C2142682|T047||CCS_10|INFANTILE FIBROSARCOMA OF PROSTATE GLAND
C2142682|T047||CCS_10|INFANTILE FIBROSARCOMA OF PROSTATE GLAND 
C2142689|T047||CCS_10|MALIGNANT SOLITARY FIBROUS TUMOR OF PROSTATE GLAND 
C2142689|T047||CCS_10|MALIGNANT SOLITARY FIBROUS TUMOR OF PROSTATE GLAND
C2168295|T047||CCS_10|LEIOMYOSARCOMA OF PROSTATE GLAND 
C2168295|T047||CCS_10|LEIOMYOSARCOMA OF PROSTATE GLAND
C2168263|T047||CCS_10|PROSTATE GLAND NEOPLASM MALIGNANT LEIOMYOSARCOMA EPITHELIOID
C2168263|T047||CCS_10|EPITHELIOID LEIOMYOSARCOMA OF PROSTATE GLAND 
C2168263|T047||CCS_10|EPITHELIOID LEIOMYOSARCOMA OF PROSTATE GLAND
C2212298|T047||CCS_10|MYXOID LEIOMYOSARCOMA OF PROSTATE GLAND 
C2212298|T047||CCS_10|MYXOID LEIOMYOSARCOMA OF PROSTATE GLAND
C1335518|T047||CCS_10|RHABDOMYOSARCOMA OF PROSTATE 
C1335518|T047||CCS_10|PROSTATE GLAND NEOPLASM MALIGNANT RHABDOMYOSARCOMA
C1335518|T047||CCS_10|RHABDOMYOSARCOMA OF PROSTATE
C1335518|T047||CCS_10|PROSTATE RHABDOMYOSARCOMA
C1335518|T047||CCS_10|RHABDOMYOSARCOMA OF THE PROSTATE
C2212299|T047||CCS_10|ADULT TYPE PLEOMORPHIC RHABDOMYOSARCOMA OF PROSTATE 
C2212299|T047||CCS_10|PROSTATE GLAND RHABDOMYOSARCOMA PLEOMORPHIC, ADULT TYPE
C2212299|T047||CCS_10|ADULT TYPE PLEOMORPHIC RHABDOMYOSARCOMA OF PROSTATE
C1335508|T047||CCS_10|PROSTATE GLAND RHABDOMYOSARCOMA EMBRYONAL
C1335508|T047||CCS_10|EMBRYONAL RHABDOMYOSARCOMA OF PROSTATE
C1335508|T047||CCS_10|EMBRYONAL RHABDOMYOSARCOMA OF PROSTATE 
C1335508|T047||CCS_10|EMBRYONAL RHABDOMYOSARCOMA OF THE PROSTATE
C1335508|T047||CCS_10|PROSTATE EMBRYONAL RHABDOMYOSARCOMA
C2018449|T047||CCS_10|SPINDLE CELL RHABDOMYOSARCOMA OF PROSTATE
C2018449|T047||CCS_10|PROSTATE GLAND RHABDOMYOSARCOMA SPINDLE CELL
C2018449|T047||CCS_10|SPINDLE CELL RHABDOMYOSARCOMA OF PROSTATE 
C2212300|T047||CCS_10|ALVEOLAR RHABDOMYOSARCOMA OF PROSTATE 
C2212300|T047||CCS_10|ALVEOLAR RHABDOMYOSARCOMA OF PROSTATE
C2212300|T047||CCS_10|PROSTATE GLAND RHABDOMYOSARCOMA ALVEOLAR
C2200364|T047||CCS_10|RHABDOMYOSARCOMA OF PROSTATE WITH GANGLIONIC DIFFERENTIATION
C2200364|T047||CCS_10|RHABDOMYOSARCOMA OF PROSTATE WITH GANGLIONIC DIFFERENTIATION 
C2200364|T047||CCS_10|PROSTATE RHABDOMYOSARCOMA WITH GANGLIONIC DIFFERENTIATION
C2212301|T047||CCS_10|ANGIOMYOSARCOMA OF PROSTATE GLAND 
C2212301|T047||CCS_10|ANGIOMYOSARCOMA OF PROSTATE GLAND
C2078063|T047||CCS_10|INTRADUCTAL PAPILLARY ADENOCARCINOMA OF PROSTATE WITH INVASION 
C2078063|T047||CCS_10|INTRADUCTAL PAPILLARY ADENOCARCINOMA OF PROSTATE WITH INVASION
C2212302|T047||CCS_10|PROSTATE GLAND RHABDOMYOSARCOMA MIXED TYPE
C2212302|T047||CCS_10|MIXED TYPE RHABDOMYOSARCOMA OF PROSTATE
C2212302|T047||CCS_10|MIXED TYPE RHABDOMYOSARCOMA OF PROSTATE 
C2212303|T047||CCS_10|EMBRYONAL CARCINOSARCOMA OF PROSTATE GLAND 
C2212303|T047||CCS_10|EMBRYONAL CARCINOSARCOMA OF PROSTATE GLAND
C2212304|T047||CCS_10|MALIGNANT MYOEPITHELIOMA OF PROSTATE GLAND
C2212304|T047||CCS_10|MALIGNANT MYOEPITHELIOMA OF PROSTATE GLAND 
C2217396|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE TNM STAGING 
C2217396|T047||CCS_10|MALIGNANT PROSTATE NEOPLASM TNM STAGING
C2217396|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE TNM STAGING
C2217396|T047||CCS_10|MALIGNANT PROSTATIC NEOPLASM TNM STAGING
C2217396|T047||CCS_10|PROSTATIC CANCER TNM STAGING
C2217396|T047||CCS_10|MALIGNANT TUMOR OF PROSTATE TNM STAGING
C2217394|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE STAGE III
C2217394|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE STAGE III 
C2217394|T047||CCS_10|MALIGNANT PROSTATIC NEOPLASM STAGE III
C2217394|T047||CCS_10|PROSTATIC CANCER STAGE III
C2217394|T047||CCS_10|MALIGNANT TUMOR OF PROSTATE STAGE III
C2217408|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE TNM STAGING HISTIOPATHIC GRADE (G) GX
C2217408|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE TNM STAGING HISTIOPATHIC GRADE (G) GX 
C2217408|T047||CCS_10|MALIGNANT PROSTATIC NEOPLASM GX
C2217408|T047||CCS_10|PROSTATIC CANCER TNM STAGING HISTIOPATHIC GRADE (G) GX
C2217408|T047||CCS_10|MALIGNANT TUMOR OF PROSTATE TNM STAGING HISTIOPATHIC GRADE (G) GX
C2217405|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE TNM STAGING HISTIOPATHIC GRADE (G) G1 
C2217405|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE TNM STAGING HISTIOPATHIC GRADE (G) G1
C2217405|T047||CCS_10|MALIGNANT PROSTATIC NEOPLASM G1
C2217405|T047||CCS_10|PROSTATIC CANCER TNM STAGING HISTIOPATHIC GRADE (G) G1
C2217405|T047||CCS_10|MALIGNANT TUMOR OF PROSTATE TNM STAGING HISTIOPATHIC GRADE (G) G1
C2217406|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE TNM STAGING HISTIOPATHIC GRADE (G) G2 
C2217406|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE TNM STAGING HISTIOPATHIC GRADE (G) G2
C2217406|T047||CCS_10|MALIGNANT PROSTATIC NEOPLASM G2
C2217406|T047||CCS_10|MALIGNANT TUMOR OF PROSTATE TNM STAGING HISTIOPATHIC GRADE (G) G2
C2217406|T047||CCS_10|PROSTATIC CANCER TNM STAGING HISTIOPATHIC GRADE (G) G2
C2217407|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE TNM STAGING HISTIOPATHIC GRADE (G) G3-4
C2217407|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE TNM STAGING HISTIOPATHIC GRADE (G) G3-4 
C2217407|T047||CCS_10|MALIGNANT PROSTATIC NEOPLASM G3-4
C2217407|T047||CCS_10|PROSTATIC CANCER TNM STAGING HISTIOPATHIC GRADE (G) G3-4
C2217407|T047||CCS_10|MALIGNANT TUMOR OF PROSTATE TNM STAGING HISTIOPATHIC GRADE (G) G3-4
C2217387|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE JEWETT STAGING SYSTEM
C2217387|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE JEWETT STAGING SYSTEM 
C2217387|T047||CCS_10|MALIGNANT PROSTATIC NEOPLASM JEWETT STAGING SYSTEM
C2217387|T047||CCS_10|MALIGNANT TUMOR OF PROSTATE JEWETT STAGING SYSTEM
C2217387|T047||CCS_10|PROSTATIC CANCER JEWETT STAGING SYSTEM
C2217388|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE JEWETT STAGING SYSTEM STAGE A 
C2217388|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE JEWETT STAGING SYSTEM STAGE A
C2217388|T047||CCS_10|MALIGNANT PROSTATIC NEOPLASM STAGE A
C2217388|T047||CCS_10|PROSTATIC CANCER JEWETT STAGING SYSTEM STAGE A
C2217388|T047||CCS_10|MALIGNANT TUMOR OF PROSTATE JEWETT STAGING SYSTEM STAGE A
C2217389|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE JEWETT STAGING SYSTEM STAGE B
C2217389|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE JEWETT STAGING SYSTEM STAGE B 
C2217389|T047||CCS_10|MALIGNANT PROSTATIC NEOPLASM STAGE B
C2217389|T047||CCS_10|PROSTATIC CANCER JEWETT STAGING SYSTEM STAGE B
C2217389|T047||CCS_10|MALIGNANT TUMOR OF PROSTATE JEWETT STAGING SYSTEM STAGE B
C2217390|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE JEWETT STAGING SYSTEM STAGE C
C2217390|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE JEWETT STAGING SYSTEM STAGE C 
C2217390|T047||CCS_10|MALIGNANT PROSTATIC NEOPLASM STAGE C
C2217390|T047||CCS_10|MALIGNANT TUMOR OF PROSTATE JEWETT STAGING SYSTEM STAGE C
C2217390|T047||CCS_10|PROSTATIC CANCER JEWETT STAGING SYSTEM STAGE C
C2217391|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE JEWETT STAGING SYSTEM STAGE D 
C2217391|T047||CCS_10|MALIGNANT NEOPLASM OF PROSTATE JEWETT STAGING SYSTEM STAGE D
C2217391|T047||CCS_10|MALIGNANT PROSTATIC NEOPLASM STAGE D
C2217391|T047||CCS_10|MALIGNANT TUMOR OF PROSTATE JEWETT STAGING SYSTEM STAGE D
C2217391|T047||CCS_10|PROSTATIC CANCER JEWETT STAGING SYSTEM STAGE D
C3469524|T047||CCS_10|PROSTATE CANCER SUSCEPTIBILITY
C3469524|T047||CCS_10|PROSTATE CANCER SUSCEPTIBILITY 
C3469524|T047||CCS_10|PROSTATE CANCER, SUSCEPTIBILITY TO
C1328504|T047||CCS_10|HORMONE REFRACTORY PROSTATE CANCER 
C1328504|T047||CCS_10|HORMONE REFRACTORY PROSTATE CANCER
C1328504|T047||CCS_10|HORMONE-REFRACTORY PROSTATE CANCER
C1328504|T047||CCS_10|PROSTATE GLAND MALIGNANT HORMONE REFRACTORY CANCER
C1328504|T047||CCS_10|HORMONE REFRACTORY PROSTATE CANCER 
C1328504|T047||CCS_10|HRPC
C3160891|T047||CCS_10|HORMONE-DEPENDENT PROSTATE CANCER
C1330959|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF PROSTATE 
C1330959|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF PROSTATE
C1330959|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF PROSTATE 
C0347001|T047||CCS_10|METASTATIC NEOPLASM TO THE PROSTATE
C0347001|T047||CCS_10|METASTASES TO PROSTATE
C0347001|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF PROSTATE
C0347001|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF PROSTATE 
C0347001|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO THE PROSTATE GLAND
C0347001|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM IN THE PROSTATE GLAND
C0347001|T047||CCS_10|CANCER METASTATIC TO PROSTATE
C0347001|T047||CCS_10|METASTASIS TO PROSTATE
C0347001|T047||CCS_10|METASTATIC TUMOR TO PROSTATE
C0347001|T047||CCS_10|METASTATIC TUMOUR TO PROSTATE
C0347001|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO PROSTATE
C0347001|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF PROSTATE 
C0347001|T047||CCS_10|METASTASES TO THE PROSTATE
C0347001|T047||CCS_10|METASTASIS TO THE PROSTATE
C0347001|T047||CCS_10|METASTATIC TUMOR TO THE PROSTATE
C1282482|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT NEOPLASM OF PROSTATE
C1282482|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT NEOPLASM OF PROSTATE 
C1282482|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOR OF PROSTATE 
C1282482|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOR OF PROSTATE
C1282482|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOUR OF PROSTATE
C4030346|T047||CCS_10|BIOPSY OF PROSTATE SHOWED CRIBRIFORM CARCINOMA 
C4030346|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA CRIBRIFORM
C4030346|T047||CCS_10|BIOPSY OF PROSTATE SHOWED CRIBRIFORM CARCINOMA
C4030340|T047||CCS_10|BIOPSY OF PROSTATE SHOWED GIANT CELL AND SPINDLE CELL CARCINOMA 
C4030340|T047||CCS_10|BIOPSY OF PROSTATE SHOWED GIANT CELL AND SPINDLE CELL CARCINOMA
C4030340|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA GIANT CELL AND SPINDLE CELL
C4030339|T047||CCS_10|BIOPSY OF PROSTATE SHOWED GIANT CELL CARCINOMA
C4030339|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA GIANT CELL
C4030339|T047||CCS_10|BIOPSY OF PROSTATE SHOWED GIANT CELL CARCINOMA 
C4030286|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT SMALL CELL TYPE 
C4030286|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT SMALL CELL TYPE
C4030304|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT FIBROSARCOMA SOLITARY FIBROUS TUMOR 
C4030304|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT FIBROSARCOMA SOLITARY FIBROUS TUMOR
C4030342|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA EPITHELIAL-MYOEPITHELIAL
C4030342|T047||CCS_10|BIOPSY OF PROSTATE SHOWED EPITHELIAL-MYOEPITHELIAL CARCINOMA
C4030342|T047||CCS_10|BIOPSY OF PROSTATE SHOWED EPITHELIAL-MYOEPITHELIAL CARCINOMA 
C4030293|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MYOSARCOMA RHABDOMYOSARCOMA MIXED TYPE
C4030293|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MYOSARCOMA RHABDOMYOSARCOMA MIXED TYPE 
C4030309|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CLEAR CELL TYPE
C4030309|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CLEAR CELL TYPE 
C4030355|T047||CCS_10|BIOPSY OF PROSTATE SHOWED BASAL CELL ADENOCARCINOMA
C4030355|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT ADENOCARCINOMA BASAL CELL
C4030355|T047||CCS_10|BIOPSY OF PROSTATE SHOWED BASAL CELL ADENOCARCINOMA 
C4030300|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MYOSARCOMA ANGIOMYOSARCOMA 
C4030300|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MYOSARCOMA ANGIOMYOSARCOMA
C4030348|T047||CCS_10|BIOPSY OF PROSTATE SHOWED CLEAR CELL ADENOCARCINOMA 
C4030348|T047||CCS_10|BIOPSY OF PROSTATE SHOWED CLEAR CELL ADENOCARCINOMA
C4030348|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT ADENOCARCINOMA CLEAR CELL
C4030333|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT ADENOCARCINOMA IN TUBULOVILLOUS ADENOMA 
C4030333|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT ADENOCARCINOMA IN TUBULOVILLOUS ADENOMA
C4030297|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MYOSARCOMA LEIOMYOSARCOMA MYXOID
C4030297|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MYOSARCOMA LEIOMYOSARCOMA MYXOID 
C4030275|T047||CCS_10|BIOPSY OF PROSTATE SHOWED SCIRRHOUS ADENOCARCINOMA 
C4030275|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT ADENOCARCINOMA SCIRRHOUS
C4030275|T047||CCS_10|BIOPSY OF PROSTATE SHOWED SCIRRHOUS ADENOCARCINOMA
C4030325|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA SMALL CELL FUSIFORM CELL
C4030325|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA SMALL CELL FUSIFORM CELL 
C4030307|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT FIBROSARCOMA FASCIAL 
C4030307|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT FIBROSARCOMA FASCIAL
C4030305|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT FIBROSARCOMA INFANTILE
C4030305|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT FIBROSARCOMA INFANTILE 
C4030302|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MARGINAL ZONE B-CELL LYMPHOMA
C4030302|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MARGINAL ZONE B-CELL LYMPHOMA 
C4030368|T047||CCS_10|BIOPSY OF PROSTATE SHOWED ACINAR CELL CYSTADENOCARCINOMA 
C4030368|T047||CCS_10|BIOPSY OF PROSTATE SHOWED ACINAR CELL CYSTADENOCARCINOMA
C4030368|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA ACINAR CELL CYSTADENOCARCINOMA
C4030295|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MYOSARCOMA RHABDOMYOSARCOMA ALVEOLAR 
C4030295|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MYOSARCOMA RHABDOMYOSARCOMA ALVEOLAR
C4030287|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT SARCOMA UNDIFFERENTIATED
C4030287|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT SARCOMA UNDIFFERENTIATED 
C4030283|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT ADENOCARCINOMA MUCINOUS
C4030283|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MUCINOUS ADENOCARCINOMA
C4030283|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MUCINOUS ADENOCARCINOMA 
C4030330|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA LARGE CELL WITH RHABDOID PHENOTYPE
C4030330|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA LARGE CELL WITH RHABDOID PHENOTYPE 
C4030288|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT SARCOMA SMALL CELL 
C4030288|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT SARCOMA SMALL CELL
C4030285|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT SPINDLE CELL TYPE 
C4030285|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT SPINDLE CELL TYPE
C4030277|T047||CCS_10|BIOPSY OF PROSTATE SHOWED PLEOMORPHIC CARCINOMA 
C4030277|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA PLEOMORPHIC
C4030277|T047||CCS_10|BIOPSY OF PROSTATE SHOWED PLEOMORPHIC CARCINOMA
C4030322|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA SQUAMOUS CELL LARGE CELL, NONKERAT 
C4030322|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA SQUAMOUS CELL LARGE CELL, NONKERAT
C4030312|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOSARCOMA 
C4030312|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOSARCOMA
C4030334|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA LARGE CELL NEUROENDOCRINE
C4030334|T047||CCS_10|BIOPSY OF PROSTATE SHOWED LARGE CELL NEUROENDOCRINE CARCINOMA 
C4030334|T047||CCS_10|BIOPSY OF PROSTATE SHOWED LARGE CELL NEUROENDOCRINE CARCINOMA
C4030298|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MYOSARCOMA LEIOMYOSARCOMA EPITHELIOID 
C4030298|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MYOSARCOMA LEIOMYOSARCOMA EPITHELIOID
C4030294|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MYOSARCOMA RHABDOMYOSARCOMA EMBRYONAL
C4030294|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MYOSARCOMA RHABDOMYOSARCOMA EMBRYONAL 
C4030271|T047||CCS_10|BIOPSY OF PROSTATE SHOWED SUPERFICIAL SPREADING ADENOCARCINOMA
C4030271|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT ADENOCARCINOMA SUPERFICIAL SPREADING
C4030271|T047||CCS_10|BIOPSY OF PROSTATE SHOWED SUPERFICIAL SPREADING ADENOCARCINOMA 
C4030267|T047||CCS_10|BIOPSY OF PROSTATE SHOWED VILLOUS ADENOCARCINOMA 
C4030267|T047||CCS_10|BIOPSY OF PROSTATE SHOWED VILLOUS ADENOCARCINOMA
C4030267|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT ADENOCARCINOMA VILLOUS
C4030323|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA SQUAMOUS CELL KERATINIZING
C4030323|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA SQUAMOUS CELL KERATINIZING 
C4030308|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT FIBROSARCOMA 
C4030308|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT FIBROSARCOMA
C4030363|T047||CCS_10|BIOPSY OF PROSTATE SHOWED ADENOCARCINOMA WITH METAPLASIA 
C4030363|T047||CCS_10|BIOPSY OF PROSTATE SHOWED ADENOCARCINOMA WITH METAPLASIA
C4030363|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT ADENOCARCINOMA WITH METAPLASIA
C4030344|T047||CCS_10|BIOPSY OF PROSTATE SHOWED DUCT CARCINOMA, DESMOPLASTIC TYPE 
C4030344|T047||CCS_10|BIOPSY OF PROSTATE SHOWED DUCT CARCINOMA, DESMOPLASTIC TYPE
C4030344|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA DUCT, DESMOPLASTIC TYPE
C4030296|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MYOSARCOMA RHABDOMYOSARCOMA
C4030296|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MYOSARCOMA RHABDOMYOSARCOMA 
C4030278|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA PAPILLARY
C4030278|T047||CCS_10|BIOPSY OF PROSTATE SHOWED PAPILLARY CARCINOMA 
C4030278|T047||CCS_10|BIOPSY OF PROSTATE SHOWED PAPILLARY CARCINOMA
C4030269|T047||CCS_10|BIOPSY OF PROSTATE SHOWED TUBULAR ADENOCARCINOMA
C4030269|T047||CCS_10|BIOPSY OF PROSTATE SHOWED TUBULAR ADENOCARCINOMA 
C4030269|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT ADENOCARCINOMA TUBULAR
C4030328|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA PSEUDOSARCOMATOUS
C4030328|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA PSEUDOSARCOMATOUS 
C4030318|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA SQUAMOUS CELL WITH HORN FORMATION
C4030318|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA SQUAMOUS CELL WITH HORN FORMATION 
C4030303|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT GIANT CELL TYPE
C4030303|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT GIANT CELL TYPE 
C4030356|T047||CCS_10|BIOPSY OF PROSTATE SHOWED ANAPLASTIC CARCINOMA 
C4030356|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA ANAPLASTIC
C4030356|T047||CCS_10|BIOPSY OF PROSTATE SHOWED ANAPLASTIC CARCINOMA
C4030331|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA EPITHELIOMA
C4030331|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA EPITHELIOMA 
C4030281|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MYOSARCOMA RHABDOMYOSARCOMA PLEOMORPHIC, ADULT TYPE
C4030281|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MYOSARCOMA RHABDOMYOSARCOMA PLEOMORPHIC, ADULT TYPE 
C4030279|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT ADENOCARCINOMA PAPILLARY
C4030279|T047||CCS_10|BIOPSY OF PROSTATE SHOWED PAPILLARY ADENOCARCINOMA
C4030279|T047||CCS_10|BIOPSY OF PROSTATE SHOWED PAPILLARY ADENOCARCINOMA 
C4030268|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA VERRUCOUS
C4030268|T047||CCS_10|BIOPSY OF PROSTATE SHOWED VERRUCOUS CARCINOMA
C4030268|T047||CCS_10|BIOPSY OF PROSTATE SHOWED VERRUCOUS CARCINOMA 
C4030301|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MYOSARCOMA
C4030301|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MYOSARCOMA 
C4030299|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MYOSARCOMA LEIOMYOSARCOMA
C4030299|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MYOSARCOMA LEIOMYOSARCOMA 
C4030292|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MYOSARCOMA RHABDOMYOSARCOMA SPINDLE CELL
C4030292|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT MYOSARCOMA RHABDOMYOSARCOMA SPINDLE CELL 
C4030291|T047||CCS_10|BIOPSY OF PROSTATE SHOWED A MALIGNANT NEOPLASM
C4030291|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT NEOPLASM 
C4030291|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT NEOPLASM
C4030290|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT SARCOMA 
C4030290|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT SARCOMA
C4030273|T047||CCS_10|BIOPSY OF PROSTATE SHOWED SPINDLE CELL SARCOMA
C4030273|T047||CCS_10|BIOPSY OF PROSTATE SHOWED SPINDLE CELL SARCOMA 
C4030273|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT SARCOMA SPINDLE CELL
C4030324|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA SQUAMOUS CELL ADENOID
C4030324|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA SQUAMOUS CELL ADENOID 
C4030317|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA TRANSITIONAL CELL MICROPAPILLARY 
C4030317|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA TRANSITIONAL CELL MICROPAPILLARY
C4030338|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA GLASSY CELL
C4030338|T047||CCS_10|BIOPSY OF PROSTATE SHOWED GLASSY CELL CARCINOMA
C4030338|T047||CCS_10|BIOPSY OF PROSTATE SHOWED GLASSY CELL CARCINOMA 
C4030276|T047||CCS_10|BIOPSY OF PROSTATE SHOWED POLYGONAL CELL CARCINOMA
C4030276|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA POLYGONAL CELL
C4030276|T047||CCS_10|BIOPSY OF PROSTATE SHOWED POLYGONAL CELL CARCINOMA 
C4030274|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA SPINDLE CELL
C4030274|T047||CCS_10|BIOPSY OF PROSTATE SHOWED SPINDLE CELL CARCINOMA
C4030274|T047||CCS_10|BIOPSY OF PROSTATE SHOWED SPINDLE CELL CARCINOMA 
C4030321|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA SQUAMOUS CELL MICROINVASIVE
C4030321|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA SQUAMOUS CELL MICROINVASIVE 
C4030313|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA WITH OSTEOCLAST-LIKE CELLS 
C4030313|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA WITH OSTEOCLAST-LIKE CELLS
C4030280|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MYOSARCOMA RHABDOMYOSARCOMA WITH GANGLIONIC DIFFERENTIATION
C4030280|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MYOSARCOMA RHABDOMYOSARCOMA WITH GANGLIONIC DIFFERENTIATION 
C4030289|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT SARCOMA GIANT CELL 
C4030289|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT SARCOMA GIANT CELL
C4030327|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA SCHNEIDERIAN 
C4030327|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA SCHNEIDERIAN
C4030311|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOSARCOMA EMBRYONAL TYPE
C4030311|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOSARCOMA EMBRYONAL TYPE 
C4030310|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOSARCOMA MYOEPITHELIOMA 
C4030310|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOSARCOMA MYOEPITHELIOMA
C4030345|T047||CCS_10|BIOPSY OF PROSTATE SHOWED DESMOPLASTIC SMALL ROUND CELL SARCOMA 
C4030345|T047||CCS_10|BIOPSY OF PROSTATE SHOWED DESMOPLASTIC SMALL ROUND CELL SARCOMA
C4030345|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT SARCOMA DESMOPLASTIC SMALL ROUND CELL
C4030272|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA SQUAMOUS CELL
C4030272|T047||CCS_10|BIOPSY OF PROSTATE SHOWED SQUAMOUS CELL CARCINOMA
C4030272|T047||CCS_10|BIOPSY OF PROSTATE SHOWED SQUAMOUS CELL CARCINOMA 
C4030270|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA TRANSITIONAL CELL
C4030270|T047||CCS_10|BIOPSY OF PROSTATE SHOWED TRANSITIONAL CELL CARCINOMA 
C4030270|T047||CCS_10|BIOPSY OF PROSTATE SHOWED TRANSITIONAL CELL CARCINOMA
C4030316|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA TRANSITIONAL CELL PAPILLARY
C4030316|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA TRANSITIONAL CELL PAPILLARY 
C4030358|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA ADENOSQUAMOUS
C4030358|T047||CCS_10|BIOPSY OF PROSTATE SHOWED ADENOSQUAMOUS CARCINOMA
C4030358|T047||CCS_10|BIOPSY OF PROSTATE SHOWED ADENOSQUAMOUS CARCINOMA 
C4030357|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT ADENOCARCINOMA ALVEOLAR
C4030357|T047||CCS_10|BIOPSY OF PROSTATE SHOWED ALVEOLAR ADENOCARCINOMA 
C4030357|T047||CCS_10|BIOPSY OF PROSTATE SHOWED ALVEOLAR ADENOCARCINOMA
C4030341|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT SARCOMA EPITHELIOID
C4030341|T047||CCS_10|BIOPSY OF PROSTATE SHOWED EPITHELIOID SARCOMA 
C4030341|T047||CCS_10|BIOPSY OF PROSTATE SHOWED EPITHELIOID SARCOMA
C4030332|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT ADENOCARCINOMA IN VILLOUS ADENOMA 
C4030332|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT ADENOCARCINOMA IN VILLOUS ADENOMA
C4030319|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA SQUAMOUS CELL SPINDLE CELL 
C4030319|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA SQUAMOUS CELL SPINDLE CELL
C4030314|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA UNDIFFERENTIATED
C4030314|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA UNDIFFERENTIATED 
C4030359|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA ADENOID CYSTIC
C4030359|T047||CCS_10|BIOPSY OF PROSTATE SHOWED ADENOID CYSTIC CARCINOMA 
C4030359|T047||CCS_10|BIOPSY OF PROSTATE SHOWED ADENOID CYSTIC CARCINOMA
C4030354|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA BASALOID
C4030354|T047||CCS_10|BIOPSY OF PROSTATE SHOWED BASALOID CARCINOMA 
C4030354|T047||CCS_10|BIOPSY OF PROSTATE SHOWED BASALOID CARCINOMA
C4030335|T047||CCS_10|BIOPSY OF PROSTATE SHOWED LARGE CELL CARCINOMA
C4030335|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA LARGE CELL
C4030335|T047||CCS_10|BIOPSY OF PROSTATE SHOWED LARGE CELL CARCINOMA 
C4030366|T047||CCS_10|BIOPSY OF PROSTATE SHOWED ADENOCARCINOMA INTRADUCTAL PAPILLARY, WITH INVASION
C4030366|T047||CCS_10|BIOPSY OF PROSTATE SHOWED ADENOCARCINOMA INTRADUCTAL PAPILLARY, WITH INVASION 
C4030284|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MEDULLARY CARCINOMA
C4030284|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA MEDULLARY
C4030284|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MEDULLARY CARCINOMA 
C4030282|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT ADENOCARCINOMA MUCIN-PRODUCING
C4030282|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MUCIN-PRODUCING ADENOCARCINOMA
C4030282|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MUCIN-PRODUCING ADENOCARCINOMA 
C4030369|T047||CCS_10|BIOPSY OF PROSTATE SHOWED ACINAR CELL CARCINOMA
C4030369|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA ACINAR CELL
C4030369|T047||CCS_10|BIOPSY OF PROSTATE SHOWED ACINAR CELL CARCINOMA 
C4030347|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA CLOACOGENIC
C4030347|T047||CCS_10|BIOPSY OF PROSTATE SHOWED CLOACOGENIC CARCINOMA
C4030347|T047||CCS_10|BIOPSY OF PROSTATE SHOWED CLOACOGENIC CARCINOMA 
C4030329|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA PAPILLARY SQUAMOUS CELL 
C4030329|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA PAPILLARY SQUAMOUS CELL
C4030320|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA SQUAMOUS CELL SMALL CELL, NONKERAT 
C4030320|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA SQUAMOUS CELL SMALL CELL, NONKERAT
C4030315|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA TRANSITIONAL CELL SPINDLE CELL
C4030315|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT CARCINOMA TRANSITIONAL CELL SPINDLE CELL 
C4030306|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT FIBROSARCOMA FIBROMYXOSARCOMA
C4030306|T047||CCS_10|BIOPSY OF PROSTATE SHOWED MALIGNANT FIBROSARCOMA FIBROMYXOSARCOMA 
C1282496|T047||CCS_10|METASTASIS FROM MALIGNANT NEOPLASM OF PROSTATE 
C1282496|T047||CCS_10|METASTASIS FROM MALIGNANT NEOPLASM OF PROSTATE
C1282496|T047||CCS_10|CANCER OF THE PROSTATE WITH METASTASIS
C1282496|T047||CCS_10|METASTATIC PROSTATE CANCER
C1282496|T047||CCS_10|METASTASIS FROM MALIGNANT TUMOR OF PROSTATE
C1282496|T047||CCS_10|METASTASIS FROM MALIGNANT TUMOR OF PROSTATE 
C1282496|T047||CCS_10|METASTASIS FROM MALIGNANT TUMOUR OF PROSTATE
C4081803|T047||CCS_10|PROSTATE CANCER METASTATIC TO EYE 
C4081803|T047||CCS_10|PROSTATE CANCER METASTATIC TO EYE
C1302530|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF PROSTATE GLAND
C1302530|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF PROSTATE GLAND 
C1302530|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF PROSTATE 
C1302530|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF PROSTATE
C1302530|T047||CCS_10|PROSTATE SQUAMOUS CELL CARCINOMA
C1302530|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE PROSTATE
C0154088|T047||CCS_10|CARCINOMA IN SITU OF PROSTATE
C0154088|T047||CCS_10|CARCINOMA IN SITU OF PROSTATE GLAND 
C0154088|T047||CCS_10|CARCINOMA IN SITU OF PROSTATE GLAND
C0154088|T047||CCS_10|CA IN SITU PROSTATE
C0154088|T047||CCS_10|CIS - CARCINOMA IN SITU OF PROSTATE
C0154088|T047||CCS_10|CANCER IN SITU OF PROSTATE
C0154088|T047||CCS_10|CIS (CARCINOMA IN SITU) OF PROSTATE
C0154088|T047||CCS_10|CARCINOMA IN SITU OF PROSTATE 
C0154088|T047||CCS_10|PIN III
C0154088|T047||CCS_10|PROSTATIC INTRAEPITHELIAL NEOPLASIA, GRADE III
C0154088|T047||CCS_10|ADENOCARCINOMA IN SITU OF PROSTATE
C0154088|T047||CCS_10|ADENOCARCINOMA IN SITU OF THE PROSTATE
C0154088|T047||CCS_10|GRADE 3 PIN
C0154088|T047||CCS_10|GRADE 3 PROSTATIC INTRAEPITHELIAL NEOPLASIA
C0154088|T047||CCS_10|GRADE III PIN
C0154088|T047||CCS_10|GRADE III PROSTATIC INTRAEPITHELIAL NEOPLASIA
C0154088|T047||CCS_10|PROSTATE ADENOCARCINOMA IN SITU
C1386259|T047||CCS_10|ENDOMETRIOID; ADENOCARCINOMA, UNSPECIFIED SITE, MALE
C1386259|T047||CCS_10|ADENOCARCINOMA; ENDOMETRIOID, UNSPECIFIED SITE, MALE
C1391907|T047||CCS_10|CARCINOMA; ENDOMETRIOID, UNSPECIFIED SITE, MALE
C1391907|T047||CCS_10|ENDOMETRIOID; CARCINOMA, UNSPECIFIED SITE, MALE
C1394298|T047||CCS_10|CYSTADENOCARCINOMA; ENDOMETRIOID, UNSPECIFIED SITE, MALE
C1394298|T047||CCS_10|ENDOMETRIOID; CYSTADENOCARCINOMA, UNSPECIFIED SITE, MALE
C0279882|T047||CCS_10|CELLULAR DIAGNOSIS, PROSTATE CANCER
C0279882|T047||CCS_10|PROSTATE CANCER CELLULAR DIAGNOSIS
C0280280|T047||CCS_10|STAGE, PROSTATE CANCER
C0280280|T047||CCS_10|PROSTATE CANCER STAGE
C1335514|T047||CCS_10|EXTRAMEDULLARY MYELOID NEOPLASM OF PROSTATE
C1335514|T047||CCS_10|EXTRAMEDULLARY MYELOID NEOPLASM OF THE PROSTATE
C1335514|T047||CCS_10|EXTRAMEDULLARY MYELOID TUMOR OF PROSTATE
C1335514|T047||CCS_10|EXTRAMEDULLARY MYELOID TUMOR OF THE PROSTATE
C1335514|T047||CCS_10|PROSTATE EXTRAMEDULLARY MYELOID NEOPLASM
C1335514|T047||CCS_10|PROSTATE EXTRAMEDULLARY MYELOID TUMOR
C1335514|T047||CCS_10|PROSTATE MYELOID SARCOMA
C1335514|T047||CCS_10|PROSTATIC CHLOROMA
C1335514|T047||CCS_10|PROSTATIC EXTRAMEDULLARY MYELOID NEOPLASM
C1335514|T047||CCS_10|PROSTATIC EXTRAMEDULLARY MYELOID TUMOR
C1335514|T047||CCS_10|PROSTATIC MYELOID SARCOMA
C0238393|T047||CCS_10|PROSTATE SARCOMA
C0238393|T047||CCS_10|SARCOMA OF PROSTATE
C0238393|T047||CCS_10|SARCOMA OF THE PROSTATE
C1334615|T047||CCS_10|MALIGNANT PHYLLODES TUMOR OF PROSTATE
C1334615|T047||CCS_10|PHYLLODES TUMOR OF THE PROSTATE
C1334615|T047||CCS_10|MALIGNANT PHYLLODES NEOPLASM OF PROSTATE
C1334615|T047||CCS_10|MALIGNANT PHYLLODES NEOPLASM OF THE PROSTATE
C1334615|T047||CCS_10|MALIGNANT PHYLLODES TUMOR OF THE PROSTATE
C1334615|T047||CCS_10|MALIGNANT PROSTATE PHYLLODES NEOPLASM
C1334615|T047||CCS_10|MALIGNANT PROSTATE PHYLLODES TUMOR
C1335512|T047||CCS_10|PRIMARY PROSTATE LYMPHOMA
C1335512|T047||CCS_10|LYMPHOMA OF PROSTATE
C1335512|T047||CCS_10|LYMPHOMA OF THE PROSTATE
C1335512|T047||CCS_10|PROSTATE LYMPHOMA
C1276489|T047||CCS_10|T3A: PROSTATE TUMOR WITH EXTRACAPSULAR EXTENSION (UNILATERAL OR BILATERAL) 
C1276489|T047||CCS_10|T3A: PROSTATE TUMOR WITH EXTRACAPSULAR EXTENSION (UNILATERAL OR BILATERAL)
C1276489|T047||CCS_10|T3A: PROSTATE TUMOUR WITH EXTRACAPSULAR EXTENSION (UNILATERAL OR BILATERAL)
C1276489|T047||CCS_10|T3A: PROSTATE TUMOR WITH EXTRACAPSULAR EXTENSION (UNILATERAL OR BILATERAL) (TUMOR STAGING)
C1720586|T047||CCS_10|EXTRAPROSTATIC EXTENSION OF TUMOR PRESENT, NON-FOCAL 
C1720586|T047||CCS_10|EXTRAPROSTATIC EXTENSION OF TUMOR PRESENT, NON-FOCAL
C1720586|T047||CCS_10|EXTRAPROSTATIC EXTENSION OF TUMOUR PRESENT, NON-FOCAL
C1300585|T047||CCS_10|SMALL CELL CARCINOMA OF PROSTATE GLAND 
C1300585|T047||CCS_10|SMALL CELL CARCINOMA OF PROSTATE GLAND
C1300585|T047||CCS_10|PROSTATE SMALL CELL NEC
C1300585|T047||CCS_10|PROSTATE SMALL CELL NEUROENDOCRINE CARCINOMA
C1300585|T047||CCS_10|OAT CELL CARCINOMA OF PROSTATE
C1300585|T047||CCS_10|SMALL CELL CARCINOMA OF PROSTATE 
C1300585|T047||CCS_10|SMALL CELL CARCINOMA OF PROSTATE
C1300585|T047||CCS_10|OAT CELL CARCINOMA OF THE PROSTATE
C1300585|T047||CCS_10|PROSTATE OAT CELL CARCINOMA
C1300585|T047||CCS_10|PROSTATE SMALL CELL CARCINOMA
C1300585|T047||CCS_10|SMALL CELL CARCINOMA OF THE PROSTATE
C1276487|T047||CCS_10|T2A: PROSTATE TUMOR INVOLVES ONE LOBE 
C1276487|T047||CCS_10|T2A: PROSTATE TUMOR INVOLVES ONE LOBE
C1276487|T047||CCS_10|T2A: PROSTATE TUMOUR INVOLVES ONE LOBE
C1276487|T047||CCS_10|T2A: PROSTATE TUMOR INVOLVES ONE LOBE (TUMOR STAGING)
C0349672|T047||CCS_10|ENDOMETRIOID CARCINOMA OF PROSTATE
C0349672|T047||CCS_10|PROSTATE GLAND MALIGNANT CARCINOMA ENDOMETRIOID
C0349672|T047||CCS_10|ENDOMETRIOID CARCINOMA OF PROSTATE 
C0349672|T047||CCS_10|ENDOMETRIOID CARCINOMA OF PROSTATE 
C0349672|T047||CCS_10|DUCTAL ADENOCARCINOMA OF PROSTATE
C0349672|T047||CCS_10|DUCTAL ADENOCARCINOMA OF THE PROSTATE
C0349672|T047||CCS_10|ENDOMETRIOID ADENOCARCINOMA OF PROSTATE
C0349672|T047||CCS_10|ENDOMETRIOID ADENOCARCINOMA OF THE PROSTATE
C0349672|T047||CCS_10|ENDOMETRIOID CARCINOMA OF THE PROSTATE
C0349672|T047||CCS_10|PROSTATE DUCTAL ADENOCARCINOMA
C0349672|T047||CCS_10|PROSTATE ENDOMETRIOID ADENOCARCINOMA
C0349672|T047||CCS_10|PROSTATE ENDOMETRIOID CARCINOMA
C0349672|T047||CCS_10|PROSTATIC ENDOMETRIOID CARCINOMA
C1276488|T047||CCS_10|T3: PROSTATE TUMOR EXTENDS THROUGH THE PROSTATIC CAPSULE 
C1276488|T047||CCS_10|T3: PROSTATE TUMOR EXTENDS THROUGH THE PROSTATIC CAPSULE
C1276488|T047||CCS_10|T3: PROSTATE TUMOUR EXTENDS THROUGH THE PROSTATIC CAPSULE
C1276488|T047||CCS_10|T3: PROSTATE TUMOR EXTENDS THROUGH THE PROSTATIC CAPSULE (TUMOR STAGING)
C1276626|T047||CCS_10|T2: TUMOR CONFINED WITHIN THE PROSTATE 
C1276626|T047||CCS_10|T2: TUMOR CONFINED WITHIN THE PROSTATE
C1276626|T047||CCS_10|T2: TUMOUR CONFINED WITHIN THE PROSTATE
C1276626|T047||CCS_10|T2: TUMOR CONFINED WITHIN THE PROSTATE (TUMOR STAGING)
C0392920|T047||CCS_10|CANCER CHEMOTHERAPY
C0392920|T047||CCS_10|CHEMOTHERAPY REGIMEN
C0392920|T047||CCS_10|CHEMOTHERAPEUTICS REGIMEN
C0392920|T047||CCS_10|CHEMOTHERAPEUTICS REGIMEN 
C0392920|T047||CCS_10|NEOPLASM/CANCER CHEMOTHERAPY
C0392920|T047||CCS_10|NEOPLASM CHEMOTHERAPY
C0392920|T047||CCS_10|CHEMOTHERAPY
C0392920|T047||CCS_10|CANCER CHEMOTHERAPY (REGIME/THERAPY)
C0392920|T047||CCS_10|CHEMOTHERAPY 
C0392920|T047||CCS_10|CANCER CHEMOTHERAPY REGIMEN
C0392920|T047||CCS_10|ANTINEOPLASTIC CHEMOTHERAPY REGIMEN 
C0392920|T047||CCS_10|ANTINEOPLASTIC CHEMOTHERAPY REGIMEN
C0392920|T047||CCS_10|NEOPLASM/CANCER PHARMACOTHERAPY
C0392920|T047||CCS_10|NEOPLASM PHARMACOTHERAPY
C0392920|T047||CCS_10|CANCER; CHEMOTHERAPY
C0392920|T047||CCS_10|CHEMOTHERAPY; CANCER
C0392920|T047||CCS_10|CHEMOTHERAPY; NEOPLASM
C0392920|T047||CCS_10|NEOPLASM; CHEMOTHERAPY
C0392920|T047||CCS_10|CHEMOTHERAPY, NOS
C0392920|T047||CCS_10|ANTINEOPLASTIC CHEMOTHERAPY REGIMEN (REGIME/THERAPY)
C0280024|T047||CCS_10|MERCAPTOPURINE/METHOTREXATE/PREDNISOLONE/VINCRISTINE
C0280024|T047||CCS_10|POMP
C0280024|T047||CCS_10|MP/MTX/PRDL/VCR
C0280024|T047||CCS_10|MERCAPTOPURINE/METHOTREXATE/PREDNISOLONE/VINCRISTINE PROTOCOL
C0280075|T047||CCS_10|MERCAPTOPURINE/METHOTREXATE/METHYLPREDNISOLONE/VINCRISTINE
C0280075|T047||CCS_10|POMP
C0280075|T047||CCS_10|MEPRDL/MP/MTX/VCR
C0280075|T047||CCS_10|MERCAPTOPURINE/METHOTREXATE/METHYLPREDNISOLONE/VINCRISTINE PROTOCOL
C0280580|T047||CCS_10|DOXORUBICIN/FLUOROURACIL
C0280580|T047||CCS_10|DOX/5-FU
C0280580|T047||CCS_10|DOXORUBICIN/FLUOROURACIL PROTOCOL
C0280593|T047||CCS_10|DOXORUBICIN/FLUOROURACIL/SEMUSTINE
C0280593|T047||CCS_10|FAME
C0280593|T047||CCS_10|DOX/5-FU/MECCNU
C0280593|T047||CCS_10|DOXORUBICIN/FLUOROURACIL/SEMUSTINE PROTOCOL
C0338272|T047||CCS_10|CYCLOPHOSPHAMIDE/LOSOXANTRONE
C0338272|T047||CCS_10|CTX/DUP-941
C2045825|T047||CCS_10|CHEMOTHERAPEUTICS REGIMEN FIRST LINE OF TREATMENT
C2045825|T047||CCS_10|CHEMOTHERAPEUTICS REGIMEN FIRST LINE OF TREATMENT 
C2045828|T047||CCS_10|CHEMOTHERAPEUTICS REGIMEN SECOND LINE OF TREATMENT
C2045828|T047||CCS_10|CHEMOTHERAPEUTICS REGIMEN SECOND LINE OF TREATMENT 
C2045827|T047||CCS_10|ORAL CHEMOTHERAPEUTICS REGIMEN
C2045827|T047||CCS_10|ORAL CHEMOTHERAPEUTICS REGIMEN 
C2045826|T047||CCS_10|INTRAVENOUS CHEMOTHERAPEUTICS REGIMEN
C2045826|T047||CCS_10|INTRAVENOUS CHEMOTHERAPEUTICS REGIMEN 
C3179010|T047||CCS_10|INDUCTION CHEMOTHERAPY
C3179010|T047||CCS_10|CHEMOTHERAPY, INDUCTION
C3179010|T047||CCS_10|CHEMOTHERAPIES, INDUCTION
C3179010|T047||CCS_10|INDUCTION CHEMOTHERAPIES
C3179010|T047||CCS_10|INDUCTION CHEMOTHERAPY 
C0374470|T047||CCS_10|CHEMO INTRALESIONAL OVER 7
C0374470|T047||CCS_10|INTRALESIONAL CHEMOTHERAPY ADMINISTRATION FOR MORE THAN 7 LESIONS
C0374470|T047||CCS_10|INTRALESIONAL CHEMOTHERAPY ADMINISTRATION FOR MORE THAN 7 LESIONS 
C0374470|T047||CCS_10|CHEMOTHERAPY ADMINISTRATION INTRALESIONAL >7
C0374470|T047||CCS_10|CHEMOTHERAPY ADMINISTRATION; INTRALESIONAL, MORE THAN 7 LESIONS
C1302181|T047||CCS_10|CHEMOTHERAPEUTICS REGIMEN CYCLE 
C1302181|T047||CCS_10|CHEMOTHERAPEUTICS REGIMEN CYCLE
C1302181|T047||CCS_10|CHEMOTHERAPY CYCLE
C1302181|T047||CCS_10|CHEMOTHERAPY CYCLE 
C1302181|T047||CCS_10|CHEMOTHERAPY CYCLE (REGIME/THERAPY)
C0413365|T047||CCS_10|INTRAVENOUS CHEMOTHERAPY
C0413365|T047||CCS_10|INTRAVENOUS CHEMOTHERAPY 
C0413365|T047||CCS_10|INTRAVENOUS CHEMOTHERAPY 
C0260835|T047||CCS_10|CHEMOTHERAPY FOLLOW-UP 
C0260835|T047||CCS_10|CHEMOTHERAPY FOLLOW-UP
C0260835|T047||CCS_10|CHEMOTHERAPY FOLLOW-UP (REGIME/THERAPY)
C0199957|T047||CCS_10|CHEMOTHERAPY ADMINISTRATION, SUBCUTANEOUS, WITH LOCAL ANESTHESIA
C0199957|T047||CCS_10|CHEMOTHERAPY ADMINISTRATION, SUBCUTANEOUS, WITH LOCAL ANAESTHESIA
C0199957|T047||CCS_10|CHEMOTHERAPY ADMINISTRATION, SUBCUTANEOUS, WITH LOCAL ANESTHESIA 
C0199957|T047||CCS_10|CHEMOTHERAPY ADMINISTRATION, SUBCUTANEOUS, WITH LOCAL ANESTHESIA (REGIME/THERAPY)
C0198526|T047||CCS_10|CHEMOTHERAPY ADMINISTRATION INTO PERITONEAL CAVITY REQUIRING PARACENTESIS
C0198526|T047||CCS_10|CHEMOTHERAPY ADMINISTRATION INTO PERITONEAL CAVITY REQUIRING PARACENTESIS 
C0198526|T047||CCS_10|CHEMOTHERAPY ADMINISTRATION INTO PERITONEAL CAVITY REQUIRING PARACENTESIS (REGIME/THERAPY)
C0189560|T047||CCS_10|CHEMOTHERAPY ADMINISTRATION INTO PLEURAL CAVITY, REQUIRING AND INCLUDING THORACENTESIS
C0189560|T047||CCS_10|CHEMOTHERAPY ADMINISTRATION INTO PLEURAL CAVITY REQUIRING THORACENTESIS 
C0189560|T047||CCS_10|CHEMOTHERAPY INTRACAVITARY
C0189560|T047||CCS_10|CHEMOTHERAPY ADMINISTRATION INTO PLEURAL CAVITY WITH THORACENTESIS
C0189560|T047||CCS_10|CHEMOTHERAPY ADMINISTRATION INTO PLEURAL CAVITY REQUIRING THORACENTESIS
C0189560|T047||CCS_10|CHEMOTHERAPY ADMINISTRATION INTO PLEURAL CAVITY REQUIRING THORACENTESIS (REGIME/THERAPY)
C0189560|T047||CCS_10|CHEMOTX ADMN PLEURAL CAVITY REQ&W/THORACNTS
C0419073|T047||CCS_10|ORAL CYTOTOXIC DRUG THERAPY
C0419073|T047||CCS_10|ORAL CHEMOTHERAPY
C0419073|T047||CCS_10|ORAL CHEMOTHERAPY 
C0419073|T047||CCS_10|ORAL CHEMOTHERAPY (REGIME/THERAPY)
C1276154|T047||CCS_10|AMBULATORY CHEMOTHERAPY 
C1276154|T047||CCS_10|AMBULATORY CHEMOTHERAPY
C1276154|T047||CCS_10|AMBULATORY CHEMOTHERAPY ADMINISTRATION 
C1276154|T047||CCS_10|CHEMOTHERAPY ADMINISTRATION AMBULATORY
C1276154|T047||CCS_10|AMBULATORY CHEMOTHERAPY ADMINISTRATION
C1276154|T047||CCS_10|AMBULATORY CHEMOTHERAPY (REGIME/THERAPY)
C3695058|T047||CCS_10|CHEMOTHERAPEUTICS REGIMEN INTRACAVITARY 
C3695058|T047||CCS_10|CHEMOTHERAPEUTICS REGIMEN INTRACAVITARY
C3665477|T047||CCS_10|CHEMOTHERAPY REGIMEN OR AGENT COMBINATION
C3665477|T047||CCS_10|COMBINATION CHEMOTHERAPY REGIMEN
C0476658|T047||CCS_10|CHEMOTHERAPY SESSION FOR NEOPLASM
C0476658|T047||CCS_10|[V]CHEMOTHERAPY SESSION FOR NEOPLASM (CONTEXT-DEPENDENT CATEGORY)
C0476658|T047||CCS_10|ENCOUNTER FOR ANTINEOPLASTIC CHEMOTHERAPY AND IMMUNOTHERAPY
C0476658|T047||CCS_10|[V]CHEMOTHERAPY SESSION FOR NEOPLASM
C0476658|T047||CCS_10|[V]CHEMOTHERAPY SESSION FOR NEOPLASM 
C0476658|T047||CCS_10|ENCOUNTER DUE TO CHEMOTHERAPY SESSION FOR NEOPLASM
C0476658|T047||CCS_10|ENCOUNTER OR ADMISSION FOR CHEMOTHERAPY
C0178200|T047||CCS_10|INJECT CA CHEMOTHER NEC
C0178200|T047||CCS_10|INJECTION OR INFUSION OF CANCER CHEMOTHERAPEUTIC SUBSTANCE
C0178200|T047||CCS_10|INJECTION OR INFUSION OF ANTINEOPLASTIC AGENT
C0374469|T047||CCS_10|INTRALESIONAL CHEMOTHERAPY ADMINISTRATION UP TO AND INCLUDING 7 LESIONS
C0374469|T047||CCS_10|INTRALESIONAL CHEMOTHERAPY ADMINISTRATION UP TO AND INCLUDING 7 LESIONS 
C0374469|T047||CCS_10|CHEMO INTRALESIONAL UP TO 7
C0374469|T047||CCS_10|CHEMOTHERAPY ADMINISTRATION INTRALESIONAL </7
C0374469|T047||CCS_10|CHEMOTHERAPY ADMINISTRATION; INTRALESIONAL, UP TO AND INCLUDING 7 LESIONS
C0374473|T047||CCS_10|CHEMOTHERAPY INTO CNS
C0374473|T047||CCS_10|CHEMOTX ADMN CNS REQ SPINAL PUNCTURE
C0374473|T047||CCS_10|CHEMOTHERAPY ADMINISTRATION, INTO CNS (EG, INTRATHECAL), REQUIRING AND INCLUDING SPINAL PUNCTURE
C0199944|T047||CCS_10|ORAL CHEMOTHERAPEUTICS REGIMEN FOR MALIGNANT NEOPLASM 
C0199944|T047||CCS_10|ORAL CHEMOTHERAPEUTICS REGIMEN FOR MALIGNANT NEOPLASM
C0199944|T047||CCS_10|CHEMOTHERAPEUTICS REGIMEN ORAL FOR MALIGNANT NEOPLASM
C0199944|T047||CCS_10|ORAL CHEMOTHERAPY FOR MALIGNANT NEOPLASM
C0199944|T047||CCS_10|ORAL CHEMOTHERAPY FOR MALIGNANT NEOPLASM 
C0199944|T047||CCS_10|ORAL CHEMOTHERAPY FOR MALIGNANT NEOPLASM (REGIME/THERAPY)
C0279023|T047||CCS_10|CHEMOSENSITIZATION/POTENTIATION
C0279023|T047||CCS_10|POTENTIATION/CHEMOSENSITIZATION
C0279023|T047||CCS_10|CHEMOSENSITIZATION
C0281488|T047||CCS_10|IN VITRO SENSITIVITY-DIRECTED CHEMOTHERAPY
C0199946|T047||CCS_10|TOPICAL CHEMOTHERAPY FOR MALIGNANT NEOPLASM 
C0199946|T047||CCS_10|TOPICAL CHEMOTHERAPY FOR MALIGNANT NEOPLASM
C0199946|T047||CCS_10|TOPICAL CHEMOTHERAPY FOR MALIGNANT NEOPLASM 
C0199946|T047||CCS_10|TOPICAL CHEMOTHERAPY FOR MALIGNANT NEOPLASM (REGIME/THERAPY)
C0189561|T047||CCS_10|PLEURODESIS WITH CANCER CHEMOTHERAPY SUBSTANCE
C0189561|T047||CCS_10|PLEURODESIS WITH CANCER CHEMOTHERAPY SUBSTANCE 
C0199942|T047||CCS_10|PERFUSION CHEMOTHERAPY FOR MALIGNANT NEOPLASM
C0199942|T047||CCS_10|PERFUSION CHEMOTHERAPY FOR MALIGNANT NEOPLASM 
C0199942|T047||CCS_10|PERFUSION CHEMOTHERAPY FOR MALIGNANT NEOPLASM 
C0199942|T047||CCS_10|PERFUSION CHEMOTHERAPY FOR MALIGNANT NEOPLASM (REGIME/THERAPY)
C0199940|T047||CCS_10|PARENTERAL CHEMOTHERAPY FOR MALIGNANT NEOPLASM
C0199940|T047||CCS_10|PARENTERAL CHEMOTHERAPY FOR MALIGNANT NEOPLASM 
C0199940|T047||CCS_10|PARENTERAL CHEMOTHERAPY FOR MALIGNANT NEOPLASM 
C0199940|T047||CCS_10|PARENTERAL CHEMOTHERAPY FOR MALIGNANT NEOPLASM (REGIME/THERAPY)
C0199943|T047||CCS_10|CHEMOTHERAPEUTICS REGIMEN INTRACAVITARY FOR MALIGNANT NEOPLASM
C0199943|T047||CCS_10|INTRACAVITARY CHEMOTHERAPEUTICS REGIMEN FOR MALIGNANT NEOPLASM 
C0199943|T047||CCS_10|INTRACAVITARY CHEMOTHERAPEUTICS REGIMEN FOR MALIGNANT NEOPLASM
C0199943|T047||CCS_10|INTRACAVITARY CHEMOTHERAPY FOR MALIGNANT NEOPLASM
C0199943|T047||CCS_10|INTRACAVITARY CHEMOTHERAPY FOR MALIGNANT NEOPLASM 
C0199943|T047||CCS_10|INTRACAVITARY CHEMOTHERAPY FOR MALIGNANT NEOPLASM (REGIME/THERAPY)
C0199941|T047||CCS_10|INTRAVENOUS CHEMOTHERAPY FOR MALIGNANT NEOPLASM 
C0199941|T047||CCS_10|INTRAVENOUS CHEMOTHERAPY FOR MALIGNANT NEOPLASM
C0199941|T047||CCS_10|CHEMOTHERAPY INTRAVENOUS FOR MALIGNANT NEOPLASM
C0199941|T047||CCS_10|INFUSION CHEMOTHERAPY FOR MALIGNANT NEOPLASM
C0199941|T047||CCS_10|INFUSION CHEMOTHERAPY FOR MALIGNANT NEOPLASM 
C0199941|T047||CCS_10|INFUSION CHEMOTHERAPY FOR MALIGNANT NEOPLASM (REGIME/THERAPY)
C0191103|T047||CCS_10|INTRAVENOUS, PUSH TECHNIQUE CHEMOTHERAPY ADMINISTRATION
C0191103|T047||CCS_10|INTRAVENOUS CHEMOTHERAPY ADMINISTRATION BY PUSH TECHNIQUE
C0191103|T047||CCS_10|INTRAVENOUS CHEMOTHERAPY ADMINISTRATION BY PUSH TECHNIQUE 
C0199945|T047||CCS_10|LOCAL CHEMOTHERAPY FOR MALIGNANT NEOPLASM 
C0199945|T047||CCS_10|LOCAL CHEMOTHERAPY FOR MALIGNANT NEOPLASM
C0199945|T047||CCS_10|LOCAL CHEMOTHERAPY FOR MALIGNANT NEOPLASM 
C0199945|T047||CCS_10|LOCAL CHEMOTHERAPY FOR MALIGNANT NEOPLASM (REGIME/THERAPY)
C0436299|T047||CCS_10|RADIOMIMETIC CHEMOTHERAPY 
C0436299|T047||CCS_10|RADIOMIMETIC CHEMOTHERAPY
C0436299|T047||CCS_10|RADIOMIMETIC CHEMOTHERAPY 
C0436299|T047||CCS_10|RADIOMIMETIC CHEMOTHERAPY (REGIME/THERAPY)
C0279512|T047||CCS_10|CYTARABINE/DAUNORUBICIN/PREDNISONE/THIOGUANINE
C0279512|T047||CCS_10|ARA-C/DNR/PRED/TG
C1521869|T047||CCS_10|CTX/IFF/VP-16
C1521869|T047||CCS_10|IFOSFAMIDE/CYCLOPHOSPHAMIDE/ETOPOSIDE
C1327770|T047||CCS_10|CCI-779/IFN-A
C1327770|T047||CCS_10|INTERFERON ALFA/TEMSIROLIMUS
C1327770|T047||CCS_10|CCI-779/INTERFERON ALFA
C1327912|T047||CCS_10|GALIXIMAB/RITUXIMAB
C1327912|T047||CCS_10|IDEC-114 MONOCLONAL ANTIBODY/RITUXIMAB
C1327912|T047||CCS_10|MOAB IDEC-114/MOAB IDEC-C2B8
C1327970|T047||CCS_10|LETROZOLE/TEMSIROLIMUS
C1327970|T047||CCS_10|CCI-779/LTZ
C1327970|T047||CCS_10|CCI-779/LETROZOLE
C1328116|T047||CCS_10|CAPTOPRIL/RECOMBINANT TISSUE PLASMINOGEN ACTIVATOR
C1328116|T047||CCS_10|CAPTOPRIL/TISSUE PLASMINOGEN ACTIVATOR
C1328116|T047||CCS_10|CPT/T-PA
C0935858|T047||CCS_10|ARA-C/ASP/DNR/MTX/PRDL/VCR
C0935858|T047||CCS_10|ASPARAGINASE/CYTARABINE/DAUNORUBICIN/METHOTREXATE/PREDNISOLONE/VINCRISTINE
C1134539|T047||CCS_10|APC8015 VACCINE/BEVACIZUMAB
C1134539|T047||CCS_10|APC8015/BEVACIZUMAB
C1134539|T047||CCS_10|APC 8015/MOAB VEGF
C1134602|T047||CCS_10|FOWLPOX VIRUS VACCINE VECTOR/GP100 ANTIGEN/INTERLEUKIN-2
C1134602|T047||CCS_10|FOWLPOX VIRUS VACCINE/GP100 ANTIGEN/INTERLEUKIN-2
C1134602|T047||CCS_10|FOWLVAC/GP100/IL-2
C0278888|T047||CCS_10|INTERLEUKIN-2/RECOMBINANT INTERFERON BETA
C0278888|T047||CCS_10|IFN-B/IL-2
C0278888|T047||CCS_10|INTERFERON BETA/INTERLEUKIN-2
C0278889|T047||CCS_10|INTERFERON GAMMA/RECOMBINANT INTERFERON BETA
C0278889|T047||CCS_10|IFN-B/IFN-G
C0278889|T047||CCS_10|INTERFERON BETA/INTERFERON GAMMA
C0279438|T047||CCS_10|FLUOROURACIL/RECOMBINANT INTERFERON BETA
C0279438|T047||CCS_10|5-FU/IFN-B
C0279438|T047||CCS_10|FLUOROURACIL/INTERFERON BETA
C0281419|T047||CCS_10|ISOTRETINOIN/RECOMBINANT INTERFERON BETA
C0281419|T047||CCS_10|13-CRA/IFN-B
C0281419|T047||CCS_10|INTERFERON BETA/ISOTRETINOIN
C0281711|T047||CCS_10|CISPLATIN/DIHYDROSPHINGOSINE
C0281711|T047||CCS_10|CDDP/SAFINGOL
C0281711|T047||CCS_10|CISPLATIN/SAFINGOL
C0393027|T047||CCS_10|ETHYNYLURACIL/FLUOROURACIL
C0393027|T047||CCS_10|ENILURACIL / 5-FU COMBINATION TABLET
C0393027|T047||CCS_10|GW776/5-FU
C0393027|T047||CCS_10|GW776/5-FLUOROURACIL
C0393027|T047||CCS_10|776C85/5-FU
C0393027|T047||CCS_10|ENILURACIL/FLUOROURACIL
C0393028|T047||CCS_10|ETHYNYLURACIL/FLUOROURACIL/LEUCOVORIN CALCIUM
C0393028|T047||CCS_10|776C85/CF/5-FU
C0393028|T047||CCS_10|ENILURACIL/FLUOROURACIL/LEUCOVORIN CALCIUM
C0796602|T047||CCS_10|FOWLPOX VIRUS VACCINE VECTOR/INTERLEUKIN-2
C0796602|T047||CCS_10|FOWLVAC/IL-2
C0796602|T047||CCS_10|FOWLPOX VIRUS VACCINE/INTERLEUKIN-2
C0796658|T047||CCS_10|FOWLPOX VIRUS VACCINE VECTOR/INTERLEUKIN-2/VACCINIA-TYROSINASE VACCINE
C0796658|T047||CCS_10|FOWLPOX VIRUS VACCINE/INTERLEUKIN-2/VACCINIA-TYROSINASE VACCINE
C0796658|T047||CCS_10|FOWLVAC/IL-2/VACTYROS
C0879332|T047||CCS_10|HER-2/NEU PEPTIDE VACCINE/MONTANIDE ISA-51
C0879332|T047||CCS_10|HER-2-NEU PEPTIDE VACCINE/MONTANIDE ISA-51
C0879332|T047||CCS_10|HER-2/ISA-51
C0879358|T047||CCS_10|HER-2/NEU PEPTIDE VACCINE/SARGRAMOSTIM
C0879358|T047||CCS_10|HER-2-NEU PEPTIDE VACCINE/SARGRAMOSTIM
C0879358|T047||CCS_10|GM-CSF/HER-2
C1831695|T047||CCS_10|CTX/DOX/MOAB VEGF/TXT
C1831695|T047||CCS_10|BEVACIZUMAB/CYCLOPHOSPHAMIDE/DOCETAXEL/DOXORUBICIN
C1831713|T047||CCS_10|CISPLATIN/DOXORUBICIN/ETOPOSIDE/IFOSFAMIDE/METHOTREXATE
C1831713|T047||CCS_10|CDDP/DOX/IFF/MTX/VP-16
C1880034|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT MALIGNANT BRAIN NEOPLASM
C1880033|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT ACUTE MYELOID LEUKEMIA
C1880060|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT PLASMA CELL MYELOMA
C1880065|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT SMALL CELL LUNG CARCINOMA
C1880051|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT MALIGNANT MESOTHELIOMA
C1880043|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT CHRONIC LYMPHOCYTIC LEUKEMIA
C1880064|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT SARCOMA
C1880052|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT MALIGNANT RENAL NEOPLASM
C1880052|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT KIDNEY CANCER
C1880055|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT NON-HODGKIN LYMPHOMA
C1880056|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT NON-SMALL CELL LUNG CARCINOMA
C1880053|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT MALIGNANT TESTICULAR NEOPLASM
C1880053|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT TESTICULAR CANCER
C1880035|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT BLADDER CARCINOMA
C1880032|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT ACUTE LYMPHOBLASTIC LEUKEMIA
C1880036|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT BREAST CARCINOMA
C1880054|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT MELANOMA
C1880044|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT COLORECTAL CARCINOMA
C1880037|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT CERVICAL CARCINOMA
C1880048|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT GASTRIC CARCINOMA
C1880058|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT MALIGNANT OVARIAN NEOPLASM
C1880050|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT MALIGNANT HEAD AND NECK NEOPLASM
C1880049|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT HODGKINS LYMPHOMA
C1880045|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT ENDOMETRIAL CARCINOMA
C1880061|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT LIVER CANCER
C1880061|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT PRIMARY MALIGNANT NEOPLASM OF LIVER
C1880046|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT ESOPHAGEAL CARCINOMA
C1880059|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT PANCREATIC CARCINOMA
C1880059|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT PANCREATIC CANCER
C1880062|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT PROSTATE CARCINOMA
C2347611|T047||CCS_10|CHEMOTHERAPY REGIMEN USED TO TREAT GESTATIONAL TROPHOBLASTIC TUMOR
C0152018|T047||CCS_10|CARCINOMA OF ESOPHAGUS
C0152018|T047||CCS_10|ESOPHAGEAL CARCINOMA
C0152018|T047||CCS_10|ESOPHAGEAL CANCER
C0152018|T047||CCS_10|CARCINOMA OF ESOPHAGUS 
C0152018|T047||CCS_10|CARCINOMA;OESOPHAGUS
C0152018|T047||CCS_10|CARCINOMA OF OESOPHAGUS
C0152018|T047||CCS_10|CARCINOMA OF OESOPHAGUS 
C0152018|T047||CCS_10|CANCER OF OESOPHAGUS
C0152018|T047||CCS_10|CARCINOMA OF ESOPHAGUS 
C0152018|T047||CCS_10|ESOPHAGEAL CANCER, NOS
C0152018|T047||CCS_10|ESOPHAGEAL CARCINOMA NOS
C0152018|T047||CCS_10|CARCINOMA OF OESOPHAGUS NOS
C0152018|T047||CCS_10|CARCINOMA OF ESOPHAGUS NOS
C0152018|T047||CCS_10|OESOPHAGEAL CARCINOMA
C0152018|T047||CCS_10|OESOPHAGEAL CARCINOMA NOS
C0152018|T047||CCS_10|CANCER OF ESOPHAGUS
C0152018|T047||CCS_10|CANCER OF THE ESOPHAGUS
C0152018|T047||CCS_10|ESOPHAGUS CARCINOMA
C0152018|T047||CCS_10|CARCINOMA OF THE ESOPHAGUS
C0152018|T047||CCS_10|CARCINOMA;ESOPHAGUS
C0152018|T047||CCS_10|CARCINOMA OF THE OESOPHAGUS
C0496775|T047||CCS_10|MALIGNANT NEOPLASM OF ABDOMINAL PART OF ESOPHAGUS
C0496775|T047||CCS_10|MALIGNANT NEOPLASM OF ABDOMINAL PART OF OESOPHAGUS
C0496775|T047||CCS_10|MALIGNANT NEOPLASM OF ABDOMINAL ESOPHAGUS
C0496775|T047||CCS_10|MALIGNANT NEOPLASM OF ABDOMINAL ESOPHAGUS 
C0496775|T047||CCS_10|MALIGNANT TUMOR OF ABDOMINAL ESOPHAGUS
C0496775|T047||CCS_10|MAL NEO ABDOMIN ESOPHAG
C0496775|T047||CCS_10|MALIGNANT NEOPLASM OF ABDOMINAL OESOPHAGUS
C0496775|T047||CCS_10|MALIGNANT TUMOR OF ABDOMINAL PART OF ESOPHAGUS
C0496775|T047||CCS_10|MALIGNANT TUMOUR OF ABDOMINAL PART OF OESOPHAGUS
C0496775|T047||CCS_10|MALIGNANT TUMOR OF ABDOMINAL PART OF ESOPHAGUS 
C0496775|T047||CCS_10|MALIGNANT NEOPLASM OF THE ABDOMINAL ESOPHAGUS
C0496775|T047||CCS_10|MALIGNANT TUMOR OF THE ABDOMINAL ESOPHAGUS
C0496773|T047||CCS_10|MALIGNANT NEOPLASM OF CERVICAL PART OF ESOPHAGUS
C0496773|T047||CCS_10|MALIGNANT NEOPLASM OF CERVICAL PART OF OESOPHAGUS
C0496773|T047||CCS_10|MALIGNANT NEOPLASM OF CERVICAL ESOPHAGUS 
C0496773|T047||CCS_10|MALIGNANT NEOPLASM OF CERVICAL ESOPHAGUS
C0496773|T047||CCS_10|MALIGNANT TUMOR OF CERVICAL ESOPHAGUS
C0496773|T047||CCS_10|MAL NEO CERVICAL ESOPHAG
C0496773|T047||CCS_10|MALIGNANT NEOPLASM OF CERVICAL OESOPHAGUS
C0496773|T047||CCS_10|MALIGNANT TUMOR OF CERVICAL PART OF ESOPHAGUS
C0496773|T047||CCS_10|MALIGNANT TUMOUR OF CERVICAL PART OF OESOPHAGUS
C0496773|T047||CCS_10|MALIGNANT TUMOR OF CERVICAL PART OF ESOPHAGUS 
C0496773|T047||CCS_10|MALIGNANT NEOPLASM OF THE CERVICAL ESOPHAGUS
C0153411|T047||CCS_10|MALIGNANT NEOPLASM OF THORACIC ESOPHAGUS
C0153411|T047||CCS_10|MALIGNANT NEOPLASM OF THORACIC PART OF ESOPHAGUS
C0153411|T047||CCS_10|MALIGNANT NEOPLASM OF THORACIC PART OF OESOPHAGUS
C0153411|T047||CCS_10|MALIGNANT NEOPLASM OF THORACIC ESOPHAGUS 
C0153411|T047||CCS_10|MALIGNANT TUMOR OF THORACIC ESOPHAGUS
C0153411|T047||CCS_10|MAL NEO THORACIC ESOPHAG
C0153411|T047||CCS_10|MALIGNANT NEOPLASM OF THORACIC OESOPHAGUS
C0153411|T047||CCS_10|MALIGNANT TUMOR OF THORACIC PART OF ESOPHAGUS
C0153411|T047||CCS_10|MALIGNANT TUMOUR OF THORACIC PART OF OESOPHAGUS
C0153411|T047||CCS_10|MALIGNANT TUMOR OF THORACIC PART OF ESOPHAGUS 
C0153411|T047||CCS_10|MALIGNANT NEOPLASM OF THE THORACIC ESOPHAGUS
C0153416|T047||CCS_10|MALIGNANT NEOPLASM OF OTHER SPECIFIED PART OF ESOPHAGUS
C0153416|T047||CCS_10|MALIGNANT NEOPLASM OF OTHER SPECIFIED PART OF OESOPHAGUS
C0153416|T047||CCS_10|MAL NEO ESOPHAGUS NEC
C0153416|T047||CCS_10|MALIGNANT NEOPLASM OF OTHER SPECIFIED PART OF ESOPHAGUS 
C0153413|T047||CCS_10|MALIGNANT NEOPLASM OF UPPER THIRD OF ESOPHAGUS
C0153413|T047||CCS_10|MALIGNANT NEOPLASM OF UPPER THIRD OF OESOPHAGUS
C0153413|T047||CCS_10|MALIGNANT NEOPLASM OF UPPER THIRD ESOPHAGUS
C0153413|T047||CCS_10|MALIGNANT NEOPLASM OF UPPER THIRD OF ESOPHAGUS 
C0153413|T047||CCS_10|MALIGNANT TUMOR OF UPPER THIRD OF ESOPHAGUS
C0153413|T047||CCS_10|MAL NEO UPPER 3RD ESOPH
C0153413|T047||CCS_10|MALIGNANT TUMOUR OF UPPER THIRD OF OESOPHAGUS
C0153413|T047||CCS_10|MALIGNANT TUMOR OF UPPER THIRD OF ESOPHAGUS 
C0153413|T047||CCS_10|MALIGNANT NEOPLASM OF PROXIMAL THIRD OF ESOPHAGUS
C0153413|T047||CCS_10|MALIGNANT NEOPLASM OF THE PROXIMAL THIRD OF THE ESOPHAGUS
C0153413|T047||CCS_10|MALIGNANT NEOPLASM OF THE UPPER THIRD OF THE ESOPHAGUS
C0153413|T047||CCS_10|MALIGNANT TUMOR OF PROXIMAL THIRD OF ESOPHAGUS
C0153413|T047||CCS_10|MALIGNANT TUMOR OF THE PROXIMAL THIRD OF THE ESOPHAGUS
C0153413|T047||CCS_10|MALIGNANT TUMOR OF THE UPPER THIRD OF THE ESOPHAGUS
C0153415|T047||CCS_10|MALIGNANT NEOPLASM OF LOWER THIRD OF ESOPHAGUS
C0153415|T047||CCS_10|MALIGNANT NEOPLASM OF LOWER THIRD OF OESOPHAGUS
C0153415|T047||CCS_10|MALIGNANT NEOPLASM OF LOWER THIRD OF ESOPHAGUS 
C0153415|T047||CCS_10|MALIGNANT TUMOR OF LOWER THIRD OF ESOPHAGUS
C0153415|T047||CCS_10|MAL NEO LOWER 3RD ESOPH
C0153415|T047||CCS_10|CA LOWER THIRD ESOPHAGUS 
C0153415|T047||CCS_10|CA LOWER THIRD ESOPHAGUS
C0153415|T047||CCS_10|CA LOWER THIRD OESOPHAGUS
C0153415|T047||CCS_10|CA LOWER THIRD OESOPHAGUS 
C0153415|T047||CCS_10|MALIGNANT TUMOUR OF LOWER THIRD OF OESOPHAGUS
C0153415|T047||CCS_10|MALIGNANT TUMOR OF LOWER THIRD OF ESOPHAGUS 
C0153415|T047||CCS_10|MALIGNANT LOWER THIRD OF ESOPHAGUS NEOPLASM
C0153415|T047||CCS_10|MALIGNANT LOWER THIRD OF ESOPHAGUS TUMOR
C0153415|T047||CCS_10|MALIGNANT LOWER THIRD OF THE ESOPHAGUS NEOPLASM
C0153415|T047||CCS_10|MALIGNANT LOWER THIRD OF THE ESOPHAGUS TUMOR
C0153415|T047||CCS_10|MALIGNANT NEOPLASM OF DISTAL THIRD OF ESOPHAGUS
C0153415|T047||CCS_10|MALIGNANT NEOPLASM OF THE DISTAL THIRD OF THE ESOPHAGUS
C0153415|T047||CCS_10|MALIGNANT NEOPLASM OF THE LOWER THIRD OF THE ESOPHAGUS
C0153415|T047||CCS_10|MALIGNANT TUMOR OF DISTAL THIRD OF ESOPHAGUS
C0153415|T047||CCS_10|MALIGNANT TUMOR OF THE DISTAL THIRD OF THE ESOPHAGUS
C0153415|T047||CCS_10|MALIGNANT TUMOR OF THE LOWER THIRD OF THE ESOPHAGUS
C0153414|T047||CCS_10|MALIGNANT NEOPLASM OF MIDDLE THIRD OF ESOPHAGUS
C0153414|T047||CCS_10|MALIGNANT NEOPLASM OF MIDDLE THIRD OF OESOPHAGUS
C0153414|T047||CCS_10|MALIGNANT NEOPLASM OF MIDDLE THIRD OF ESOPHAGUS 
C0153414|T047||CCS_10|MALIGNANT TUMOR OF MIDDLE THIRD OF ESOPHAGUS
C0153414|T047||CCS_10|MAL NEO MIDDLE 3RD ESOPH
C0153414|T047||CCS_10|CA MIDDLE THIRD ESOPHAGUS 
C0153414|T047||CCS_10|CA MIDDLE THIRD OESOPHAGUS
C0153414|T047||CCS_10|CA MIDDLE THIRD OESOPHAGUS 
C0153414|T047||CCS_10|CA MIDDLE THIRD ESOPHAGUS
C0153414|T047||CCS_10|MALIGNANT TUMOUR OF MIDDLE THIRD OF OESOPHAGUS
C0153414|T047||CCS_10|MALIGNANT TUMOR OF MIDDLE THIRD OF ESOPHAGUS 
C0153414|T047||CCS_10|MALIGNANT MIDDLE THIRD OF ESOPHAGUS NEOPLASM
C0153414|T047||CCS_10|MALIGNANT MIDDLE THIRD OF ESOPHAGUS TUMOR
C0153414|T047||CCS_10|MALIGNANT MIDDLE THIRD OF THE ESOPHAGUS NEOPLASM
C0153414|T047||CCS_10|MALIGNANT MIDDLE THIRD OF THE ESOPHAGUS TUMOR
C0153414|T047||CCS_10|MALIGNANT NEOPLASM OF THE MIDDLE THIRD OF THE ESOPHAGUS
C0153414|T047||CCS_10|MALIGNANT TUMOR OF THE MIDDLE THIRD OF THE ESOPHAGUS
C0546837|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS
C0546837|T047||CCS_10|CANCER OF ESOPHAGUS
C0546837|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS, UNSPECIFIED
C0546837|T047||CCS_10|ESOPHAGUS, UNSPECIFIED
C0546837|T047||CCS_10|MALIGNANT NEOPLASM OF OESOPHAGUS
C0546837|T047||CCS_10|MALIGNANT NEOPLASM OF OESOPHAGUS, UNSPECIFIED
C0546837|T047||CCS_10|OESOPHAGUS, UNSPECIFIED
C0546837|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS 
C0546837|T047||CCS_10|ESOPHAGEAL CANCER
C0546837|T047||CCS_10|ESOPHAGEAL CANCER 
C0546837|T047||CCS_10|MALIGNANT ESOPHAGEAL NEOPLASM
C0546837|T047||CCS_10|CA ESOPHAGUS
C0546837|T047||CCS_10|OESOPHAGEAL NEOPLASMS MALIGNANT
C0546837|T047||CCS_10|CANCER, ESOPHAGEAL
C0546837|T047||CCS_10|CANCERS, ESOPHAGEAL
C0546837|T047||CCS_10|ESOPHAGEAL CANCERS
C0546837|T047||CCS_10|CANCERS, ESOPHAGUS
C0546837|T047||CCS_10|ESOPHAGUS CANCERS
C0546837|T047||CCS_10|MALIGNANT TUMOR OF ESOPHAGUS
C0546837|T047||CCS_10|MAL NEO ESOPHAGUS NOS
C0546837|T047||CCS_10|CANCER, ESOPHAGUS
C0546837|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS, UNSPECIFIED SITE
C0546837|T047||CCS_10|OESOPHAGEAL CANCER
C0546837|T047||CCS_10|MALIGNANT NEOPLASM OF OESOPHAGUS NOS
C0546837|T047||CCS_10|CA ESOPHAGUS NOS 
C0546837|T047||CCS_10|CA ESOPHAGUS NOS
C0546837|T047||CCS_10|(MALIGNANT NEOPLASM OF OESOPHAGUS NOS OR OESOPHAGEAL CANCER
C0546837|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS NOS
C0546837|T047||CCS_10|CA OESOPHAGUS NOS
C0546837|T047||CCS_10|CA OESOPHAGUS NOS 
C0546837|T047||CCS_10|CA - CANCER OF ESOPHAGUS
C0546837|T047||CCS_10|CA - CANCER OF OESOPHAGUS
C0546837|T047||CCS_10|CANCER OF OESOPHAGUS
C0546837|T047||CCS_10|MALIGNANT TUMOUR OF OESOPHAGUS
C0546837|T047||CCS_10|MALIGNANT TUMOUR OF OESOPHAGUS 
C0546837|T047||CCS_10|(MALIGNANT NEOPLASM OF ESOPHAGUS NOS OR ESOPHAGEAL CANCER
C0546837|T047||CCS_10|(MALIGNANT NEOPLASM OF OESOPHAGUS NOS OR OESOPHAGEAL CANCER 
C0546837|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS NOS 
C0546837|T047||CCS_10|ESOPHAGUS--CANCER
C0546837|T047||CCS_10|-- ESOPHAGEAL CANCER
C0546837|T047||CCS_10|OESOPHAGEAL CANCER NOS
C0546837|T047||CCS_10|ESOPHAGEAL CANCER NOS
C0546837|T047||CCS_10|ESOPHAGUS CANCER
C0546837|T047||CCS_10|CANCER OF THE ESOPHAGUS
C0546837|T047||CCS_10|CA OESOPHAGUS
C0546837|T047||CCS_10|MALIGNANT TUMOR OF ESOPHAGUS 
C0546837|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS, NOS
C0546837|T047||CCS_10|MALIGNANT ESOPHAGEAL TUMOR
C0546837|T047||CCS_10|MALIGNANT ESOPHAGUS TUMOR
C0546837|T047||CCS_10|MALIGNANT NEOPLASM OF THE ESOPHAGUS
C0546837|T047||CCS_10|MALIGNANT TUMOR OF THE ESOPHAGUS
C0546837|T047||CCS_10|ESOPHAGEAL NEOPLASMS MALIGNANT
C0546837|T047||CCS_10|NEOPLASM MALIG;ESOPHAGUS
C0546837|T047||CCS_10|NEOPLASM MALIG;OESOPHAGUS
C0546837|T047||CCS_10|MALIGNANT NEOSPLASM OF THE ESOPHAGUS
C0546837|T047||CCS_10|MALIGNANT NEOSPLASM OF THE OESOPHAGUS
C0496776|T047||CCS_10|MALIGNANT NEOPLASM OVERLAPPING ESOPHAGUS SITE
C0496776|T047||CCS_10|MALIGNANT NEOPLASM OVERLAPPING OESOPHAGUS SITE
C0496776|T047||CCS_10|OVERLAPPING LESION OF ESOPHAGUS
C0496776|T047||CCS_10|OVERLAPPING LESION OF OESOPHAGUS
C0496776|T047||CCS_10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF ESOPHAGUS
C0496776|T047||CCS_10|ESOPHAGEAL NEOPLASM MALIGNANT OVERLAPPING SITES OF ESOPHAGUS
C0496776|T047||CCS_10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF ESOPHAGUS 
C0279628|T047||CCS_10|ADENOCARCINOMA OF ESOPHAGUS 
C0279628|T047||CCS_10|ADENOCARCINOMA OF ESOPHAGUS
C0279628|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA
C0279628|T047||CCS_10|ADENOCARCINOMA - ESOPHAGUS
C0279628|T047||CCS_10|ADENOCARCINOMA OF THE ESOPHAGUS
C0279628|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA NOS
C0279628|T047||CCS_10|OESOPHAGEAL ADENOCARCINOMA
C0279628|T047||CCS_10|OESOPHAGEAL ADENOCARCINOMA NOS
C0279628|T047||CCS_10|ADENOCARCINOMA OF OESOPHAGUS
C0279628|T047||CCS_10|ADENOCARCINOMA OF ESOPHAGUS 
C0279628|T047||CCS_10|ESOPHAGEAL CANCER, ADENOCARCINOMA
C0279628|T047||CCS_10|ESOPHAGUS CANCER, ADENOCARCINOMA
C0279628|T047||CCS_10|ESOPHAGUS ADENOCARCINOMA
C0854762|T047||CCS_10|OESOPHAGEAL ADENOCARCINOMA RECURRENT
C0854762|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA RECURRENT
C0854762|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA, RECURRENT
C0854762|T047||CCS_10|RECURRENT ADENOCARCINOMA OF ESOPHAGUS
C0854762|T047||CCS_10|RECURRENT ADENOCARCINOMA OF THE ESOPHAGUS
C0854762|T047||CCS_10|RECURRENT ESOPHAGEAL ADENOCARCINOMA
C0854762|T047||CCS_10|RECURRENT ESOPHAGUS ADENOCARCINOMA
C0854762|T047||CCS_10|RELAPSED ADENOCARCINOMA OF ESOPHAGUS
C0854762|T047||CCS_10|RELAPSED ADENOCARCINOMA OF THE ESOPHAGUS
C0854762|T047||CCS_10|RELAPSED ESOPHAGEAL ADENOCARCINOMA
C0854762|T047||CCS_10|RELAPSED ESOPHAGUS ADENOCARCINOMA
C0854764|T047||CCS_10|ADENOCARCINOMA IN SITU OF ESOPHAGUS 
C0854764|T047||CCS_10|ADENOCARCINOMA IN SITU OF ESOPHAGUS
C0854764|T047||CCS_10|OESOPHAGEAL ADENOCARCINOMA STAGE 0
C0854764|T047||CCS_10|STAGE 0 ESOPHAGEAL ADENOCARCINOMA AJCC V7
C0854764|T047||CCS_10|STAGE 0 ESOPHAGEAL ADENOCARCINOMA
C0854764|T047||CCS_10|OESOPHAGEAL ADENOCARCINOMA SITE UNSPECIFIED STAGE 0
C0854764|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA IN SITU
C0854764|T047||CCS_10|OESOPHAGEAL ADENOCARCINOMA SITE UNSPECIFIED IN SITU
C0854764|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA SITE UNSPECIFIED STAGE 0
C0854764|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA STAGE 0
C0854764|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA SITE UNSPECIFIED IN SITU
C0854764|T047||CCS_10|OESOPHAGEAL ADENOCARCINOMA IN SITU
C0854764|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA, STAGE 0
C0854764|T047||CCS_10|ADENOCARCINOMA IN SITU OF THE ESOPHAGUS
C0854764|T047||CCS_10|ESOPHAGUS ADENOCARCINOMA IN SITU
C0854764|T047||CCS_10|STAGE 0 ADENOCARCINOMA OF ESOPHAGUS
C0854764|T047||CCS_10|STAGE 0 ADENOCARCINOMA OF THE ESOPHAGUS
C0854764|T047||CCS_10|STAGE 0 ESOPHAGUS ADENOCARCINOMA
C0854765|T047||CCS_10|OESOPHAGEAL ADENOCARCINOMA STAGE I
C0854765|T047||CCS_10|STAGE I ESOPHAGEAL ADENOCARCINOMA AJCC V7
C0854765|T047||CCS_10|STAGE I ESOPHAGEAL ADENOCARCINOMA
C0854765|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA SITE UNSPECIFIED STAGE I
C0854765|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA STAGE I
C0854765|T047||CCS_10|OESOPHAGEAL ADENOCARCINOMA SITE UNSPECIFIED STAGE I
C0854765|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA, STAGE I
C0854765|T047||CCS_10|STAGE I ADENOCARCINOMA OF ESOPHAGUS
C0854765|T047||CCS_10|STAGE I ADENOCARCINOMA OF THE ESOPHAGUS
C0854765|T047||CCS_10|STAGE I ESOPHAGUS ADENOCARCINOMA
C0854763|T047||CCS_10|OESOPHAGEAL ADENOCARCINOMA STAGE II
C0854763|T047||CCS_10|STAGE II ESOPHAGEAL ADENOCARCINOMA AJCC V7
C0854763|T047||CCS_10|STAGE II ESOPHAGEAL ADENOCARCINOMA
C0854763|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA SITE UNSPECIFIED STAGE II
C0854763|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA STAGE II
C0854763|T047||CCS_10|OESOPHAGEAL ADENOCARCINOMA SITE UNSPECIFIED STAGE II
C0854763|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA, STAGE II
C0854763|T047||CCS_10|STAGE II ADENOCARCINOMA OF ESOPHAGUS
C0854763|T047||CCS_10|STAGE II ADENOCARCINOMA OF THE ESOPHAGUS
C0854763|T047||CCS_10|STAGE II ESOPHAGUS ADENOCARCINOMA
C0854766|T047||CCS_10|OESOPHAGEAL ADENOCARCINOMA STAGE III
C0854766|T047||CCS_10|STAGE III ESOPHAGEAL ADENOCARCINOMA AJCC V7
C0854766|T047||CCS_10|STAGE III ESOPHAGEAL ADENOCARCINOMA
C0854766|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA STAGE III
C0854766|T047||CCS_10|OESOPHAGEAL ADENOCARCINOMA SITE UNSPECIFIED STAGE III
C0854766|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA SITE UNSPECIFIED STAGE III
C0854766|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA, STAGE III
C0854766|T047||CCS_10|STAGE III ADENOCARCINOMA OF ESOPHAGUS
C0854766|T047||CCS_10|STAGE III ADENOCARCINOMA OF THE ESOPHAGUS
C0854766|T047||CCS_10|STAGE III ESOPHAGUS ADENOCARCINOMA
C1142347|T047||CCS_10|OESOPHAGEAL ADENOCARCINOMA STAGE IV
C1142347|T047||CCS_10|STAGE IV ESOPHAGEAL ADENOCARCINOMA AJCC V7
C1142347|T047||CCS_10|STAGE IV ESOPHAGEAL ADENOCARCINOMA
C1142347|T047||CCS_10|OESOPHAGEAL ADENOCARCINOMA METASTATIC
C1142347|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA METASTATIC
C1142347|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA SITE UNSPECIFIED STAGE IV
C1142347|T047||CCS_10|OESOPHAGEAL ADENOCARCINOMA SITE UNSPECIFIED STAGE IV
C1142347|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA STAGE IV
C1142347|T047||CCS_10|ESOPHAGEAL ADENOCARCINOMA, STAGE IV
C1142347|T047||CCS_10|METASTATIC ADENOCARCINOMA OF ESOPHAGUS
C1142347|T047||CCS_10|METASTATIC ADENOCARCINOMA OF THE ESOPHAGUS
C1142347|T047||CCS_10|METASTATIC ESOPHAGEAL ADENOCARCINOMA
C1142347|T047||CCS_10|METASTATIC ESOPHAGUS ADENOCARCINOMA
C1142347|T047||CCS_10|STAGE IV ADENOCARCINOMA OF ESOPHAGUS
C1142347|T047||CCS_10|STAGE IV ADENOCARCINOMA OF THE ESOPHAGUS
C1142347|T047||CCS_10|STAGE IV ESOPHAGUS ADENOCARCINOMA
C0854761|T047||CCS_10|OESOPHAGEAL CARCINOMA RECURRENT
C0854761|T047||CCS_10|RECURRENT ESOPHAGEAL CANCER
C0854761|T047||CCS_10|RECURRENT ESOPHAGEAL CARCINOMA
C0854761|T047||CCS_10|OESOPHAGEAL CARCINOMA SITE UNSPECIFIED RECURRENT
C0854761|T047||CCS_10|ESOPHAGEAL CARCINOMA RECURRENT
C0854761|T047||CCS_10|ESOPHAGEAL CARCINOMA SITE UNSPECIFIED RECURRENT
C0854761|T047||CCS_10|ESOPHAGEAL CANCER, RECURRENT
C0854761|T047||CCS_10|ESOPHAGUS CANCER, RECURRENT
C0854761|T047||CCS_10|ESOPHAGEAL CARCINOMA, RECURRENT
C0854761|T047||CCS_10|RECURRENT CANCER OF ESOPHAGUS
C0854761|T047||CCS_10|RECURRENT CANCER OF THE ESOPHAGUS
C0854761|T047||CCS_10|RECURRENT CARCINOMA OF ESOPHAGUS
C0854761|T047||CCS_10|RECURRENT CARCINOMA OF THE ESOPHAGUS
C0854761|T047||CCS_10|RECURRENT ESOPHAGUS CANCER
C0854761|T047||CCS_10|RELAPSED CANCER OF ESOPHAGUS
C0854761|T047||CCS_10|RELAPSED CANCER OF THE ESOPHAGUS
C0854761|T047||CCS_10|RELAPSED CARCINOMA OF ESOPHAGUS
C0854761|T047||CCS_10|RELAPSED CARCINOMA OF THE ESOPHAGUS
C0854761|T047||CCS_10|RELAPSED ESOPHAGEAL CANCER
C0854761|T047||CCS_10|RELAPSED ESOPHAGUS CARCINOMA
C0154059|T047||CCS_10|ESOPHAGUS
C0154059|T047||CCS_10|CARCINOMA IN SITU OF ESOPHAGUS
C0154059|T047||CCS_10|CARCINOMA IN SITU OF OESOPHAGUS
C0154059|T047||CCS_10|OESOPHAGUS
C0154059|T047||CCS_10|CARCINOMA IN SITU OF ESOPHAGUS 
C0154059|T047||CCS_10|CA IN SITU ESOPHAGUS
C0154059|T047||CCS_10|ESOPHAGEAL CARCINOMA IN SITU AJCC V7
C0154059|T047||CCS_10|SEVERE ESOPHAGEAL DYSPLASIA AJCC V7
C0154059|T047||CCS_10|SEVERE ESOPHAGEAL DYSPLASIA
C0154059|T047||CCS_10|STAGE 0 ESOPHAGEAL CANCER AJCC V7
C0154059|T047||CCS_10|ESOPHAGEAL CARCINOMA IN SITU
C0154059|T047||CCS_10|STAGE 0 ESOPHAGEAL CANCER
C0154059|T047||CCS_10|CARCINOMA IN SITU OF ESOPHAGUS NOS
C0154059|T047||CCS_10|CARCINOMA IN SITU OF OESOPHAGUS NOS
C0154059|T047||CCS_10|CARCINOMA IN SITU OF ESOPHAGUS NOS 
C0154059|T047||CCS_10|STAGE 0 ESOPHAGEAL CARCINOMA IN SITU
C0154059|T047||CCS_10|CANCER IN SITU OF ESOPHAGUS
C0154059|T047||CCS_10|CANCER IN SITU OF OESOPHAGUS
C0154059|T047||CCS_10|OESOPHAGEAL CARCINOMA NOS STAGE 0
C0154059|T047||CCS_10|ESOPHAGEAL CARCINOMA STAGE 0
C0154059|T047||CCS_10|ESOPHAGEAL CARCINOMA SITE UNSPECIFIED STAGE 0
C0154059|T047||CCS_10|OESOPHAGEAL CARCINOMA SITE UNSPECIFIED STAGE 0
C0154059|T047||CCS_10|OESOPHAGEAL CARCINOMA IN SITU
C0154059|T047||CCS_10|OESOPHAGEAL CARCINOMA STAGE 0
C0154059|T047||CCS_10|ESOPHAGEAL CARCINOMA NOS STAGE 0
C0154059|T047||CCS_10|SEVERE OESOPHAGEAL DYSPLASIA
C0154059|T047||CCS_10|CARCINOMA IN SITU OF ESOPHAGUS 
C0154059|T047||CCS_10|SEVERE ESOPHAGEAL DYSPLASIA 
C0154059|T047||CCS_10|ESOPHAGEAL CANCER, STAGE 0
C0154059|T047||CCS_10|ESOPHAGUS CANCER, STAGE 0
C0154059|T047||CCS_10|CARCINOMA IN SITU OF ESOPHAGUS, NOS
C0854769|T047||CCS_10|OESOPHAGEAL SQUAMOUS CELL CARCINOMA RECURRENT
C0854769|T047||CCS_10|ESOPHAGEAL SQUAMOUS CELL CARCINOMA SITE UNSPECIFIED RECURRENT
C0854769|T047||CCS_10|ESOPHAGEAL SQUAMOUS CELL CARCINOMA RECURRENT
C0854769|T047||CCS_10|OESOPHAGEAL SQUAMOUS CELL CARCINOMA SITE UNSPECIFIED RECURRENT
C0854769|T047||CCS_10|RECURRENT ESOPHAGEAL SQUAMOUS CELL CARCINOMA
C0854769|T047||CCS_10|RECURRENT SQUAMOUS CELL CARCINOMA OF ESOPHAGUS
C0854769|T047||CCS_10|RECURRENT SQUAMOUS CELL CARCINOMA OF THE ESOPHAGUS
C0854770|T047||CCS_10|SQUAMOUS CELL CARCINOMA IN SITU OF ESOPHAGUS 
C0854770|T047||CCS_10|SQUAMOUS CELL CARCINOMA IN SITU OF ESOPHAGUS
C0854770|T047||CCS_10|OESOPHAGEAL SQUAMOUS CELL CARCINOMA STAGE 0
C0854770|T047||CCS_10|STAGE 0 ESOPHAGEAL SQUAMOUS CELL CARCINOMA AJCC V7
C0854770|T047||CCS_10|STAGE 0 ESOPHAGEAL SQUAMOUS CELL CARCINOMA
C0854770|T047||CCS_10|OESOPHAGEAL SQUAMOUS CELL CARCINOMA IN SITU
C0854770|T047||CCS_10|ESOPHAGEAL SQUAMOUS CELL CARCINOMA IN SITU
C0854770|T047||CCS_10|ESOPHAGEAL SQUAMOUS CELL CARCINOMA STAGE 0
C0854770|T047||CCS_10|ESOPHAGUS SQUAMOUS CELL CARCINOMA IN SITU
C0854770|T047||CCS_10|SQUAMOUS CELL CARCINOMA IN SITU OF THE ESOPHAGUS
C0854770|T047||CCS_10|STAGE 0 ESOPHAGUS SQUAMOUS CELL CARCINOMA
C0854770|T047||CCS_10|STAGE 0 SQUAMOUS CELL CARCINOMA OF ESOPHAGUS
C0854770|T047||CCS_10|STAGE 0 SQUAMOUS CELL CARCINOMA OF THE ESOPHAGUS
C0854771|T047||CCS_10|OESOPHAGEAL SQUAMOUS CELL CARCINOMA STAGE I
C0854771|T047||CCS_10|STAGE I ESOPHAGEAL SQUAMOUS CELL CARCINOMA AJCC V7
C0854771|T047||CCS_10|STAGE I ESOPHAGEAL SQUAMOUS CELL CARCINOMA
C0854771|T047||CCS_10|ESOPHAGEAL SQUAMOUS CELL CARCINOMA SITE UNSPECIFIED STAGE I
C0854771|T047||CCS_10|ESOPHAGEAL SQUAMOUS CELL CARCINOMA STAGE I
C0854771|T047||CCS_10|OESOPHAGEAL SQUAMOUS CELL CARCINOMA SITE UNSPECIFIED STAGE I
C0854771|T047||CCS_10|STAGE I ESOPHAGUS SQUAMOUS CELL CARCINOMA
C0854771|T047||CCS_10|STAGE I SQUAMOUS CELL CARCINOMA OF ESOPHAGUS
C0854771|T047||CCS_10|STAGE I SQUAMOUS CELL CARCINOMA OF THE ESOPHAGUS
C0854772|T047||CCS_10|OESOPHAGEAL SQUAMOUS CELL CARCINOMA STAGE II
C0854772|T047||CCS_10|STAGE II ESOPHAGEAL SQUAMOUS CELL CARCINOMA AJCC V7
C0854772|T047||CCS_10|STAGE II ESOPHAGEAL SQUAMOUS CELL CARCINOMA
C0854772|T047||CCS_10|ESOPHAGEAL SQUAMOUS CELL CARCINOMA SITE UNSPECIFIED STAGE II
C0854772|T047||CCS_10|OESOPHAGEAL SQUAMOUS CELL CARCINOMA SITE UNSPECIFIED STAGE II
C0854772|T047||CCS_10|ESOPHAGEAL SQUAMOUS CELL CARCINOMA STAGE II
C0854772|T047||CCS_10|STAGE II ESOPHAGUS SQUAMOUS CELL CARCINOMA
C0854772|T047||CCS_10|STAGE II SQUAMOUS CELL CARCINOMA OF ESOPHAGUS
C0854772|T047||CCS_10|STAGE II SQUAMOUS CELL CARCINOMA OF THE ESOPHAGUS
C0854773|T047||CCS_10|OESOPHAGEAL SQUAMOUS CELL CARCINOMA STAGE III
C0854773|T047||CCS_10|STAGE III ESOPHAGEAL SQUAMOUS CELL CARCINOMA AJCC V7
C0854773|T047||CCS_10|STAGE III ESOPHAGEAL SQUAMOUS CELL CARCINOMA
C0854773|T047||CCS_10|ESOPHAGEAL SQUAMOUS CELL CARCINOMA STAGE III
C0854773|T047||CCS_10|STAGE III ESOPHAGUS SQUAMOUS CELL CARCINOMA
C0854773|T047||CCS_10|STAGE III SQUAMOUS CELL CARCINOMA OF ESOPHAGUS
C0854773|T047||CCS_10|STAGE III SQUAMOUS CELL CARCINOMA OF THE ESOPHAGUS
C1142025|T047||CCS_10|OESOPHAGEAL SQUAMOUS CELL CARCINOMA STAGE IV
C1142025|T047||CCS_10|STAGE IV ESOPHAGEAL SQUAMOUS CELL CARCINOMA AJCC V7
C1142025|T047||CCS_10|STAGE IV ESOPHAGEAL SQUAMOUS CELL CARCINOMA
C1142025|T047||CCS_10|OESOPHAGEAL SQUAMOUS CELL CARCINOMA METASTATIC
C1142025|T047||CCS_10|OESOPHAGEAL SQUAMOUS CELL CARCINOMA SITE UNSPECIFIED STAGE IV
C1142025|T047||CCS_10|ESOPHAGEAL SQUAMOUS CELL CARCINOMA METASTATIC
C1142025|T047||CCS_10|ESOPHAGEAL SQUAMOUS CELL CARCINOMA SITE UNSPECIFIED STAGE IV
C1142025|T047||CCS_10|ESOPHAGEAL SQUAMOUS CELL CARCINOMA STAGE IV
C1142025|T047||CCS_10|METASTATIC ESOPHAGEAL SQUAMOUS CELL CARCINOMA
C1142025|T047||CCS_10|METASTATIC ESOPHAGUS SQUAMOUS CELL CARCINOMA
C1142025|T047||CCS_10|METASTATIC SQUAMOUS CELL CARCINOMA OF ESOPHAGUS
C1142025|T047||CCS_10|METASTATIC SQUAMOUS CELL CARCINOMA OF THE ESOPHAGUS
C1142025|T047||CCS_10|STAGE IV ESOPHAGUS SQUAMOUS CELL CARCINOMA
C1142025|T047||CCS_10|STAGE IV SQUAMOUS CELL CARCINOMA OF ESOPHAGUS
C1142025|T047||CCS_10|STAGE IV SQUAMOUS CELL CARCINOMA OF THE ESOPHAGUS
C0278562|T047||CCS_10|STAGE IV ESOPHAGEAL CANCER AJCC V7
C0278562|T047||CCS_10|STAGE IV ESOPHAGEAL CANCER
C0278562|T047||CCS_10|OESOPHAGEAL CANCER METASTATIC
C0278562|T047||CCS_10|OESOPHAGEAL NEOPLASM METASTATIC
C0278562|T047||CCS_10|ESOPHAGEAL NEOPLASM METASTATIC
C0278562|T047||CCS_10|ESOPHAGEAL CANCER METASTATIC
C0278562|T047||CCS_10|ESOPHAGEAL CANCER, METASTATIC
C0278562|T047||CCS_10|ESOPHAGEAL CANCER, STAGE IV
C0278562|T047||CCS_10|ESOPHAGUS CANCER, METASTATIC
C0278562|T047||CCS_10|ESOPHAGUS CANCER, STAGE IV
C0278562|T047||CCS_10|METASTATIC ESOPHAGEAL CANCER
C0279626|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF ESOPHAGUS
C0279626|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF ESOPHAGUS 
C0279626|T047||CCS_10|ESCC
C0279626|T047||CCS_10|ESOPHAGEAL SQUAMOUS CELL CARCINOMA
C0279626|T047||CCS_10|SQUAMOUS CELL CAR. - ESOPHAGUS
C0279626|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE ESOPHAGUS
C0279626|T047||CCS_10|OESOPHAGEAL SQUAMOUS CELL CARCINOMA STAGE UNSPECIFIED
C0279626|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF OESOPHAGUS
C0279626|T047||CCS_10|ESOPHAGEAL SQUAMOUS CELL CARCINOMA STAGE UNSPECIFIED
C0279626|T047||CCS_10|OESOPHAGEAL SQUAMOUS CELL CARCINOMA NOS
C0279626|T047||CCS_10|ESOPHAGEAL SQUAMOUS CELL CARCINOMA NOS
C0279626|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF ESOPHAGUS NOS
C0279626|T047||CCS_10|OESOPHAGEAL EPIDERMOID CARCINOMA NOS
C0279626|T047||CCS_10|OESOPHAGEAL SQUAMOUS CELL CARCINOMA
C0279626|T047||CCS_10|ESOPHAGEAL EPIDERMOID CARCINOMA NOS
C0279626|T047||CCS_10|SCC - SQUAMOUS CELL CARCINOMA OF ESOPHAGUS
C0279626|T047||CCS_10|SCC - SQUAMOUS CELL CARCINOMA OF OESOPHAGUS
C0279626|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF ESOPHAGUS 
C0279626|T047||CCS_10|ESOPHAGEAL CANCER, SQUAMOUS CELL
C0279626|T047||CCS_10|ESOPHAGUS CANCER, SQUAMOUS CELL
C0279626|T047||CCS_10|SQUAMOUS CELL ESOPHAGEAL CANCER
C0279626|T047||CCS_10|SQUAMOUS CELL ESOPHAGUS CANCER
C0279626|T047||CCS_10|ESOPHAGEAL EPIDERMOID CARCINOMA
C0279626|T047||CCS_10|ESOPHAGEAL SCC
C0279626|T047||CCS_10|ESOPHAGUS SCC
C0279626|T047||CCS_10|ESOPHAGUS SQUAMOUS CELL CARCINOMA
C0279626|T047||CCS_10|SCC OF ESOPHAGUS
C0279626|T047||CCS_10|SCC OF THE ESOPHAGUS
C2204789|T047||CCS_10|MALIGNANT SMALL CELL NEOPLASM OF ESOPHAGUS 
C2204789|T047||CCS_10|MALIGNANT SMALL CELL NEOPLASM OF ESOPHAGUS
C2011363|T047||CCS_10|GIANT CELL TYPE NEOPLASM OF ESOPHAGUS
C2011363|T047||CCS_10|GIANT CELL TYPE NEOPLASM OF ESOPHAGUS 
C2018647|T047||CCS_10|SPINDLE CELL TYPE NEOPLASM OF ESOPHAGUS 
C2018647|T047||CCS_10|SPINDLE CELL TYPE NEOPLASM OF ESOPHAGUS
C2075606|T047||CCS_10|CLEAR CELL TYPE NEOPLASM OF ESOPHAGUS 
C2075606|T047||CCS_10|CLEAR CELL TYPE NEOPLASM OF ESOPHAGUS
C2204810|T047||CCS_10|MYOSARCOMA OF ESOPHAGUS
C2204810|T047||CCS_10|MYOSARCOMA OF ESOPHAGUS 
C2204823|T047||CCS_10|MALIGNANT PLASMACYTOMA OF ESOPHAGUS 
C2204823|T047||CCS_10|MALIGNANT PLASMACYTOMA OF ESOPHAGUS
C2204825|T047||CCS_10|MALIGNANT MASTOCYTOSIS OF ESOPHAGUS
C2204825|T047||CCS_10|MALIGNANT MASTOCYTOSIS OF ESOPHAGUS 
C1333466|T047||CCS_10|SARCOMA OF ESOPHAGUS 
C1333466|T047||CCS_10|SARCOMA OF ESOPHAGUS
C1333466|T047||CCS_10|ESOPHAGEAL SARCOMA
C1333466|T047||CCS_10|ESOPHAGUS SARCOMA
C1333466|T047||CCS_10|SARCOMA OF THE ESOPHAGUS
C1333466|T047||CCS_10|SARCOMA, ESOPHAGUS
C2216771|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS STAGING 
C2216771|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS STAGING
C2216771|T047||CCS_10|MALIGNANT ESOPHAGEAL NEOPLASM STAGING
C2216771|T047||CCS_10|MALIGNANT TUMOR OF ESOPHAGUS STAGING
C2216771|T047||CCS_10|ESOPHAGEAL CANCER STAGING
C2062505|T047||CCS_10|MALIGNANT LYMPHOMA OF ESOPHAGUS 
C2062505|T047||CCS_10|MALIGNANT LYMPHOMA OF ESOPHAGUS
C1333453|T047||CCS_10|ESOPHAGEAL KAPOSI SARCOMA
C1333453|T047||CCS_10|ESOPHAGEAL KAPOSI'S SARCOMA
C1333453|T047||CCS_10|KAPOSI'S SARCOMA OF ESOPHAGUS 
C1333453|T047||CCS_10|KAPOSI'S SARCOMA OF ESOPHAGUS
C1333453|T047||CCS_10|ESOPHAGUS KAPOSI'S SARCOMA
C1333453|T047||CCS_10|KAPOSI'S SARCOMA OF THE ESOPHAGUS
C1333463|T047||CCS_10|NEUROFIBROMA OF ESOPHAGUS
C1333463|T047||CCS_10|NEUROFIBROMA OF ESOPHAGUS 
C1333463|T047||CCS_10|ESOPHAGEAL NEUROFIBROMA
C1333463|T047||CCS_10|ESOPHAGUS NEUROFIBROMA
C1333463|T047||CCS_10|NEUROFIBROMA OF THE ESOPHAGUS
C2007067|T047||CCS_10|CARCINOSARCOMA OF ESOPHAGUS 
C2007067|T047||CCS_10|CARCINOSARCOMA OF ESOPHAGUS
C1333444|T047||CCS_10|MALIGNANT CARCINOID TUMOR OF ESOPHAGUS 
C1333444|T047||CCS_10|MALIGNANT CARCINOID TUMOR OF ESOPHAGUS
C1333444|T047||CCS_10|ESOPHAGEAL NEUROENDOCRINE TUMOR G1
C1333444|T047||CCS_10|ESOPHAGEAL NET G1 (CARCINOID)
C1333444|T047||CCS_10|ESOPHAGEAL CARCINOID TUMOR
C1333444|T047||CCS_10|ESOPHAGEAL NEUROENDOCRINE TUMOR G1 (CARCINOID)
C1333444|T047||CCS_10|ESOPHAGEAL NET G1
C1333444|T047||CCS_10|CARCINOID TUMOR OF ESOPHAGUS
C1333444|T047||CCS_10|CARCINOID TUMOR OF THE ESOPHAGUS
C2204829|T047||CCS_10|BALLOON CELL MELANOMA OF ESOPHAGUS 
C2204829|T047||CCS_10|BALLOON CELL MELANOMA OF ESOPHAGUS
C2063891|T047||CCS_10|MELANOMA OF SKIN OF ESOPHAGUS
C2063891|T047||CCS_10|MELANOMA OF SKIN OF ESOPHAGUS 
C2984901|T047||CCS_10|MALIGNANT ESOPHAGEAL PERIPHERAL NERVE SHEATH TUMOR
C2216772|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS TNM STAGING
C2216772|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS TNM STAGING 
C2216772|T047||CCS_10|ESOPHAGEAL CANCER TNM STAGING
C2216772|T047||CCS_10|MALIGNANT TUMOR OF ESOPHAGUS TNM STAGING
C2216783|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS TNM STAGING REGIONAL LYMPH NODES (N) 
C2216783|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS TNM STAGING REGIONAL LYMPH NODES (N)
C2216783|T047||CCS_10|MALIGNANT ESOPHAGEAL NEOPLASM TNM STAGING OF REGIONAL LYMPH NODES (N)
C2216783|T047||CCS_10|ESOPHAGEAL CANCER TNM STAGING REGIONAL LYMPH NODES (N)
C2216783|T047||CCS_10|MALIGNANT TUMOR OF ESOPHAGUS TNM STAGING REGIONAL LYMPH NODES (N)
C2216784|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS TNM STAGING REGIONAL LYMPH NODES (N) N0 
C2216784|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS TNM STAGING REGIONAL LYMPH NODES (N) N0
C2216784|T047||CCS_10|MALIGNANT ESOPHAGEAL NEOPLASM N0
C2216784|T047||CCS_10|ESOPHAGEAL CANCER TNM STAGING REGIONAL LYMPH NODES (N) N0
C2216784|T047||CCS_10|MALIGNANT TUMOR OF ESOPHAGUS TNM STAGING REGIONAL LYMPH NODES (N) N0
C2216785|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS TNM STAGING REGIONAL LYMPH NODES (N) N1 
C2216785|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS TNM STAGING REGIONAL LYMPH NODES (N) N1
C2216785|T047||CCS_10|MALIGNANT ESOPHAGEAL NEOPLASM N1
C2216785|T047||CCS_10|MALIGNANT TUMOR OF ESOPHAGUS TNM STAGING REGIONAL LYMPH NODES (N) N1
C2216785|T047||CCS_10|ESOPHAGEAL CANCER TNM STAGING REGIONAL LYMPH NODES (N) N1
C2216776|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS TNM STAGING DISTANT METASTASIS (M) 
C2216776|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS TNM STAGING DISTANT METASTASIS (M)
C2216776|T047||CCS_10|MALIGNANT ESOPHAGEAL NEOPLASM TNM STAGING OF DISTANT METASTASIS (M)
C2216776|T047||CCS_10|MALIGNANT TUMOR OF ESOPHAGUS TNM STAGING DISTANT METASTASIS (M)
C2216776|T047||CCS_10|ESOPHAGEAL CANCER TNM STAGING DISTANT METASTASIS (M)
C2216775|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS TNM STAGING DISTAL METASTASIS (M) M1B
C2216775|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS TNM STAGING DISTAL METASTASIS (M) M1B 
C2216775|T047||CCS_10|MALIGNANT ESOPHAGEAL NEOPLASM M1B
C2216775|T047||CCS_10|MALIGNANT TUMOR OF ESOPHAGUS TNM STAGING DISTAL METASTASIS (M) M1B
C2216775|T047||CCS_10|ESOPHAGEAL CANCER TNM STAGING DISTAL METASTASIS (M) M1B
C2216773|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS TNM STAGING DISTAL METASTASIS (M) M0 
C2216773|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS TNM STAGING DISTAL METASTASIS (M) M0
C2216773|T047||CCS_10|MALIGNANT ESOPHAGEAL NEOPLASM M0
C2216773|T047||CCS_10|MALIGNANT TUMOR OF ESOPHAGUS TNM STAGING DISTAL METASTASIS (M) M0
C2216773|T047||CCS_10|ESOPHAGEAL CANCER TNM STAGING DISTAL METASTASIS (M) M0
C2216774|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS TNM STAGING DISTAL METASTASIS (M) M1A
C2216774|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS TNM STAGING DISTAL METASTASIS (M) M1A 
C2216774|T047||CCS_10|MALIGNANT ESOPHAGEAL NEOPLASM M1A
C2216774|T047||CCS_10|ESOPHAGEAL CANCER TNM STAGING DISTAL METASTASIS (M) M1A
C2216774|T047||CCS_10|MALIGNANT TUMOR OF ESOPHAGUS TNM STAGING DISTAL METASTASIS (M) M1A
C3165092|T047||CCS_10|LEIOMYOSARCOMA OF LOWER ESOPHAGUS
C3165092|T047||CCS_10|LEIOMYOSARCOMA OF LOWER ESOPHAGUS 
C3165092|T047||CCS_10|LEIOMYOSARCOMA OF LOWER OESOPHAGUS
C3165092|T047||CCS_10|MALIGNANT NEOPLASM MYOSARCOMA LEIOMYOSARCOMA LOWER ESOPHAGUS
C3165092|T047||CCS_10|LEIOMYOSARCOMA OF LOWER ESOPHAGUS 
C3165036|T047||CCS_10|LYMPHOMA OF LOWER ESOPHAGUS 
C3165036|T047||CCS_10|LYMPHOMA OF LOWER ESOPHAGUS
C3165036|T047||CCS_10|LYMPHOMA OF LOWER OESOPHAGUS
C3165036|T047||CCS_10|ESOPHAGEAL MALIGNANT LYMPHOMA OF LOWER ESOPHAGUS
C3165036|T047||CCS_10|LYMPHOMA OF LOWER ESOPHAGUS 
C2111603|T047||CCS_10|LARGE CELL CARCINOMA OF ESOPHAGUS 
C2111603|T047||CCS_10|LARGE CELL CARCINOMA OF ESOPHAGUS
C2111715|T047||CCS_10|LARGE CELL NEUROENDOCRINE CARCINOMA OF ESOPHAGUS
C2111715|T047||CCS_10|LARGE CELL NEUROENDOCRINE CARCINOMA OF ESOPHAGUS 
C2111604|T047||CCS_10|LARGE CELL CARCINOMA OF ESOPHAGUS WITH RHABDOID PHENOTYPE 
C2111604|T047||CCS_10|LARGE CELL CARCINOMA OF ESOPHAGUS WITH RHABDOID PHENOTYPE
C2012076|T047||CCS_10|GLASSY CELL CARCINOMA OF ESOPHAGUS 
C2012076|T047||CCS_10|GLASSY CELL CARCINOMA OF ESOPHAGUS
C2188058|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF ESOPHAGUS 
C2188058|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF ESOPHAGUS
C2188058|T047||CCS_10|ESOPHAGEAL UNDIFFERENTIATED CARCINOMA
C2009877|T047||CCS_10|FUSIFORM TYPE SMALL CELL CARCINOMA OF ESOPHAGUS 
C2009877|T047||CCS_10|FUSIFORM TYPE SMALL CELL CARCINOMA OF ESOPHAGUS
C2037374|T047||CCS_10|SUPERFICIAL SPREADING MELANOMA OF ESOPHAGUS
C2037374|T047||CCS_10|SUPERFICIAL SPREADING MELANOMA OF ESOPHAGUS 
C2204836|T047||CCS_10|MIXED EPITHELIOID AND SPINDLE CELL MELANOMA OF ESOPHAGUS 
C2204836|T047||CCS_10|MIXED EPITHELIOID AND SPINDLE CELL MELANOMA OF ESOPHAGUS
C2063886|T047||CCS_10|ADENOSQUAMOUS CARCINOMA OF ESOPHAGUS
C2063886|T047||CCS_10|ADENOSQUAMOUS CARCINOMA OF ESOPHAGUS 
C2063886|T047||CCS_10|ESOPHAGEAL ADENOSQUAMOUS CARCINOMA
C1333441|T047||CCS_10|ADENOID CYSTIC CARCINOMA OF ESOPHAGUS
C1333441|T047||CCS_10|ADENOID CYSTIC CARCINOMA OF ESOPHAGUS 
C1333441|T047||CCS_10|ESOPHAGEAL ADENOID CYSTIC CARCINOMA
C1333441|T047||CCS_10|ESOPHAGUS ADENOID CYSTIC CARCINOMA
C1333441|T047||CCS_10|ADENOID CYSTIC CARCINOMA OF THE ESOPHAGUS
C1333441|T047||CCS_10|ADENOID CYSTIC CARCINOMA, ESOPHAGUS
C1333441|T047||CCS_10|ADENOID CYSTIC ESOPHAGUS CARCINOMA
C1333461|T047||CCS_10|MUCOEPIDERMOID CARCINOMA OF ESOPHAGUS
C1333461|T047||CCS_10|MUCOEPIDERMOID CARCINOMA OF ESOPHAGUS 
C1333461|T047||CCS_10|ESOPHAGEAL MUCOEPIDERMOID CARCINOMA
C1333461|T047||CCS_10|MUCOEPIDERMOID CARCINOMA OF THE ESOPHAGUS
C1333461|T047||CCS_10|MUCOEPIDERMOID ESOPHAGEAL CARCINOMA
C1333461|T047||CCS_10|MUCOEPIDERMOID ESOPHAGUS CARCINOMA
C2237936|T047||CCS_10|X-RAY UGI BA SWALLOW- ESOPHAGEAL MASS MALIGNANT NEOPLASM ___
C2237936|T047||CCS_10|BARIUM SWALLOW: MALIGNANT NEOPLASM OF ESOPHAGUS
C2237936|T047||CCS_10|BARIUM SWALLOW: MALIGNANT NEOPLASM OF ESOPHAGUS 
C2204790|T047||CCS_10|MALIGNANT EPITHELIOMA OF ESOPHAGUS 
C2204790|T047||CCS_10|MALIGNANT EPITHELIOMA OF ESOPHAGUS
C2204834|T047||CCS_10|EPITHELIOID CELL MELANOMA OF ESOPHAGUS 
C2204834|T047||CCS_10|EPITHELIOID CELL MELANOMA OF ESOPHAGUS
C1282473|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT NEOPLASM OF ESOPHAGUS
C1282473|T047||CCS_10|ESOPHAGEAL MALIGNANT NEOPLASM, LOCAL RECURRENCE
C1282473|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT NEOPLASM OF ESOPHAGUS 
C1282473|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOR OF ESOPHAGUS 
C1282473|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOR OF ESOPHAGUS
C1282473|T047||CCS_10|LOCAL RECURRENCE OF MALIGNANT TUMOUR OF OESOPHAGUS
C0349048|T047||CCS_10|MALIGNANT NEOPLASM, OVERLAPPING LESION OF ESOPHAGUS
C0349048|T047||CCS_10|MALIGNANT NEOPLASM, OVERLAPPING LESION OF OESOPHAGUS
C0349048|T047||CCS_10|MALIGNANT NEOPLASM, OVERLAPPING LESION OF ESOPHAGUS 
C0349048|T047||CCS_10|OVERLAPPING MALIGNANT NEOPLASM OF ESOPHAGUS 
C0349048|T047||CCS_10|OVERLAPPING MALIGNANT NEOPLASM OF ESOPHAGUS
C0349048|T047||CCS_10|OVERLAPPING MALIGNANT NEOPLASM OF OESOPHAGUS
C0346619|T047||CCS_10|MALIGNANT NEOPLASM OF CARDIOESOPHAGEAL JUNCTION OF STOMACH
C0346619|T047||CCS_10|MALIGNANT NEOPLASM OF GASTRO-ESOPHAGEAL JUNCTION
C0346619|T047||CCS_10|MALIGNANT NEOPLASM OF CARDIOESOPHAGEAL JUNCTION OF STOMACH 
C0346619|T047||CCS_10|ESOPHAGEAL NEOPLASM MALIGNANT CARDIOESOPHAGEAL JUNCTION OF STOMACH
C0346619|T047||CCS_10|MALIGNANT NEOPLASM OF CARDIO-ESOPHAGEAL JUNCTION OF STOMACH
C0346619|T047||CCS_10|MALIGNANT NEOPLASM OF CARDIO-OESOPHAGEAL JUNCTION OF STOMACH
C0346619|T047||CCS_10|MALIGNANT NEOPLASM OF GASTRO-OESOPHAGEAL JUNCTION
C0346619|T047||CCS_10|MALIGNANT NEOPLASM OF CARDIOESOPHAGEAL JUNCTION OF STOMACH 
C1300083|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF OESOPHAGUS
C1300083|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF ESOPHAGUS 
C1300083|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF ESOPHAGUS
C1300083|T047||CCS_10|PRIMARY MALIGNANT NEOPLASM OF ESOPHAGUS 
C1300083|T047||CCS_10|ESOPHAGEAL MALIGNANT NEOPLASM PRIMARY
C0686055|T047||CCS_10|METASTATIC NEOPLASM TO THE ESOPHAGUS
C0686055|T047||CCS_10|METASTASES TO OESOPHAGUS
C0686055|T047||CCS_10|ESOPHAGEAL MALIGNANT NEOPLASM SECONDARY
C0686055|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF ESOPHAGUS
C0686055|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF ESOPHAGUS 
C0686055|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO THE ESOPHAGUS
C0686055|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM IN THE ESOPHAGUS
C0686055|T047||CCS_10|CANCER METASTATIC TO ESOPHAGUS
C0686055|T047||CCS_10|METASTASES TO ESOPHAGUS
C0686055|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO ESOPHAGUS
C0686055|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF ESOPHAGUS 
C0686055|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF OESOPHAGUS
C0686055|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO OESOPHAGUS
C0686055|T047||CCS_10|METASTATIC MALIGNANT NEOPLASM TO ESOPHAGUS, NOS
C0686055|T047||CCS_10|SECONDARY MALIGNANT NEOPLASM OF ESOPHAGUS, NOS
C0686055|T047||CCS_10|ESOPHAGEAL METASTASIS
C0686055|T047||CCS_10|METASTASES TO THE ESOPHAGUS
C0686055|T047||CCS_10|METASTASIS TO ESOPHAGUS
C0686055|T047||CCS_10|METASTASIS TO THE ESOPHAGUS
C0686055|T047||CCS_10|METASTATIC TUMOR TO THE ESOPHAGUS
C4065138|T047||CCS_10|ESOPHAGOSCOPY MASS MALIGNANT NEOPLASM
C4065138|T047||CCS_10|ESOPHAGOSCOPY MASS MALIGNANT NEOPLASM 
C0346618|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS, STOMACH, AND DUODENUM
C0346618|T047||CCS_10|DIGESTIVE NEOPLASM MALIGNANT OF ESOPHAGUS, STOMACH, AND DUODENUM
C0346618|T047||CCS_10|MALIGNANT NEOPLASM OF ESOPHAGUS, STOMACH, AND DUODENUM 
C0346618|T047||CCS_10|MALIGNANT TUMOR OF ESOPHAGUS, STOMACH AND DUODENUM
C0346618|T047||CCS_10|MALIGNANT TUMOUR OF OESOPHAGUS, STOMACH AND DUODENUM
C0346618|T047||CCS_10|MALIGNANT TUMOR OF ESOPHAGUS, STOMACH AND DUODENUM 
C0279865|T047||CCS_10|CELLULAR DIAGNOSIS, ESOPHAGEAL CANCER
C0279865|T047||CCS_10|ESOPHAGEAL CANCER, CELLULAR DIAGNOSIS
C0279865|T047||CCS_10|ESOPHAGUS CANCER CELLULAR DIAGNOSIS
C0280257|T047||CCS_10|STAGE, ESOPHAGEAL CANCER
C0280257|T047||CCS_10|ESOPHAGEAL CANCER, STAGE
C1333459|T047||CCS_10|PRIMARY ESOPHAGEAL LYMPHOMA
C1333459|T047||CCS_10|ESOPHAGEAL LYMPHOMA
C1333459|T047||CCS_10|ESOPHAGUS LYMPHOMA
C1333459|T047||CCS_10|LYMPHOMA OF ESOPHAGUS
C1333459|T047||CCS_10|LYMPHOMA OF THE ESOPHAGUS
C1334579|T047||CCS_10|MALIGNANT ESOPHAGEAL NEOPLASM BY TOPOGRAPHIC REGION
C1333460|T047||CCS_10|ESOPHAGEAL MELANOMA
C1333460|T047||CCS_10|ESOPHAGUS MELANOMA
C1333460|T047||CCS_10|MELANOMA OF ESOPHAGUS
C1333460|T047||CCS_10|MELANOMA OF THE ESOPHAGUS
C1334578|T047||CCS_10|MALIGNANT ESOPHAGEAL NEOPLASM BY ANATOMIC REGION
C0585126|T047||CCS_10|PERFORATED CARCINOMA OF ESOPHAGUS 
C0585126|T047||CCS_10|ESOPHAGEAL NEOPLASM MALIGNANT CARCINOMA, PERFORATED
C0585126|T047||CCS_10|PERFORATED CARCINOMA OF ESOPHAGUS
C0585126|T047||CCS_10|PERFORATED CARCINOMA OF OESOPHAGUS
C0585126|T047||CCS_10|PERFORATED CARCINOMA OF ESOPHAGUS 
C1276562|T047||CCS_10|T3: ESOPHAGEAL TUMOR INVADES ADVENTITIA 
C1276562|T047||CCS_10|T3: ESOPHAGEAL TUMOR INVADES ADVENTITIA
C1276562|T047||CCS_10|T3: OESOPHAGEAL TUMOUR INVADES ADVENTITIA
C1276562|T047||CCS_10|T3: ESOPHAGEAL TUMOR INVADES ADVENTITIA (TUMOR STAGING)
C2204817|T047||CCS_10|ANGIOIMMUNOBLASTIC T-CELL LYMPHOMA OF ESOPHAGUS
C2204817|T047||CCS_10|ANGIOIMMUNOBLASTIC T-CELL LYMPHOMA OF ESOPHAGUS 
C2204817|T047||CCS_10|ANGIOIMMUNOBLASTIC LYMPHADENOPATHY WITH DYSPROTEINEMIA (AILD) OF ESOPHAGUS
C2204821|T047||CCS_10|NK/T-CELL LYMPHOMA OF ESOPHAGUS
C2204821|T047||CCS_10|NK/T-CELL LYMPHOMA OF ESOPHAGUS 
C2113687|T047||CCS_10|PRECURSOR CELL LYMPHOBLASTIC LYMPHOMA OF ESOPHAGUS 
C2113687|T047||CCS_10|PRECURSOR CELL LYMPHOBLASTIC LYMPHOMA OF ESOPHAGUS
C2204826|T047||CCS_10|MAST CELL SARCOMA OF ESOPHAGUS 
C2204826|T047||CCS_10|MAST CELL SARCOMA OF ESOPHAGUS
C2113618|T047||CCS_10|PRECURSOR B-CELL LYMPHOBLASTIC LYMPHOMA OF ESOPHAGUS
C2113618|T047||CCS_10|PRECURSOR B-CELL LYMPHOBLASTIC LYMPHOMA OF ESOPHAGUS 
C2204822|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF ESOPHAGUS
C2204822|T047||CCS_10|MALIGNANT HISTIOCYTOSIS OF ESOPHAGUS 
C2204837|T047||CCS_10|SEZARY SYNDROME OF ESOPHAGUS
C2204837|T047||CCS_10|SEZARY SYNDROME OF ESOPHAGUS 
C2204815|T047||CCS_10|MARGINAL ZONE B-CELL LYMPHOMA OF ESOPHAGUS
C2204815|T047||CCS_10|MARGINAL ZONE B-CELL LYMPHOMA OF ESOPHAGUS 
C2113758|T047||CCS_10|PRECURSOR T-CELL LYMPHOBLASTIC LYMPHOMA OF ESOPHAGUS 
C2113758|T047||CCS_10|PRECURSOR T-CELL LYMPHOBLASTIC LYMPHOMA OF ESOPHAGUS
C2204816|T047||CCS_10|MATURE T-CELL LYMPHOMA OF ESOPHAGUS
C2204816|T047||CCS_10|MATURE T-CELL LYMPHOMA OF ESOPHAGUS 
C0345819|T047||CCS_10|GASTRIC MALIGNANT CARCINOMA LESSER CURVE
C0345819|T047||CCS_10|CARCINOMA OF LESSER CURVE OF STOMACH 
C0345819|T047||CCS_10|CARCINOMA OF LESSER CURVE OF STOMACH
C0345819|T047||CCS_10|CARCINOMA OF LESSER CURVE OF STOMACH 
C0153423|T047||CCS_10|MALIGNANT NEOPLASM OF GREATER CURVATURE OF STOMACH, UNSPECIFIED
C0153423|T047||CCS_10|GREATER CURVATURE OF STOMACH, UNSPECIFIED
C0153423|T047||CCS_10|MALIGNANT NEOPLASM OF GREATER CURVATURE OF STOMACH
C0153423|T047||CCS_10|MALIGNANT NEOPLASM OF GREATER CURVATURE OF STOMACH 
C0153423|T047||CCS_10|MALIGNANT TUMOR OF GREATER CURVATURE OF STOMACH
C0153423|T047||CCS_10|MAL NEO STOM GREAT CURV
C0153423|T047||CCS_10|MALIGNANT NEOPLASM OF GREATER CURVATURE OF STOMACH, UNSP
C0153423|T047||CCS_10|CA GREATER CURVATURE - STOMACH
C0153423|T047||CCS_10|MALIGNANT NEOPLASM OF GREATER CURVE OF STOMACH UNSPECIFIED
C0153423|T047||CCS_10|CA GREATER CURVATURE - STOMACH 
C0153423|T047||CCS_10|MALIGNANT NEOPLASM OF GREATER CURVE OF STOMACH UNSPECIFIED 
C0153423|T047||CCS_10|MALIGNANT TUMOR OF GREATER CURVE OF STOMACH
C0153423|T047||CCS_10|MALIGNANT TUMOUR OF GREATER CURVE OF STOMACH
C0153423|T047||CCS_10|MALIGNANT TUMOR OF GREATER CURVE OF STOMACH 
C0153423|T047||CCS_10|MALIGNANT NEOPLASM OF GREATER CURVATURE OF STOMACH, NOS
C0699791|T047||CCS_10|CANCER OF STOMACH
C0699791|T047||CCS_10|CARCINOMA OF STOMACH 
C0699791|T047||CCS_10|CARCINOMA OF STOMACH
C0699791|T047||CCS_10|GASTRIC CARCINOMA
C0699791|T047||CCS_10|CARCINOMA;STOMACH
C0699791|T047||CCS_10|GASTRIC CANCER
C0699791|T047||CCS_10|STOMACH CANCER
C0699791|T047||CCS_10|CARCINOMA OF STOMACH 
C0699791|T047||CCS_10|GASTRIC CANCER, NOS
C0699791|T047||CCS_10|CARCINOMA GASTRIC
C0699791|T047||CCS_10|CARCINOMA STOMACH
C0699791|T047||CCS_10|STOMACH CARCINOMA
C0699791|T047||CCS_10|STOMACH (GASTRIC) CANCER
C0699791|T047||CCS_10|CANCER OF THE STOMACH
C0699791|T047||CCS_10|CARCINOMA OF THE STOMACH
C2204845|T047||CCS_10|MALIGNANT EPITHELIOMA OF STOMACH 
C2204845|T047||CCS_10|MALIGNANT EPITHELIOMA OF STOMACH
C2111678|T047||CCS_10|LARGE CELL CARCINOMA OF STOMACH 
C2111678|T047||CCS_10|LARGE CELL CARCINOMA OF STOMACH
C2012116|T047||CCS_10|GLASSY CELL CARCINOMA OF STOMACH 
C2012116|T047||CCS_10|GLASSY CELL CARCINOMA OF STOMACH
C1336858|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF STOMACH
C1336858|T047||CCS_10|ANAPLASTIC CARCINOMA OF STOMACH 
C1336858|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF STOMACH 
C1336858|T047||CCS_10|ANAPLASTIC CARCINOMA OF STOMACH
C1336858|T047||CCS_10|UNDIFFERENTIATED GASTRIC CARCINOMA
C1336858|T047||CCS_10|ANAPLASTIC CARCINOMA OF THE STOMACH
C1336858|T047||CCS_10|ANAPLASTIC GASTRIC CARCINOMA
C1336858|T047||CCS_10|UNDIFFERENTIATED CARCINOMA OF THE STOMACH
C2082464|T047||CCS_10|PLEOMORPHIC CARCINOMA OF STOMACH
C2082464|T047||CCS_10|PLEOMORPHIC CARCINOMA OF STOMACH 
C2011266|T047||CCS_10|GIANT CELL CARCINOMA OF STOMACH 
C2011266|T047||CCS_10|GIANT CELL CARCINOMA OF STOMACH
C2018406|T047||CCS_10|SPINDLE CELL CARCINOMA OF STOMACH 
C2018406|T047||CCS_10|SPINDLE CELL CARCINOMA OF STOMACH
C2011231|T047||CCS_10|GIANT CELL AND SPINDLE CELL CARCINOMA OF STOMACH
C2011231|T047||CCS_10|GIANT CELL AND SPINDLE CELL CARCINOMA OF STOMACH 
C2142936|T047||CCS_10|PSEUDOSARCOMATOUS CARCINOMA OF STOMACH
C2142936|T047||CCS_10|PSEUDOSARCOMATOUS CARCINOMA OF STOMACH 
C2111818|T047||CCS_10|POLYGONAL CELL CARCINOMA OF STOMACH
C2111818|T047||CCS_10|POLYGONAL CELL CARCINOMA OF STOMACH 
C2010505|T047||CCS_10|CARCINOMA OF STOMACH WITH OSTEOCLAST-LIKE GIANT CELLS
C2010505|T047||CCS_10|CARCINOMA OF STOMACH WITH OSTEOCLAST-LIKE GIANT CELLS 
C2010505|T047||CCS_10|GASTRIC CARCINOMA WITH OSTEOCLAST-LIKE GIANT CELLS
C2033236|T047||CCS_10|PAPILLARY CARCINOMA OF STOMACH 
C2033236|T047||CCS_10|PAPILLARY CARCINOMA OF STOMACH
C2189366|T047||CCS_10|VERRUCOUS CARCINOMA OF STOMACH
C2189366|T047||CCS_10|VERRUCOUS CARCINOMA OF STOMACH 
C2010501|T047||CCS_10|DIFFUSE CARCINOMA OF STOMACH 
C2010501|T047||CCS_10|DIFFUSE CARCINOMA OF STOMACH
C2010503|T047||CCS_10|PARIETAL CELL CARCINOMA OF STOMACH 
C2010503|T047||CCS_10|PARIETAL CELL CARCINOMA OF STOMACH
C2017458|T047||CCS_10|SOLID CARCINOMA OF STOMACH
C2017458|T047||CCS_10|SOLID CARCINOMA OF STOMACH 
C2010504|T047||CCS_10|CARCINOMA SIMPLEX OF STOMACH 
C2010504|T047||CCS_10|CARCINOMA SIMPLEX OF STOMACH
C2010502|T047||CCS_10|NEUROENDOCRINE CARCINOMA OF STOMACH 
C2010502|T047||CCS_10|NEUROENDOCRINE CARCINOMA OF STOMACH
C2204850|T047||CCS_10|MEDULLARY CARCINOMA OF STOMACH
C2204850|T047||CCS_10|MEDULLARY CARCINOMA OF STOMACH 
C2204851|T047||CCS_10|EPITHELIAL-MYOEPITHELIAL CARCINOMA OF STOMACH 
C2204851|T047||CCS_10|EPITHELIAL-MYOEPITHELIAL CARCINOMA OF STOMACH
C2064167|T047||CCS_10|SIGNET RING CELL CARCINOMA OF STOMACH
C2064167|T047||CCS_10|SIGNET RING CELL CARCINOMA OF STOMACH 
C2064167|T047||CCS_10|GASTRIC SIGNET RING CELL CARCINOMA
C1333761|T047||CCS_10|ADENOSQUAMOUS CARCINOMA OF STOMACH 
C1333761|T047||CCS_10|ADENOSQUAMOUS CARCINOMA OF STOMACH
C1333761|T047||CCS_10|GASTRIC ADENOSQUAMOUS CARCINOMA
C1333761|T047||CCS_10|ADENOSQUAMOUS CARCINOMA OF THE STOMACH
C1333789|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF STOMACH 
C1333789|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF STOMACH
C1333789|T047||CCS_10|GASTRIC SQUAMOUS CELL CARCINOMA
C1333789|T047||CCS_10|SQUAMOUS CELL CARCINOMA OF THE STOMACH
C1333788|T047||CCS_10|SMALL CELL CARCINOMA OF STOMACH 
C1333788|T047||CCS_10|SMALL CELL CARCINOMA OF STOMACH
C1333788|T047||CCS_10|GASTRIC SMALL CELL CARCINOMA
C1333788|T047||CCS_10|GASTRIC SMALL CELL NEUROENDOCRINE CARCINOMA
C1333788|T047||CCS_10|OAT CELL CARCINOMA OF STOMACH
C1333788|T047||CCS_10|GASTRIC OAT CELL CARCINOMA
C1333788|T047||CCS_10|OAT CELL CARCINOMA OF THE STOMACH
C1333788|T047||CCS_10|SMALL CELL CARCINOMA OF THE STOMACH
C2983703|T047||CCS_10|GASTRIC CARCINOMA BY AJCC V6 STAGE
C2984086|T047||CCS_10|GASTRIC CARCINOMA BY AJCC V7 STAGE
C3272409|T047||CCS_10|GASTRIC NEUROENDOCRINE CARCINOMA
C3272409|T047||CCS_10|GASTRIC NEC
C3272411|T047||CCS_10|GASTRIC MIXED ADENONEUROENDOCRINE CARCINOMA
C3272411|T047||CCS_10|GASTRIC MANEC
C0345804|T047||CCS_10|GASTRIC MALIGNANT CARCINOMA BODY
C0345804|T047||CCS_10|CARCINOMA OF BODY OF STOMACH 
C0345804|T047||CCS_10|CARCINOMA OF BODY OF STOMACH
C0345804|T047||CCS_10|CARCINOMA OF BODY OF STOMACH 
C0345804|T047||CCS_10|GASTRIC BODY CANCER
C0345804|T047||CCS_10|GASTRIC BODY CARCINOMA
C0345804|T047||CCS_10|CANCER OF BODY OF STOMACH
C0345804|T047||CCS_10|CANCER OF GASTRIC BODY
C0345804|T047||CCS_10|CANCER OF THE BODY OF THE STOMACH
C0345804|T047||CCS_10|CANCER OF THE GASTRIC BODY
C0345804|T047||CCS_10|CARCINOMA OF GASTRIC BODY
C0345804|T047||CCS_10|CARCINOMA OF THE BODY OF THE STOMACH
C0345804|T047||CCS_10|CARCINOMA OF THE GASTRIC BODY
C0345814|T047||CCS_10|GASTRIC MALIGNANT CARCINOMA PYLORUS
C0345814|T047||CCS_10|CARCINOMA OF PYLORUS 
C0345814|T047||CCS_10|CARCINOMA OF PYLORUS
C0345814|T047||CCS_10|PYLORIC CARCINOMA
C0345814|T047||CCS_10|CARCINOMA OF PYLORUS 
C0345809|T047||CCS_10|GASTRIC MALIGNANT CARCINOMA PYLORIC ANTRUM
C0345809|T047||CCS_10|CARCINOMA OF PYLORIC ANTRUM
C0345809|T047||CCS_10|CARCINOMA OF PYLORIC ANTRUM 
C0345809|T047||CCS_10|CARCINOMA OF PYLORIC ANTRUM 
C0345794|T047||CCS_10|GASTRIC MALIGNANT CARCINOMA CARDIA
C0345794|T047||CCS_10|CARCINOMA OF CARDIA
C0345794|T047||CCS_10|CARCINOMA OF CARDIA 
C0345794|T047||CCS_10|CARCINOMA OF CARDIA 
C0345799|T047||CCS_10|CARCINOMA OF FUNDUS OF STOMACH
C0345799|T047||CCS_10|CARCINOMA OF FUNDUS OF STOMACH 
C0345799|T047||CCS_10|GASTRIC MALIGNANT CARCINOMA FUNDUS
C0345799|T047||CCS_10|CARCINOMA OF FUNDUS OF STOMACH 
C0345799|T047||CCS_10|GASTRIC FUNDUS CANCER
C0345799|T047||CCS_10|GASTRIC FUNDUS CARCINOMA
C0345799|T047||CCS_10|CANCER OF FUNDUS OF STOMACH
C0345799|T047||CCS_10|CANCER OF GASTRIC FUNDUS
C0345799|T047||CCS_10|CANCER OF THE FUNDUS OF THE STOMACH
C0345799|T047||CCS_10|CANCER OF THE GASTRIC FUNDUS
C0345799|T047||CCS_10|CARCINOMA OF GASTRIC FUNDUS
C0345799|T047||CCS_10|CARCINOMA OF THE FUNDUS OF THE STOMACH
C0345799|T047||CCS_10|CARCINOMA OF THE GASTRIC FUNDUS
C0740488|T047||CCS_10|GASTRIC MALIGNANT CARCINOMA GREATER CURVE
C0740488|T047||CCS_10|CARCINOMA OF GREATER CURVE OF STOMACH 
C0740488|T047||CCS_10|CARCINOMA OF GREATER CURVE OF STOMACH
C0740488|T047||CCS_10|CARCINOMA OF GREATER CURVE OF STOMACH 
C0349530|T047||CCS_10|EARLY GASTRIC CANCER
C0349530|T047||CCS_10|GASTRIC NEOPLASM MALIGNANT EARLY CANCER
C0349530|T047||CCS_10|EARLY GASTRIC CANCER 
C0349530|T047||CCS_10|EGC - EARLY GASTRIC CANCER
C0349530|T047||CCS_10|EARLY GASTRIC CANCER 
C0349530|T047||CCS_10|MICROINVASIVE GASTRIC CANCER
C0349530|T047||CCS_10|SUPERFICIAL GASTRIC CANCER
C0349530|T047||CCS_10|SUPERFICIAL SPREADING GASTRIC CANCER
C0349530|T047||CCS_10|SURFACE GASTRIC CANCER
C0349531|T047||CCS_10|LATE GASTRIC CANCER 
C0349531|T047||CCS_10|LATE GASTRIC CANCER
C0349531|T047||CCS_10|GASTRIC NEOPLASM MALIGNANT LATE CANCER
C0349531|T047||CCS_10|LGC - LATE GASTRIC CANCER
C0349531|T047||CCS_10|LATE GASTRIC CANCER 
C3899661|T047||CCS_10|CHILDHOOD GASTRIC CARCINOMA
C0280253|T047||CCS_10|STAGE, GASTRIC CANCER
C0280253|T047||CCS_10|GASTRIC CANCER STAGE
C0280253|T047||CCS_10|STOMACH CANCER STAGE
C0279889|T047||CCS_10|CELLULAR DIAGNOSIS, GASTRIC CANCER
C0279889|T047||CCS_10|GASTRIC CANCER CELLULAR DIAGNOSIS
C0279889|T047||CCS_10|STOMACH CANCER CELLULAR DIAGNOSIS
C1333763|T047||CCS_10|GASTRIC CARDIA CANCER
C1333763|T047||CCS_10|GASTRIC CARDIA CARCINOMA
C1333763|T047||CCS_10|CANCER OF GASTRIC CARDIA
C1333763|T047||CCS_10|CANCER OF THE GASTRIC CARDIA
C1333763|T047||CCS_10|CARCINOMA OF CARDIA OF STOMACH
C1333763|T047||CCS_10|CARCINOMA OF GASTRIC CARDIA
C1333763|T047||CCS_10|CARCINOMA OF THE CARDIA OF THE STOMACH
C1333763|T047||CCS_10|CARCINOMA OF THE GASTRIC CARDIA
C0278502|T047||CCS_10|GASTRIC CANCER RECURRENT
C0278502|T047||CCS_10|RECURRENT GASTRIC CARCINOMA
C0278502|T047||CCS_10|RECURRENT GASTRIC CANCER
C0278502|T047||CCS_10|STOMACH CANCER RECURRENT
C0278502|T047||CCS_10|GASTRIC CARCINOMA RECURRENT
C0278502|T047||CCS_10|STOMACH CARCINOMA RECURRENT
C0278502|T047||CCS_10|GASTRIC CANCER, RECURRENT
C0278502|T047||CCS_10|STOMACH CANCER, RECURRENT
C0278502|T047||CCS_10|GASTRIC CARCINOMA, RECURRENT
C0278502|T047||CCS_10|RECURRENT CANCER OF STOMACH
C0278502|T047||CCS_10|RECURRENT CANCER OF THE STOMACH
C0278502|T047||CCS_10|RECURRENT CARCINOMA OF STOMACH
C0278502|T047||CCS_10|RECURRENT CARCINOMA OF THE STOMACH
C0278502|T047||CCS_10|RECURRENT STOMACH CANCER
C0278502|T047||CCS_10|RECURRENT STOMACH CARCINOMA
C1333787|T047||CCS_10|GASTRIC PYLORUS CANCER
C1333787|T047||CCS_10|GASTRIC PYLORUS CARCINOMA
C1333787|T047||CCS_10|CANCER OF GASTRIC PYLORUS
C1333787|T047||CCS_10|CANCER OF PYLORUS OF STOMACH
C1333787|T047||CCS_10|CANCER OF THE GASTRIC PYLORUS
C1333787|T047||CCS_10|CANCER OF THE PYLORUS OF THE STOMACH
C1333787|T047||CCS_10|CARCINOMA OF GASTRIC PYLORUS
C1333787|T047||CCS_10|CARCINOMA OF PYLORUS OF STOMACH
C1333787|T047||CCS_10|CARCINOMA OF THE GASTRIC PYLORUS
C1333787|T047||CCS_10|CARCINOMA OF THE PYLORUS OF THE STOMACH
C0278701|T047||CCS_10|GASTRIC ADENOCARCINOMA
C0278701|T047||CCS_10|ADENOCARCINOMA OF STOMACH
C0278701|T047||CCS_10|ADENOCARCINOMA OF STOMACH 
C0278701|T047||CCS_10|ADENOCARCINOMA GASTRIC
C0278701|T047||CCS_10|ADENOCARCINOMA - STOMACH
C0278701|T047||CCS_10|ADENOCARCINOMA OF THE STOMACH
C0278701|T047||CCS_10|CANCER OF STOMACH, ADENOCARCINOMA
C0278701|T047||CCS_10|ADENOCARCINOMA OF STOMACH 
C0278701|T047||CCS_10|GASTRIC CANCER, ADENOCARCINOMA
C0278701|T047||CCS_10|STOMACH CANCER, ADENOCARCINOMA
C0278701|T047||CCS_10|STOMACH, ADENOCARCINOMA OF THE
C0278701|T047||CCS_10|STOMACH ADENOCARCINOMA
C0809960|T047|15|CCS_10|CANCER OF RECTUM AND ANUS|CANCER OF RECTUM AND ANUS
C0809962|T047|18|CCS_10|CANCER OF OTHER GI ORGANS; PERITONEUM|CANCER OF OTHER GI ORGANS; PERITONEUM
