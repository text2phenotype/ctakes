C0524909|T047|61977001|SNOMEDCT_US|HEPATITIS B, CHRONIC|CHRONIC TYPE B VIRAL HEPATITIS (DISORDER)
C0744831|T047|266539002|SNOMEDCT_US|CHRONIC ACTIVE HEPATITIS B|CHRONIC ACTIVE HEPATITIS B
C0276612|T047|50167007|SNOMEDCT_US|CHRONIC ACTIVE TYPE B VIRAL HEPATITIS|CHRONIC ACTIVE TYPE B VIRAL HEPATITIS (DISORDER)
C0276613|T047|38662009|SNOMEDCT_US|CHRONIC PERSISTENT TYPE B VIRAL HEPATITIS|CHRONIC PERSISTENT TYPE B VIRAL HEPATITIS (DISORDER)
C0744833|T047||SNOMEDCT_US|HEPATITIS B CHRONIC PERSISTENT INFECTION
C1827079|T047|424340000|SNOMEDCT_US|HEPATIC COMA DUE TO CHRONIC HEPATITIS B|CHRONIC HEPATITIS B WITH HEPATIC COMA
C2074982|T047||SNOMEDCT_US|CHRONIC VIRAL HEPATITIS DELTA INFECTION WITH HEPATITIS B 
C2118427|T047||SNOMEDCT_US|ACUTE HEPATITIS D INFECTION WITH CHRONIC HEPATITIS B
C2074977|T047||SNOMEDCT_US|CHRONIC HEPATITIS B INFECTION WITH FULMINANT HEPATIC FAILURE
C2074978|T047||SNOMEDCT_US|CHRONIC HEPATITIS B INFECTION WITH HEPATIC COMA
C4075603|T047|713966008|SNOMEDCT_US|OCCULT CHRONIC TYPE B VIRAL HEPATITIS|OCCULT CHRONIC TYPE B VIRAL HEPATITIS (DISORDER)
C0375002|T047||SNOMEDCT_US|CHRONIC VIRAL HEPATITIS B WITH HEPATIC COMA WITHOUT HEPATITIS DELTA
C0375003|T047||SNOMEDCT_US|CHRONIC VIRAL HEPATITIS B WITH HEPATIC COMA WITH HEPATITIS DELTA
C0375007|T047||SNOMEDCT_US|CHRONIC VIRAL HEPATITIS B WITHOUT MENTION OF HEPATIC COMA WITH HEPATITIS DELTA
C0276612|T047|50167007|SNOMEDCT_US|CHRONIC ACTIVE TYPE HEPATITIS B VIRUS |CHRONIC ACTIVE TYPE B VIRAL HEPATITIS (DISORDER)
C0276612|T047|50167007|SNOMEDCT_US|CHRONIC ACTIVE TYPE HEPATITIS B VIRUS|CHRONIC ACTIVE TYPE B VIRAL HEPATITIS (DISORDER)
C0276612|T047|50167007|SNOMEDCT_US|HEPATITIS B VIRUS - CHRONIC ACTIVE|CHRONIC ACTIVE TYPE B VIRAL HEPATITIS (DISORDER)
C0276612|T047|50167007|SNOMEDCT_US|CHRONIC ACTIVE TYPE B VIRAL HEPATITIS|CHRONIC ACTIVE TYPE B VIRAL HEPATITIS (DISORDER)
C0276612|T047|50167007|SNOMEDCT_US|CHRONIC ACTIVE TYPE B VIRAL HEPATITIS |CHRONIC ACTIVE TYPE B VIRAL HEPATITIS (DISORDER)
C0276613|T047|38662009|SNOMEDCT_US|CHRONIC PERSISTENT TYPE B VIRAL HEPATITIS |CHRONIC PERSISTENT TYPE B VIRAL HEPATITIS (DISORDER)
C0276613|T047|38662009|SNOMEDCT_US|CHRONIC PERSISTENT TYPE B VIRAL HEPATITIS|CHRONIC PERSISTENT TYPE B VIRAL HEPATITIS (DISORDER)
C0276613|T047|38662009|SNOMEDCT_US|HEPATITIS B VIRUS - CHRONIC PERSISTENT|CHRONIC PERSISTENT TYPE B VIRAL HEPATITIS (DISORDER)
C0276613|T047|38662009|SNOMEDCT_US|CHRONIC IMMUNE TOLERANT HEPATITIS B|CHRONIC PERSISTENT TYPE B VIRAL HEPATITIS (DISORDER)
C0276613|T047|38662009|SNOMEDCT_US|CHRONIC PERSISTENT TYPE B VIRAL HEPATITIS |CHRONIC PERSISTENT TYPE B VIRAL HEPATITIS (DISORDER)
C0276614|T047|1116000|SNOMEDCT_US|CHRONIC AGGRESSIVE TYPE B VIRAL HEPATITIS |CHRONIC AGGRESSIVE TYPE B VIRAL HEPATITIS (DISORDER)
C0276614|T047|1116000|SNOMEDCT_US|CHRONIC AGGRESSIVE TYPE B VIRAL HEPATITIS|CHRONIC AGGRESSIVE TYPE B VIRAL HEPATITIS (DISORDER)
C0276614|T047|1116000|SNOMEDCT_US|HEPATITIS B VIRUS - CHRONIC AGGRESSIVE TYPE|CHRONIC AGGRESSIVE TYPE B VIRAL HEPATITIS (DISORDER)
C0276614|T047|1116000|SNOMEDCT_US|CHRONIC AGGRESSIVE TYPE B VIRAL HEPATITIS |CHRONIC AGGRESSIVE TYPE B VIRAL HEPATITIS (DISORDER)
C0276610|T047|186639003|SNOMEDCT_US|CHRONIC VIRAL HEPATITIS B WITHOUT DELTA-AGENT|CHRONIC VIRAL HEPATITIS B WITHOUT DELTA-AGENT (DISORDER)
C0276610|T047|186639003|SNOMEDCT_US|CHRONIC VIRAL HEPATITIS B WITHOUT DELTA-AGENT |CHRONIC VIRAL HEPATITIS B WITHOUT DELTA-AGENT (DISORDER)
C0524909|T047|61977001|SNOMEDCT_US|HEPATITIS B, CHRONIC|CHRONIC TYPE B VIRAL HEPATITIS (DISORDER)
C0524909|T047|61977001|SNOMEDCT_US|CHRONIC VIRAL HEPATITIS B INFECTION|CHRONIC TYPE B VIRAL HEPATITIS (DISORDER)
C0524909|T047|61977001|SNOMEDCT_US|CHRONIC HEPATITIS B INFECTION |CHRONIC TYPE B VIRAL HEPATITIS (DISORDER)
C0524909|T047|61977001|SNOMEDCT_US|CHRONIC HEPATITIS B INFECTION|CHRONIC TYPE B VIRAL HEPATITIS (DISORDER)
C0524909|T047|61977001|SNOMEDCT_US|CHRONIC HEPATITIS, B VIRUS|CHRONIC TYPE B VIRAL HEPATITIS (DISORDER)
C0524909|T047|61977001|SNOMEDCT_US|CHRONIC (VIRAL) HEPATITIS B|CHRONIC TYPE B VIRAL HEPATITIS (DISORDER)
C0524909|T047|61977001|SNOMEDCT_US|CHRONIC HEPATITIS B|CHRONIC TYPE B VIRAL HEPATITIS (DISORDER)
C0524909|T047|61977001|SNOMEDCT_US|HEPATITIS B, CHRONIC [DISEASE/FINDING]|CHRONIC TYPE B VIRAL HEPATITIS (DISORDER)
C0524909|T047|61977001|SNOMEDCT_US|CHRONIC TYPE B VIRAL HEPATITIS|CHRONIC TYPE B VIRAL HEPATITIS (DISORDER)
C0524909|T047|61977001|SNOMEDCT_US|CHRONIC VIRAL HEPATITIS B|CHRONIC TYPE B VIRAL HEPATITIS (DISORDER)
C0524909|T047|61977001|SNOMEDCT_US|CHRONIC TYPE B VIRAL HEPATITIS |CHRONIC TYPE B VIRAL HEPATITIS (DISORDER)
C0524909|T047|61977001|SNOMEDCT_US|HEPATITIS; VIRUS, CHRONIC, TYPE B|CHRONIC TYPE B VIRAL HEPATITIS (DISORDER)
C0400918|T047|235869004|SNOMEDCT_US|CHRONIC VIRAL HEPATITIS B WITH DELTA-AGENT|CHRONIC VIRAL HEPATITIS B WITH HEPATITIS D (DISORDER)
C0400918|T047|235869004|SNOMEDCT_US|CHRONIC VIRAL HEPATITIS B INFECTION WITH HEPATITIS DELTA|CHRONIC VIRAL HEPATITIS B WITH HEPATITIS D (DISORDER)
C0400918|T047|235869004|SNOMEDCT_US|CHRONIC HEPATITIS B INFECTION WITH HEPATITIS DELTA|CHRONIC VIRAL HEPATITIS B WITH HEPATITIS D (DISORDER)
C0400918|T047|235869004|SNOMEDCT_US|CHRONIC HEPATITIS, B VIRUS WITH HEPATITIS DELTA|CHRONIC VIRAL HEPATITIS B WITH HEPATITIS D (DISORDER)
C0400918|T047|235869004|SNOMEDCT_US|CHRONIC HEPATITIS B INFECTION WITH HEPATITIS DELTA |CHRONIC VIRAL HEPATITIS B WITH HEPATITIS D (DISORDER)
C0400918|T047|235869004|SNOMEDCT_US|CHRONIC VIRAL HEPATITIS B WITH HEPATITIS D|CHRONIC VIRAL HEPATITIS B WITH HEPATITIS D (DISORDER)
C0400918|T047|235869004|SNOMEDCT_US|CHRONIC VIRAL HEPATITIS B WITH HEPATITIS D |CHRONIC VIRAL HEPATITIS B WITH HEPATITIS D (DISORDER)
C0400918|T047|235869004|SNOMEDCT_US|HEPATITIS; VIRUS, CHRONIC, TYPE B, WITH DELTA-AGENT|CHRONIC VIRAL HEPATITIS B WITH HEPATITIS D (DISORDER)
C2074978|T047||SNOMEDCT_US|CHRONIC HEPATITIS, B VIRUS WITH HEPATIC COMA
C2074978|T047||SNOMEDCT_US|CHRONIC VIRAL HEPATITIS B INFECTION WITH HEPATIC COMA
C2074978|T047||SNOMEDCT_US|CHRONIC HEPATITIS B INFECTION WITH HEPATIC COMA
C2074978|T047||SNOMEDCT_US|CHRONIC HEPATITIS B INFECTION WITH HEPATIC COMA 
C2074976|T047||SNOMEDCT_US|CHRONIC HEPATITIS B INFECTION WITH COMA WITH HEPATITIS DELTA 
C2074976|T047||SNOMEDCT_US|CHRONIC HEPATITIS B INFECTION WITH COMA WITH HEPATITIS DELTA
C2074976|T047||SNOMEDCT_US|CHRONIC HEPATITIS, B VIRUS COMA WITH HEPATITIS DELTA
C2074976|T047||SNOMEDCT_US|CHRONIC VIRAL HEPATITIS B INFECTION WITH COMA WITH HEPATITIS DELTA
C2074977|T047||SNOMEDCT_US|CHRONIC VIRAL HEPATITIS B INFECTION WITH FULMINANT HEPATIC FAILURE
C2074977|T047||SNOMEDCT_US|CHRONIC HEPATITIS B INFECTION WITH FULMINANT HEPATIC FAILURE 
C2074977|T047||SNOMEDCT_US|CHRONIC HEPATITIS B INFECTION WITH FULMINANT HEPATIC FAILURE
C2074977|T047||SNOMEDCT_US|CHRONIC HEPATITIS, B VIRUS WITH FULMINANT HEPATIC FAILURE
C3838179|T047||SNOMEDCT_US|HEPATITIS, B VIRUS - CHRONIC WITHOUT HEPATITIS DELTA
C3838179|T047||SNOMEDCT_US|CHRONIC HEPATITIS, B VIRUS WITHOUT HEPATITIS DELTA 
C3838179|T047||SNOMEDCT_US|CHRONIC HEPATITIS, B VIRUS WITHOUT HEPATITIS DELTA
C4075603|T047|713966008|SNOMEDCT_US|OCCULT CHRONIC TYPE B VIRAL HEPATITIS |OCCULT CHRONIC TYPE B VIRAL HEPATITIS (DISORDER)
C4075603|T047|713966008|SNOMEDCT_US|OCCULT CHRONIC TYPE B VIRAL HEPATITIS|OCCULT CHRONIC TYPE B VIRAL HEPATITIS (DISORDER)
C4075603|T047|713966008|SNOMEDCT_US|OCCULT HEPATITIS B INFECTION|OCCULT CHRONIC TYPE B VIRAL HEPATITIS (DISORDER)
C1827079|T047|424340000|SNOMEDCT_US|CHRONIC VIRAL HEPATITIS B WITH HEPATIC COMA|CHRONIC HEPATITIS B WITH HEPATIC COMA
C1827079|T047|424340000|SNOMEDCT_US|HEPATIC COMA DUE TO CHRONIC HEPATITIS B |CHRONIC HEPATITIS B WITH HEPATIC COMA
C1827079|T047|424340000|SNOMEDCT_US|CHRONIC HEPATITIS B WITH HEPATIC COMA|CHRONIC HEPATITIS B WITH HEPATIC COMA
C1827079|T047|424340000|SNOMEDCT_US|HEPATIC COMA DUE TO CHRONIC HEPATITIS B|CHRONIC HEPATITIS B WITH HEPATIC COMA
C1827079|T047|424340000|SNOMEDCT_US|CHRONIC HEPATITIS B WITH HEPATIC COMA |CHRONIC HEPATITIS B WITH HEPATIC COMA
C0494789|T047||SNOMEDCT_US|CHRONIC ACTIVE HEPATITIS, NOT ELSEWHERE CLASSIFIED
C0494787|T047||SNOMEDCT_US|CHRONIC PERSISTENT HEPATITIS, NOT ELSEWHERE CLASSIFIED
C4041189|T047|153091000119109|SNOMEDCT_US|HEPATIC COMA DUE TO CHRONIC HEPATITIS B WITH DELTA AGENT |HEPATIC COMA DUE TO CHRONIC HEPATITIS B WITH DELTA AGENT (DISORDER)
C4041189|T047|153091000119109|SNOMEDCT_US|HEPATIC COMA DUE TO CHRONIC HEPATITIS B WITH DELTA AGENT|HEPATIC COMA DUE TO CHRONIC HEPATITIS B WITH DELTA AGENT (DISORDER)
C2074981|T047||SNOMEDCT_US|CHRONIC HEPATITIS D INFECTION WITH CHRONIC HEPATITIS B 
C2074981|T047||SNOMEDCT_US|CHRONIC HEPATITIS, DELTA VIRUS WITH CHRONIC HEPATITIS B
C2074981|T047||SNOMEDCT_US|CHRONIC HEPATITIS D INFECTION WITH CHRONIC HEPATITIS B
C2074983|T047||SNOMEDCT_US|CHRONIC HEPATITIS D INFECTION WITH HEPATITIS B CARRIER STATE 
C2074983|T047||SNOMEDCT_US|CHRONIC HEPATITIS, DELTA VIRUS WITH CARRIER STATE HEPATITIS B
C2074983|T047||SNOMEDCT_US|CHRONIC HEPATITIS D INFECTION WITH HEPATITIS B CARRIER STATE
C0375002|T047||SNOMEDCT_US|HPT B CHRN COMA WO DLTA
C0375002|T047||SNOMEDCT_US|CHRONIC VIRAL HEPATITIS B WITH HEPATIC COMA WITHOUT HEPATITIS DELTA
C0375002|T047||SNOMEDCT_US|VIRAL HEPATITIS B WITH HEPATIC COMA, CHRONIC, WITHOUT MENTION OF HEPATITIS DELTA
C0375003|T047||SNOMEDCT_US|HPT B CHRN COMA W DLTA
C0375003|T047||SNOMEDCT_US|CHRONIC VIRAL HEPATITIS B WITH HEPATIC COMA WITH HEPATITIS DELTA
C0375007|T047||SNOMEDCT_US|HPT B CHRN WO CM W DLTA
C0375007|T047||SNOMEDCT_US|CHRONIC VIRAL HEPATITIS B WITHOUT MENTION OF HEPATIC COMA WITH HEPATITIS DELTA
