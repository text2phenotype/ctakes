C2229883|T034||LNC|TIBC
C2229883|T034||LNC|SERUM TOTAL IRON BINDING CAPACITY (TIBC)
C0036835|T034|LP32077-7|LNC|SERUM TOTAL IRON-BINDING CAPACITY RESULT|IRON BINDING CAPACITY.TOTAL
C0036835|T034|LP32077-7|LNC|TIBC|IRON BINDING CAPACITY.TOTAL
C0036835|T034|LP32077-7|LNC|SERUM TOTAL IRON-BINDING CAPACITY RESULT|IRON BINDING CAPACITY.TOTAL
