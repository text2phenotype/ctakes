C0364639|T034|2498-4|LNC|IRON[MASS/VOLUME] IN SERUM OR PLASMA|IRON SERPL-MCNC
C0428578|T034||LNC|IRON LEVEL RESULT
C0364639|T034|2498-4|LNC|IRON [MASS/VOLUME] IN SERUM OR PLASMA|IRON SERPL-MCNC
C0364639|T034|2498-4|LNC|IRON SERPL-MCNC|IRON SERPL-MCNC
C0364639|T034|2498-4|LNC|IRON:MCNC:PT:SER/PLAS:QN|IRON SERPL-MCNC
C0364639|T034|2498-4|LNC|IRON:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|IRON SERPL-MCNC
C0853169|T034||LNC|BLOOD IRON MEASUREMENT
C0853169|T034||LNC|BLOOD IRON
C1318312|T034||LNC|SERUM IRON
C1318312|T034||LNC|SERUM IRON MEASUREMENT 
C1318312|T034||LNC|SERUM IRON LEVEL
C1318312|T034||LNC|(SERUM IRON TESTS) OR (SERUM IRON LEVEL) 
C1318312|T034||LNC|(SERUM IRON TESTS) OR (SERUM IRON LEVEL)
C1318312|T034||LNC|SERUM IRON: [TESTS] OR [LEVEL] 
C1318312|T034||LNC|SERUM IRON: [TESTS] OR [LEVEL]
C1277709|T034|MTHU023012|LNC|IRON SATURATION|TRANSFERRIN SATURATION
C1272108|T034||LNC|PLASMA IRON LEVEL
C0302583|T034||LNC|IRON|IRON
