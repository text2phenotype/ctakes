C0033707|T034||LNC|PROTIME
C0033707|T034||LNC|PROTHROMBIN TIME
C0033707|T034||LNC|PROTHROMBIN TIME ASSAY
C0151872|T034||LNC|PROTHROMBIN TIME INCREASED
C0482694|T034|5902-2|LNC|COAGULATION TISSUE FACTOR INDUCED:TIME:PT:PPP:QN:COAG|COAGULATION TISSUE FACTOR INDUCED:TIME:POINT IN TIME:PLATELET POOR PLASMA:QUANTITATIVE:COAGULATION ASSAY
C0482694|T034|5902-2|LNC|COAGULATION TISSUE FACTOR INDUCED|COAGULATION TISSUE FACTOR INDUCED:TIME:POINT IN TIME:PLATELET POOR PLASMA:QUANTITATIVE:COAGULATION ASSAY
C0482694|T034|5902-2|LNC|COAGULATION TIME|COAGULATION TISSUE FACTOR INDUCED:TIME:POINT IN TIME:PLATELET POOR PLASMA:QUANTITATIVE:COAGULATION ASSAY
C0482694|T034|5902-2|LNC|LOINC 5902-2|COAGULATION TISSUE FACTOR INDUCED:TIME:POINT IN TIME:PLATELET POOR PLASMA:QUANTITATIVE:COAGULATION ASSAY
C0482694|T034|5902-2|LNC|LNC 5902-2|COAGULATION TISSUE FACTOR INDUCED:TIME:POINT IN TIME:PLATELET POOR PLASMA:QUANTITATIVE:COAGULATION ASSAY
C0482694|T034|5902-2|LNC|5902-2|COAGULATION TISSUE FACTOR INDUCED:TIME:POINT IN TIME:PLATELET POOR PLASMA:QUANTITATIVE:COAGULATION ASSAY
C0482694|T034|5902-2|LNC|PROTHROMBIN TIME|COAGULATION TISSUE FACTOR INDUCED:TIME:POINT IN TIME:PLATELET POOR PLASMA:QUANTITATIVE:COAGULATION ASSAY
C0236453|T034||LNC|PLASMA PATIENT PROTHROMBIN TEST
C0033707|T034||LNC|PROTHROMBIN TIME
C0033707|T034||LNC|PROTHROMBIN TIMES
C0033707|T034||LNC|TIME, PROTHROMBIN
C0033707|T034||LNC|TIMES, PROTHROMBIN
C0033707|T034||LNC|PROTHROMBIN TIME (PT)
# C0033707|T034||LNC|PT
C0033707|T034||LNC|PROTHROMBIN TIME TEST
C0033707|T034||LNC|PROTHROMBIN TIME (PT) 
C0033707|T034||LNC|TEST;PROTHROMBIN TIME
C0033707|T034||LNC|PROTHROMBIN TIME ASSAY
C0033707|T034||LNC|PT ASSAY
C0033707|T034||LNC|PROTIME
C0033707|T034||LNC|PTT - PROTHROMBIN TIME
C0033707|T034||LNC|QUICK ONE STAGE PROTHROMBIN TIME
C0033707|T034||LNC|PT - PROTHROMBIN TIME
C0033707|T034||LNC|PROTHROMBIN TIME 
C0033707|T034||LNC|ONE STAGE PROTHROMBIN TIME
C0033707|T034||LNC|ONE STAGE PROTHROMBIN TIME 
C0033707|T034||LNC|PRO-THROMBIN TIME
C0033707|T034||LNC|PROTHROMBIN TEST
C0033707|T034||LNC|PLASMA PROTHROMBIN TEST
C1271785|T034||LNC|PROTHROMBIN TIME - REFERENCE
C1271785|T034||LNC|PROTHROMBIN TIME - REFERENCE 
C0373814|T034||LNC|PROTHROMBIN TIME; SUBSTITUTION, PLASMA FRACTIONS, EACH
C0373814|T034||LNC|PROTHROMBIN TIME ASSAY; SUBSTITUTION, PLASMA FRACTIONS, EACH
C0373814|T034||LNC|PROTHROMBIN TIME SUBSTITUTION PLASMA FRCTJ EACH
C0373814|T034||LNC|PROTHROMBIN TEST
C4027891|T034||LNC|PROTHROMBIN TIME IN PLATELET-POOR PLASMA BY COAGULATION ASSAY
C4027891|T034||LNC|PROTHROMBIN TIME (PT) IN PLATELET-POOR PLASMA BY COAGULATION ASSAY
C4027891|T034||LNC|PROTHROMBIN TIME IN PLATELET-POOR PLASMA BY COAGULATION ASSAY 
C4027892|T034||LNC|PROTHROMBIN TIME (PT) IN CAPILLARY BLOOD 
C4027892|T034||LNC|PROTHROMBIN TIME (PT) IN CAPILLARY BLOOD
C0151872|T034||LNC|PROLONGED PROTHROMBIN TIME
C0151872|T034||LNC|PROTHROMBIN TIME INC
C0151872|T034||LNC|PT INC
C0151872|T034||LNC|PROTHROMBIN LEVEL INCREASED
C0151872|T034||LNC|PROTHROMBIN TIME PROLONGED
C0151872|T034||LNC|PT PROLONGED
C0151872|T034||LNC|PROTHROMBIN TIME INCREASED
C0151872|T034||LNC|COAGULATION FACTOR II LEVEL INCREASED
C0151872|T034||LNC|PROTHROMBIN INCREASED
C0151872|T034||LNC|PT INCREASED
C0151872|T034||LNC|PROLONGED; PROTHROMBIN TIME
C0151872|T034||LNC|PROTHROMBIN TIME; PROLONGED
C0151872|T034||LNC|PROTHROMBIN TIME INCREASED 
C0151872|T034||LNC|ABNORMAL OR PROLONGED PROTHROMBIN TIME
C0151872|T034||LNC|ABNORMAL OR PROLONGED PT
C3670570|T034||LNC|OSPT INCREASED
C3670570|T034||LNC|ONE STAGE PROTHROMBIN TIME INCREASED
C3670570|T034||LNC|ONE STAGE PROTHROMBIN TIME INCREASED 
C3670543|T034||LNC|THROMBOTEST PROLONGED
C3670543|T034||LNC|PIVKA TEST PROLONGED
C3670543|T034||LNC|THROMBOTEST PROLONGED 
C0482694|T034|5902-2|LNC|COAGULATION TISSUE FACTOR INDUCED:TIME:PT:PPP:QN:COAG|COAGULATION TISSUE FACTOR INDUCED:TIME:POINT IN TIME:PLATELET POOR PLASMA:QUANTITATIVE:COAGULATION ASSAY
C0482694|T034|5902-2|LNC|COAGULATION TISSUE FACTOR INDUCED:TIME:POINT IN TIME:PLATELET POOR PLASMA:QUANTITATIVE:COAGULATION ASSAY|COAGULATION TISSUE FACTOR INDUCED:TIME:POINT IN TIME:PLATELET POOR PLASMA:QUANTITATIVE:COAGULATION ASSAY
C0482694|T034|5902-2|LNC|PROTHROMBIN TIME|COAGULATION TISSUE FACTOR INDUCED:TIME:POINT IN TIME:PLATELET POOR PLASMA:QUANTITATIVE:COAGULATION ASSAY
C0482694|T034|5902-2|LNC|PROTHROMBIN TIME (PT)|COAGULATION TISSUE FACTOR INDUCED:TIME:POINT IN TIME:PLATELET POOR PLASMA:QUANTITATIVE:COAGULATION ASSAY
