C0019151|T047|123049003|SNOMEDCT_US|HEPATIC ENCEPHALOPATHY|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C3266165|T047|449901005|SNOMEDCT_US|HEPATIC ENCEPHALOPATHY IN FULMINANT HEPATIC FAILURE|HEPATIC ENCEPHALOPATHY IN FULMINANT HEPATIC FAILURE (DISORDER)
C2729507|T047||SNOMEDCT_US|HEPATIC ENCEPHALOPATHY WITH COMA
C3888788|T047||SNOMEDCT_US|MINIMAL HEPATIC ENCEPHALOPATHY
C4024937|T047||SNOMEDCT_US|CHRONIC HEPATIC ENCEPHALOPATHY
C3889995|T047||SNOMEDCT_US|CDISC SDTM WEST HAVEN HEPATIC ENCEPHALOPATHY GRADE TERMINOLOGY
C3890564|T047||SNOMEDCT_US|WEST HAVEN HEPATIC ENCEPHALOPATHY GRADE
C4086961|T047||SNOMEDCT_US|WEST HAVEN CRITERIA - WEST HAVEN HEPATIC ENCEPHALOPATHY GRADE
C3151062|T047||SNOMEDCT_US|INFECTIONS, RECURRENT, WITH ENCEPHALOPATHY, HEPATIC DYSFUNCTION, AND CARDIOVASCULAR MALFORMATIONS
C3889290|T047||SNOMEDCT_US|WEST HAVEN HEPATIC ENCEPHALOPATHY GRADE 3
C3889292|T047||SNOMEDCT_US|WEST HAVEN HEPATIC ENCEPHALOPATHY GRADE 1
C3889293|T047||SNOMEDCT_US|WEST HAVEN HEPATIC ENCEPHALOPATHY GRADE 4
C3889824|T047||SNOMEDCT_US|WEST HAVEN HEPATIC ENCEPHALOPATHY GRADE 2
C3890401|T047||SNOMEDCT_US|WEST HAVEN HEPATIC ENCEPHALOPATHY GRADE 0
C4016797|T047||SNOMEDCT_US|INFECTIONS, RECURRENT, ASSOCIATED WITH ENCEPHALOPATHY, HEPATIC DYSFUNCTION, AND CARDIOVASCULAR MALFORMATIONS
C4086072|T047||SNOMEDCT_US|CDISC CLINICAL CLASSIFICATION WEST HAVEN CRITERIA TEST CODE TERMINOLOGY
C4086073|T047||SNOMEDCT_US|CDISC CLINICAL CLASSIFICATION WEST HAVEN CRITERIA TEST NAME TERMINOLOGY
C0019151|T047|123049003|SNOMEDCT_US|ENCEPHALOPATHIES, HEPATIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|ENCEPHALOPATHIES, PORTOSYSTEMIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|HEPATIC ENCEPHALOPATHIES|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|HEPATIC ENCEPHALOPATHY|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|PORTOSYSTEMIC ENCEPHALOPATHIES|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|ENCEPH HEPATOCEREBRAL|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|ENCEPH PORTAL SYSTEMIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|HEPATIC ENCEPH|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|PORTOSYSTEMIC ENCEPH|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|ENCEPH PORTOSYSTEMIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|PORTAL SYSTEMIC ENCEPH|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|HEPATOCEREBRAL ENCEPH|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|ENCEPH HEPATIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|HEPATIC ENCEPHALOPATHY |HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|HEPATOCEREBRAL ENCEPHALOPATHY -RETIRED-|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|ENCEPHALOPATHIES, HEPATOCEREBRAL|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|HEPATOCEREBRAL ENCEPHALOPATHIES|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|ENCEPHALOPATHIES, PORTAL-SYSTEMIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|PORTAL SYSTEMIC ENCEPHALOPATHY|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|PORTAL-SYSTEMIC ENCEPHALOPATHIES|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|HEPATIC ENCEPHALOPATHY NOS|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|PORTOSYSTEMIC ENCEPHALOPATHY|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|ENCEPHALOPATHY, HEPATOCEREBRAL|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|HEPATOCEREBRAL ENCEPHALOPATHY|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|HEPATIC ENCEPHALOPATHY [DISEASE/FINDING]|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|PORTAL-SYSTEMIC ENCEPHALOPATHY|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|ENCEPHALOPATHY, HEPATIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|ENCEPHALOPATHY, PORTAL-SYSTEMIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|ENCEPHALOPATHY, PORTOSYSTEMIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|HEPATIC COMA/ENCEPHALOPATHY|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|ENCEPHALOPATHY, PORTAL SYSTEMIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|GAUSTAD'S SYNDROME|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|PORTAL SYSTEMIC ENCEPHALOPATHY |HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|TRANSIENT HEPATARGY SYNDROME|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|ENCEPHALOPATHY - HEPATIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|HEPATOCEREBRAL ENCEPHALOPATHY |HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|ENCEPHALOPATHY HEPATIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|HE - HEPATIC ENCEPHALOPATHY|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|HEPATIC ENCEPHALOPATHY |HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|ENCEPHALOPATHY; HEPATIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|ENCEPHALOPATHY; PORTOSYSTEMIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|HEPATIC; ENCEPHALOPATHY|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T047|123049003|SNOMEDCT_US|PORTOSYSTEMIC; ENCEPHALOPATHY|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C2729507|T047||SNOMEDCT_US|HEPATIC ENCEPHALOPATHY WITH COMA 
C2729507|T047||SNOMEDCT_US|HEPATIC ENCEPHALOPATHY WITH COMA
C0019147|T047|72836002|SNOMEDCT_US|COMAS, HEPATIC|HEPATIC COMA (DISORDER)
C0019147|T047|72836002|SNOMEDCT_US|HEPATIC COMAS|HEPATIC COMA (DISORDER)
C0019147|T047|72836002|SNOMEDCT_US|COMA, HEPATIC|HEPATIC COMA (DISORDER)
C0019147|T047|72836002|SNOMEDCT_US|HEPATIC COMA|HEPATIC COMA (DISORDER)
C0019147|T047|72836002|SNOMEDCT_US|COMA HEPATIC|HEPATIC COMA (DISORDER)
C0019147|T047|72836002|SNOMEDCT_US|HEPATIC COMA NOS|HEPATIC COMA (DISORDER)
C0019147|T047|72836002|SNOMEDCT_US|COMA;HEPATIC|HEPATIC COMA (DISORDER)
C0019147|T047|72836002|SNOMEDCT_US|HEPATIC COMA |HEPATIC COMA (DISORDER)
C0019147|T047|72836002|SNOMEDCT_US|HEPATOCEREBRAL INTOXICATION|HEPATIC COMA (DISORDER)
C0019147|T047|72836002|SNOMEDCT_US|COMA; HEPATIC|HEPATIC COMA (DISORDER)
C0019147|T047|72836002|SNOMEDCT_US|HEPATIC; COMA|HEPATIC COMA (DISORDER)
C3266165|T047|449901005|SNOMEDCT_US|HEPATIC ENCEPHALOPATHY IN FULMINANT HEPATIC FAILURE|HEPATIC ENCEPHALOPATHY IN FULMINANT HEPATIC FAILURE (DISORDER)
C3266165|T047|449901005|SNOMEDCT_US|HEPATIC ENCEPHALOPATHY IN FULMINANT HEPATIC FAILURE |HEPATIC ENCEPHALOPATHY IN FULMINANT HEPATIC FAILURE (DISORDER)
C0751198|T047||SNOMEDCT_US|HEPATIC STUPORS
C0751198|T047||SNOMEDCT_US|STUPOR, HEPATIC
C0751198|T047||SNOMEDCT_US|STUPORS, HEPATIC
C0751198|T047||SNOMEDCT_US|HEPATIC STUPOR
C1836797|T047||SNOMEDCT_US|GENETIC DEFICIENCY, WOULD NOT BE RELATED TO CIRRHOSIS
C1836797|T047||SNOMEDCT_US|HEPATOENCEPHALOPATHY, EARLY FATAL PROGRESSIVE
C4024937|T047||SNOMEDCT_US|CHRONIC HEPATIC ENCEPHALOPATHY
C3888788|T047||SNOMEDCT_US|MINIMAL HEPATIC ENCEPHALOPATHY
C3889824|T047||SNOMEDCT_US|WEST HAVEN HEPATIC ENCEPHALOPATHY GRADE 2
C3890401|T047||SNOMEDCT_US|WEST HAVEN HEPATIC ENCEPHALOPATHY GRADE 0
C3889292|T047||SNOMEDCT_US|WEST HAVEN HEPATIC ENCEPHALOPATHY GRADE 1
C3889290|T047||SNOMEDCT_US|WEST HAVEN HEPATIC ENCEPHALOPATHY GRADE 3
C3889293|T047||SNOMEDCT_US|WEST HAVEN HEPATIC ENCEPHALOPATHY GRADE 4
