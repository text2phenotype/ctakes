C0005910|T034|6063|MEDCIN|BODY WEIGHT|WEIGHT (PHYSICAL FINDING)
C0944911|T034||MEDCIN|BODY WEIGHT:MASS:POINT IN TIME:^PATIENT:QUANTITATIVE
C0005910|T034|6063|MEDCIN|BODY WEIGHT|WEIGHT (PHYSICAL FINDING)
C0005910|T034|6063|MEDCIN|WEIGHT, BODY|WEIGHT (PHYSICAL FINDING)
C0005910|T034|6063|MEDCIN|WEIGHTS, BODY|WEIGHT (PHYSICAL FINDING)
C0005910|T034|6063|MEDCIN|WEIGHT|WEIGHT (PHYSICAL FINDING)
C0005910|T034|6063|MEDCIN|WEIGHT (PHYSICAL FINDING)|WEIGHT (PHYSICAL FINDING)
C0005910|T034|6063|MEDCIN|BODY WEIGHT [DISEASE/FINDING]|WEIGHT (PHYSICAL FINDING)
C0005910|T034|6063|MEDCIN|BODY WEIGHT - OBSERVATION|WEIGHT (PHYSICAL FINDING)
C0005910|T034|6063|MEDCIN|BODY WEIGHT (OBSERVABLE ENTITY)|WEIGHT (PHYSICAL FINDING)
C0005910|T034|6063|MEDCIN|BW|WEIGHT (PHYSICAL FINDING)
C0005910|T034|6063|MEDCIN|BODY WEIGHT, NOS|WEIGHT (PHYSICAL FINDING)
C0005910|T034|6063|MEDCIN|BODY WEIGHT [DUP] (OBSERVABLE ENTITY)|WEIGHT (PHYSICAL FINDING)
C0005910|T034|6063|MEDCIN|WEIGHT (BODY)|WEIGHT (PHYSICAL FINDING)
C2709005|T034||MEDCIN|DRY BODY WEIGHT
C2709005|T034||MEDCIN|DRY WEIGHT
C2709005|T034||MEDCIN|DRY BODY WEIGHT (OBSERVABLE ENTITY)
C1439839|T034|268429|MEDCIN|DRY WEIGHT (PHYSICAL FINDING)|DRY WEIGHT
C1439839|T034|268429|MEDCIN|DRY WEIGHT|DRY WEIGHT
C2266789|T034|293332|MEDCIN|WEIGHT RECORDED|WEIGHT WAS RECORDED
C2266789|T034|293332|MEDCIN|WEIGHT RECORDED (PHYSICAL FINDING)|WEIGHT WAS RECORDED
C1303013|T034||MEDCIN|BASELINE WEIGHT (OBSERVABLE ENTITY)
C1303013|T034||MEDCIN|BASELINE WEIGHT
C0424662|T034||MEDCIN|REFERENCE WEIGHT
C0424662|T034||MEDCIN|REFERENCE WEIGHT (OBSERVABLE ENTITY)
C3645728|T034|297539|MEDCIN|WEIGHT OBTAINED FROM PRIOR MEDICAL RECORD (___ LBS) (PHYSICAL FINDING)|WEIGHT OBTAINED FROM PRIOR MEDICAL RECORD (___ LBS) (PHYSICAL FINDING)
C3645728|T034|297539|MEDCIN|WEIGHT OBTAINED FROM PRIOR MEDICAL RECORD (___ LBS)|WEIGHT OBTAINED FROM PRIOR MEDICAL RECORD (___ LBS) (PHYSICAL FINDING)
C3834630|T034|297812|MEDCIN|WEIGHT WITH CLOTHES (PHYSICAL FINDING)|WEIGHT WITH CLOTHES (PHYSICAL FINDING)
C3834630|T034|297812|MEDCIN|WEIGHT WITH CLOTHES|WEIGHT WITH CLOTHES (PHYSICAL FINDING)
C3834629|T034|297813|MEDCIN|WEIGHT WITHOUT CLOTHES (PHYSICAL FINDING)|WEIGHT WITHOUT CLOTHES (PHYSICAL FINDING)
C3834629|T034|297813|MEDCIN|WEIGHT WITHOUT CLOTHES|WEIGHT WITHOUT CLOTHES (PHYSICAL FINDING)
C3834631|T034|297862|MEDCIN|WEIGHT AT INITIAL ENCOUNTER ___|WEIGHT AT INITIAL ENCOUNTER ___ (PHYSICAL FINDING)
C3834631|T034|297862|MEDCIN|WEIGHT AT INITIAL ENCOUNTER ___ (PHYSICAL FINDING)|WEIGHT AT INITIAL ENCOUNTER ___ (PHYSICAL FINDING)
C4032003|T034|298347|MEDCIN|ANTEPARTUM WEIGHT (___LBS)|ANTEPARTUM WEIGHT (___LBS)
C4032003|T034|298347|MEDCIN|ANTEPARTUM WEIGHT|ANTEPARTUM WEIGHT (___LBS)
C4032003|T034|298347|MEDCIN|ANTEPARTUM WEIGHT (PHYSICAL FINDING)|ANTEPARTUM WEIGHT (___LBS)
C4027960|T034|298305|MEDCIN|WEIGHT POST-SURGERY (___ LBS)|POST-SURGERY WEIGHT (PHYSICAL FINDING)
C4027960|T034|298305|MEDCIN|POST-SURGERY WEIGHT (PHYSICAL FINDING)|POST-SURGERY WEIGHT (PHYSICAL FINDING)
C4027960|T034|298305|MEDCIN|POST-SURGERY WEIGHT|POST-SURGERY WEIGHT (PHYSICAL FINDING)
C4027367|T034|298300|MEDCIN|WEIGHT PRE-SURGERY (___ LBS)|WEIGHT PRE-SURGERY (___ LBS) (PHYSICAL FINDING)
C4027367|T034|298300|MEDCIN|WEIGHT PRE-SURGERY (___ LBS) (PHYSICAL FINDING)|WEIGHT PRE-SURGERY (___ LBS) (PHYSICAL FINDING)
C1827199|T034||MEDCIN|BODY WEIGHT WITHOUT SHOES
C1827199|T034||MEDCIN|BODY WEIGHT WITHOUT SHOES (OBSERVABLE ENTITY)
C1828456|T034||MEDCIN|BODY WEIGHT WITH SHOES (OBSERVABLE ENTITY)
C1828456|T034||MEDCIN|BODY WEIGHT WITH SHOES
C0944911|T034||MEDCIN|BODY WEIGHT:MASS:POINT IN TIME:^PATIENT:QUANTITATIVE
C0944911|T034||MEDCIN|BODY WEIGHT:MASS:PT:^PATIENT:QN
C0944911|T034||MEDCIN|WEIGHT
C0944911|T034||MEDCIN|BODY WEIGHT
