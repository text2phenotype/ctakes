C0001899|T034||LNC|ALANINE TRANSAMINASE
C0201836|T034||LNC|ALANINE AMINOTRANSFERASE MEASUREMENT
C2257651|T034||LNC|L-ALANINE:2-OXOGLUTARATE AMINOTRANSFERASE ACTIVITY
C0001899|T034||LNC|ALANINE 2 OXOGLUTARATE AMINOTRANSFERASE
C0001899|T034||LNC|ALANINE AMINOTRANSFERASE
C0001899|T034||LNC|AMINOTRANSFERASE, ALANINE
C0001899|T034||LNC|AMINOTRANSFERASE, ALANINE-2-OXOGLUTARATE
C0001899|T034||LNC|GLUTAMIC ALANINE TRANSAMINASE
C0001899|T034||LNC|GLUTAMIC PYRUVIC TRANSAMINASE
C0001899|T034||LNC|GLUTAMIC-PYRUVIC TRANSAMINASE
C0001899|T034||LNC|TRANSAMINASE, GLUTAMIC-ALANINE
C0001899|T034||LNC|TRANSAMINASE, GLUTAMIC-PYRUVIC
C0001899|T034||LNC|L-ALANINE:2-OXOGLUTARATE AMINOTRANSFERASE
C0001899|T034||LNC|ALANINE TRANSAMINASE
C0001899|T034||LNC|TRANSAMINASE, ALANINE
C0001899|T034||LNC|GLUTAMIC-ALANINE TRANSAMINASE
C0001899|T034||LNC|ALANINE TRANSAMINASE [CHEMICAL/INGREDIENT]
C0001899|T034||LNC|ALANINE-2-OXOGLUTARATE AMINOTRANSFERASE
C0001899|T034||LNC|GPT
C0001899|T034||LNC|ALAT - ALANINE AMINOTRANSFERASE
C0001899|T034||LNC|ALT - ALANINE AMINOTRANSFERASE
C0001899|T034||LNC|GLUTAMATE PYRUVATE TRANSAMINASE
C0001899|T034||LNC|ALANINE AMINOTRANSFERASE 
C1980933|T034|LP44699-4|LNC|ALANINE AMINOTRANSFERASE &#X7C; BLD-SER-PLAS|ALANINE AMINOTRANSFERASE &#X7C; BLD-SER-PLAS
C1980938|T034|LP62238-8|LNC|ALANINE AMINOTRANSFERASE.MACROMOLECULAR &#X7C; BLD-SER-PLAS|ALANINE AMINOTRANSFERASE.MACROMOLECULAR &#X7C; BLD-SER-PLAS
C0376147|T034||LNC|SGPT
C0376147|T034||LNC|SGPT - GLUTAMATE PYRUVATE TRANSAMINASE
C0376147|T034||LNC|ALT
C0376147|T034||LNC|SERUM GLUTAMATE PYRUVATE TRANSAMINASE
C0376147|T034||LNC|ALANINE TRANSFERASE
C0376147|T034||LNC|SGPT (ALT)
C3887708|T034||LNC|GLUTAMATE PYRUVATE TRANSAMINASE 1
C3887708|T034||LNC|GLUTAMIC--ALANINE TRANSAMINASE 1
C3887708|T034||LNC|GLUTAMIC-PYRUVATE TRANSAMINASE
C3887708|T034||LNC|GPT 1
C3887708|T034||LNC|GLUTAMIC--PYRUVIC TRANSAMINASE 1
C3887708|T034||LNC|ALANINE AMINOTRANSFERASE 1
C3887708|T034||LNC|EC 2.6.1.2
C3887708|T034||LNC|ALANINE AMINOTRANSFERASE 1, HUMAN
C3887708|T034||LNC|ALANINE AMINOTRANSFERASE
C3887708|T034||LNC|GLUTAMIC-ALANINE TRANSAMINASE
C3887708|T034||LNC|GLUTAMIC-PYRUVIC TRANSAMINASE
C3887708|T034||LNC|GPT
C3887708|T034||LNC|AAT1
C3887708|T034||LNC|GPT1
C3887708|T034||LNC|ALT1
C0201836|T034||LNC|ALANINE AMINOTRANSFERASE MEASUREMENT
C0201836|T034||LNC|ALANINE AMINOTRANSFERASE
C0201836|T034||LNC|ALT
C0201836|T034||LNC|TRANSFERASE; ALANINE AMINO (ALT) (SGPT)
C0201836|T034||LNC|TEST;ALANINE AMINOTRANSFERASE
C0201836|T034||LNC|TRANSFERASE ALANINE AMINO ALT SGPT
C0201836|T034||LNC|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T034||LNC|MEASUREMENT OF ALANINE AMINO TRANSFERASE
C0201836|T034||LNC|LIVER ENZYME (SGPT), LEVEL
C0201836|T034||LNC|ALANINE AMINO (ALT) (SGPT)
C0201836|T034||LNC|SGPT
C0201836|T034||LNC|GLUTAMIC-PYRUVATE TRANSAMINASE
C0201836|T034||LNC|GPT
C0201836|T034||LNC|GPT MEASUREMENT
C0201836|T034||LNC|GLUTAMIC PYRUVATE TRANSAMINASE MEASUREMENT
C0201836|T034||LNC|SGPT MEASUREMENT
C0201836|T034||LNC|ALT MEASUREMENT
C0201836|T034||LNC|ALANINE AMINOTRANSFERASE MEASUREMENT 
C0201836|T034||LNC|ALANINE AMINOTRANSFERASE TEST
C1883008|T034||LNC|SERUM ALANINE AMINOTRANSFERASE MEASUREMENT
C1883008|T034||LNC|SERUM SGPT MEASUREMENT
C1883008|T034||LNC|SERUM ALANINE TRANSAMINASE MEASUREMENT
C1883008|T034||LNC|SERUM ALANINE AMINOTRANSFERASE MEASUREMENT 
C1883008|T034||LNC|ALT (SGPT) LEVEL
C0428324|T034||LNC|ALANINE TRANSAMINASE LEVEL
C0428324|T034||LNC|ALANINE TRANSAMINASE LEVEL 
C0428325|T034||LNC|ALT/SGPT SERUM LEVEL
C0428325|T034||LNC|ALT/SGPT SERUM LEVEL 
C0523461|T034||LNC|I BELIEVE THIS IS THE STANDARD METHOD BUT NOT 100%
C0523461|T034||LNC|ALANINE AMINOTRANSFERASE (ALT) MEASUREMENT, METHOD WITH PYRIDOXAL-5'-PHOSPHATE
C0523461|T034||LNC|ALANINE AMINOTRANSFERASE MEASUREMENT, METHOD WITH PYRIDOXAL-5'-PHOSPHATE 
C0523461|T034||LNC|ALANINE AMINOTRANSFERASE (ALT) MEASUREMENT, METHOD WITH PYRIDOXAL-5'-PHOSPHATE 
C0523461|T034||LNC|ALANINE AMINOTRANSFERASE MEASUREMENT, METHOD WITH PYRIDOXAL-5'-PHOSPHATE
C0523461|T034||LNC|ALT MEASUREMENT, METHOD WITH PYRIDOXAL-5'-PHOSPHATE
C0523462|T034||LNC|ALT MEASUREMENT, METHOD WITHOUT PYRIDOXAL-5'-PHOSPHATE 
C0523462|T034||LNC|ALANINE AMINOTRANSFERASE (ALT) MEASUREMENT, METHOD WITHOUT PYRIDOXAL-5'-PHOSPHATE
C0523462|T034||LNC|ALANINE AMINOTRANSFERASE MEASUREMENT, METHOD WITHOUT PYRIDOXAL-5'-PHOSPHATE 
C0523462|T034||LNC|ALANINE AMINOTRANSFERASE MEASUREMENT, METHOD WITHOUT PYRIDOXAL-5'-PHOSPHATE
C0523462|T034||LNC|ALANINE AMINOTRANSFERASE (ALT) MEASUREMENT, METHOD WITHOUT PYRIDOXAL-5'-PHOSPHATE 
C0523462|T034||LNC|ALT MEASUREMENT, METHOD WITHOUT PYRIDOXAL-5'-PHOSPHATE
C0428326|T034||LNC|SERUM GLUTAMIC OXALOACETIC TRANSAMINASE (SGPT) - BLOOD MEASUREMENT 
C0428326|T034||LNC|SERUM GLUTAMIC OXALOACETIC TRANSAMINASE (SGPT) - BLOOD MEASUREMENT
C0428326|T034||LNC|SGPT - BLOOD MEASUREMENT 
C0428326|T034||LNC|SGPT - BLOOD LEVEL
C0428326|T034||LNC|SGPT - BLOOD MEASUREMENT
C0428327|T034||LNC|ALT - BLOOD MEASUREMENT 
C0428327|T034||LNC|ALANINE AMINOTRANSFERASE (ALT) - BLOOD MEASUREMENT
C0428327|T034||LNC|LIVER ENZYMES (& BLOOD LEVEL [ALT] OR [SGPT])
C0428327|T034||LNC|LIVER ENZYMES (& BLOOD LEVEL [ALT] OR [SGPT]) 
C0428327|T034||LNC|SGPT - BLOOD LEVEL
C0428327|T034||LNC|ALT - BLOOD LEVEL
C0428327|T034||LNC|ALANINE AMINOTRANSFERASE - BLOOD MEASUREMENT
C0428327|T034||LNC|ALANINE AMINOTRANSFERASE (ALT) - BLOOD MEASUREMENT 
C0428327|T034||LNC|ALANINE AMINOTRANSFERASE - BLOOD MEASUREMENT 
C0428327|T034||LNC|ALT - BLOOD MEASUREMENT
C0428327|T034||LNC|ALT BLOOD MEASUREMENT