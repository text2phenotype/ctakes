#CUI|TUI|CODE|SAB|STR|PREF_TEXT|TS|STT|ISPREF
C0004886|T129|3055-2365|CSP|Bacillus Calmette Guerin vaccine||S|VCW|Y
C0004886|T121|3055-2365|CSP|Bacillus Calmette Guerin vaccine||S|VCW|Y
C0004886|T129|3055-2365|CSP|BCG vaccine||P|VC|Y
C0004886|T121|3055-2365|CSP|BCG vaccine||P|VC|Y
C0004886|T129|19|CVX|Bacillus Calmette-Guerin vaccine||S|VCW|Y
C0004886|T121|19|CVX|Bacillus Calmette-Guerin vaccine||S|VCW|Y
C0004886|T129|19|CVX|BCG||S|PF|N
C0004886|T121|19|CVX|BCG||S|PF|N
C0004886|T129|19|HL7V2.5|BCG||S|PF|N
C0004886|T121|19|HL7V2.5|BCG||S|PF|N
C0004886|T129|19|HL7V3.0|BCG||S|PF|N
C0004886|T121|19|HL7V3.0|BCG||S|PF|N
C0004886|T129|sh88000480|LCH_NW|BCG vaccines||P|VO|Y
C0004886|T121|sh88000480|LCH_NW|BCG vaccines||P|VO|Y
C0004886|T129|133312|MEDCIN|BCG vaccine, live, attenuated for tuberculosis (percutaneous use)||S|PF|Y
C0004886|T121|133312|MEDCIN|BCG vaccine, live, attenuated for tuberculosis (percutaneous use)||S|PF|Y
C0004886|T129|133312|MEDCIN|BCG vaccine, live, attenuated for tuberculosis (percutaneous use) (medication)||S|PF|Y
C0004886|T121|133312|MEDCIN|BCG vaccine, live, attenuated for tuberculosis (percutaneous use) (medication)||S|PF|Y
C0004886|T129|133312|MEDCIN|live attenuated BCG vaccine for tuberculosis (percutaneous use)||S|VW|Y
C0004886|T121|133312|MEDCIN|live attenuated BCG vaccine for tuberculosis (percutaneous use)||S|VW|Y
C0004886|T129|133313|MEDCIN|BCG vaccine, live, attenuated for bladder cancer (intravesical)||S|PF|Y
C0004886|T121|133313|MEDCIN|BCG vaccine, live, attenuated for bladder cancer (intravesical)||S|PF|Y
C0004886|T129|133313|MEDCIN|BCG vaccine, live, attenuated for bladder cancer (intravesical) (medication)||S|PF|Y
C0004886|T121|133313|MEDCIN|BCG vaccine, live, attenuated for bladder cancer (intravesical) (medication)||S|PF|Y
C0004886|T129|133313|MEDCIN|live attenuated BCG vaccine for bladder cancer (intravesical)||S|VW|Y
C0004886|T121|133313|MEDCIN|live attenuated BCG vaccine for bladder cancer (intravesical)||S|VW|Y
C0004886|T129|44458|MEDCIN|BCG vaccine, live, attenuated||S|PF|Y
C0004886|T121|44458|MEDCIN|BCG vaccine, live, attenuated||S|PF|Y
C0004886|T129|44458|MEDCIN|BCG vaccine, live, attenuated (medication)||S|PF|Y
C0004886|T121|44458|MEDCIN|BCG vaccine, live, attenuated (medication)||S|PF|Y
C0004886|T129|44458|MEDCIN|live attenuated BCG vaccine||S|VW|Y
C0004886|T121|44458|MEDCIN|live attenuated BCG vaccine||S|VW|Y
C0004886|T129|178022|MMSL|BCG Vaccine||P|PF|N
C0004886|T121|178022|MMSL|BCG Vaccine||P|PF|N
C0004886|T129|D001500|MSH|Bacillus Calmette Guerin Vaccine||S|VW|Y
C0004886|T121|D001500|MSH|Bacillus Calmette Guerin Vaccine||S|VW|Y
C0004886|T129|D001500|MSH|BCG Vaccine||P|PF|N
C0004886|T121|D001500|MSH|BCG Vaccine||P|PF|N
C0004886|T129|D001500|MSH|Calmette Guerin Bacillus Vaccine||S|PF|Y
C0004886|T121|D001500|MSH|Calmette Guerin Bacillus Vaccine||S|PF|Y
C0004886|T129|D001500|MSH|Calmette Vaccine||S|VO|Y
C0004886|T121|D001500|MSH|Calmette Vaccine||S|VO|Y
C0004886|T129|D001500|MSH|Calmette's Vaccine||S|PF|Y
C0004886|T121|D001500|MSH|Calmette's Vaccine||S|PF|Y
C0004886|T129|D001500|MSH|Calmettes Vaccine||S|VO|Y
C0004886|T121|D001500|MSH|Calmettes Vaccine||S|VO|Y
C0004886|T129|D001500|MSH|Vaccine, BCG||P|VW|Y
C0004886|T121|D001500|MSH|Vaccine, BCG||P|VW|Y
C0004886|T129|D001500|MSH|Vaccine, Calmette's||S|VW|Y
C0004886|T121|D001500|MSH|Vaccine, Calmette's||S|VW|Y
C0004886|T129|U001728|MTH|BCG Vaccine||P|PF|Y
C0004886|T121|U001728|MTH|BCG Vaccine||P|PF|Y
C0004886|T129|C298|NCI|Bacille Calmette-Guerin Live||S|PF|Y
C0004886|T121|C298|NCI|Bacille Calmette-Guerin Live||S|PF|Y
C0004886|T129|C298|NCI|Bacillius Calmette-Guerin Vaccine||S|PF|Y
C0004886|T121|C298|NCI|Bacillius Calmette-Guerin Vaccine||S|PF|Y
C0004886|T129|C298|NCI|Bacillus Calmette-Guerin||S|PF|Y
C0004886|T121|C298|NCI|Bacillus Calmette-Guerin||S|PF|Y
C0004886|T129|C298|NCI|BCG||S|PF|Y
C0004886|T121|C298|NCI|BCG||S|PF|Y
C0004886|T129|C298|NCI|BCG (Pasteur)||S|PF|Y
C0004886|T121|C298|NCI|BCG (Pasteur)||S|PF|Y
C0004886|T129|C298|NCI|BCG Vaccine||P|PF|N
C0004886|T121|C298|NCI|BCG Vaccine||P|PF|N
C0004886|T129|C298|NCI|Live Intravesical BCG||S|PF|Y
C0004886|T121|C298|NCI|Live Intravesical BCG||S|PF|Y
C0004886|T129|C298|NCI|Mycobacterium bovis (Strain BCG)||S|PF|Y
C0004886|T121|C298|NCI|Mycobacterium bovis (Strain BCG)||S|PF|Y
C0004886|T129|00495|NCI_DCP|Bacillus Calmette-Guerin||S|PF|N
C0004886|T121|00495|NCI_DCP|Bacillus Calmette-Guerin||S|PF|N
C0004886|T129|NSC0007817|NCI_DTP|Bacillus Calmette-Guerin||S|PF|N
C0004886|T121|NSC0007817|NCI_DTP|Bacillus Calmette-Guerin||S|PF|N
C0004886|T129|CDR0000044581|NCI_NCI-GLOSS|Bacillus Calmette Guerin||S|VO|Y
C0004886|T121|CDR0000044581|NCI_NCI-GLOSS|Bacillus Calmette Guerin||S|VO|Y
C0004886|T129|CDR0000045987|NCI_NCI-GLOSS|BCG||S|PF|N
C0004886|T121|CDR0000045987|NCI_NCI-GLOSS|BCG||S|PF|N
C0004886|T129|N0000010507|NDFRT|Bacillus Calmette Guerin Vaccine||S|VW|N
C0004886|T121|N0000010507|NDFRT|Bacillus Calmette Guerin Vaccine||S|VW|N
C0004886|T129|N0000010507|NDFRT|BCG Vaccine||P|PF|N
C0004886|T121|N0000010507|NDFRT|BCG Vaccine||P|PF|N
C0004886|T129|N0000010507|NDFRT|BCG Vaccine [Chemical/Ingredient]||S|PF|Y
C0004886|T121|N0000010507|NDFRT|BCG Vaccine [Chemical/Ingredient]||S|PF|Y
C0004886|T129|N0000010507|NDFRT|Calmette Guerin Bacillus Vaccine||S|PF|N
C0004886|T121|N0000010507|NDFRT|Calmette Guerin Bacillus Vaccine||S|PF|N
C0004886|T129|N0000010507|NDFRT|Calmette's Vaccine||S|PF|N
C0004886|T121|N0000010507|NDFRT|Calmette's Vaccine||S|PF|N
C0004886|T129|N0000147189|NDFRT|BACILLUS CALMETTE-GUERIN VACCINE||S|VCW|N
C0004886|T121|N0000147189|NDFRT|BACILLUS CALMETTE-GUERIN VACCINE||S|VCW|N
C0004886|T129|N0000147717|NDFRT|BCG VACCINE||P|VC|N
C0004886|T121|N0000147717|NDFRT|BCG VACCINE||P|VC|N
C0004886|T129|1344|RXNORM|BCG Vaccine||P|PF|N
C0004886|T121|1344|RXNORM|BCG Vaccine||P|PF|N
C0004886|T129|255701000|SNOMEDCT_US|BCG vaccine||P|VC|N
C0004886|T121|255701000|SNOMEDCT_US|BCG vaccine||P|VC|N
C0004886|T129|255701000|SNOMEDCT_US|BCG vaccine (substance)||S|PF|N
C0004886|T121|255701000|SNOMEDCT_US|BCG vaccine (substance)||S|PF|N
C0004886|T129|396419007|SNOMEDCT_US|Bacillus Calmette-Guérin vaccine||S|VO|Y
C0004886|T129|396419007|SNOMEDCT_US|Bacillus Calmette-Guerin vaccine||S|VCW|N
C0004886|T121|396419007|SNOMEDCT_US|Bacillus Calmette-Guérin vaccine||S|VO|Y
C0004886|T121|396419007|SNOMEDCT_US|Bacillus Calmette-Guerin vaccine||S|VCW|N
C0004886|T129|396419007|SNOMEDCT_US|BCG vaccine||P|VC|N
C0004886|T121|396419007|SNOMEDCT_US|BCG vaccine||P|VC|N
C0004886|T129|396419007|SNOMEDCT_US|BCG vaccine (substance)||S|PF|Y
C0004886|T121|396419007|SNOMEDCT_US|BCG vaccine (substance)||S|PF|Y
C0004886|T129|418268006|SNOMEDCT_US|Attenuated Bacillus Calmette Guerin||S|PF|Y
C0004886|T121|418268006|SNOMEDCT_US|Attenuated Bacillus Calmette Guerin||S|PF|Y
C0004886|T129|418268006|SNOMEDCT_US|Attenuated Bacillus Calmette Guerin (product)||S|PF|Y
C0004886|T121|418268006|SNOMEDCT_US|Attenuated Bacillus Calmette Guerin (product)||S|PF|Y
C0004886|T129|418571002|SNOMEDCT_US|Attenuated Bacillus Calmette Guerin||S|PF|N
C0004886|T121|418571002|SNOMEDCT_US|Attenuated Bacillus Calmette Guerin||S|PF|N
C0004886|T129|418571002|SNOMEDCT_US|Attenuated Bacillus Calmette Guerin (substance)||S|PF|Y
C0004886|T121|418571002|SNOMEDCT_US|Attenuated Bacillus Calmette Guerin (substance)||S|PF|Y
C0004886|T129|76685007|SNOMEDCT_US|Bacillus Calmette-Guérin vaccine||S|VO|N
C0004886|T129|76685007|SNOMEDCT_US|Bacillus Calmette-Guerin vaccine||S|VCW|N
C0004886|T121|76685007|SNOMEDCT_US|Bacillus Calmette-Guérin vaccine||S|VO|N
C0004886|T121|76685007|SNOMEDCT_US|Bacillus Calmette-Guerin vaccine||S|VCW|N
C0004886|T129|76685007|SNOMEDCT_US|BCG vaccine||P|VC|N
C0004886|T121|76685007|SNOMEDCT_US|BCG vaccine||P|VC|N
C0004886|T129|76685007|SNOMEDCT_US|BCG vaccine (product)||S|PF|Y
C0004886|T121|76685007|SNOMEDCT_US|BCG vaccine (product)||S|PF|Y
C0004886|T129|76685007|SNOMEDCT_US|BCG vaccine (substance)||S|PF|N
C0004886|T121|76685007|SNOMEDCT_US|BCG vaccine (substance)||S|PF|N
C0004886|T129|4018895|VANDF|BACILLUS CALMETTE-GUERIN VACCINE||S|VCW|Y
C0004886|T121|4018895|VANDF|BACILLUS CALMETTE-GUERIN VACCINE||S|VCW|Y
C0004886|T129|4019624|VANDF|BCG VACCINE||P|VC|Y
C0004886|T121|4019624|VANDF|BCG VACCINE||P|VC|Y
C0006044|T121|27|CVX|botulinum antitoxin||P|VC|N
C0006044|T121|27|CVX|botulinum antitoxin||P|VC|Y
C0006044|T129|27|CVX|botulinum antitoxin||P|VC|N
C0006044|T129|27|CVX|botulinum antitoxin||P|VC|Y
C0006044|T109|27|CVX|botulinum antitoxin||P|VC|N
C0006044|T109|27|CVX|botulinum antitoxin||P|VC|Y
C0006044|T121|27|HL7V2.5|botulinum antitoxin||P|VC|N
C0006044|T129|27|HL7V2.5|botulinum antitoxin||P|VC|N
C0006044|T109|27|HL7V2.5|botulinum antitoxin||P|VC|N
C0006044|T121|27|HL7V3.0|botulinum antitoxin||P|VC|N
C0006044|T129|27|HL7V3.0|botulinum antitoxin||P|VC|N
C0006044|T109|27|HL7V3.0|botulinum antitoxin||P|VC|N
C0006044|T121|40117|MEDCIN|botulism antitoxin||S|VC|N
C0006044|T129|40117|MEDCIN|botulism antitoxin||S|VC|N
C0006044|T109|40117|MEDCIN|botulism antitoxin||S|VC|N
C0006044|T121|40117|MEDCIN|botulism antitoxin (medication)||S|PF|Y
C0006044|T129|40117|MEDCIN|botulism antitoxin (medication)||S|PF|Y
C0006044|T109|40117|MEDCIN|botulism antitoxin (medication)||S|PF|Y
C0006044|T121|18704|MMSL|botulism antitoxin||S|VC|N
C0006044|T129|18704|MMSL|botulism antitoxin||S|VC|N
C0006044|T109|18704|MMSL|botulism antitoxin||S|VC|N
C0006044|T121|46487|MMSL|Botulism Antitoxin||S|PF|N
C0006044|T129|46487|MMSL|Botulism Antitoxin||S|PF|N
C0006044|T109|46487|MMSL|Botulism Antitoxin||S|PF|N
C0006044|T121|d04856|MMSL|botulism antitoxin||S|VC|Y
C0006044|T129|d04856|MMSL|botulism antitoxin||S|VC|Y
C0006044|T109|d04856|MMSL|botulism antitoxin||S|VC|Y
C0006044|T121|D001904|MSH|Antitoxin, Botulinum||P|VW|Y
C0006044|T129|D001904|MSH|Antitoxin, Botulinum||P|VW|Y
C0006044|T109|D001904|MSH|Antitoxin, Botulinum||P|VW|Y
C0006044|T121|D001904|MSH|Antitoxin, Botulism||S|VW|Y
C0006044|T129|D001904|MSH|Antitoxin, Botulism||S|VW|Y
C0006044|T109|D001904|MSH|Antitoxin, Botulism||S|VW|Y
C0006044|T121|D001904|MSH|Botulinum Antitoxin||P|PF|N
C0006044|T129|D001904|MSH|Botulinum Antitoxin||P|PF|N
C0006044|T109|D001904|MSH|Botulinum Antitoxin||P|PF|N
C0006044|T121|D001904|MSH|Botulism Antitoxin||S|PF|Y
C0006044|T129|D001904|MSH|Botulism Antitoxin||S|PF|Y
C0006044|T109|D001904|MSH|Botulism Antitoxin||S|PF|Y
C0006044|T121|NOCODE|MTH|Botulinum Antitoxin||P|PF|Y
C0006044|T129|NOCODE|MTH|Botulinum Antitoxin||P|PF|Y
C0006044|T109|NOCODE|MTH|Botulinum Antitoxin||P|PF|Y
C0006044|T121|N0000022498|NDFRT|BOTULISM ANTITOXIN||S|VC|N
C0006044|T129|N0000022498|NDFRT|BOTULISM ANTITOXIN||S|VC|N
C0006044|T109|N0000022498|NDFRT|BOTULISM ANTITOXIN||S|VC|N
C0006044|T121|N0000169329|NDFRT|Botulinum Antitoxin||P|PF|N
C0006044|T129|N0000169329|NDFRT|Botulinum Antitoxin||P|PF|N
C0006044|T109|N0000169329|NDFRT|Botulinum Antitoxin||P|PF|N
C0006044|T121|N0000169329|NDFRT|Botulinum Antitoxin [Chemical/Ingredient]||S|PF|Y
C0006044|T129|N0000169329|NDFRT|Botulinum Antitoxin [Chemical/Ingredient]||S|PF|Y
C0006044|T109|N0000169329|NDFRT|Botulinum Antitoxin [Chemical/Ingredient]||S|PF|Y
C0006044|T121|N0000169329|NDFRT|Botulism Antitoxin||S|PF|N
C0006044|T129|N0000169329|NDFRT|Botulism Antitoxin||S|PF|N
C0006044|T109|N0000169329|NDFRT|Botulism Antitoxin||S|PF|N
C0006044|T121|385336006|SNOMEDCT_US|Botulinum antitoxin||P|VC|Y
C0006044|T129|385336006|SNOMEDCT_US|Botulinum antitoxin||P|VC|Y
C0006044|T109|385336006|SNOMEDCT_US|Botulinum antitoxin||P|VC|Y
C0006044|T121|385336006|SNOMEDCT_US|Botulinum antitoxin (substance)||S|PF|Y
C0006044|T129|385336006|SNOMEDCT_US|Botulinum antitoxin (substance)||S|PF|Y
C0006044|T109|385336006|SNOMEDCT_US|Botulinum antitoxin (substance)||S|PF|Y
C0006044|T121|385336006|SNOMEDCT_US|Botulism antitoxin||S|VC|N
C0006044|T129|385336006|SNOMEDCT_US|Botulism antitoxin||S|VC|N
C0006044|T109|385336006|SNOMEDCT_US|Botulism antitoxin||S|VC|N
C0006044|T121|86080005|SNOMEDCT_US|Botulinum antitoxin||P|VC|N
C0006044|T129|86080005|SNOMEDCT_US|Botulinum antitoxin||P|VC|N
C0006044|T109|86080005|SNOMEDCT_US|Botulinum antitoxin||P|VC|N
C0006044|T121|86080005|SNOMEDCT_US|Botulism antitoxin||S|VC|Y
C0006044|T129|86080005|SNOMEDCT_US|Botulism antitoxin||S|VC|Y
C0006044|T109|86080005|SNOMEDCT_US|Botulism antitoxin||S|VC|Y
C0006044|T121|86080005|SNOMEDCT_US|Botulism antitoxin (product)||S|PF|Y
C0006044|T129|86080005|SNOMEDCT_US|Botulism antitoxin (product)||S|PF|Y
C0006044|T109|86080005|SNOMEDCT_US|Botulism antitoxin (product)||S|PF|Y
C0006044|T121|86080005|SNOMEDCT_US|Botulism antitoxin (substance)||S|PF|Y
C0006044|T129|86080005|SNOMEDCT_US|Botulism antitoxin (substance)||S|PF|Y
C0006044|T109|86080005|SNOMEDCT_US|Botulism antitoxin (substance)||S|PF|Y
C0006044|T121|4019149|VANDF|BOTULISM ANTITOXIN||S|VC|Y
C0006044|T129|4019149|VANDF|BOTULISM ANTITOXIN||S|VC|Y
C0006044|T109|4019149|VANDF|BOTULISM ANTITOXIN||S|VC|Y
C0008359|T121|90625|CPT|Cholera vaccine||P|VC|N
C0008359|T129|90625|CPT|Cholera vaccine||P|VC|N
C0008359|T121|3055-6111|CSP|cholera vaccine||P|VC|N
C0008359|T129|3055-6111|CSP|cholera vaccine||P|VC|N
C0008359|T121|26|CVX|cholera||S|VC|N
C0008359|T129|26|CVX|cholera||S|VC|N
C0008359|T121|26|CVX|cholera vaccine||P|VC|N
C0008359|T129|26|CVX|cholera vaccine||P|VC|N
C0008359|T121|26|HL7V2.5|cholera||S|VC|Y
C0008359|T129|26|HL7V2.5|cholera||S|VC|Y
C0008359|T121|26|HL7V3.0|Cholera||S|PF|Y
C0008359|T129|26|HL7V3.0|Cholera||S|PF|Y
C0008359|T121|40143|MEDCIN|cholera vaccine||P|VC|N
C0008359|T129|40143|MEDCIN|cholera vaccine||P|VC|N
C0008359|T121|40143|MEDCIN|cholera vaccine (medication)||S|PF|Y
C0008359|T129|40143|MEDCIN|cholera vaccine (medication)||S|PF|Y
C0008359|T121|4377|MMSL|Cholera Vaccine||P|PF|N
C0008359|T129|4377|MMSL|Cholera Vaccine||P|PF|N
C0008359|T121|d01154|MMSL|cholera vaccine||P|VC|Y
C0008359|T129|d01154|MMSL|cholera vaccine||P|VC|Y
C0008359|T121|D022121|MSH|Cholera Vaccines||P|VO|Y
C0008359|T129|D022121|MSH|Cholera Vaccines||P|VO|Y
C0008359|T121|D022121|MSH|Vaccines, Cholera||P|VO|Y
C0008359|T129|D022121|MSH|Vaccines, Cholera||P|VO|Y
C0008359|T121|U001808|MTH|Cholera Vaccine||P|PF|Y
C0008359|T129|U001808|MTH|Cholera Vaccine||P|PF|Y
C0008359|T121|N0000170887|NDFRT|Cholera Vaccines||P|VO|N
C0008359|T129|N0000170887|NDFRT|Cholera Vaccines||P|VO|N
C0008359|T121|N0000170887|NDFRT|Cholera Vaccines [Chemical/Ingredient]||S|PF|Y
C0008359|T129|N0000170887|NDFRT|Cholera Vaccines [Chemical/Ingredient]||S|PF|Y
C0008359|T121|2427|RXNORM|Cholera Vaccine||P|PF|N
C0008359|T129|2427|RXNORM|Cholera Vaccine||P|PF|N
C0008359|T121|35736007|SNOMEDCT_US|Cholera vaccine||P|VC|Y
C0008359|T129|35736007|SNOMEDCT_US|Cholera vaccine||P|VC|Y
C0008359|T121|35736007|SNOMEDCT_US|Cholera vaccine (product)||S|PF|Y
C0008359|T129|35736007|SNOMEDCT_US|Cholera vaccine (product)||S|PF|Y
C0008359|T121|35736007|SNOMEDCT_US|Cholera vaccine (substance)||S|PF|N
C0008359|T129|35736007|SNOMEDCT_US|Cholera vaccine (substance)||S|PF|N
C0008359|T121|35736007|SNOMEDCT_US|Cholera vaccines||P|VO|Y
C0008359|T129|35736007|SNOMEDCT_US|Cholera vaccines||P|VO|Y
C0008359|T121|396422009|SNOMEDCT_US|Cholera vaccine||P|VC|N
C0008359|T129|396422009|SNOMEDCT_US|Cholera vaccine||P|VC|N
C0008359|T121|396422009|SNOMEDCT_US|Cholera vaccine (substance)||S|PF|Y
C0008359|T129|396422009|SNOMEDCT_US|Cholera vaccine (substance)||S|PF|Y
C0012547|T121|12|CVX|diphtheria antitoxin||P|VC|N
C0012547|T129|12|CVX|diphtheria antitoxin||P|VC|N
C0012547|T116|12|CVX|diphtheria antitoxin||P|VC|N
C0012547|T121|12|HL7V2.5|diphtheria antitoxin||P|VC|N
C0012547|T129|12|HL7V2.5|diphtheria antitoxin||P|VC|N
C0012547|T116|12|HL7V2.5|diphtheria antitoxin||P|VC|N
C0012547|T121|12|HL7V3.0|diphtheria antitoxin||P|VC|N
C0012547|T129|12|HL7V3.0|diphtheria antitoxin||P|VC|N
C0012547|T116|12|HL7V3.0|diphtheria antitoxin||P|VC|N
C0012547|T121|sh85038154|LCH_NW|Diphtheria antitoxin||P|VC|N
C0012547|T129|sh85038154|LCH_NW|Diphtheria antitoxin||P|VC|N
C0012547|T116|sh85038154|LCH_NW|Diphtheria antitoxin||P|VC|N
C0012547|T121|40136|MEDCIN|diphtheria antitoxin||P|VC|N
C0012547|T129|40136|MEDCIN|diphtheria antitoxin||P|VC|N
C0012547|T116|40136|MEDCIN|diphtheria antitoxin||P|VC|N
C0012547|T121|40136|MEDCIN|diphtheria antitoxin (medication)||S|PF|Y
C0012547|T129|40136|MEDCIN|diphtheria antitoxin (medication)||S|PF|Y
C0012547|T116|40136|MEDCIN|diphtheria antitoxin (medication)||S|PF|Y
C0012547|T121|1701|MMSL|Diphtheria Antitoxin||P|PF|N
C0012547|T129|1701|MMSL|Diphtheria Antitoxin||P|PF|N
C0012547|T116|1701|MMSL|Diphtheria Antitoxin||P|PF|N
C0012547|T121|4615|MMSL|diphtheria antitoxin||P|VC|N
C0012547|T129|4615|MMSL|diphtheria antitoxin||P|VC|N
C0012547|T116|4615|MMSL|diphtheria antitoxin||P|VC|N
C0012547|T121|d01142|MMSL|diphtheria antitoxin||P|VC|Y
C0012547|T129|d01142|MMSL|diphtheria antitoxin||P|VC|Y
C0012547|T116|d01142|MMSL|diphtheria antitoxin||P|VC|Y
C0012547|T121|D004166|MSH|Antitoxin, Diphtheria||P|VW|Y
C0012547|T129|D004166|MSH|Antitoxin, Diphtheria||P|VW|Y
C0012547|T116|D004166|MSH|Antitoxin, Diphtheria||P|VW|Y
C0012547|T121|D004166|MSH|Diphtheria Antitoxin||P|PF|N
C0012547|T129|D004166|MSH|Diphtheria Antitoxin||P|PF|N
C0012547|T116|D004166|MSH|Diphtheria Antitoxin||P|PF|N
C0012547|T121|NOCODE|MTH|Diphtheria Antitoxin||P|PF|Y
C0012547|T129|NOCODE|MTH|Diphtheria Antitoxin||P|PF|Y
C0012547|T116|NOCODE|MTH|Diphtheria Antitoxin||P|PF|Y
C0012547|T121|N0000004696|NDFRT|Diphtheria Antitoxin||P|PF|N
C0012547|T129|N0000004696|NDFRT|Diphtheria Antitoxin||P|PF|N
C0012547|T116|N0000004696|NDFRT|Diphtheria Antitoxin||P|PF|N
C0012547|T121|N0000004696|NDFRT|Diphtheria Antitoxin [Chemical/Ingredient]||S|PF|Y
C0012547|T129|N0000004696|NDFRT|Diphtheria Antitoxin [Chemical/Ingredient]||S|PF|Y
C0012547|T116|N0000004696|NDFRT|Diphtheria Antitoxin [Chemical/Ingredient]||S|PF|Y
C0012547|T121|N0000020115|NDFRT|DIPHTHERIA ANTITOXIN||P|VC|N
C0012547|T129|N0000020115|NDFRT|DIPHTHERIA ANTITOXIN||P|VC|N
C0012547|T116|N0000020115|NDFRT|DIPHTHERIA ANTITOXIN||P|VC|N
C0012547|T121|3510|RXNORM|Diphtheria Antitoxin||P|PF|N
C0012547|T129|3510|RXNORM|Diphtheria Antitoxin||P|PF|N
C0012547|T116|3510|RXNORM|Diphtheria Antitoxin||P|PF|N
C0012547|T121|412175006|SNOMEDCT_US|Diphtheria antitoxin||P|VC|N
C0012547|T129|412175006|SNOMEDCT_US|Diphtheria antitoxin||P|VC|N
C0012547|T116|412175006|SNOMEDCT_US|Diphtheria antitoxin||P|VC|N
C0012547|T121|412175006|SNOMEDCT_US|Diphtheria antitoxin (substance)||S|PF|Y
C0012547|T129|412175006|SNOMEDCT_US|Diphtheria antitoxin (substance)||S|PF|Y
C0012547|T116|412175006|SNOMEDCT_US|Diphtheria antitoxin (substance)||S|PF|Y
C0012547|T121|412175006|SNOMEDCT_US|Diphtheria immunoglobulin||S|PF|Y
C0012547|T129|412175006|SNOMEDCT_US|Diphtheria immunoglobulin||S|PF|Y
C0012547|T116|412175006|SNOMEDCT_US|Diphtheria immunoglobulin||S|PF|Y
C0012547|T121|412175006|SNOMEDCT_US|Diptheria antitoxin||P|VO|Y
C0012547|T129|412175006|SNOMEDCT_US|Diptheria antitoxin||P|VO|Y
C0012547|T116|412175006|SNOMEDCT_US|Diptheria antitoxin||P|VO|Y
C0012547|T121|412175006|SNOMEDCT_US|Diptheria antitoxin (substance)||S|VO|Y
C0012547|T129|412175006|SNOMEDCT_US|Diptheria antitoxin (substance)||S|VO|Y
C0012547|T116|412175006|SNOMEDCT_US|Diptheria antitoxin (substance)||S|VO|Y
C0012547|T121|412175006|SNOMEDCT_US|Diptheria immunoglobulin||S|VO|Y
C0012547|T129|412175006|SNOMEDCT_US|Diptheria immunoglobulin||S|VO|Y
C0012547|T116|412175006|SNOMEDCT_US|Diptheria immunoglobulin||S|VO|Y
C0012547|T121|77048008|SNOMEDCT_US|Dip/ser||S|PF|Y
C0012547|T129|77048008|SNOMEDCT_US|Dip/ser||S|PF|Y
C0012547|T116|77048008|SNOMEDCT_US|Dip/ser||S|PF|Y
C0012547|T121|77048008|SNOMEDCT_US|Diphtheria antitoxin||P|VC|Y
C0012547|T129|77048008|SNOMEDCT_US|Diphtheria antitoxin||P|VC|Y
C0012547|T116|77048008|SNOMEDCT_US|Diphtheria antitoxin||P|VC|Y
C0012547|T121|77048008|SNOMEDCT_US|Diphtheria antitoxin (product)||S|PF|Y
C0012547|T129|77048008|SNOMEDCT_US|Diphtheria antitoxin (product)||S|PF|Y
C0012547|T116|77048008|SNOMEDCT_US|Diphtheria antitoxin (product)||S|PF|Y
C0012547|T121|77048008|SNOMEDCT_US|Diphtheria antitoxin (substance)||S|PF|N
C0012547|T129|77048008|SNOMEDCT_US|Diphtheria antitoxin (substance)||S|PF|N
C0012547|T116|77048008|SNOMEDCT_US|Diphtheria antitoxin (substance)||S|PF|N
C0012547|T121|4022109|VANDF|DIPHTHERIA ANTITOXIN||P|VC|Y
C0012547|T129|4022109|VANDF|DIPHTHERIA ANTITOXIN||P|VC|Y
C0012547|T116|4022109|VANDF|DIPHTHERIA ANTITOXIN||P|VC|Y
C0012559|T121|01|CVX|diphtheria, tetanus toxoids and pertussis vaccine||S|PF|Y
C0012559|T129|01|CVX|diphtheria, tetanus toxoids and pertussis vaccine||S|PF|Y
C0012559|T121|01|CVX|DTP||S|PF|N
C0012559|T129|01|CVX|DTP||S|PF|N
C0012559|T121|79263|GS|DTP Vaccine||S|PF|Y
C0012559|T129|79263|GS|DTP Vaccine||S|PF|Y
C0012559|T121|01|HL7V2.5|DTP||S|PF|N
C0012559|T129|01|HL7V2.5|DTP||S|PF|N
C0012559|T121|1|HL7V3.0|DTP||S|PF|Y
C0012559|T129|1|HL7V3.0|DTP||S|PF|Y
C0012559|T121|436|MMSL|DTP Vaccine||S|PF|N
C0012559|T129|436|MMSL|DTP Vaccine||S|PF|N
C0012559|T121|7421|MMSL|diphtheria, pertussis, tetanus vaccine||P|VCW|Y
C0012559|T129|7421|MMSL|diphtheria, pertussis, tetanus vaccine||P|VCW|Y
C0012559|T121|NOCODE|MTH|Diphtheria-Tetanus-Pertussis Vaccine||P|PF|Y
C0012559|T129|NOCODE|MTH|Diphtheria-Tetanus-Pertussis Vaccine||P|PF|Y
C0012559|T121|421245007|SNOMEDCT_US|Diphtheria + pertussis + tetanus vaccine||P|VCW|Y
C0012559|T129|421245007|SNOMEDCT_US|Diphtheria + pertussis + tetanus vaccine||P|VCW|Y
C0012559|T121|421245007|SNOMEDCT_US|Diphtheria + pertussis + tetanus vaccine (product)||S|PF|Y
C0012559|T129|421245007|SNOMEDCT_US|Diphtheria + pertussis + tetanus vaccine (product)||S|PF|Y
C0012559|T121|421245007|SNOMEDCT_US|Diphtheria and tetanus toxoids with pertussis, combined vaccine||S|PF|Y
C0012559|T129|421245007|SNOMEDCT_US|Diphtheria and tetanus toxoids with pertussis, combined vaccine||S|PF|Y
C0012559|T121|421245007|SNOMEDCT_US|Diptheria + pertussis + tetanus vaccine||P|VO|Y
C0012559|T129|421245007|SNOMEDCT_US|Diptheria + pertussis + tetanus vaccine||P|VO|Y
C0012559|T121|421245007|SNOMEDCT_US|Diptheria + pertussis + tetanus vaccine (product)||S|VO|Y
C0012559|T129|421245007|SNOMEDCT_US|Diptheria + pertussis + tetanus vaccine (product)||S|VO|Y
C0012559|T121|421245007|SNOMEDCT_US|DPT - Diphtheria + pertussis + tetanus vaccine||S|PF|Y
C0012559|T129|421245007|SNOMEDCT_US|DPT - Diphtheria + pertussis + tetanus vaccine||S|PF|Y
C0012559|T121|421245007|SNOMEDCT_US|DTP - Diphtheria + tetanus + pertussis vaccine||S|PF|Y
C0012559|T129|421245007|SNOMEDCT_US|DTP - Diphtheria + tetanus + pertussis vaccine||S|PF|Y
C0012559|T121|54667003|SNOMEDCT_US|Diphtheria and tetanus toxoids with pertussis, combined vaccine||S|PF|N
C0012559|T129|54667003|SNOMEDCT_US|Diphtheria and tetanus toxoids with pertussis, combined vaccine||S|PF|N
C0012559|T121|54667003|SNOMEDCT_US|Diphtheria and tetanus toxoids with pertussis, combined vaccine (product)||S|PF|Y
C0012559|T129|54667003|SNOMEDCT_US|Diphtheria and tetanus toxoids with pertussis, combined vaccine (product)||S|PF|Y
C0012559|T121|54667003|SNOMEDCT_US|Diphtheria and tetanus toxoids with pertussis, combined vaccine (substance)||S|PF|Y
C0012559|T129|54667003|SNOMEDCT_US|Diphtheria and tetanus toxoids with pertussis, combined vaccine (substance)||S|PF|Y
C0012559|T121|54667003|SNOMEDCT_US|Diphtheria+tetanus+pertussis vaccine||P|VC|Y
C0012559|T129|54667003|SNOMEDCT_US|Diphtheria+tetanus+pertussis vaccine||P|VC|Y
C0012559|T121|54667003|SNOMEDCT_US|DPT||S|PF|Y
C0012559|T129|54667003|SNOMEDCT_US|DPT||S|PF|Y
C0012559|T121|54667003|SNOMEDCT_US|DTP||S|PF|N
C0012559|T129|54667003|SNOMEDCT_US|DTP||S|PF|N
C0025010|T121|3060-1063|CSP|measles vaccine||P|VC|Y
C0025010|T129|3060-1063|CSP|measles vaccine||P|VC|Y
C0025010|T121|05|CVX|measles||S|PF|N
C0025010|T129|05|CVX|measles||S|PF|N
C0025010|T121|05|CVX|measles virus vaccine||S|PF|N
C0025010|T129|05|CVX|measles virus vaccine||S|PF|N
C0025010|T121|05|HL7V2.5|measles||S|PF|N
C0025010|T129|05|HL7V2.5|measles||S|PF|N
C0025010|T121|5|HL7V3.0|measles||S|PF|Y
C0025010|T129|5|HL7V3.0|measles||S|PF|Y
C0025010|T121|sh85082698|LCH_NW|Measles vaccine||P|VC|N
C0025010|T129|sh85082698|LCH_NW|Measles vaccine||P|VC|N
C0025010|T121|7408|MMSL|measles virus vaccine||S|PF|N
C0025010|T129|7408|MMSL|measles virus vaccine||S|PF|N
C0025010|T121|d01159|MMSL|measles virus vaccine||S|PF|Y
C0025010|T129|d01159|MMSL|measles virus vaccine||S|PF|Y
C0025010|T121|D008458|MSH|Measles Vaccine||P|PF|N
C0025010|T129|D008458|MSH|Measles Vaccine||P|PF|N
C0025010|T121|D008458|MSH|Vaccine, Measles||P|VW|Y
C0025010|T129|D008458|MSH|Vaccine, Measles||P|VW|Y
C0025010|T121|NOCODE|MTH|Measles Vaccine||P|PF|Y
C0025010|T129|NOCODE|MTH|Measles Vaccine||P|PF|Y
C0025010|T121|N0000170910|NDFRT|Measles Vaccine||P|PF|N
C0025010|T129|N0000170910|NDFRT|Measles Vaccine||P|PF|N
C0025010|T121|N0000170910|NDFRT|Measles Vaccine [Chemical/Ingredient]||S|PF|Y
C0025010|T129|N0000170910|NDFRT|Measles Vaccine [Chemical/Ingredient]||S|PF|Y
C0025010|T121|6669|RXNORM|Measles Vaccine||P|PF|N
C0025010|T129|6669|RXNORM|Measles Vaccine||P|PF|N
C0025010|T121|386012008|SNOMEDCT_US|Measles live virus vaccine||S|PF|N
C0025010|T129|386012008|SNOMEDCT_US|Measles live virus vaccine||S|PF|N
C0025010|T121|386012008|SNOMEDCT_US|Measles vaccine||P|VC|Y
C0025010|T129|386012008|SNOMEDCT_US|Measles vaccine||P|VC|Y
C0025010|T121|386012008|SNOMEDCT_US|Measles vaccine (product)||S|PF|Y
C0025010|T129|386012008|SNOMEDCT_US|Measles vaccine (product)||S|PF|Y
C0025010|T121|386012008|SNOMEDCT_US|Rubeola virus vaccine||S|PF|Y
C0025010|T129|386012008|SNOMEDCT_US|Rubeola virus vaccine||S|PF|Y
C0025010|T121|396427003|SNOMEDCT_US|Measles live virus vaccine||S|PF|Y
C0025010|T129|396427003|SNOMEDCT_US|Measles live virus vaccine||S|PF|Y
C0025010|T121|396427003|SNOMEDCT_US|Measles vaccine||P|VC|N
C0025010|T129|396427003|SNOMEDCT_US|Measles vaccine||P|VC|N
C0025010|T121|396427003|SNOMEDCT_US|Measles vaccine (substance)||S|PF|Y
C0025010|T129|396427003|SNOMEDCT_US|Measles vaccine (substance)||S|PF|Y
C0025010|T121|396427003|SNOMEDCT_US|Rubeola virus vaccine||S|PF|N
C0025010|T129|396427003|SNOMEDCT_US|Rubeola virus vaccine||S|PF|N
C0025010|T121|396428008|SNOMEDCT_US|Measles live virus vaccine||S|PF|N
C0025010|T129|396428008|SNOMEDCT_US|Measles live virus vaccine||S|PF|N
C0025010|T121|396428008|SNOMEDCT_US|Measles live virus vaccine (substance)||S|PF|Y
C0025010|T129|396428008|SNOMEDCT_US|Measles live virus vaccine (substance)||S|PF|Y
C0025010|T121|87939007|SNOMEDCT_US|Measles live virus vaccine||S|PF|N
C0025010|T129|87939007|SNOMEDCT_US|Measles live virus vaccine||S|PF|N
C0025010|T121|87939007|SNOMEDCT_US|Measles live virus vaccine (product)||S|PF|Y
C0025010|T129|87939007|SNOMEDCT_US|Measles live virus vaccine (product)||S|PF|Y
C0025010|T121|87939007|SNOMEDCT_US|Measles live virus vaccine (substance)||S|PF|N
C0025010|T129|87939007|SNOMEDCT_US|Measles live virus vaccine (substance)||S|PF|N
C0025010|T121|87939007|SNOMEDCT_US|Rubeola virus vaccine||S|PF|N
C0025010|T129|87939007|SNOMEDCT_US|Rubeola virus vaccine||S|PF|N
C0026782|T121|07|CVX|mumps||S|PF|N
C0026782|T129|07|CVX|mumps||S|PF|N
C0026782|T121|07|CVX|mumps virus vaccine||S|PF|N
C0026782|T129|07|CVX|mumps virus vaccine||S|PF|N
C0026782|T121|07|HL7V2.5|mumps||S|PF|N
C0026782|T129|07|HL7V2.5|mumps||S|PF|N
C0026782|T121|7|HL7V3.0|mumps||S|PF|Y
C0026782|T129|7|HL7V3.0|mumps||S|PF|Y
C0026782|T121|40150|MEDCIN|vaccines viral mumps, live||S|PF|Y
C0026782|T129|40150|MEDCIN|vaccines viral mumps, live||S|PF|Y
C0026782|T121|40150|MEDCIN|vaccines viral mumps, live (medication)||S|PF|Y
C0026782|T129|40150|MEDCIN|vaccines viral mumps, live (medication)||S|PF|Y
C0026782|T121|7418|MMSL|mumps virus vaccine, live||S|VCW|Y
C0026782|T129|7418|MMSL|mumps virus vaccine, live||S|VCW|Y
C0026782|T121|d01161|MMSL|mumps virus vaccine||S|PF|Y
C0026782|T129|d01161|MMSL|mumps virus vaccine||S|PF|Y
C0026782|T121|D009108|MSH|Mumps Vaccine||P|PF|N
C0026782|T129|D009108|MSH|Mumps Vaccine||P|PF|N
C0026782|T121|D009108|MSH|Vaccine, Mumps||P|VW|Y
C0026782|T129|D009108|MSH|Vaccine, Mumps||P|VW|Y
C0026782|T121|NOCODE|MTH|Mumps Vaccine||P|PF|Y
C0026782|T129|NOCODE|MTH|Mumps Vaccine||P|PF|Y
C0026782|T121|N0000146322|NDFRT|MUMPS VIRUS VACCINE,LIVE||S|VCW|N
C0026782|T129|N0000146322|NDFRT|MUMPS VIRUS VACCINE,LIVE||S|VCW|N
C0026782|T121|N0000170898|NDFRT|Mumps Vaccine||P|PF|N
C0026782|T129|N0000170898|NDFRT|Mumps Vaccine||P|PF|N
C0026782|T121|N0000170898|NDFRT|Mumps Vaccine [Chemical/Ingredient]||S|PF|Y
C0026782|T129|N0000170898|NDFRT|Mumps Vaccine [Chemical/Ingredient]||S|PF|Y
C0026782|T121|763656|RXNORM|Mumps Vaccine||P|PF|N
C0026782|T129|763656|RXNORM|Mumps Vaccine||P|PF|N
C0026782|T121|396431009|SNOMEDCT_US|Mumps vaccine||P|VC|Y
C0026782|T129|396431009|SNOMEDCT_US|Mumps vaccine||P|VC|Y
C0026782|T121|396431009|SNOMEDCT_US|Mumps vaccine (substance)||S|PF|Y
C0026782|T129|396431009|SNOMEDCT_US|Mumps vaccine (substance)||S|PF|Y
C0026782|T121|90043005|SNOMEDCT_US|Mumps live virus vaccine||S|PF|Y
C0026782|T129|90043005|SNOMEDCT_US|Mumps live virus vaccine||S|PF|Y
C0026782|T121|90043005|SNOMEDCT_US|Mumps live virus vaccine (product)||S|PF|Y
C0026782|T129|90043005|SNOMEDCT_US|Mumps live virus vaccine (product)||S|PF|Y
C0026782|T121|90043005|SNOMEDCT_US|Mumps live virus vaccine (substance)||S|PF|Y
C0026782|T129|90043005|SNOMEDCT_US|Mumps live virus vaccine (substance)||S|PF|Y
C0026782|T121|90043005|SNOMEDCT_US|Mumps vaccine||P|VC|N
C0026782|T129|90043005|SNOMEDCT_US|Mumps vaccine||P|VC|N
C0026782|T121|4017972|VANDF|MUMPS VIRUS VACCINE,LIVE||S|VCW|Y
C0026782|T129|4017972|VANDF|MUMPS VIRUS VACCINE,LIVE||S|VCW|Y
C0031237|T121|3055-7984|CSP|pertussis vaccine||P|VC|N
C0031237|T129|3055-7984|CSP|pertussis vaccine||P|VC|N
C0031237|T121|11|CVX|pertussis||S|VC|N
C0031237|T129|11|CVX|pertussis||S|VC|N
C0031237|T121|11|CVX|pertussis vaccine||P|VC|Y
C0031237|T129|11|CVX|pertussis vaccine||P|VC|Y
C0031237|T121|11|HL7V2.5|pertussis||S|VC|N
C0031237|T129|11|HL7V2.5|pertussis||S|VC|N
C0031237|T121|11|HL7V3.0|pertussis||S|VC|Y
C0031237|T129|11|HL7V3.0|pertussis||S|VC|Y
C0031237|T121|LA10493-7|LNC|Pertussis||S|PF|Y
C0031237|T129|LA10493-7|LNC|Pertussis||S|PF|Y
C0031237|T121|461|MEDLINEPLUS|Pertussis||S|PF|N
C0031237|T129|461|MEDLINEPLUS|Pertussis||S|PF|N
C0031237|T121|D010567|MSH|Pertussis Vaccine||P|PF|N
C0031237|T129|D010567|MSH|Pertussis Vaccine||P|PF|N
C0031237|T121|D010567|MSH|Vaccine, Pertussis||P|VW|Y
C0031237|T129|D010567|MSH|Vaccine, Pertussis||P|VW|Y
C0031237|T121|NOCODE|MTH|Pertussis Vaccine||P|PF|Y
C0031237|T129|NOCODE|MTH|Pertussis Vaccine||P|PF|Y
C0031237|T121|N0000005258|NDFRT|Pertussis Vaccine||P|PF|N
C0031237|T129|N0000005258|NDFRT|Pertussis Vaccine||P|PF|N
C0031237|T121|N0000005258|NDFRT|Pertussis Vaccine [Chemical/Ingredient]||S|PF|Y
C0031237|T129|N0000005258|NDFRT|Pertussis Vaccine [Chemical/Ingredient]||S|PF|Y
C0031237|T121|N0000146177|NDFRT|PERTUSSIS VACCINE||P|VC|N
C0031237|T129|N0000146177|NDFRT|PERTUSSIS VACCINE||P|VC|N
C0031237|T121|8080|RXNORM|Pertussis Vaccine||P|PF|N
C0031237|T129|8080|RXNORM|Pertussis Vaccine||P|PF|N
C0031237|T121|396433007|SNOMEDCT_US|Pertussis vaccine||P|VC|Y
C0031237|T129|396433007|SNOMEDCT_US|Pertussis vaccine||P|VC|Y
C0031237|T121|396433007|SNOMEDCT_US|Pertussis vaccine (substance)||S|PF|Y
C0031237|T129|396433007|SNOMEDCT_US|Pertussis vaccine (substance)||S|PF|Y
C0031237|T121|61602008|SNOMEDCT_US|Pertussis vaccine||P|VC|N
C0031237|T129|61602008|SNOMEDCT_US|Pertussis vaccine||P|VC|N
C0031237|T121|61602008|SNOMEDCT_US|Pertussis vaccine (product)||S|PF|Y
C0031237|T129|61602008|SNOMEDCT_US|Pertussis vaccine (product)||S|PF|Y
C0031237|T121|61602008|SNOMEDCT_US|Pertussis vaccine (substance)||S|PF|N
C0031237|T129|61602008|SNOMEDCT_US|Pertussis vaccine (substance)||S|PF|N
C0031237|T121|61602008|SNOMEDCT_US|Whooping-cough vaccine||S|PF|Y
C0031237|T129|61602008|SNOMEDCT_US|Whooping-cough vaccine||S|PF|Y
C0031237|T121|4017817|VANDF|PERTUSSIS VACCINE||P|VC|Y
C0031237|T129|4017817|VANDF|PERTUSSIS VACCINE||P|VC|Y
C0032066|T121|23|CVX|plague||S|PF|N
C0032066|T129|23|CVX|plague||S|PF|N
C0032066|T121|23|CVX|plague vaccine||P|VC|N
C0032066|T129|23|CVX|plague vaccine||P|VC|N
C0032066|T121|23|HL7V2.5|plague||S|PF|N
C0032066|T129|23|HL7V2.5|plague||S|PF|N
C0032066|T121|23|HL7V3.0|plague||S|PF|Y
C0032066|T129|23|HL7V3.0|plague||S|PF|Y
C0032066|T121|sh85102598|LCH_NW|Plague vaccines||P|VO|Y
C0032066|T129|sh85102598|LCH_NW|Plague vaccines||P|VO|Y
C0032066|T121|40151|MEDCIN|plague vaccine||P|VC|N
C0032066|T129|40151|MEDCIN|plague vaccine||P|VC|N
C0032066|T121|40151|MEDCIN|plague vaccine (medication)||S|PF|Y
C0032066|T129|40151|MEDCIN|plague vaccine (medication)||S|PF|Y
C0032066|T121|5982|MMSL|Plague Vaccine||P|PF|N
C0032066|T129|5982|MMSL|Plague Vaccine||P|PF|N
C0032066|T121|d01155|MMSL|plague vaccine||P|VC|Y
C0032066|T129|d01155|MMSL|plague vaccine||P|VC|Y
C0032066|T121|D010931|MSH|Plague Vaccine||P|PF|N
C0032066|T129|D010931|MSH|Plague Vaccine||P|PF|N
C0032066|T121|D010931|MSH|Vaccine, Plague||P|VW|Y
C0032066|T129|D010931|MSH|Vaccine, Plague||P|VW|Y
C0032066|T121|U002172|MTH|Plague Vaccine||P|PF|Y
C0032066|T129|U002172|MTH|Plague Vaccine||P|PF|Y
C0032066|T121|N0000005307|NDFRT|Plague Vaccine||P|PF|N
C0032066|T129|N0000005307|NDFRT|Plague Vaccine||P|PF|N
C0032066|T121|N0000005307|NDFRT|Plague Vaccine [Chemical/Ingredient]||S|PF|Y
C0032066|T129|N0000005307|NDFRT|Plague Vaccine [Chemical/Ingredient]||S|PF|Y
C0032066|T121|N0000022466|NDFRT|PLAGUE VACCINE||P|VC|N
C0032066|T129|N0000022466|NDFRT|PLAGUE VACCINE||P|VC|N
C0032066|T121|11866009|SNOMEDCT_US|Plague vaccine||P|VC|Y
C0032066|T129|11866009|SNOMEDCT_US|Plague vaccine||P|VC|Y
C0032066|T121|11866009|SNOMEDCT_US|Plague vaccine (product)||S|PF|Y
C0032066|T129|11866009|SNOMEDCT_US|Plague vaccine (product)||S|PF|Y
C0032066|T121|11866009|SNOMEDCT_US|Plague vaccine (substance)||S|PF|N
C0032066|T129|11866009|SNOMEDCT_US|Plague vaccine (substance)||S|PF|N
C0032066|T121|412477009|SNOMEDCT_US|Plague vaccine||P|VC|N
C0032066|T129|412477009|SNOMEDCT_US|Plague vaccine||P|VC|N
C0032066|T121|412477009|SNOMEDCT_US|Plague vaccine (substance)||S|PF|Y
C0032066|T129|412477009|SNOMEDCT_US|Plague vaccine (substance)||S|PF|Y
C0032066|T121|4018881|VANDF|PLAGUE VACCINE||P|VC|Y
C0032066|T129|4018881|VANDF|PLAGUE VACCINE||P|VC|Y
C0032375|T109|02|CVX|OPV||S|PF|N
C0032375|T129|02|CVX|OPV||S|PF|N
C0032375|T121|02|CVX|OPV||S|PF|N
C0032375|T109|02|CVX|poliovirus vaccine, live, oral||S|PF|Y
C0032375|T129|02|CVX|poliovirus vaccine, live, oral||S|PF|Y
C0032375|T121|02|CVX|poliovirus vaccine, live, oral||S|PF|Y
C0032375|T109|02|HL7V2.5|OPV||S|PF|N
C0032375|T129|02|HL7V2.5|OPV||S|PF|N
C0032375|T121|02|HL7V2.5|OPV||S|PF|N
C0032375|T109|2|HL7V3.0|OPV||S|PF|N
C0032375|T129|2|HL7V3.0|OPV||S|PF|N
C0032375|T121|2|HL7V3.0|OPV||S|PF|N
C0032375|T109|sh85104278|LCH_NW|Poliomyelitis vaccine, Oral||S|PF|Y
C0032375|T129|sh85104278|LCH_NW|Poliomyelitis vaccine, Oral||S|PF|Y
C0032375|T121|sh85104278|LCH_NW|Poliomyelitis vaccine, Oral||S|PF|Y
C0032375|T109|D011055|MSH|Oral Poliovirus Vaccine||P|PF|N
C0032375|T129|D011055|MSH|Oral Poliovirus Vaccine||P|PF|N
C0032375|T121|D011055|MSH|Oral Poliovirus Vaccine||P|PF|N
C0032375|T109|D011055|MSH|Poliovirus Vaccine, Oral||P|VW|Y
C0032375|T129|D011055|MSH|Poliovirus Vaccine, Oral||P|VW|Y
C0032375|T121|D011055|MSH|Poliovirus Vaccine, Oral||P|VW|Y
C0032375|T109|D011055|MSH|Sabin Vaccine||S|PF|Y
C0032375|T129|D011055|MSH|Sabin Vaccine||S|PF|Y
C0032375|T121|D011055|MSH|Sabin Vaccine||S|PF|Y
C0032375|T109|D011055|MSH|Vaccine, Oral Poliovirus||P|VW|Y
C0032375|T129|D011055|MSH|Vaccine, Oral Poliovirus||P|VW|Y
C0032375|T121|D011055|MSH|Vaccine, Oral Poliovirus||P|VW|Y
C0032375|T109|D011055|MSH|Vaccine, Sabin||S|VW|Y
C0032375|T129|D011055|MSH|Vaccine, Sabin||S|VW|Y
C0032375|T121|D011055|MSH|Vaccine, Sabin||S|VW|Y
C0032375|T109|NOCODE|MTH|Oral Poliovirus Vaccine||P|PF|Y
C0032375|T129|NOCODE|MTH|Oral Poliovirus Vaccine||P|PF|Y
C0032375|T121|NOCODE|MTH|Oral Poliovirus Vaccine||P|PF|Y
C0032375|T109|C96401|NCI|OPV||S|PF|N
C0032375|T129|C96401|NCI|OPV||S|PF|N
C0032375|T121|C96401|NCI|OPV||S|PF|N
C0032375|T109|C96401|NCI|Oral Polio Vaccine||S|PF|Y
C0032375|T129|C96401|NCI|Oral Polio Vaccine||S|PF|Y
C0032375|T121|C96401|NCI|Oral Polio Vaccine||S|PF|Y
C0032375|T109|C96401|NCI_NICHD|Oral Polio Vaccine||S|PF|N
C0032375|T129|C96401|NCI_NICHD|Oral Polio Vaccine||S|PF|N
C0032375|T121|C96401|NCI_NICHD|Oral Polio Vaccine||S|PF|N
C0032375|T109|N0000170901|NDFRT|Poliovirus Vaccine, Oral||P|VW|N
C0032375|T129|N0000170901|NDFRT|Poliovirus Vaccine, Oral||P|VW|N
C0032375|T121|N0000170901|NDFRT|Poliovirus Vaccine, Oral||P|VW|N
C0032375|T109|N0000170901|NDFRT|Poliovirus Vaccine, Oral [Chemical/Ingredient]||S|PF|Y
C0032375|T129|N0000170901|NDFRT|Poliovirus Vaccine, Oral [Chemical/Ingredient]||S|PF|Y
C0032375|T121|N0000170901|NDFRT|Poliovirus Vaccine, Oral [Chemical/Ingredient]||S|PF|Y
C0032375|T109|N0000170901|NDFRT|Sabin Vaccine||S|PF|N
C0032375|T129|N0000170901|NDFRT|Sabin Vaccine||S|PF|N
C0032375|T121|N0000170901|NDFRT|Sabin Vaccine||S|PF|N
C0032375|T109|111164008|SNOMEDCT_US|OPV||S|PF|Y
C0032375|T129|111164008|SNOMEDCT_US|OPV||S|PF|Y
C0032375|T121|111164008|SNOMEDCT_US|OPV||S|PF|Y
C0032375|T109|111164008|SNOMEDCT_US|Sabin vaccine||S|VC|Y
C0032375|T129|111164008|SNOMEDCT_US|Sabin vaccine||S|VC|Y
C0032375|T121|111164008|SNOMEDCT_US|Sabin vaccine||S|VC|Y
C0032375|T109|111164008|SNOMEDCT_US|TOPV||S|PF|Y
C0032375|T129|111164008|SNOMEDCT_US|TOPV||S|PF|Y
C0032375|T121|111164008|SNOMEDCT_US|TOPV||S|PF|Y
C0032375|T109|125690004|SNOMEDCT_US|OPV||S|PF|N
C0032375|T129|125690004|SNOMEDCT_US|OPV||S|PF|N
C0032375|T121|125690004|SNOMEDCT_US|OPV||S|PF|N
C0032375|T109|125690004|SNOMEDCT_US|Pol/Vac (oral)||S|PF|N
C0032375|T129|125690004|SNOMEDCT_US|Pol/Vac (oral)||S|PF|N
C0032375|T121|125690004|SNOMEDCT_US|Pol/Vac (oral)||S|PF|N
C0032375|T109|125690004|SNOMEDCT_US|Sabin vaccine||S|VC|N
C0032375|T129|125690004|SNOMEDCT_US|Sabin vaccine||S|VC|N
C0032375|T121|125690004|SNOMEDCT_US|Sabin vaccine||S|VC|N
C0032375|T109|268590009|SNOMEDCT_US|Oral polio vaccine||S|VC|Y
C0032375|T129|268590009|SNOMEDCT_US|Oral polio vaccine||S|VC|Y
C0032375|T121|268590009|SNOMEDCT_US|Oral polio vaccine||S|VC|Y
C0032375|T109|396436004|SNOMEDCT_US|OPV||S|PF|N
C0032375|T129|396436004|SNOMEDCT_US|OPV||S|PF|N
C0032375|T121|396436004|SNOMEDCT_US|OPV||S|PF|N
C0032375|T109|396436004|SNOMEDCT_US|Pol/Vac (oral)||S|PF|Y
C0032375|T129|396436004|SNOMEDCT_US|Pol/Vac (oral)||S|PF|Y
C0032375|T121|396436004|SNOMEDCT_US|Pol/Vac (oral)||S|PF|Y
C0032375|T109|396436004|SNOMEDCT_US|Sabin vaccine||S|VC|N
C0032375|T129|396436004|SNOMEDCT_US|Sabin vaccine||S|VC|N
C0032375|T121|396436004|SNOMEDCT_US|Sabin vaccine||S|VC|N
C0035923|T121|06|CVX|rubella||S|PF|N
C0035923|T116|06|CVX|rubella||S|PF|N
C0035923|T129|06|CVX|rubella||S|PF|N
C0035923|T121|06|CVX|rubella virus vaccine||P|VC|N
C0035923|T116|06|CVX|rubella virus vaccine||P|VC|N
C0035923|T129|06|CVX|rubella virus vaccine||P|VC|N
C0035923|T121|06|HL7V2.5|rubella||S|PF|N
C0035923|T116|06|HL7V2.5|rubella||S|PF|N
C0035923|T129|06|HL7V2.5|rubella||S|PF|N
C0035923|T121|6|HL7V3.0|rubella||S|PF|Y
C0035923|T116|6|HL7V3.0|rubella||S|PF|Y
C0035923|T129|6|HL7V3.0|rubella||S|PF|Y
C0035923|T121|sh85115674|LCH_NW|Rubella vaccines||S|VO|Y
C0035923|T116|sh85115674|LCH_NW|Rubella vaccines||S|VO|Y
C0035923|T129|sh85115674|LCH_NW|Rubella vaccines||S|VO|Y
C0035923|T121|7419|MMSL|rubella virus vaccine||P|VC|N
C0035923|T116|7419|MMSL|rubella virus vaccine||P|VC|N
C0035923|T129|7419|MMSL|rubella virus vaccine||P|VC|N
C0035923|T121|d01160|MMSL|rubella virus vaccine||P|VC|Y
C0035923|T116|d01160|MMSL|rubella virus vaccine||P|VC|Y
C0035923|T129|d01160|MMSL|rubella virus vaccine||P|VC|Y
C0035923|T121|D012411|MSH|Rubella Vaccine||S|PF|Y
C0035923|T116|D012411|MSH|Rubella Vaccine||S|PF|Y
C0035923|T129|D012411|MSH|Rubella Vaccine||S|PF|Y
C0035923|T121|D012411|MSH|Vaccine, Rubella||S|VW|Y
C0035923|T116|D012411|MSH|Vaccine, Rubella||S|VW|Y
C0035923|T129|D012411|MSH|Vaccine, Rubella||S|VW|Y
C0035923|T121|NOCODE|MTH|Rubella virus vaccine||P|PF|Y
C0035923|T116|NOCODE|MTH|Rubella virus vaccine||P|PF|Y
C0035923|T129|NOCODE|MTH|Rubella virus vaccine||P|PF|Y
C0035923|T121|N0000146325|NDFRT|RUBELLA VIRUS VACCINE,LIVE||S|PF|N
C0035923|T116|N0000146325|NDFRT|RUBELLA VIRUS VACCINE,LIVE||S|PF|N
C0035923|T129|N0000146325|NDFRT|RUBELLA VIRUS VACCINE,LIVE||S|PF|N
C0035923|T121|N0000170894|NDFRT|Rubella Vaccine||S|PF|N
C0035923|T116|N0000170894|NDFRT|Rubella Vaccine||S|PF|N
C0035923|T129|N0000170894|NDFRT|Rubella Vaccine||S|PF|N
C0035923|T121|N0000170894|NDFRT|Rubella Vaccine [Chemical/Ingredient]||S|PF|Y
C0035923|T116|N0000170894|NDFRT|Rubella Vaccine [Chemical/Ingredient]||S|PF|Y
C0035923|T129|N0000170894|NDFRT|Rubella Vaccine [Chemical/Ingredient]||S|PF|Y
C0035923|T121|9486|RXNORM|Rubella virus vaccine||P|PF|N
C0035923|T116|9486|RXNORM|Rubella virus vaccine||P|PF|N
C0035923|T129|9486|RXNORM|Rubella virus vaccine||P|PF|N
C0035923|T121|386013003|SNOMEDCT_US|German measles vaccine||S|PF|Y
C0035923|T116|386013003|SNOMEDCT_US|German measles vaccine||S|PF|Y
C0035923|T129|386013003|SNOMEDCT_US|German measles vaccine||S|PF|Y
C0035923|T121|386013003|SNOMEDCT_US|Rubella vaccine||S|VC|Y
C0035923|T116|386013003|SNOMEDCT_US|Rubella vaccine||S|VC|Y
C0035923|T129|386013003|SNOMEDCT_US|Rubella vaccine||S|VC|Y
C0035923|T121|386013003|SNOMEDCT_US|Rubella vaccine (product)||S|PF|Y
C0035923|T116|386013003|SNOMEDCT_US|Rubella vaccine (product)||S|PF|Y
C0035923|T129|386013003|SNOMEDCT_US|Rubella vaccine (product)||S|PF|Y
C0035923|T121|396438003|SNOMEDCT_US|German measles vaccine||S|PF|N
C0035923|T116|396438003|SNOMEDCT_US|German measles vaccine||S|PF|N
C0035923|T129|396438003|SNOMEDCT_US|German measles vaccine||S|PF|N
C0035923|T121|396438003|SNOMEDCT_US|Rubella vaccine||S|VC|N
C0035923|T116|396438003|SNOMEDCT_US|Rubella vaccine||S|VC|N
C0035923|T129|396438003|SNOMEDCT_US|Rubella vaccine||S|VC|N
C0035923|T121|396438003|SNOMEDCT_US|Rubella vaccine (substance)||S|PF|Y
C0035923|T116|396438003|SNOMEDCT_US|Rubella vaccine (substance)||S|PF|Y
C0035923|T129|396438003|SNOMEDCT_US|Rubella vaccine (substance)||S|PF|Y
C0035923|T121|5524008|SNOMEDCT_US|German measles virus vaccine||S|PF|Y
C0035923|T116|5524008|SNOMEDCT_US|German measles virus vaccine||S|PF|Y
C0035923|T129|5524008|SNOMEDCT_US|German measles virus vaccine||S|PF|Y
C0035923|T121|5524008|SNOMEDCT_US|Rubella live virus vaccine||S|VCW|Y
C0035923|T116|5524008|SNOMEDCT_US|Rubella live virus vaccine||S|VCW|Y
C0035923|T129|5524008|SNOMEDCT_US|Rubella live virus vaccine||S|VCW|Y
C0035923|T121|5524008|SNOMEDCT_US|Rubella live virus vaccine (product)||S|PF|Y
C0035923|T116|5524008|SNOMEDCT_US|Rubella live virus vaccine (product)||S|PF|Y
C0035923|T129|5524008|SNOMEDCT_US|Rubella live virus vaccine (product)||S|PF|Y
C0035923|T121|5524008|SNOMEDCT_US|Rubella live virus vaccine (substance)||S|PF|Y
C0035923|T116|5524008|SNOMEDCT_US|Rubella live virus vaccine (substance)||S|PF|Y
C0035923|T129|5524008|SNOMEDCT_US|Rubella live virus vaccine (substance)||S|PF|Y
C0035923|T121|5524008|SNOMEDCT_US|Rubella vaccine||S|VC|N
C0035923|T116|5524008|SNOMEDCT_US|Rubella vaccine||S|VC|N
C0035923|T129|5524008|SNOMEDCT_US|Rubella vaccine||S|VC|N
C0035923|T121|5524008|SNOMEDCT_US|Rubella virus vaccine||P|PF|N
C0035923|T116|5524008|SNOMEDCT_US|Rubella virus vaccine||P|PF|N
C0035923|T129|5524008|SNOMEDCT_US|Rubella virus vaccine||P|PF|N
C0035923|T121|4017976|VANDF|RUBELLA VIRUS VACCINE,LIVE||S|PF|Y
C0035923|T116|4017976|VANDF|RUBELLA VIRUS VACCINE,LIVE||S|PF|Y
C0035923|T129|4017976|VANDF|RUBELLA VIRUS VACCINE,LIVE||S|PF|Y
C0037355|T121|5003-0043|CSP|smallpox vaccine||P|VC|N
C0037355|T129|5003-0043|CSP|smallpox vaccine||P|VC|N
C0037355|T121|75|CVX|vaccinia (smallpox)||S|PF|Y
C0037355|T129|75|CVX|vaccinia (smallpox)||S|PF|Y
C0037355|T121|75|CVX|vaccinia (smallpox) vaccine||S|PF|Y
C0037355|T129|75|CVX|vaccinia (smallpox) vaccine||S|PF|Y
C0037355|T121|75|HL7V2.5|smallpox||S|PF|N
C0037355|T129|75|HL7V2.5|smallpox||S|PF|N
C0037355|T121|75|HL7V3.0|smallpox||S|PF|Y
C0037355|T129|75|HL7V3.0|smallpox||S|PF|Y
C0037355|T121|sh85123618|LCH_NW|Smallpox vaccine||P|VC|N
C0037355|T129|sh85123618|LCH_NW|Smallpox vaccine||P|VC|N
C0037355|T121|40157|MEDCIN|smallpox vaccine||P|VC|N
C0037355|T129|40157|MEDCIN|smallpox vaccine||P|VC|N
C0037355|T121|40157|MEDCIN|smallpox vaccine (medication)||S|PF|Y
C0037355|T129|40157|MEDCIN|smallpox vaccine (medication)||S|PF|Y
C0037355|T121|40157|MEDCIN|vaccines viral smallpox||S|PF|Y
C0037355|T129|40157|MEDCIN|vaccines viral smallpox||S|PF|Y
C0037355|T121|d04831|MMSL|smallpox vaccine||P|VC|Y
C0037355|T129|d04831|MMSL|smallpox vaccine||P|VC|Y
C0037355|T121|D012900|MSH|Smallpox Vaccine||P|PF|N
C0037355|T129|D012900|MSH|Smallpox Vaccine||P|PF|N
C0037355|T121|D012900|MSH|Vaccine, Smallpox||P|VW|Y
C0037355|T129|D012900|MSH|Vaccine, Smallpox||P|VW|Y
C0037355|T121|NOCODE|MTH|Smallpox Vaccine||P|PF|Y
C0037355|T129|NOCODE|MTH|Smallpox Vaccine||P|PF|Y
C0037355|T121|N0000010563|NDFRT|Smallpox Vaccine||P|PF|N
C0037355|T129|N0000010563|NDFRT|Smallpox Vaccine||P|PF|N
C0037355|T121|N0000010563|NDFRT|Smallpox Vaccine [Chemical/Ingredient]||S|PF|Y
C0037355|T129|N0000010563|NDFRT|Smallpox Vaccine [Chemical/Ingredient]||S|PF|Y
C0037355|T121|N0000023075|NDFRT|SMALLPOX VACCINE||P|VC|N
C0037355|T129|N0000023075|NDFRT|SMALLPOX VACCINE||P|VC|N
C0037355|T121|9835|RXNORM|Smallpox Vaccine||P|PF|N
C0037355|T129|9835|RXNORM|Smallpox Vaccine||P|PF|N
C0037355|T121|33234009|SNOMEDCT_US|Smallpox vaccine||P|VC|Y
C0037355|T129|33234009|SNOMEDCT_US|Smallpox vaccine||P|VC|Y
C0037355|T121|33234009|SNOMEDCT_US|Smallpox vaccine (product)||S|PF|Y
C0037355|T129|33234009|SNOMEDCT_US|Smallpox vaccine (product)||S|PF|Y
C0037355|T121|33234009|SNOMEDCT_US|Smallpox vaccine (substance)||S|PF|N
C0037355|T129|33234009|SNOMEDCT_US|Smallpox vaccine (substance)||S|PF|N
C0037355|T121|33234009|SNOMEDCT_US|Var/Vac||S|PF|Y
C0037355|T129|33234009|SNOMEDCT_US|Var/Vac||S|PF|Y
C0037355|T121|396439006|SNOMEDCT_US|Smallpox vaccine||P|VC|N
C0037355|T129|396439006|SNOMEDCT_US|Smallpox vaccine||P|VC|N
C0037355|T121|396439006|SNOMEDCT_US|Smallpox vaccine (substance)||S|PF|Y
C0037355|T129|396439006|SNOMEDCT_US|Smallpox vaccine (substance)||S|PF|Y
C0037355|T121|396439006|SNOMEDCT_US|Var/Vac||S|PF|N
C0037355|T129|396439006|SNOMEDCT_US|Var/Vac||S|PF|N
C0037355|T121|4021502|VANDF|SMALLPOX VACCINE||P|VC|Y
C0037355|T129|4021502|VANDF|SMALLPOX VACCINE||P|VC|Y
C0051981|T121|65|CVX|leprosy||S|PF|N
C0051981|T129|65|CVX|leprosy||S|PF|N
C0051981|T121|65|CVX|leprosy vaccine||S|PF|Y
C0051981|T129|65|CVX|leprosy vaccine||S|PF|Y
C0051981|T121|65|HL7V2.5|leprosy||S|PF|N
C0051981|T129|65|HL7V2.5|leprosy||S|PF|N
C0051981|T121|65|HL7V3.0|leprosy||S|PF|Y
C0051981|T129|65|HL7V3.0|leprosy||S|PF|Y
C0051981|T121|5360|MEDLINEPLUS|Leprosy||S|VC|Y
C0051981|T129|5360|MEDLINEPLUS|Leprosy||S|VC|Y
C0051981|T121|C060596|MSH|anti-leprosy vaccine||P|PF|N
C0051981|T129|C060596|MSH|anti-leprosy vaccine||P|PF|N
C0051981|T121|C060596|MSH|antileprosy vaccine||S|PF|Y
C0051981|T129|C060596|MSH|antileprosy vaccine||S|PF|Y
C0051981|T121|NOCODE|MTH|anti-leprosy vaccine||P|PF|Y
C0051981|T129|NOCODE|MTH|anti-leprosy vaccine||P|PF|Y
C0062525|T116|90371|CPT|Human hepatitis B immune globulin||S|VCW|Y
C0062525|T129|90371|CPT|Human hepatitis B immune globulin||S|VCW|Y
C0062525|T121|90371|CPT|Human hepatitis B immune globulin||S|VCW|Y
C0062525|T116|30|CVX|HBIG||S|PF|N
C0062525|T129|30|CVX|HBIG||S|PF|N
C0062525|T121|30|CVX|HBIG||S|PF|N
C0062525|T116|30|CVX|hepatitis B immune globulin||P|PF|N
C0062525|T129|30|CVX|hepatitis B immune globulin||P|PF|N
C0062525|T121|30|CVX|hepatitis B immune globulin||P|PF|N
C0062525|T116|30|HL7V2.5|HBIG||S|PF|N
C0062525|T129|30|HL7V2.5|HBIG||S|PF|N
C0062525|T121|30|HL7V2.5|HBIG||S|PF|N
C0062525|T116|30|HL7V3.0|HBIG||S|PF|N
C0062525|T129|30|HL7V3.0|HBIG||S|PF|N
C0062525|T121|30|HL7V3.0|HBIG||S|PF|N
C0062525|T116|133255|MEDCIN|globulin, hepatitis B immune (human) for intramuscular use||S|VW|Y
C0062525|T129|133255|MEDCIN|globulin, hepatitis B immune (human) for intramuscular use||S|VW|Y
C0062525|T121|133255|MEDCIN|globulin, hepatitis B immune (human) for intramuscular use||S|VW|Y
C0062525|T116|133255|MEDCIN|human hepatitis B immune globulin for intramuscular use||S|PF|Y
C0062525|T129|133255|MEDCIN|human hepatitis B immune globulin for intramuscular use||S|PF|Y
C0062525|T121|133255|MEDCIN|human hepatitis B immune globulin for intramuscular use||S|PF|Y
C0062525|T116|133255|MEDCIN|human hepatitis B immune globulin for intramuscular use (medication)||S|PF|Y
C0062525|T129|133255|MEDCIN|human hepatitis B immune globulin for intramuscular use (medication)||S|PF|Y
C0062525|T121|133255|MEDCIN|human hepatitis B immune globulin for intramuscular use (medication)||S|PF|Y
C0062525|T116|48433|MEDCIN|globulin, hepatitis B immune (human)||S|VCW|Y
C0062525|T129|48433|MEDCIN|globulin, hepatitis B immune (human)||S|VCW|Y
C0062525|T121|48433|MEDCIN|globulin, hepatitis B immune (human)||S|VCW|Y
C0062525|T116|48433|MEDCIN|human hepatitis B immune globulin||S|VCW|Y
C0062525|T129|48433|MEDCIN|human hepatitis B immune globulin||S|VCW|Y
C0062525|T121|48433|MEDCIN|human hepatitis B immune globulin||S|VCW|Y
C0062525|T116|48433|MEDCIN|human hepatitis B immune globulin (medication)||S|PF|Y
C0062525|T129|48433|MEDCIN|human hepatitis B immune globulin (medication)||S|PF|Y
C0062525|T121|48433|MEDCIN|human hepatitis B immune globulin (medication)||S|PF|Y
C0062525|T116|7404|MMSL|hepatitis B immune globulin||P|PF|N
C0062525|T129|7404|MMSL|hepatitis B immune globulin||P|PF|N
C0062525|T121|7404|MMSL|hepatitis B immune globulin||P|PF|N
C0062525|T116|d01136|MMSL|hepatitis B immune globulin||P|PF|N
C0062525|T129|d01136|MMSL|hepatitis B immune globulin||P|PF|N
C0062525|T121|d01136|MMSL|hepatitis B immune globulin||P|PF|N
C0062525|T116|C045213|MSH|HBIG||S|PF|N
C0062525|T129|C045213|MSH|HBIG||S|PF|N
C0062525|T121|C045213|MSH|HBIG||S|PF|N
C0062525|T116|C045213|MSH|hepatitis B hyperimmune globulin||S|PF|Y
C0062525|T129|C045213|MSH|hepatitis B hyperimmune globulin||S|PF|Y
C0062525|T121|C045213|MSH|hepatitis B hyperimmune globulin||S|PF|Y
C0062525|T116|NOCODE|MTH|hepatitis B immune globulin||P|PF|Y
C0062525|T129|NOCODE|MTH|hepatitis B immune globulin||P|PF|Y
C0062525|T121|NOCODE|MTH|hepatitis B immune globulin||P|PF|Y
C0062525|T116|XII270YC6M|MTHSPL|HUMAN HEPATITIS B VIRUS IMMUNE GLOBULIN||S|PF|Y
C0062525|T116|XII270YC6M|MTHSPL|Human Hepatitis B Virus Immune Globulin||S|VC|Y
C0062525|T129|XII270YC6M|MTHSPL|HUMAN HEPATITIS B VIRUS IMMUNE GLOBULIN||S|PF|Y
C0062525|T129|XII270YC6M|MTHSPL|Human Hepatitis B Virus Immune Globulin||S|VC|Y
C0062525|T121|XII270YC6M|MTHSPL|HUMAN HEPATITIS B VIRUS IMMUNE GLOBULIN||S|PF|Y
C0062525|T121|XII270YC6M|MTHSPL|Human Hepatitis B Virus Immune Globulin||S|VC|Y
C0062525|T116|C80827|NCI|Human Hepatitis B Virus Immune Globulin||S|VC|N
C0062525|T129|C80827|NCI|Human Hepatitis B Virus Immune Globulin||S|VC|N
C0062525|T121|C80827|NCI|Human Hepatitis B Virus Immune Globulin||S|VC|N
C0062525|T116|XII270YC6M|NCI_FDA|HUMAN HEPATITIS B VIRUS IMMUNE GLOBULIN||S|PF|N
C0062525|T129|XII270YC6M|NCI_FDA|HUMAN HEPATITIS B VIRUS IMMUNE GLOBULIN||S|PF|N
C0062525|T121|XII270YC6M|NCI_FDA|HUMAN HEPATITIS B VIRUS IMMUNE GLOBULIN||S|PF|N
C0062525|T116|N0000146326|NDFRT|HEPATITIS B IMMUNE GLOBULIN||P|VC|N
C0062525|T129|N0000146326|NDFRT|HEPATITIS B IMMUNE GLOBULIN||P|VC|N
C0062525|T121|N0000146326|NDFRT|HEPATITIS B IMMUNE GLOBULIN||P|VC|N
C0062525|T116|N0000146328|NDFRT|HEPATITIS B IMMUNE GLOBULIN,HUMAN||S|VC|N
C0062525|T129|N0000146328|NDFRT|HEPATITIS B IMMUNE GLOBULIN,HUMAN||S|VC|N
C0062525|T121|N0000146328|NDFRT|HEPATITIS B IMMUNE GLOBULIN,HUMAN||S|VC|N
C0062525|T116|N0000179149|NDFRT|HBIG||S|PF|N
C0062525|T129|N0000179149|NDFRT|HBIG||S|PF|N
C0062525|T121|N0000179149|NDFRT|HBIG||S|PF|N
C0062525|T116|N0000179149|NDFRT|hepatitis B hyperimmune globulin||S|PF|N
C0062525|T129|N0000179149|NDFRT|hepatitis B hyperimmune globulin||S|PF|N
C0062525|T121|N0000179149|NDFRT|hepatitis B hyperimmune globulin||S|PF|N
C0062525|T116|N0000179149|NDFRT|hepatitis B hyperimmune globulin [Chemical/Ingredient]||S|PF|Y
C0062525|T129|N0000179149|NDFRT|hepatitis B hyperimmune globulin [Chemical/Ingredient]||S|PF|Y
C0062525|T121|N0000179149|NDFRT|hepatitis B hyperimmune globulin [Chemical/Ingredient]||S|PF|Y
C0062525|T116|26744|RXNORM|hepatitis B immune globulin||P|PF|N
C0062525|T129|26744|RXNORM|hepatitis B immune globulin||P|PF|N
C0062525|T121|26744|RXNORM|hepatitis B immune globulin||P|PF|N
C0062525|T116|170456004|SNOMEDCT_US|Anti-Hepatitis B immunoglob.||S|PF|Y
C0062525|T129|170456004|SNOMEDCT_US|Anti-Hepatitis B immunoglob.||S|PF|Y
C0062525|T121|170456004|SNOMEDCT_US|Anti-Hepatitis B immunoglob.||S|PF|Y
C0062525|T116|275846008|SNOMEDCT_US|Hepatitis B immunoglobulin||S|PF|N
C0062525|T129|275846008|SNOMEDCT_US|Hepatitis B immunoglobulin||S|PF|N
C0062525|T121|275846008|SNOMEDCT_US|Hepatitis B immunoglobulin||S|PF|N
C0062525|T116|275846008|SNOMEDCT_US|Hepatitis B immunoglobulin (substance)||S|PF|Y
C0062525|T129|275846008|SNOMEDCT_US|Hepatitis B immunoglobulin (substance)||S|PF|Y
C0062525|T121|275846008|SNOMEDCT_US|Hepatitis B immunoglobulin (substance)||S|PF|Y
C0062525|T116|9542007|SNOMEDCT_US|Antihepatitis B immunoglobulin||S|PF|Y
C0062525|T129|9542007|SNOMEDCT_US|Antihepatitis B immunoglobulin||S|PF|Y
C0062525|T121|9542007|SNOMEDCT_US|Antihepatitis B immunoglobulin||S|PF|Y
C0062525|T116|9542007|SNOMEDCT_US|HBIG||S|PF|Y
C0062525|T129|9542007|SNOMEDCT_US|HBIG||S|PF|Y
C0062525|T121|9542007|SNOMEDCT_US|HBIG||S|PF|Y
C0062525|T116|9542007|SNOMEDCT_US|Hepatitis B immune globulin (human)||S|PF|Y
C0062525|T129|9542007|SNOMEDCT_US|Hepatitis B immune globulin (human)||S|PF|Y
C0062525|T121|9542007|SNOMEDCT_US|Hepatitis B immune globulin (human)||S|PF|Y
C0062525|T116|9542007|SNOMEDCT_US|Hepatitis B immune globulin (human) (product)||S|PF|Y
C0062525|T129|9542007|SNOMEDCT_US|Hepatitis B immune globulin (human) (product)||S|PF|Y
C0062525|T121|9542007|SNOMEDCT_US|Hepatitis B immune globulin (human) (product)||S|PF|Y
C0062525|T116|9542007|SNOMEDCT_US|Hepatitis B immune globulin (human) (substance)||S|PF|Y
C0062525|T129|9542007|SNOMEDCT_US|Hepatitis B immune globulin (human) (substance)||S|PF|Y
C0062525|T121|9542007|SNOMEDCT_US|Hepatitis B immune globulin (human) (substance)||S|PF|Y
C0062525|T116|9542007|SNOMEDCT_US|Hepatitis B immunoglobulin||S|PF|Y
C0062525|T129|9542007|SNOMEDCT_US|Hepatitis B immunoglobulin||S|PF|Y
C0062525|T121|9542007|SNOMEDCT_US|Hepatitis B immunoglobulin||S|PF|Y
C0062525|T116|4017979|VANDF|HEPATITIS B IMMUNE GLOBULIN||P|VC|Y
C0062525|T129|4017979|VANDF|HEPATITIS B IMMUNE GLOBULIN||P|VC|Y
C0062525|T121|4017979|VANDF|HEPATITIS B IMMUNE GLOBULIN||P|VC|Y
C0062525|T116|4017981|VANDF|HEPATITIS B IMMUNE GLOBULIN,HUMAN||S|VC|Y
C0062525|T129|4017981|VANDF|HEPATITIS B IMMUNE GLOBULIN,HUMAN||S|VC|Y
C0062525|T121|4017981|VANDF|HEPATITIS B IMMUNE GLOBULIN,HUMAN||S|VC|Y
C0065828|T121|90707|CPT|Live measles, mumps and rubella virus vaccine||S|VO|Y
C0065828|T129|90707|CPT|Live measles, mumps and rubella virus vaccine||S|VO|Y
C0065828|T121|03|CVX|measles, mumps and rubella virus vaccine||S|VO|Y
C0065828|T129|03|CVX|measles, mumps and rubella virus vaccine||S|VO|Y
C0065828|T121|03|CVX|MMR||S|PF|N
C0065828|T129|03|CVX|MMR||S|PF|N
C0065828|T121|03|HL7V2.5|MMR||S|PF|N
C0065828|T129|03|HL7V2.5|MMR||S|PF|N
C0065828|T121|3|HL7V3.0|MMR||S|PF|N
C0065828|T129|3|HL7V3.0|MMR||S|PF|N
C0065828|T121|sh2005000940|LCH_NW|MMR vaccine||S|VC|N
C0065828|T129|sh2005000940|LCH_NW|MMR vaccine||S|VC|N
C0065828|T121|d03007|MMSL|measles/mumps/rubella virus vaccine||S|PF|Y
C0065828|T129|d03007|MMSL|measles/mumps/rubella virus vaccine||S|PF|Y
C0065828|T121|D022542|MSH|Measles Mumps Rubella Vaccine||P|VO|N
C0065828|T129|D022542|MSH|Measles Mumps Rubella Vaccine||P|VO|N
C0065828|T121|D022542|MSH|Measles-Mumps-Rubella Vaccine||P|PF|N
C0065828|T129|D022542|MSH|Measles-Mumps-Rubella Vaccine||P|PF|N
C0065828|T121|D022542|MSH|Measles, Mumps, Rubella Vaccine||P|VO|Y
C0065828|T129|D022542|MSH|Measles, Mumps, Rubella Vaccine||P|VO|Y
C0065828|T121|D022542|MSH|MMR Vaccine||S|PF|Y
C0065828|T129|D022542|MSH|MMR Vaccine||S|PF|Y
C0065828|T121|D022542|MSH|Mumps Measles Rubella Vaccine||P|VW|Y
C0065828|T129|D022542|MSH|Mumps Measles Rubella Vaccine||P|VW|Y
C0065828|T121|D022542|MSH|Mumps-Measles-Rubella Vaccine||P|VW|Y
C0065828|T129|D022542|MSH|Mumps-Measles-Rubella Vaccine||P|VW|Y
C0065828|T121|D022542|MSH|Vaccine, Measles-Mumps-Rubella||P|VW|Y
C0065828|T129|D022542|MSH|Vaccine, Measles-Mumps-Rubella||P|VW|Y
C0065828|T121|D022542|MSH|Vaccine, MMR||S|VW|Y
C0065828|T129|D022542|MSH|Vaccine, MMR||S|VW|Y
C0065828|T121|D022542|MSH|Vaccine, Mumps-Measles-Rubella||P|VW|Y
C0065828|T129|D022542|MSH|Vaccine, Mumps-Measles-Rubella||P|VW|Y
C0065828|T121|NOCODE|MTH|Measles-Mumps-Rubella Vaccine||P|PF|Y
C0065828|T129|NOCODE|MTH|Measles-Mumps-Rubella Vaccine||P|PF|Y
C0065828|T121|C96403|NCI|M-M-R II||S|PF|Y
C0065828|T129|C96403|NCI|M-M-R II||S|PF|Y
C0065828|T121|C96403|NCI|Measles Mumps Rubella Vaccine||P|VO|Y
C0065828|T129|C96403|NCI|Measles Mumps Rubella Vaccine||P|VO|Y
C0065828|T121|C96403|NCI|Measles, Mumps and Rubella Virus Vaccine, Live||S|VO|Y
C0065828|T129|C96403|NCI|Measles, Mumps and Rubella Virus Vaccine, Live||S|VO|Y
C0065828|T121|C96403|NCI|Measles, Mumps, and Rubella Vaccine||P|VO|Y
C0065828|T129|C96403|NCI|Measles, Mumps, and Rubella Vaccine||P|VO|Y
C0065828|T121|C96403|NCI|Measles/Mumps/Rubella Vaccine||P|VO|Y
C0065828|T129|C96403|NCI|Measles/Mumps/Rubella Vaccine||P|VO|Y
C0065828|T121|C96403|NCI|MMR Vaccine||S|PF|N
C0065828|T129|C96403|NCI|MMR Vaccine||S|PF|N
C0065828|T121|C96403|NCI_NICHD|Measles Mumps Rubella Vaccine||P|VO|N
C0065828|T129|C96403|NCI_NICHD|Measles Mumps Rubella Vaccine||P|VO|N
C0065828|T121|C96403|NCI_NICHD|Measles/Mumps/Rubella Vaccine||P|VO|N
C0065828|T129|C96403|NCI_NICHD|Measles/Mumps/Rubella Vaccine||P|VO|N
C0065828|T121|C96403|NCI_NICHD|MMR||S|PF|Y
C0065828|T129|C96403|NCI_NICHD|MMR||S|PF|Y
C0065828|T121|N0000022440|NDFRT|MEASLES/MUMPS/RUBELLA VIRUS VACCINE,LIVE||S|PF|N
C0065828|T129|N0000022440|NDFRT|MEASLES/MUMPS/RUBELLA VIRUS VACCINE,LIVE||S|PF|N
C0065828|T121|N0000170911|NDFRT|Measles-Mumps-Rubella Vaccine||P|PF|N
C0065828|T129|N0000170911|NDFRT|Measles-Mumps-Rubella Vaccine||P|PF|N
C0065828|T121|N0000170911|NDFRT|Measles-Mumps-Rubella Vaccine [Chemical/Ingredient]||S|PF|Y
C0065828|T129|N0000170911|NDFRT|Measles-Mumps-Rubella Vaccine [Chemical/Ingredient]||S|PF|Y
C0065828|T121|N0000170911|NDFRT|Measles, Mumps, Rubella Vaccine||P|VO|N
C0065828|T129|N0000170911|NDFRT|Measles, Mumps, Rubella Vaccine||P|VO|N
C0065828|T121|N0000170911|NDFRT|MMR Vaccine||S|PF|N
C0065828|T129|N0000170911|NDFRT|MMR Vaccine||S|PF|N
C0065828|T121|N0000170911|NDFRT|Mumps-Measles-Rubella Vaccine||P|VW|N
C0065828|T129|N0000170911|NDFRT|Mumps-Measles-Rubella Vaccine||P|VW|N
C0065828|T121|396429000|SNOMEDCT_US|Measles, mumps and rubella vaccine||P|VO|Y
C0065828|T129|396429000|SNOMEDCT_US|Measles, mumps and rubella vaccine||P|VO|Y
C0065828|T121|396429000|SNOMEDCT_US|Measles, mumps and rubella vaccine (substance)||S|PF|Y
C0065828|T129|396429000|SNOMEDCT_US|Measles, mumps and rubella vaccine (substance)||S|PF|Y
C0065828|T121|396429000|SNOMEDCT_US|MMR vaccine||S|VC|Y
C0065828|T129|396429000|SNOMEDCT_US|MMR vaccine||S|VC|Y
C0065828|T121|61153008|SNOMEDCT_US|Measles + Mumps + Rubella vaccine||P|VC|Y
C0065828|T129|61153008|SNOMEDCT_US|Measles + Mumps + Rubella vaccine||P|VC|Y
C0065828|T121|61153008|SNOMEDCT_US|Measles, mumps and rubella vaccine||P|VO|N
C0065828|T129|61153008|SNOMEDCT_US|Measles, mumps and rubella vaccine||P|VO|N
C0065828|T121|61153008|SNOMEDCT_US|Measles, mumps and rubella vaccine (product)||S|PF|Y
C0065828|T129|61153008|SNOMEDCT_US|Measles, mumps and rubella vaccine (product)||S|PF|Y
C0065828|T121|61153008|SNOMEDCT_US|Measles, mumps and rubella vaccine (substance)||S|PF|N
C0065828|T129|61153008|SNOMEDCT_US|Measles, mumps and rubella vaccine (substance)||S|PF|N
C0065828|T121|61153008|SNOMEDCT_US|Measles/mumps/rubella vaccine||P|VC|Y
C0065828|T129|61153008|SNOMEDCT_US|Measles/mumps/rubella vaccine||P|VC|Y
C0065828|T121|4017978|VANDF|MEASLES/MUMPS/RUBELLA VIRUS VACCINE,LIVE||S|PF|Y
C0065828|T129|4017978|VANDF|MEASLES/MUMPS/RUBELLA VIRUS VACCINE,LIVE||S|PF|Y
C0065829|T121|94|CVX|measles, mumps, rubella, and varicella virus vaccine||S|VO|Y
C0065829|T129|94|CVX|measles, mumps, rubella, and varicella virus vaccine||S|VO|Y
C0065829|T121|94|CVX|MMRV||S|PF|N
C0065829|T129|94|CVX|MMRV||S|PF|N
C0065829|T121|94|HL7V2.5|MMRV||S|PF|N
C0065829|T129|94|HL7V2.5|MMRV||S|PF|N
C0065829|T121|94|HL7V3.0|MMRV||S|PF|Y
C0065829|T129|94|HL7V3.0|MMRV||S|PF|Y
C0065829|T121|d05645|MMSL|measles/mumps/rubella/varicella virus vaccine||S|PF|Y
C0065829|T129|d05645|MMSL|measles/mumps/rubella/varicella virus vaccine||S|PF|Y
C0065829|T121|C050102|MSH|measles, mumps, rubella, varicella vaccine||P|PF|Y
C0065829|T129|C050102|MSH|measles, mumps, rubella, varicella vaccine||P|PF|Y
C0065829|T121|C050102|MSH|MMRV vaccine||S|PF|Y
C0065829|T129|C050102|MSH|MMRV vaccine||S|PF|Y
C0065829|T121|419550004|SNOMEDCT_US|Measles + mumps + rubella + varicella vaccine||P|VC|Y
C0065829|T129|419550004|SNOMEDCT_US|Measles + mumps + rubella + varicella vaccine||P|VC|Y
C0065829|T121|419550004|SNOMEDCT_US|Measles + mumps + rubella + varicella vaccine (product)||S|PF|Y
C0065829|T129|419550004|SNOMEDCT_US|Measles + mumps + rubella + varicella vaccine (product)||S|PF|Y
C0078048|T121|21|CVX|varicella||S|PF|N
C0078048|T129|21|CVX|varicella||S|PF|N
C0078048|T121|21|CVX|varicella virus vaccine||S|VC|N
C0078048|T129|21|CVX|varicella virus vaccine||S|VC|N
C0078048|T121|21|HL7V2.5|Varicella||S|VC|Y
C0078048|T129|21|HL7V2.5|Varicella||S|VC|Y
C0078048|T121|21|HL7V3.0|varicella||S|PF|Y
C0078048|T129|21|HL7V3.0|varicella||S|PF|Y
C0078048|T121|d03832|MMSL|varicella virus vaccine||S|VC|Y
C0078048|T129|d03832|MMSL|varicella virus vaccine||S|VC|Y
C0078048|T121|D019433|MSH|Chickenpox Vaccine||P|PF|N
C0078048|T129|D019433|MSH|Chickenpox Vaccine||P|PF|N
C0078048|T121|D019433|MSH|Oka Varicella Vaccine||S|PF|Y
C0078048|T129|D019433|MSH|Oka Varicella Vaccine||S|PF|Y
C0078048|T121|D019433|MSH|Vaccine, Chickenpox||P|VW|Y
C0078048|T129|D019433|MSH|Vaccine, Chickenpox||P|VW|Y
C0078048|T121|D019433|MSH|Vaccine, Oka Varicella||S|VW|Y
C0078048|T129|D019433|MSH|Vaccine, Oka Varicella||S|VW|Y
C0078048|T121|D019433|MSH|Vaccine, Varicella||S|VW|Y
C0078048|T129|D019433|MSH|Vaccine, Varicella||S|VW|Y
C0078048|T121|D019433|MSH|Varicella Vaccine||S|PF|Y
C0078048|T129|D019433|MSH|Varicella Vaccine||S|PF|Y
C0078048|T121|D019433|MSH|Varicella Vaccine, Oka||S|VW|Y
C0078048|T129|D019433|MSH|Varicella Vaccine, Oka||S|VW|Y
C0078048|T121|NOCODE|MTH|Chickenpox Vaccine||P|PF|Y
C0078048|T129|NOCODE|MTH|Chickenpox Vaccine||P|PF|Y
C0078048|T121|N0000170905|NDFRT|Chickenpox Vaccine||P|PF|N
C0078048|T129|N0000170905|NDFRT|Chickenpox Vaccine||P|PF|N
C0078048|T121|N0000170905|NDFRT|Chickenpox Vaccine [Chemical/Ingredient]||S|PF|Y
C0078048|T129|N0000170905|NDFRT|Chickenpox Vaccine [Chemical/Ingredient]||S|PF|Y
C0078048|T121|N0000170905|NDFRT|Oka Varicella Vaccine||S|PF|N
C0078048|T129|N0000170905|NDFRT|Oka Varicella Vaccine||S|PF|N
C0078048|T121|N0000170905|NDFRT|Varicella Vaccine||S|PF|N
C0078048|T129|N0000170905|NDFRT|Varicella Vaccine||S|PF|N
C0078048|T121|108729007|SNOMEDCT_US|Varicella vaccine||S|VC|Y
C0078048|T129|108729007|SNOMEDCT_US|Varicella vaccine||S|VC|Y
C0078048|T121|108729007|SNOMEDCT_US|Varicella virus vaccine||S|PF|Y
C0078048|T129|108729007|SNOMEDCT_US|Varicella virus vaccine||S|PF|Y
C0078048|T121|108729007|SNOMEDCT_US|Varicella virus vaccine (product)||S|PF|Y
C0078048|T129|108729007|SNOMEDCT_US|Varicella virus vaccine (product)||S|PF|Y
C0078048|T121|108729007|SNOMEDCT_US|Varicella virus vaccine (substance)||S|PF|N
C0078048|T129|108729007|SNOMEDCT_US|Varicella virus vaccine (substance)||S|PF|N
C0078048|T121|396442000|SNOMEDCT_US|Varicella virus vaccine||S|PF|N
C0078048|T129|396442000|SNOMEDCT_US|Varicella virus vaccine||S|PF|N
C0078048|T121|396442000|SNOMEDCT_US|Varicella virus vaccine (substance)||S|PF|Y
C0078048|T129|396442000|SNOMEDCT_US|Varicella virus vaccine (substance)||S|PF|Y
C0078049|T121|90396|CPT|Human varicella-zoster immune globulin||S|VC|Y
C0078049|T116|90396|CPT|Human varicella-zoster immune globulin||S|VC|Y
C0078049|T129|90396|CPT|Human varicella-zoster immune globulin||S|VC|Y
C0078049|T121|36|CVX|varicella zoster immune globulin||P|VO|N
C0078049|T116|36|CVX|varicella zoster immune globulin||P|VO|N
C0078049|T129|36|CVX|varicella zoster immune globulin||P|VO|N
C0078049|T121|36|CVX|VZIG||S|PF|N
C0078049|T116|36|CVX|VZIG||S|PF|N
C0078049|T129|36|CVX|VZIG||S|PF|N
C0078049|T121|36|HL7V2.5|VZIG||S|PF|N
C0078049|T116|36|HL7V2.5|VZIG||S|PF|N
C0078049|T129|36|HL7V2.5|VZIG||S|PF|N
C0078049|T121|36|HL7V3.0|VZIG||S|PF|N
C0078049|T116|36|HL7V3.0|VZIG||S|PF|N
C0078049|T129|36|HL7V3.0|VZIG||S|PF|N
C0078049|T121|3142|MMSL|Varicella Zoster Immune Globulin||P|VC|Y
C0078049|T116|3142|MMSL|Varicella Zoster Immune Globulin||P|VC|Y
C0078049|T129|3142|MMSL|Varicella Zoster Immune Globulin||P|VC|Y
C0078049|T121|5666|MMSL|varicella-zoster immune globulin||P|PF|N
C0078049|T116|5666|MMSL|varicella-zoster immune globulin||P|PF|N
C0078049|T129|5666|MMSL|varicella-zoster immune globulin||P|PF|N
C0078049|T121|d01138|MMSL|varicella zoster immune globulin||P|VO|Y
C0078049|T116|d01138|MMSL|varicella zoster immune globulin||P|VO|Y
C0078049|T129|d01138|MMSL|varicella zoster immune globulin||P|VO|Y
C0078049|T121|C030799|MSH|varicella-zoster immune globulin||P|PF|N
C0078049|T116|C030799|MSH|varicella-zoster immune globulin||P|PF|N
C0078049|T129|C030799|MSH|varicella-zoster immune globulin||P|PF|N
C0078049|T121|C030799|MSH|varicellon||S|PF|Y
C0078049|T116|C030799|MSH|varicellon||S|PF|Y
C0078049|T129|C030799|MSH|varicellon||S|PF|Y
C0078049|T121|C030799|MSH|VZIG||S|PF|N
C0078049|T116|C030799|MSH|VZIG||S|PF|N
C0078049|T129|C030799|MSH|VZIG||S|PF|N
C0078049|T121|NOCODE|MTH|varicella-zoster immune globulin||P|PF|Y
C0078049|T116|NOCODE|MTH|varicella-zoster immune globulin||P|PF|Y
C0078049|T129|NOCODE|MTH|varicella-zoster immune globulin||P|PF|Y
C0078049|T121|33T61IWL27|MTHSPL|HUMAN VARICELLA-ZOSTER IMMUNE GLOBULIN||S|PF|Y
C0078049|T116|33T61IWL27|MTHSPL|HUMAN VARICELLA-ZOSTER IMMUNE GLOBULIN||S|PF|Y
C0078049|T129|33T61IWL27|MTHSPL|HUMAN VARICELLA-ZOSTER IMMUNE GLOBULIN||S|PF|Y
C0078049|T121|C123431|NCI|Human Varicella Zoster Immune Globulin||S|VC|Y
C0078049|T116|C123431|NCI|Human Varicella Zoster Immune Globulin||S|VC|Y
C0078049|T129|C123431|NCI|Human Varicella Zoster Immune Globulin||S|VC|Y
C0078049|T121|C123431|NCI|Human Varicella-Zoster Immune Globulin||S|VC|Y
C0078049|T116|C123431|NCI|Human Varicella-Zoster Immune Globulin||S|VC|Y
C0078049|T129|C123431|NCI|Human Varicella-Zoster Immune Globulin||S|VC|Y
C0078049|T121|C123431|NCI|Varicella Zoster Immune Globulin Human||S|VCW|Y
C0078049|T116|C123431|NCI|Varicella Zoster Immune Globulin Human||S|VCW|Y
C0078049|T129|C123431|NCI|Varicella Zoster Immune Globulin Human||S|VCW|Y
C0078049|T121|C123431|NCI|VZIG Vaccine||S|PF|Y
C0078049|T116|C123431|NCI|VZIG Vaccine||S|PF|Y
C0078049|T129|C123431|NCI|VZIG Vaccine||S|PF|Y
C0078049|T121|33T61IWL27|NCI_FDA|HUMAN VARICELLA-ZOSTER IMMUNE GLOBULIN||S|PF|N
C0078049|T116|33T61IWL27|NCI_FDA|HUMAN VARICELLA-ZOSTER IMMUNE GLOBULIN||S|PF|N
C0078049|T129|33T61IWL27|NCI_FDA|HUMAN VARICELLA-ZOSTER IMMUNE GLOBULIN||S|PF|N
C0078049|T121|N0000020895|NDFRT|VARICELLA ZOSTER IMMUNE GLOBULIN||P|VC|N
C0078049|T116|N0000020895|NDFRT|VARICELLA ZOSTER IMMUNE GLOBULIN||P|VC|N
C0078049|T129|N0000020895|NDFRT|VARICELLA ZOSTER IMMUNE GLOBULIN||P|VC|N
C0078049|T121|N0000147358|NDFRT|VARICELLA ZOSTER IMMUNE GLOBULIN (HUMAN)||S|VW|N
C0078049|T116|N0000147358|NDFRT|VARICELLA ZOSTER IMMUNE GLOBULIN (HUMAN)||S|VW|N
C0078049|T129|N0000147358|NDFRT|VARICELLA ZOSTER IMMUNE GLOBULIN (HUMAN)||S|VW|N
C0078049|T121|N0000179279|NDFRT|varicella-zoster immune globulin||P|PF|N
C0078049|T116|N0000179279|NDFRT|varicella-zoster immune globulin||P|PF|N
C0078049|T129|N0000179279|NDFRT|varicella-zoster immune globulin||P|PF|N
C0078049|T121|N0000179279|NDFRT|varicella-zoster immune globulin [Chemical/Ingredient]||S|PF|Y
C0078049|T116|N0000179279|NDFRT|varicella-zoster immune globulin [Chemical/Ingredient]||S|PF|Y
C0078049|T129|N0000179279|NDFRT|varicella-zoster immune globulin [Chemical/Ingredient]||S|PF|Y
C0078049|T121|N0000179279|NDFRT|varicellon||S|PF|N
C0078049|T116|N0000179279|NDFRT|varicellon||S|PF|N
C0078049|T129|N0000179279|NDFRT|varicellon||S|PF|N
C0078049|T121|N0000179279|NDFRT|VZIG||S|PF|N
C0078049|T116|N0000179279|NDFRT|VZIG||S|PF|N
C0078049|T129|N0000179279|NDFRT|VZIG||S|PF|N
C0078049|T121|39385|RXNORM|varicella-zoster immune globulin||P|PF|N
C0078049|T116|39385|RXNORM|varicella-zoster immune globulin||P|PF|N
C0078049|T129|39385|RXNORM|varicella-zoster immune globulin||P|PF|N
C0078049|T121|147707008|SNOMEDCT_US|Anti-varic-Zoster immunoglob (& injection)||S|PF|N
C0078049|T116|147707008|SNOMEDCT_US|Anti-varic-Zoster immunoglob (& injection)||S|PF|N
C0078049|T129|147707008|SNOMEDCT_US|Anti-varic-Zoster immunoglob (& injection)||S|PF|N
C0078049|T121|147707008|SNOMEDCT_US|Anti-varic-Zoster immunoglob (& injection) (procedure)||S|PF|N
C0078049|T116|147707008|SNOMEDCT_US|Anti-varic-Zoster immunoglob (& injection) (procedure)||S|PF|N
C0078049|T129|147707008|SNOMEDCT_US|Anti-varic-Zoster immunoglob (& injection) (procedure)||S|PF|N
C0078049|T121|170455000|SNOMEDCT_US|Anti-varic-Zoster immunoglob||S|VO|Y
C0078049|T116|170455000|SNOMEDCT_US|Anti-varic-Zoster immunoglob||S|VO|Y
C0078049|T129|170455000|SNOMEDCT_US|Anti-varic-Zoster immunoglob||S|VO|Y
C0078049|T121|170455000|SNOMEDCT_US|Anti-varic-Zoster immunoglob (& injection)||S|PF|Y
C0078049|T121|170455000|SNOMEDCT_US|Anti-varic-Zoster immunoglob (& injection)||S|PF|N
C0078049|T116|170455000|SNOMEDCT_US|Anti-varic-Zoster immunoglob (& injection)||S|PF|Y
C0078049|T116|170455000|SNOMEDCT_US|Anti-varic-Zoster immunoglob (& injection)||S|PF|N
C0078049|T129|170455000|SNOMEDCT_US|Anti-varic-Zoster immunoglob (& injection)||S|PF|Y
C0078049|T129|170455000|SNOMEDCT_US|Anti-varic-Zoster immunoglob (& injection)||S|PF|N
C0078049|T121|170455000|SNOMEDCT_US|Anti-varic-Zoster immunoglob (& injection) (procedure)||S|PF|Y
C0078049|T116|170455000|SNOMEDCT_US|Anti-varic-Zoster immunoglob (& injection) (procedure)||S|PF|Y
C0078049|T129|170455000|SNOMEDCT_US|Anti-varic-Zoster immunoglob (& injection) (procedure)||S|PF|Y
C0078049|T121|170455000|SNOMEDCT_US|Anti-varic-Zoster immunoglob.||S|PF|Y
C0078049|T116|170455000|SNOMEDCT_US|Anti-varic-Zoster immunoglob.||S|PF|Y
C0078049|T129|170455000|SNOMEDCT_US|Anti-varic-Zoster immunoglob.||S|PF|Y
C0078049|T121|62294009|SNOMEDCT_US|Anti-varicella-zoster immunoglobulin||S|PF|Y
C0078049|T116|62294009|SNOMEDCT_US|Anti-varicella-zoster immunoglobulin||S|PF|Y
C0078049|T129|62294009|SNOMEDCT_US|Anti-varicella-zoster immunoglobulin||S|PF|Y
C0078049|T121|62294009|SNOMEDCT_US|Varicella immunoglobulin||S|PF|Y
C0078049|T116|62294009|SNOMEDCT_US|Varicella immunoglobulin||S|PF|Y
C0078049|T129|62294009|SNOMEDCT_US|Varicella immunoglobulin||S|PF|Y
C0078049|T121|62294009|SNOMEDCT_US|Varicella-zoster immune globulin||P|VC|Y
C0078049|T116|62294009|SNOMEDCT_US|Varicella-zoster immune globulin||P|VC|Y
C0078049|T129|62294009|SNOMEDCT_US|Varicella-zoster immune globulin||P|VC|Y
C0078049|T121|62294009|SNOMEDCT_US|Varicella-zoster immune globulin (product)||S|PF|Y
C0078049|T116|62294009|SNOMEDCT_US|Varicella-zoster immune globulin (product)||S|PF|Y
C0078049|T129|62294009|SNOMEDCT_US|Varicella-zoster immune globulin (product)||S|PF|Y
C0078049|T121|62294009|SNOMEDCT_US|Varicella-zoster immune globulin (substance)||S|PF|Y
C0078049|T116|62294009|SNOMEDCT_US|Varicella-zoster immune globulin (substance)||S|PF|Y
C0078049|T129|62294009|SNOMEDCT_US|Varicella-zoster immune globulin (substance)||S|PF|Y
C0078049|T121|62294009|SNOMEDCT_US|Varicella-zoster immunoglobulin||S|PF|Y
C0078049|T116|62294009|SNOMEDCT_US|Varicella-zoster immunoglobulin||S|PF|Y
C0078049|T129|62294009|SNOMEDCT_US|Varicella-zoster immunoglobulin||S|PF|Y
C0078049|T121|62294009|SNOMEDCT_US|VZIG||S|PF|Y
C0078049|T116|62294009|SNOMEDCT_US|VZIG||S|PF|Y
C0078049|T129|62294009|SNOMEDCT_US|VZIG||S|PF|Y
C0078049|T121|62294009|SNOMEDCT_US|ZIG - Zoster immune globulin||S|PF|Y
C0078049|T116|62294009|SNOMEDCT_US|ZIG - Zoster immune globulin||S|PF|Y
C0078049|T129|62294009|SNOMEDCT_US|ZIG - Zoster immune globulin||S|PF|Y
C0078049|T121|62294009|SNOMEDCT_US|Zoster immune globulin||S|PF|Y
C0078049|T116|62294009|SNOMEDCT_US|Zoster immune globulin||S|PF|Y
C0078049|T129|62294009|SNOMEDCT_US|Zoster immune globulin||S|PF|Y
C0078049|T121|4019100|VANDF|VARICELLA ZOSTER IMMUNE GLOBULIN (HUMAN)||S|VW|Y
C0078049|T116|4019100|VANDF|VARICELLA ZOSTER IMMUNE GLOBULIN (HUMAN)||S|VW|Y
C0078049|T129|4019100|VANDF|VARICELLA ZOSTER IMMUNE GLOBULIN (HUMAN)||S|VW|Y
C0078049|T121|4022890|VANDF|VARICELLA ZOSTER IMMUNE GLOBULIN||P|VC|Y
C0078049|T116|4022890|VANDF|VARICELLA ZOSTER IMMUNE GLOBULIN||P|VC|Y
C0078049|T129|4022890|VANDF|VARICELLA ZOSTER IMMUNE GLOBULIN||P|VC|Y
C0085297|T121|87|CVX|IGIV||S|PF|N
C0085297|T116|87|CVX|IGIV||S|PF|N
C0085297|T129|87|CVX|IGIV||S|PF|N
C0085297|T121|87|CVX|immune globulin, intravenous||S|VC|Y
C0085297|T116|87|CVX|immune globulin, intravenous||S|VC|Y
C0085297|T129|87|CVX|immune globulin, intravenous||S|VC|Y
C0085297|T121|87|HL7V2.5|IGIV||S|PF|N
C0085297|T116|87|HL7V2.5|IGIV||S|PF|N
C0085297|T129|87|HL7V2.5|IGIV||S|PF|N
C0085297|T121|87|HL7V3.0|IGIV||S|PF|Y
C0085297|T116|87|HL7V3.0|IGIV||S|PF|Y
C0085297|T129|87|HL7V3.0|IGIV||S|PF|Y
C0085297|T121|42500|MMSL|Immune Globulin, Intravenous||S|PF|N
C0085297|T116|42500|MMSL|Immune Globulin, Intravenous||S|PF|N
C0085297|T129|42500|MMSL|Immune Globulin, Intravenous||S|PF|N
C0085297|T121|d01133|MMSL|immune globulin intravenous||S|VC|Y
C0085297|T116|d01133|MMSL|immune globulin intravenous||S|VC|Y
C0085297|T129|d01133|MMSL|immune globulin intravenous||S|VC|Y
C0085297|T121|D016756|MSH|Antibodies, Intravenous||S|VW|Y
C0085297|T116|D016756|MSH|Antibodies, Intravenous||S|VW|Y
C0085297|T129|D016756|MSH|Antibodies, Intravenous||S|VW|Y
C0085297|T121|D016756|MSH|IG IV||S|PF|Y
C0085297|T116|D016756|MSH|IG IV||S|PF|Y
C0085297|T129|D016756|MSH|IG IV||S|PF|Y
C0085297|T121|D016756|MSH|IGIV||S|PF|N
C0085297|T116|D016756|MSH|IGIV||S|PF|N
C0085297|T129|D016756|MSH|IGIV||S|PF|N
C0085297|T121|D016756|MSH|Immune Globulin, Intravenous||S|PF|Y
C0085297|T116|D016756|MSH|Immune Globulin, Intravenous||S|PF|Y
C0085297|T129|D016756|MSH|Immune Globulin, Intravenous||S|PF|Y
C0085297|T121|D016756|MSH|Immunoglobulins, Intravenous||P|PF|N
C0085297|T116|D016756|MSH|Immunoglobulins, Intravenous||P|PF|N
C0085297|T129|D016756|MSH|Immunoglobulins, Intravenous||P|PF|N
C0085297|T121|D016756|MSH|Immunoglobulins, IV||S|VW|Y
C0085297|T116|D016756|MSH|Immunoglobulins, IV||S|VW|Y
C0085297|T129|D016756|MSH|Immunoglobulins, IV||S|VW|Y
C0085297|T121|D016756|MSH|Intravenous Antibodies||S|PF|Y
C0085297|T116|D016756|MSH|Intravenous Antibodies||S|PF|Y
C0085297|T129|D016756|MSH|Intravenous Antibodies||S|PF|Y
C0085297|T121|D016756|MSH|Intravenous IG||S|PF|Y
C0085297|T116|D016756|MSH|Intravenous IG||S|PF|Y
C0085297|T129|D016756|MSH|Intravenous IG||S|PF|Y
C0085297|T121|D016756|MSH|Intravenous Immune Globulin||S|VW|Y
C0085297|T116|D016756|MSH|Intravenous Immune Globulin||S|VW|Y
C0085297|T129|D016756|MSH|Intravenous Immune Globulin||S|VW|Y
C0085297|T121|D016756|MSH|Intravenous Immunoglobulins||P|VW|Y
C0085297|T116|D016756|MSH|Intravenous Immunoglobulins||P|VW|Y
C0085297|T129|D016756|MSH|Intravenous Immunoglobulins||P|VW|Y
C0085297|T121|D016756|MSH|IV IG||S|VW|Y
C0085297|T116|D016756|MSH|IV IG||S|VW|Y
C0085297|T129|D016756|MSH|IV IG||S|VW|Y
C0085297|T121|D016756|MSH|IV Immunoglobulins||S|PF|Y
C0085297|T116|D016756|MSH|IV Immunoglobulins||S|PF|Y
C0085297|T129|D016756|MSH|IV Immunoglobulins||S|PF|Y
C0085297|T121|D016756|MSH|IVIG||S|PF|Y
C0085297|T116|D016756|MSH|IVIG||S|PF|Y
C0085297|T129|D016756|MSH|IVIG||S|PF|Y
C0085297|T121|NOCODE|MTH|Immunoglobulins, Intravenous||P|PF|Y
C0085297|T116|NOCODE|MTH|Immunoglobulins, Intravenous||P|PF|Y
C0085297|T129|NOCODE|MTH|Immunoglobulins, Intravenous||P|PF|Y
C0085297|T121|C121331|NCI|Gamma Globulin Therapy||S|PF|Y
C0085297|T116|C121331|NCI|Gamma Globulin Therapy||S|PF|Y
C0085297|T129|C121331|NCI|Gamma Globulin Therapy||S|PF|Y
C0085297|T121|C121331|NCI|Immune Globulin Therapy||S|PF|Y
C0085297|T116|C121331|NCI|Immune Globulin Therapy||S|PF|Y
C0085297|T129|C121331|NCI|Immune Globulin Therapy||S|PF|Y
C0085297|T121|C121331|NCI|Intravenous Immunoglobulin Therapy||S|PF|Y
C0085297|T116|C121331|NCI|Intravenous Immunoglobulin Therapy||S|PF|Y
C0085297|T129|C121331|NCI|Intravenous Immunoglobulin Therapy||S|PF|Y
C0085297|T121|C121331|NCI|IVIG Therapy||S|PF|Y
C0085297|T116|C121331|NCI|IVIG Therapy||S|PF|Y
C0085297|T129|C121331|NCI|IVIG Therapy||S|PF|Y
C0085297|T121|C121331|NCI_NICHD|Gamma Globulin||S|PF|Y
C0085297|T116|C121331|NCI_NICHD|Gamma Globulin||S|PF|Y
C0085297|T129|C121331|NCI_NICHD|Gamma Globulin||S|PF|Y
C0085297|T121|C121331|NCI_NICHD|Immune Globulin||S|PF|Y
C0085297|T116|C121331|NCI_NICHD|Immune Globulin||S|PF|Y
C0085297|T129|C121331|NCI_NICHD|Immune Globulin||S|PF|Y
C0085297|T121|C121331|NCI_NICHD|Intravenous Immunoglobulin||P|VO|Y
C0085297|T116|C121331|NCI_NICHD|Intravenous Immunoglobulin||P|VO|Y
C0085297|T129|C121331|NCI_NICHD|Intravenous Immunoglobulin||P|VO|Y
C0085297|T121|C121331|NCI_NICHD|IVIG||S|PF|N
C0085297|T116|C121331|NCI_NICHD|IVIG||S|PF|N
C0085297|T129|C121331|NCI_NICHD|IVIG||S|PF|N
C0085297|T121|N0000007401|NDFRT|Antibodies, Intravenous||S|VW|N
C0085297|T116|N0000007401|NDFRT|Antibodies, Intravenous||S|VW|N
C0085297|T129|N0000007401|NDFRT|Antibodies, Intravenous||S|VW|N
C0085297|T121|N0000007401|NDFRT|Immune Globulin, Intravenous||S|PF|N
C0085297|T116|N0000007401|NDFRT|Immune Globulin, Intravenous||S|PF|N
C0085297|T129|N0000007401|NDFRT|Immune Globulin, Intravenous||S|PF|N
C0085297|T121|N0000007401|NDFRT|Immunoglobulins, Intravenous||P|PF|N
C0085297|T116|N0000007401|NDFRT|Immunoglobulins, Intravenous||P|PF|N
C0085297|T129|N0000007401|NDFRT|Immunoglobulins, Intravenous||P|PF|N
C0085297|T121|N0000007401|NDFRT|Immunoglobulins, Intravenous [Chemical/Ingredient]||S|PF|Y
C0085297|T116|N0000007401|NDFRT|Immunoglobulins, Intravenous [Chemical/Ingredient]||S|PF|Y
C0085297|T129|N0000007401|NDFRT|Immunoglobulins, Intravenous [Chemical/Ingredient]||S|PF|Y
C0085297|T121|N0000007401|NDFRT|Intravenous Antibodies||S|PF|N
C0085297|T116|N0000007401|NDFRT|Intravenous Antibodies||S|PF|N
C0085297|T129|N0000007401|NDFRT|Intravenous Antibodies||S|PF|N
C0085297|T121|N0000007401|NDFRT|Intravenous IG||S|PF|N
C0085297|T116|N0000007401|NDFRT|Intravenous IG||S|PF|N
C0085297|T129|N0000007401|NDFRT|Intravenous IG||S|PF|N
C0085297|T121|N0000007401|NDFRT|Intravenous Immunoglobulins||P|VW|N
C0085297|T116|N0000007401|NDFRT|Intravenous Immunoglobulins||P|VW|N
C0085297|T129|N0000007401|NDFRT|Intravenous Immunoglobulins||P|VW|N
C0085297|T121|N0000007401|NDFRT|IV Immunoglobulins||S|PF|N
C0085297|T116|N0000007401|NDFRT|IV Immunoglobulins||S|PF|N
C0085297|T129|N0000007401|NDFRT|IV Immunoglobulins||S|PF|N
C0085297|T121|N0000007401|NDFRT|IVIG||S|PF|N
C0085297|T116|N0000007401|NDFRT|IVIG||S|PF|N
C0085297|T129|N0000007401|NDFRT|IVIG||S|PF|N
C0085297|T121|N0000146387|NDFRT|GLOBULIN,IMMUNE (IV)||S|PF|N
C0085297|T116|N0000146387|NDFRT|GLOBULIN,IMMUNE (IV)||S|PF|N
C0085297|T129|N0000146387|NDFRT|GLOBULIN,IMMUNE (IV)||S|PF|N
C0085297|T121|CDR0000040109|PDQ|Immune Globulin Intravenous||S|VO|Y
C0085297|T116|CDR0000040109|PDQ|Immune Globulin Intravenous||S|VO|Y
C0085297|T129|CDR0000040109|PDQ|Immune Globulin Intravenous||S|VO|Y
C0085297|T121|CDR0000040109|PDQ|Immune Globulin IV||S|VCW|Y
C0085297|T116|CDR0000040109|PDQ|Immune Globulin IV||S|VCW|Y
C0085297|T129|CDR0000040109|PDQ|Immune Globulin IV||S|VCW|Y
C0085297|T121|42386|RXNORM|Immunoglobulins, Intravenous||P|PF|N
C0085297|T116|42386|RXNORM|Immunoglobulins, Intravenous||P|PF|N
C0085297|T129|42386|RXNORM|Immunoglobulins, Intravenous||P|PF|N
C0085297|T121|34245000|SNOMEDCT_US|IGIV||S|PF|N
C0085297|T116|34245000|SNOMEDCT_US|IGIV||S|PF|N
C0085297|T129|34245000|SNOMEDCT_US|IGIV||S|PF|N
C0085297|T121|34245000|SNOMEDCT_US|Immune globulin IV||S|VCW|Y
C0085297|T116|34245000|SNOMEDCT_US|Immune globulin IV||S|VCW|Y
C0085297|T129|34245000|SNOMEDCT_US|Immune globulin IV||S|VCW|Y
C0085297|T121|34245000|SNOMEDCT_US|Immune globulin IV (product)||S|PF|Y
C0085297|T116|34245000|SNOMEDCT_US|Immune globulin IV (product)||S|PF|Y
C0085297|T129|34245000|SNOMEDCT_US|Immune globulin IV (product)||S|PF|Y
C0085297|T121|34245000|SNOMEDCT_US|Immune globulin IV (substance)||S|PF|Y
C0085297|T116|34245000|SNOMEDCT_US|Immune globulin IV (substance)||S|PF|Y
C0085297|T129|34245000|SNOMEDCT_US|Immune globulin IV (substance)||S|PF|Y
C0085297|T121|350344000|SNOMEDCT_US|Intravenous immunoglobulin||P|VO|Y
C0085297|T116|350344000|SNOMEDCT_US|Intravenous immunoglobulin||P|VO|Y
C0085297|T129|350344000|SNOMEDCT_US|Intravenous immunoglobulin||P|VO|Y
C0085297|T121|350344000|SNOMEDCT_US|Intravenous immunoglobulin (product)||S|PF|Y
C0085297|T116|350344000|SNOMEDCT_US|Intravenous immunoglobulin (product)||S|PF|Y
C0085297|T129|350344000|SNOMEDCT_US|Intravenous immunoglobulin (product)||S|PF|Y
C0085297|T121|350344000|SNOMEDCT_US|Intravenous immunoglobulin (substance)||S|PF|Y
C0085297|T116|350344000|SNOMEDCT_US|Intravenous immunoglobulin (substance)||S|PF|Y
C0085297|T129|350344000|SNOMEDCT_US|Intravenous immunoglobulin (substance)||S|PF|Y
C0085297|T121|4018045|VANDF|GLOBULIN,IMMUNE (IV)||S|PF|Y
C0085297|T116|4018045|VANDF|GLOBULIN,IMMUNE (IV)||S|PF|Y
C0085297|T129|4018045|VANDF|GLOBULIN,IMMUNE (IV)||S|PF|Y
C0086413|T121|3059-5000|CSP|HIV vaccine||P|VC|Y
C0086413|T129|3059-5000|CSP|HIV vaccine||P|VC|Y
C0086413|T121|61|CVX|HIV||S|PF|N
C0086413|T129|61|CVX|HIV||S|PF|N
C0086413|T121|61|CVX|human immunodeficiency virus vaccine||S|PF|Y
C0086413|T129|61|CVX|human immunodeficiency virus vaccine||S|PF|Y
C0086413|T121|61|HL7V2.5|HIV||S|PF|N
C0086413|T129|61|HL7V2.5|HIV||S|PF|N
C0086413|T121|61|HL7V3.0|HIV||S|PF|N
C0086413|T129|61|HL7V3.0|HIV||S|PF|N
C0086413|T121|LP183501-8|LNC|HIV||S|PF|Y
C0086413|T129|LP183501-8|LNC|HIV||S|PF|Y
C0086413|T121|D016915|MSH|HIV Vaccines||P|VO|Y
C0086413|T129|D016915|MSH|HIV Vaccines||P|VO|Y
C0086413|T121|NOCODE|MTH|HIV Vaccine||P|PF|Y
C0086413|T129|NOCODE|MTH|HIV Vaccine||P|PF|Y
C0086413|T121|C1325|NCI|HIV Vaccine||P|PF|N
C0086413|T129|C1325|NCI|HIV Vaccine||P|PF|N
C0086413|T121|C1325|NCI|HIV/AIDS Vaccines||S|PF|Y
C0086413|T129|C1325|NCI|HIV/AIDS Vaccines||S|PF|Y
C0206255|T121|3058-4206|CSP|malaria vaccine||P|VO|N
C0206255|T129|3058-4206|CSP|malaria vaccine||P|VO|N
C0206255|T121|67|CVX|malaria||S|PF|N
C0206255|T129|67|CVX|malaria||S|PF|N
C0206255|T121|67|CVX|malaria vaccine||P|VO|Y
C0206255|T129|67|CVX|malaria vaccine||P|VO|Y
C0206255|T121|67|HL7V2.5|malaria||S|PF|N
C0206255|T129|67|HL7V2.5|malaria||S|PF|N
C0206255|T121|67|HL7V3.0|malaria||S|PF|Y
C0206255|T129|67|HL7V3.0|malaria||S|PF|Y
C0206255|T121|sh86005372|LCH_NW|Malaria vaccine||P|VO|Y
C0206255|T129|sh86005372|LCH_NW|Malaria vaccine||P|VO|Y
C0206255|T121|D017780|MSH|Malaria Vaccines||P|PF|N
C0206255|T129|D017780|MSH|Malaria Vaccines||P|PF|N
C0206255|T121|D017780|MSH|Malarial Vaccines||S|PF|Y
C0206255|T129|D017780|MSH|Malarial Vaccines||S|PF|Y
C0206255|T121|D017780|MSH|Vaccines, Malaria||P|VW|Y
C0206255|T129|D017780|MSH|Vaccines, Malaria||P|VW|Y
C0206255|T121|D017780|MSH|Vaccines, Malarial||S|VW|Y
C0206255|T129|D017780|MSH|Vaccines, Malarial||S|VW|Y
C0206255|T121|NOCODE|MTH|Malaria Vaccines||P|PF|Y
C0206255|T129|NOCODE|MTH|Malaria Vaccines||P|PF|Y
C0206255|T121|N0000170878|NDFRT|Malaria Vaccines||P|PF|N
C0206255|T129|N0000170878|NDFRT|Malaria Vaccines||P|PF|N
C0206255|T121|N0000170878|NDFRT|Malaria Vaccines [Chemical/Ingredient]||S|PF|Y
C0206255|T129|N0000170878|NDFRT|Malaria Vaccines [Chemical/Ingredient]||S|PF|Y
C0206255|T121|N0000170878|NDFRT|Malarial Vaccines||S|PF|N
C0206255|T129|N0000170878|NDFRT|Malarial Vaccines||S|PF|N
C0301508|T121|3059-1698|CSP|yellow fever vaccine||P|VC|N
C0301508|T129|3059-1698|CSP|yellow fever vaccine||P|VC|N
C0301508|T121|3100-3104|CSP|yellow fever vaccine||P|VC|N
C0301508|T129|3100-3104|CSP|yellow fever vaccine||P|VC|N
C0301508|T121|37|CVX|yellow fever||S|PF|N
C0301508|T129|37|CVX|yellow fever||S|PF|N
C0301508|T121|37|CVX|yellow fever vaccine||P|VC|N
C0301508|T129|37|CVX|yellow fever vaccine||P|VC|N
C0301508|T121|37|HL7V2.5|yellow fever||S|PF|N
C0301508|T129|37|HL7V2.5|yellow fever||S|PF|N
C0301508|T121|37|HL7V3.0|yellow fever||S|PF|Y
C0301508|T129|37|HL7V3.0|yellow fever||S|PF|Y
C0301508|T121|sh85149095|LCH_NW|Yellow fever vaccine||P|VC|N
C0301508|T129|sh85149095|LCH_NW|Yellow fever vaccine||P|VC|N
C0301508|T121|44445|MEDCIN|vaccines viral yellow fever||S|PF|Y
C0301508|T129|44445|MEDCIN|vaccines viral yellow fever||S|PF|Y
C0301508|T121|44445|MEDCIN|yellow fever vaccine||P|VC|N
C0301508|T129|44445|MEDCIN|yellow fever vaccine||P|VC|N
C0301508|T121|44445|MEDCIN|yellow fever vaccine (medication)||S|PF|Y
C0301508|T129|44445|MEDCIN|yellow fever vaccine (medication)||S|PF|Y
C0301508|T121|d01165|MMSL|yellow fever vaccine||P|VC|Y
C0301508|T129|d01165|MMSL|yellow fever vaccine||P|VC|Y
C0301508|T121|D022341|MSH|Fever Vaccine, Yellow||P|VW|Y
C0301508|T129|D022341|MSH|Fever Vaccine, Yellow||P|VW|Y
C0301508|T121|D022341|MSH|Vaccine, Yellow Fever||P|VW|Y
C0301508|T129|D022341|MSH|Vaccine, Yellow Fever||P|VW|Y
C0301508|T121|D022341|MSH|Yellow Fever Vaccine||P|PF|N
C0301508|T129|D022341|MSH|Yellow Fever Vaccine||P|PF|N
C0301508|T121|NOCODE|MTH|Yellow Fever Vaccine||P|PF|Y
C0301508|T129|NOCODE|MTH|Yellow Fever Vaccine||P|PF|Y
C0301508|T121|C96396|NCI|Yellow Fever Vaccine||P|PF|N
C0301508|T129|C96396|NCI|Yellow Fever Vaccine||P|PF|N
C0301508|T121|C96396|NCI_NICHD|Yellow Fever Vaccine||P|PF|N
C0301508|T129|C96396|NCI_NICHD|Yellow Fever Vaccine||P|PF|N
C0301508|T121|N0000005680|NDFRT|Yellow Fever Vaccine||P|PF|N
C0301508|T129|N0000005680|NDFRT|Yellow Fever Vaccine||P|PF|N
C0301508|T121|N0000005680|NDFRT|Yellow Fever Vaccine [Chemical/Ingredient]||S|PF|Y
C0301508|T129|N0000005680|NDFRT|Yellow Fever Vaccine [Chemical/Ingredient]||S|PF|Y
C0301508|T121|N0000146121|NDFRT|YELLOW FEVER VACCINE||P|VC|N
C0301508|T129|N0000146121|NDFRT|YELLOW FEVER VACCINE||P|VC|N
C0301508|T121|89890|RXNORM|Yellow Fever Vaccine||P|PF|N
C0301508|T129|89890|RXNORM|Yellow Fever Vaccine||P|PF|N
C0301508|T121|396444004|SNOMEDCT_US|Yellow fever vaccine||P|VC|Y
C0301508|T129|396444004|SNOMEDCT_US|Yellow fever vaccine||P|VC|Y
C0301508|T121|396444004|SNOMEDCT_US|Yellow fever vaccine (substance)||S|PF|Y
C0301508|T129|396444004|SNOMEDCT_US|Yellow fever vaccine (substance)||S|PF|Y
C0301508|T121|56844000|SNOMEDCT_US|Yellow fever vaccine||P|VC|N
C0301508|T129|56844000|SNOMEDCT_US|Yellow fever vaccine||P|VC|N
C0301508|T121|56844000|SNOMEDCT_US|Yellow fever vaccine (product)||S|PF|Y
C0301508|T129|56844000|SNOMEDCT_US|Yellow fever vaccine (product)||S|PF|Y
C0301508|T121|56844000|SNOMEDCT_US|Yellow fever vaccine (substance)||S|PF|N
C0301508|T129|56844000|SNOMEDCT_US|Yellow fever vaccine (substance)||S|PF|N
C0301508|T121|56844000|SNOMEDCT_US|Yellow fever vaccine product||S|VO|Y
C0301508|T129|56844000|SNOMEDCT_US|Yellow fever vaccine product||S|VO|Y
C0301508|T121|4017755|VANDF|YELLOW FEVER VACCINE||P|VC|Y
C0301508|T129|4017755|VANDF|YELLOW FEVER VACCINE||P|VC|Y
C0305060|T121|09|CVX|Td (adult), adsorbed||S|PF|Y
C0305060|T116|09|CVX|Td (adult), adsorbed||S|PF|Y
C0305060|T129|09|CVX|Td (adult), adsorbed||S|PF|Y
C0305060|T121|09|CVX|tetanus and diphtheria toxoids, adsorbed, for adult use||P|VO|Y
C0305060|T116|09|CVX|tetanus and diphtheria toxoids, adsorbed, for adult use||P|VO|Y
C0305060|T129|09|CVX|tetanus and diphtheria toxoids, adsorbed, for adult use||P|VO|Y
C0305060|T121|09|HL7V2.5|Td (adult)||S|PF|N
C0305060|T116|09|HL7V2.5|Td (adult)||S|PF|N
C0305060|T129|09|HL7V2.5|Td (adult)||S|PF|N
C0305060|T121|9|HL7V3.0|Td (adult)||S|PF|Y
C0305060|T116|9|HL7V3.0|Td (adult)||S|PF|Y
C0305060|T129|9|HL7V3.0|Td (adult)||S|PF|Y
C0305060|T121|NOCODE|MTH|Tetanus and diphtheria toxoid adsorbed for adult use||P|PF|Y
C0305060|T116|NOCODE|MTH|Tetanus and diphtheria toxoid adsorbed for adult use||P|PF|Y
C0305060|T129|NOCODE|MTH|Tetanus and diphtheria toxoid adsorbed for adult use||P|PF|Y
C0305060|T121|C96405|NCI|Td||S|PF|N
C0305060|T116|C96405|NCI|Td||S|PF|N
C0305060|T129|C96405|NCI|Td||S|PF|N
C0305060|T121|C96405|NCI|Tetanus and Diphtheria Toxoids Adsorbed||S|PF|Y
C0305060|T116|C96405|NCI|Tetanus and Diphtheria Toxoids Adsorbed||S|PF|Y
C0305060|T129|C96405|NCI|Tetanus and Diphtheria Toxoids Adsorbed||S|PF|Y
C0305060|T121|C96405|NCI|Tetanus and Diphtheria Toxoids Adsorbed for Adult Use||P|VO|Y
C0305060|T116|C96405|NCI|Tetanus and Diphtheria Toxoids Adsorbed for Adult Use||P|VO|Y
C0305060|T129|C96405|NCI|Tetanus and Diphtheria Toxoids Adsorbed for Adult Use||P|VO|Y
C0305060|T121|C96405|NCI_NICHD|Td||S|PF|Y
C0305060|T116|C96405|NCI_NICHD|Td||S|PF|Y
C0305060|T129|C96405|NCI_NICHD|Td||S|PF|Y
C0305060|T121|C96405|NCI_NICHD|Tetanus and Diphtheria Toxoids Adsorbed||S|PF|N
C0305060|T116|C96405|NCI_NICHD|Tetanus and Diphtheria Toxoids Adsorbed||S|PF|N
C0305060|T129|C96405|NCI_NICHD|Tetanus and Diphtheria Toxoids Adsorbed||S|PF|N
C0305060|T121|59999009|SNOMEDCT_US|TD||S|VC|Y
C0305060|T116|59999009|SNOMEDCT_US|TD||S|VC|Y
C0305060|T129|59999009|SNOMEDCT_US|TD||S|VC|Y
C0305060|T121|59999009|SNOMEDCT_US|TD toxoid||S|PF|Y
C0305060|T116|59999009|SNOMEDCT_US|TD toxoid||S|PF|Y
C0305060|T129|59999009|SNOMEDCT_US|TD toxoid||S|PF|Y
C0305060|T121|59999009|SNOMEDCT_US|Tetanus and diphtheria toxoid adsorbed for adult use||P|PF|N
C0305060|T116|59999009|SNOMEDCT_US|Tetanus and diphtheria toxoid adsorbed for adult use||P|PF|N
C0305060|T129|59999009|SNOMEDCT_US|Tetanus and diphtheria toxoid adsorbed for adult use||P|PF|N
C0305060|T121|59999009|SNOMEDCT_US|Tetanus and diphtheria toxoid adsorbed for adult use (product)||S|PF|Y
C0305060|T116|59999009|SNOMEDCT_US|Tetanus and diphtheria toxoid adsorbed for adult use (product)||S|PF|Y
C0305060|T129|59999009|SNOMEDCT_US|Tetanus and diphtheria toxoid adsorbed for adult use (product)||S|PF|Y
C0305060|T121|59999009|SNOMEDCT_US|Tetanus and diphtheria toxoid adsorbed for adult use (substance)||S|PF|Y
C0305060|T116|59999009|SNOMEDCT_US|Tetanus and diphtheria toxoid adsorbed for adult use (substance)||S|PF|Y
C0305060|T129|59999009|SNOMEDCT_US|Tetanus and diphtheria toxoid adsorbed for adult use (substance)||S|PF|Y
C0305062|T129|1554-6078|CSP|tetanus toxoid||S|VC|N
C0305062|T116|1554-6078|CSP|tetanus toxoid||S|VC|N
C0305062|T121|1554-6078|CSP|tetanus toxoid||S|VC|N
C0305062|T129|35|CVX|tetanus toxoid, adsorbed||S|VC|N
C0305062|T129|35|CVX|tetanus toxoid, adsorbed||S|VC|Y
C0305062|T116|35|CVX|tetanus toxoid, adsorbed||S|VC|N
C0305062|T116|35|CVX|tetanus toxoid, adsorbed||S|VC|Y
C0305062|T121|35|CVX|tetanus toxoid, adsorbed||S|VC|N
C0305062|T121|35|CVX|tetanus toxoid, adsorbed||S|VC|Y
C0305062|T129|35|HL7V2.5|tetanus toxoid||S|VC|N
C0305062|T116|35|HL7V2.5|tetanus toxoid||S|VC|N
C0305062|T121|35|HL7V2.5|tetanus toxoid||S|VC|N
C0305062|T129|35|HL7V3.0|tetanus toxoid||S|VC|N
C0305062|T116|35|HL7V3.0|tetanus toxoid||S|VC|N
C0305062|T121|35|HL7V3.0|tetanus toxoid||S|VC|N
C0305062|T129|LA10510-8|LNC|Tetanus||S|VC|Y
C0305062|T116|LA10510-8|LNC|Tetanus||S|VC|Y
C0305062|T121|LA10510-8|LNC|Tetanus||S|VC|Y
C0305062|T129|40141|MEDCIN|tetanus toxoid||S|VC|N
C0305062|T116|40141|MEDCIN|tetanus toxoid||S|VC|N
C0305062|T121|40141|MEDCIN|tetanus toxoid||S|VC|N
C0305062|T129|40141|MEDCIN|tetanus toxoid (medication)||S|PF|Y
C0305062|T116|40141|MEDCIN|tetanus toxoid (medication)||S|PF|Y
C0305062|T121|40141|MEDCIN|tetanus toxoid (medication)||S|PF|Y
C0305062|T129|11718|MMSL|Tetanus Toxoid||S|PF|N
C0305062|T116|11718|MMSL|Tetanus Toxoid||S|PF|N
C0305062|T121|11718|MMSL|Tetanus Toxoid||S|PF|N
C0305062|T129|2014|MMSL|Tetanus Toxoid Adsorbed||S|VC|Y
C0305062|T116|2014|MMSL|Tetanus Toxoid Adsorbed||S|VC|Y
C0305062|T121|2014|MMSL|Tetanus Toxoid Adsorbed||S|VC|Y
C0305062|T129|5556|MMSL|tetanus||S|PF|Y
C0305062|T116|5556|MMSL|tetanus||S|PF|Y
C0305062|T121|5556|MMSL|tetanus||S|PF|Y
C0305062|T129|5558|MMSL|tetanus toxoid||S|VC|N
C0305062|T116|5558|MMSL|tetanus toxoid||S|VC|N
C0305062|T121|5558|MMSL|tetanus toxoid||S|VC|N
C0305062|T129|d01168|MMSL|tetanus toxoid||S|VC|Y
C0305062|T116|d01168|MMSL|tetanus toxoid||S|VC|Y
C0305062|T121|d01168|MMSL|tetanus toxoid||S|VC|Y
C0305062|T129|D013745|MSH|Tetanus Toxoid||S|PF|Y
C0305062|T116|D013745|MSH|Tetanus Toxoid||S|PF|Y
C0305062|T121|D013745|MSH|Tetanus Toxoid||S|PF|Y
C0305062|T129|D013745|MSH|Toxoid, Tetanus||S|VW|Y
C0305062|T116|D013745|MSH|Toxoid, Tetanus||S|VW|Y
C0305062|T121|D013745|MSH|Toxoid, Tetanus||S|VW|Y
C0305062|T129|NOCODE|MTH|tetanus toxoid vaccine, inactivated||P|PF|Y
C0305062|T116|NOCODE|MTH|tetanus toxoid vaccine, inactivated||P|PF|Y
C0305062|T121|NOCODE|MTH|tetanus toxoid vaccine, inactivated||P|PF|Y
C0305062|T129|751E8J54VM|MTHSPL|CLOSTRIDIUM TETANI||S|PF|Y
C0305062|T116|751E8J54VM|MTHSPL|CLOSTRIDIUM TETANI||S|PF|Y
C0305062|T121|751E8J54VM|MTHSPL|CLOSTRIDIUM TETANI||S|PF|Y
C0305062|T129|K3W1N8YP13|MTHSPL|CLOSTRIDIUM TETANI TOXOID ANTIGEN (FORMALDEHYDE INACTIVATED)||S|PF|Y
C0305062|T116|K3W1N8YP13|MTHSPL|CLOSTRIDIUM TETANI TOXOID ANTIGEN (FORMALDEHYDE INACTIVATED)||S|PF|Y
C0305062|T121|K3W1N8YP13|MTHSPL|CLOSTRIDIUM TETANI TOXOID ANTIGEN (FORMALDEHYDE INACTIVATED)||S|PF|Y
C0305062|T129|C2660|NCI|Tetanus Toxoid||S|PF|N
C0305062|T116|C2660|NCI|Tetanus Toxoid||S|PF|N
C0305062|T121|C2660|NCI|Tetanus Toxoid||S|PF|N
C0305062|T129|C2660|NCI|Tetanus Toxoid Vaccine||S|PF|Y
C0305062|T116|C2660|NCI|Tetanus Toxoid Vaccine||S|PF|Y
C0305062|T121|C2660|NCI|Tetanus Toxoid Vaccine||S|PF|Y
C0305062|T129|C77704|NCI|Clostridium tetani Toxoid Antigen (Formaldehyde Inactivated)||S|VC|Y
C0305062|T116|C77704|NCI|Clostridium tetani Toxoid Antigen (Formaldehyde Inactivated)||S|VC|Y
C0305062|T121|C77704|NCI|Clostridium tetani Toxoid Antigen (Formaldehyde Inactivated)||S|VC|Y
C0305062|T129|C77704|NCI|Clostridium tetani Toxoid Antigen, A||S|PF|Y
C0305062|T116|C77704|NCI|Clostridium tetani Toxoid Antigen, A||S|PF|Y
C0305062|T121|C77704|NCI|Clostridium tetani Toxoid Antigen, A||S|PF|Y
C0305062|T129|C77704|NCI|Tetanus Toxoid||S|PF|N
C0305062|T116|C77704|NCI|Tetanus Toxoid||S|PF|N
C0305062|T121|C77704|NCI|Tetanus Toxoid||S|PF|N
C0305062|T129|TCGA|NCI|Tetanus Toxoid Vaccine||S|PF|N
C0305062|T116|TCGA|NCI|Tetanus Toxoid Vaccine||S|PF|N
C0305062|T121|TCGA|NCI|Tetanus Toxoid Vaccine||S|PF|N
C0305062|T129|K3W1N8YP13|NCI_FDA|CLOSTRIDIUM TETANI TOXOID ANTIGEN (FORMALDEHYDE INACTIVATED)||S|PF|N
C0305062|T116|K3W1N8YP13|NCI_FDA|CLOSTRIDIUM TETANI TOXOID ANTIGEN (FORMALDEHYDE INACTIVATED)||S|PF|N
C0305062|T121|K3W1N8YP13|NCI_FDA|CLOSTRIDIUM TETANI TOXOID ANTIGEN (FORMALDEHYDE INACTIVATED)||S|PF|N
C0305062|T129|CDR0000045064|NCI_NCI-GLOSS|tetanus toxoid||S|VC|N
C0305062|T116|CDR0000045064|NCI_NCI-GLOSS|tetanus toxoid||S|VC|N
C0305062|T121|CDR0000045064|NCI_NCI-GLOSS|tetanus toxoid||S|VC|N
C0305062|T129|C2660|NCI_NICHD|Tetanus Toxoid Vaccine||S|PF|N
C0305062|T116|C2660|NCI_NICHD|Tetanus Toxoid Vaccine||S|PF|N
C0305062|T121|C2660|NCI_NICHD|Tetanus Toxoid Vaccine||S|PF|N
C0305062|T129|C2660|NCI_NICHD|TT||S|PF|Y
C0305062|T116|C2660|NCI_NICHD|TT||S|PF|Y
C0305062|T121|C2660|NCI_NICHD|TT||S|PF|Y
C0305062|T129|N0000005564|NDFRT|Tetanus Toxoid||S|PF|N
C0305062|T116|N0000005564|NDFRT|Tetanus Toxoid||S|PF|N
C0305062|T121|N0000005564|NDFRT|Tetanus Toxoid||S|PF|N
C0305062|T129|N0000005564|NDFRT|Tetanus Toxoid [Chemical/Ingredient]||S|PF|Y
C0305062|T116|N0000005564|NDFRT|Tetanus Toxoid [Chemical/Ingredient]||S|PF|Y
C0305062|T121|N0000005564|NDFRT|Tetanus Toxoid [Chemical/Ingredient]||S|PF|Y
C0305062|T129|N0000146118|NDFRT|TETANUS TOXOID ADSORBED||S|VC|N
C0305062|T116|N0000146118|NDFRT|TETANUS TOXOID ADSORBED||S|VC|N
C0305062|T121|N0000146118|NDFRT|TETANUS TOXOID ADSORBED||S|VC|N
C0305062|T129|N0000146120|NDFRT|TETANUS TOXOID||S|VC|N
C0305062|T116|N0000146120|NDFRT|TETANUS TOXOID||S|VC|N
C0305062|T121|N0000146120|NDFRT|TETANUS TOXOID||S|VC|N
C0305062|T129|CDR0000038508|PDQ|tetanus toxoid||S|VC|N
C0305062|T116|CDR0000038508|PDQ|tetanus toxoid||S|VC|N
C0305062|T121|CDR0000038508|PDQ|tetanus toxoid||S|VC|N
C0305062|T129|CDR0000038508|PDQ|TETTOX||S|PF|Y
C0305062|T116|CDR0000038508|PDQ|TETTOX||S|PF|Y
C0305062|T121|CDR0000038508|PDQ|TETTOX||S|PF|Y
C0305062|T129|798306|RXNORM|tetanus toxoid vaccine, inactivated||P|PF|N
C0305062|T116|798306|RXNORM|tetanus toxoid vaccine, inactivated||P|PF|N
C0305062|T121|798306|RXNORM|tetanus toxoid vaccine, inactivated||P|PF|N
C0305062|T129|333621002|SNOMEDCT_US|Tetanus toxoids||S|VO|Y
C0305062|T116|333621002|SNOMEDCT_US|Tetanus toxoids||S|VO|Y
C0305062|T121|333621002|SNOMEDCT_US|Tetanus toxoids||S|VO|Y
C0305062|T129|396412003|SNOMEDCT_US|Tetanus toxoid||S|VC|Y
C0305062|T116|396412003|SNOMEDCT_US|Tetanus toxoid||S|VC|Y
C0305062|T121|396412003|SNOMEDCT_US|Tetanus toxoid||S|VC|Y
C0305062|T129|396412003|SNOMEDCT_US|Tetanus toxoid (substance)||S|PF|Y
C0305062|T116|396412003|SNOMEDCT_US|Tetanus toxoid (substance)||S|PF|Y
C0305062|T121|396412003|SNOMEDCT_US|Tetanus toxoid (substance)||S|PF|Y
C0305062|T129|58098008|SNOMEDCT_US|Tetanus toxoid adsorbed||S|PF|Y
C0305062|T116|58098008|SNOMEDCT_US|Tetanus toxoid adsorbed||S|PF|Y
C0305062|T121|58098008|SNOMEDCT_US|Tetanus toxoid adsorbed||S|PF|Y
C0305062|T129|58098008|SNOMEDCT_US|Tetanus toxoid adsorbed (product)||S|PF|Y
C0305062|T116|58098008|SNOMEDCT_US|Tetanus toxoid adsorbed (product)||S|PF|Y
C0305062|T121|58098008|SNOMEDCT_US|Tetanus toxoid adsorbed (product)||S|PF|Y
C0305062|T129|58098008|SNOMEDCT_US|Tetanus toxoid adsorbed (substance)||S|PF|Y
C0305062|T116|58098008|SNOMEDCT_US|Tetanus toxoid adsorbed (substance)||S|PF|Y
C0305062|T121|58098008|SNOMEDCT_US|Tetanus toxoid adsorbed (substance)||S|PF|Y
C0305062|T129|4017752|VANDF|TETANUS TOXOID ADSORBED||S|VC|Y
C0305062|T116|4017752|VANDF|TETANUS TOXOID ADSORBED||S|VC|Y
C0305062|T121|4017752|VANDF|TETANUS TOXOID ADSORBED||S|VC|Y
C0305062|T129|4017754|VANDF|TETANUS TOXOID||S|VC|Y
C0305062|T116|4017754|VANDF|TETANUS TOXOID||S|VC|Y
C0305062|T121|4017754|VANDF|TETANUS TOXOID||S|VC|Y
C0310756|T121|69|CVX|parainfluenza-3||S|PF|N
C0310756|T116|69|CVX|parainfluenza-3||S|PF|N
C0310756|T129|69|CVX|parainfluenza-3||S|PF|N
C0310756|T121|69|CVX|parainfluenza-3 virus vaccine||S|PF|Y
C0310756|T116|69|CVX|parainfluenza-3 virus vaccine||S|PF|Y
C0310756|T129|69|CVX|parainfluenza-3 virus vaccine||S|PF|Y
C0310756|T121|69|HL7V2.5|parainfluenza-3||S|PF|N
C0310756|T116|69|HL7V2.5|parainfluenza-3||S|PF|N
C0310756|T129|69|HL7V2.5|parainfluenza-3||S|PF|N
C0310756|T121|69|HL7V3.0|parainfluenza-3||S|PF|Y
C0310756|T116|69|HL7V3.0|parainfluenza-3||S|PF|Y
C0310756|T129|69|HL7V3.0|parainfluenza-3||S|PF|Y
C0310756|T121|82867008|SNOMEDCT_US|Parainfluenza 3 vaccine||P|PF|N
C0310756|T116|82867008|SNOMEDCT_US|Parainfluenza 3 vaccine||P|PF|N
C0310756|T129|82867008|SNOMEDCT_US|Parainfluenza 3 vaccine||P|PF|N
C0310756|T121|82867008|SNOMEDCT_US|Parainfluenza 3 vaccine (product)||S|PF|N
C0310756|T116|82867008|SNOMEDCT_US|Parainfluenza 3 vaccine (product)||S|PF|N
C0310756|T129|82867008|SNOMEDCT_US|Parainfluenza 3 vaccine (product)||S|PF|N
C0310756|T121|82867008|SNOMEDCT_US|Parainfluenza 3 vaccine (substance)||S|PF|Y
C0310756|T116|82867008|SNOMEDCT_US|Parainfluenza 3 vaccine (substance)||S|PF|Y
C0310756|T129|82867008|SNOMEDCT_US|Parainfluenza 3 vaccine (substance)||S|PF|Y
C0310756|T121|348721000009102|SNOMEDCT_VET|Parainfluenza 3 vaccine||P|PF|Y
C0310756|T116|348721000009102|SNOMEDCT_VET|Parainfluenza 3 vaccine||P|PF|Y
C0310756|T129|348721000009102|SNOMEDCT_VET|Parainfluenza 3 vaccine||P|PF|Y
C0310756|T121|348721000009102|SNOMEDCT_VET|Parainfluenza 3 vaccine (product)||S|PF|Y
C0310756|T116|348721000009102|SNOMEDCT_VET|Parainfluenza 3 vaccine (product)||S|PF|Y
C0310756|T129|348721000009102|SNOMEDCT_VET|Parainfluenza 3 vaccine (product)||S|PF|Y
C0358297|T121|90581|CPT|Anthrax vaccine||P|VO|N
C0358297|T129|90581|CPT|Anthrax vaccine||P|VO|N
C0358297|T121|5003-0003|CSP|anthrax vaccine||P|VO|N
C0358297|T129|5003-0003|CSP|anthrax vaccine||P|VO|N
C0358297|T121|24|CVX|anthrax||S|VC|N
C0358297|T129|24|CVX|anthrax||S|VC|N
C0358297|T121|24|CVX|anthrax vaccine||P|VO|Y
C0358297|T129|24|CVX|anthrax vaccine||P|VO|Y
C0358297|T121|24|HL7V2.5|anthrax||S|VC|Y
C0358297|T129|24|HL7V2.5|anthrax||S|VC|Y
C0358297|T121|24|HL7V3.0|Anthrax||S|PF|Y
C0358297|T129|24|HL7V3.0|Anthrax||S|PF|Y
C0358297|T121|308541|MEDCIN|Anthrax vaccine||P|VO|N
C0358297|T129|308541|MEDCIN|Anthrax vaccine||P|VO|N
C0358297|T121|308541|MEDCIN|anthrax vaccine (medication)||S|PF|Y
C0358297|T129|308541|MEDCIN|anthrax vaccine (medication)||S|PF|Y
C0358297|T121|D022122|MSH|Anthrax Vaccines||P|PF|N
C0358297|T129|D022122|MSH|Anthrax Vaccines||P|PF|N
C0358297|T121|D022122|MSH|Vaccines, Anthrax||P|VW|Y
C0358297|T129|D022122|MSH|Vaccines, Anthrax||P|VW|Y
C0358297|T121|NOCODE|MTH|Anthrax Vaccines||P|PF|Y
C0358297|T129|NOCODE|MTH|Anthrax Vaccines||P|PF|Y
C0358297|T121|N0000023074|NDFRT|ANTHRAX VACCINE||P|VO|N
C0358297|T129|N0000023074|NDFRT|ANTHRAX VACCINE||P|VO|N
C0358297|T121|N0000170890|NDFRT|Anthrax Vaccines||P|PF|N
C0358297|T129|N0000170890|NDFRT|Anthrax Vaccines||P|PF|N
C0358297|T121|N0000170890|NDFRT|Anthrax Vaccines [Chemical/Ingredient]||S|PF|Y
C0358297|T129|N0000170890|NDFRT|Anthrax Vaccines [Chemical/Ingredient]||S|PF|Y
C0358297|T121|N0000170890|NDFRT|Vaccines, Anthrax||P|VW|N
C0358297|T129|N0000170890|NDFRT|Vaccines, Anthrax||P|VW|N
C0358297|T121|333521006|SNOMEDCT_US|Anthrax vaccine||P|VO|Y
C0358297|T129|333521006|SNOMEDCT_US|Anthrax vaccine||P|VO|Y
C0358297|T121|333521006|SNOMEDCT_US|Anthrax vaccine (product)||S|PF|Y
C0358297|T129|333521006|SNOMEDCT_US|Anthrax vaccine (product)||S|PF|Y
C0358297|T121|333521006|SNOMEDCT_US|Anthrax vaccine (substance)||S|PF|N
C0358297|T129|333521006|SNOMEDCT_US|Anthrax vaccine (substance)||S|PF|N
C0358297|T121|396420001|SNOMEDCT_US|Anthrax vaccine||P|VO|N
C0358297|T129|396420001|SNOMEDCT_US|Anthrax vaccine||P|VO|N
C0358297|T121|396420001|SNOMEDCT_US|Anthrax vaccine (substance)||S|PF|Y
C0358297|T129|396420001|SNOMEDCT_US|Anthrax vaccine (substance)||S|PF|Y
C0358297|T121|4021501|VANDF|ANTHRAX VACCINE||P|VO|Y
C0358297|T129|4021501|VANDF|ANTHRAX VACCINE||P|VO|Y
C0359940|T121|90690|CPT|TYPHOID VACCINE LIVE ORAL||P|VCW|Y
C0359940|T129|90690|CPT|TYPHOID VACCINE LIVE ORAL||P|VCW|Y
C0359940|T116|90690|CPT|TYPHOID VACCINE LIVE ORAL||P|VCW|Y
C0359940|T121|90690|CPT|TYPHOID VACCINE ORAL||S|PF|Y
C0359940|T129|90690|CPT|TYPHOID VACCINE ORAL||S|PF|Y
C0359940|T116|90690|CPT|TYPHOID VACCINE ORAL||S|PF|Y
C0359940|T121|90690|CPT|Typhoid vaccine, live, oral||P|VW|Y
C0359940|T129|90690|CPT|Typhoid vaccine, live, oral||P|VW|Y
C0359940|T116|90690|CPT|Typhoid vaccine, live, oral||P|VW|Y
C0359940|T121|25|CVX|typhoid vaccine, live, oral||P|VCW|Y
C0359940|T129|25|CVX|typhoid vaccine, live, oral||P|VCW|Y
C0359940|T116|25|CVX|typhoid vaccine, live, oral||P|VCW|Y
C0359940|T121|25|CVX|typhoid, oral||S|PF|N
C0359940|T129|25|CVX|typhoid, oral||S|PF|N
C0359940|T116|25|CVX|typhoid, oral||S|PF|N
C0359940|T121|90690|HCPT|Typhoid vaccine oral||S|VC|Y
C0359940|T129|90690|HCPT|Typhoid vaccine oral||S|VC|Y
C0359940|T116|90690|HCPT|Typhoid vaccine oral||S|VC|Y
C0359940|T121|25|HL7V2.5|typhoid, oral||S|PF|N
C0359940|T129|25|HL7V2.5|typhoid, oral||S|PF|N
C0359940|T116|25|HL7V2.5|typhoid, oral||S|PF|N
C0359940|T121|25|HL7V3.0|typhoid, oral||S|PF|Y
C0359940|T129|25|HL7V3.0|typhoid, oral||S|PF|Y
C0359940|T116|25|HL7V3.0|typhoid, oral||S|PF|Y
C0359940|T121|133295|MEDCIN|typhoid vaccine live, oral||P|VCW|Y
C0359940|T129|133295|MEDCIN|typhoid vaccine live, oral||P|VCW|Y
C0359940|T116|133295|MEDCIN|typhoid vaccine live, oral||P|VCW|Y
C0359940|T121|133295|MEDCIN|typhoid vaccine live, oral (medication)||S|PF|Y
C0359940|T129|133295|MEDCIN|typhoid vaccine live, oral (medication)||S|PF|Y
C0359940|T116|133295|MEDCIN|typhoid vaccine live, oral (medication)||S|PF|Y
C0359940|T121|346696005|SNOMEDCT_US|Typhoid live oral vaccine||P|PF|Y
C0359940|T129|346696005|SNOMEDCT_US|Typhoid live oral vaccine||P|PF|Y
C0359940|T116|346696005|SNOMEDCT_US|Typhoid live oral vaccine||P|PF|Y
C0359940|T121|346696005|SNOMEDCT_US|Typhoid live oral vaccine (product)||S|PF|Y
C0359940|T129|346696005|SNOMEDCT_US|Typhoid live oral vaccine (product)||S|PF|Y
C0359940|T116|346696005|SNOMEDCT_US|Typhoid live oral vaccine (product)||S|PF|Y
C0359940|T121|346696005|SNOMEDCT_US|Typhoid live oral vaccine (substance)||S|PF|Y
C0359940|T129|346696005|SNOMEDCT_US|Typhoid live oral vaccine (substance)||S|PF|Y
C0359940|T116|346696005|SNOMEDCT_US|Typhoid live oral vaccine (substance)||S|PF|Y
C0360506|T121|86|CVX|IG||S|PF|N
C0360506|T116|86|CVX|IG||S|PF|N
C0360506|T129|86|CVX|IG||S|PF|N
C0360506|T121|86|CVX|immune globulin, intramuscular||S|VO|Y
C0360506|T116|86|CVX|immune globulin, intramuscular||S|VO|Y
C0360506|T129|86|CVX|immune globulin, intramuscular||S|VO|Y
C0360506|T121|86|HL7V2.5|IG||S|PF|N
C0360506|T116|86|HL7V2.5|IG||S|PF|N
C0360506|T129|86|HL7V2.5|IG||S|PF|N
C0360506|T121|86|HL7V3.0|IG||S|PF|Y
C0360506|T116|86|HL7V3.0|IG||S|PF|Y
C0360506|T129|86|HL7V3.0|IG||S|PF|Y
C0360506|T121|d01135|MMSL|immune globulin intramuscular||S|PF|Y
C0360506|T116|d01135|MMSL|immune globulin intramuscular||S|PF|Y
C0360506|T129|d01135|MMSL|immune globulin intramuscular||S|PF|Y
C0360506|T121|NOCODE|MTH|Intramuscular immunoglobulin||P|PF|Y
C0360506|T116|NOCODE|MTH|Intramuscular immunoglobulin||P|PF|Y
C0360506|T129|NOCODE|MTH|Intramuscular immunoglobulin||P|PF|Y
C0360506|T121|N0000146386|NDFRT|GLOBULIN,IMMUNE (IM)||S|VCW|N
C0360506|T116|N0000146386|NDFRT|GLOBULIN,IMMUNE (IM)||S|VCW|N
C0360506|T129|N0000146386|NDFRT|GLOBULIN,IMMUNE (IM)||S|VCW|N
C0360506|T121|108067|RXNORM|Intramuscular immunoglobulin||P|PF|N
C0360506|T116|108067|RXNORM|Intramuscular immunoglobulin||P|PF|N
C0360506|T129|108067|RXNORM|Intramuscular immunoglobulin||P|PF|N
C0360506|T121|350343006|SNOMEDCT_US|Intramuscular immunoglobulin||P|PF|N
C0360506|T116|350343006|SNOMEDCT_US|Intramuscular immunoglobulin||P|PF|N
C0360506|T129|350343006|SNOMEDCT_US|Intramuscular immunoglobulin||P|PF|N
C0360506|T121|350343006|SNOMEDCT_US|Intramuscular immunoglobulin (product)||S|PF|Y
C0360506|T116|350343006|SNOMEDCT_US|Intramuscular immunoglobulin (product)||S|PF|Y
C0360506|T129|350343006|SNOMEDCT_US|Intramuscular immunoglobulin (product)||S|PF|Y
C0360506|T121|350343006|SNOMEDCT_US|Intramuscular immunoglobulin (substance)||S|PF|Y
C0360506|T116|350343006|SNOMEDCT_US|Intramuscular immunoglobulin (substance)||S|PF|Y
C0360506|T129|350343006|SNOMEDCT_US|Intramuscular immunoglobulin (substance)||S|PF|Y
C0360506|T121|36763003|SNOMEDCT_US|IGIM||S|PF|Y
C0360506|T116|36763003|SNOMEDCT_US|IGIM||S|PF|Y
C0360506|T129|36763003|SNOMEDCT_US|IGIM||S|PF|Y
C0360506|T121|36763003|SNOMEDCT_US|Immune globulin IM||S|PF|Y
C0360506|T116|36763003|SNOMEDCT_US|Immune globulin IM||S|PF|Y
C0360506|T129|36763003|SNOMEDCT_US|Immune globulin IM||S|PF|Y
C0360506|T121|36763003|SNOMEDCT_US|Immune globulin IM (product)||S|PF|Y
C0360506|T116|36763003|SNOMEDCT_US|Immune globulin IM (product)||S|PF|Y
C0360506|T129|36763003|SNOMEDCT_US|Immune globulin IM (product)||S|PF|Y
C0360506|T121|36763003|SNOMEDCT_US|Immune globulin IM (substance)||S|PF|Y
C0360506|T116|36763003|SNOMEDCT_US|Immune globulin IM (substance)||S|PF|Y
C0360506|T129|36763003|SNOMEDCT_US|Immune globulin IM (substance)||S|PF|Y
C0360506|T121|4018044|VANDF|GLOBULIN,IMMUNE (IM)||S|VCW|Y
C0360506|T116|4018044|VANDF|GLOBULIN,IMMUNE (IM)||S|VCW|Y
C0360506|T129|4018044|VANDF|GLOBULIN,IMMUNE (IM)||S|VCW|Y
C0388013|T116|71|CVX|respiratory syncytial virus immune globulin, intravenous||P|VO|Y
C0388013|T121|71|CVX|respiratory syncytial virus immune globulin, intravenous||P|VO|Y
C0388013|T129|71|CVX|respiratory syncytial virus immune globulin, intravenous||P|VO|Y
C0388013|T116|71|CVX|RSV-IGIV||S|PF|N
C0388013|T121|71|CVX|RSV-IGIV||S|PF|N
C0388013|T129|71|CVX|RSV-IGIV||S|PF|N
C0388013|T116|71|HL7V2.5|RSV-IGIV||S|PF|N
C0388013|T121|71|HL7V2.5|RSV-IGIV||S|PF|N
C0388013|T129|71|HL7V2.5|RSV-IGIV||S|PF|N
C0388013|T116|71|HL7V3.0|RSV-IGIV||S|PF|N
C0388013|T121|71|HL7V3.0|RSV-IGIV||S|PF|N
C0388013|T129|71|HL7V3.0|RSV-IGIV||S|PF|N
C0388013|T116|5419|MMSL|respiratory syncytial virus immunoglobulin||S|VC|Y
C0388013|T121|5419|MMSL|respiratory syncytial virus immunoglobulin||S|VC|Y
C0388013|T129|5419|MMSL|respiratory syncytial virus immunoglobulin||S|VC|Y
C0388013|T116|d03881|MMSL|respiratory syncytial virus immune globulin||S|VC|Y
C0388013|T121|d03881|MMSL|respiratory syncytial virus immune globulin||S|VC|Y
C0388013|T129|d03881|MMSL|respiratory syncytial virus immune globulin||S|VC|Y
C0388013|T116|C098685|MSH|respiratory syncytial virus immune globulin intravenous||P|PF|Y
C0388013|T121|C098685|MSH|respiratory syncytial virus immune globulin intravenous||P|PF|Y
C0388013|T129|C098685|MSH|respiratory syncytial virus immune globulin intravenous||P|PF|Y
C0388013|T116|C098685|MSH|RSV-IGIV||S|PF|Y
C0388013|T121|C098685|MSH|RSV-IGIV||S|PF|Y
C0388013|T129|C098685|MSH|RSV-IGIV||S|PF|Y
C0388013|T116|78I1W13C3D|MTHSPL|RESPIRATORY SYNCYTIAL VIRUS IMMUNE GLOBULIN INTRAVENOUS (HUMAN)||S|PF|Y
C0388013|T121|78I1W13C3D|MTHSPL|RESPIRATORY SYNCYTIAL VIRUS IMMUNE GLOBULIN INTRAVENOUS (HUMAN)||S|PF|Y
C0388013|T129|78I1W13C3D|MTHSPL|RESPIRATORY SYNCYTIAL VIRUS IMMUNE GLOBULIN INTRAVENOUS (HUMAN)||S|PF|Y
C0388013|T116|119246|RXNORM|respiratory syncytial virus immune globulin intravenous||P|PF|N
C0388013|T121|119246|RXNORM|respiratory syncytial virus immune globulin intravenous||P|PF|N
C0388013|T129|119246|RXNORM|respiratory syncytial virus immune globulin intravenous||P|PF|N
C0388013|T116|108723008|SNOMEDCT_US|Respiratory syncytial virus immune globulin||S|PF|Y
C0388013|T121|108723008|SNOMEDCT_US|Respiratory syncytial virus immune globulin||S|PF|Y
C0388013|T129|108723008|SNOMEDCT_US|Respiratory syncytial virus immune globulin||S|PF|Y
C0388013|T116|108723008|SNOMEDCT_US|Respiratory syncytial virus immune globulin (product)||S|PF|Y
C0388013|T121|108723008|SNOMEDCT_US|Respiratory syncytial virus immune globulin (product)||S|PF|Y
C0388013|T129|108723008|SNOMEDCT_US|Respiratory syncytial virus immune globulin (product)||S|PF|Y
C0388013|T116|108723008|SNOMEDCT_US|Respiratory syncytial virus immune globulin (substance)||S|PF|Y
C0388013|T121|108723008|SNOMEDCT_US|Respiratory syncytial virus immune globulin (substance)||S|PF|Y
C0388013|T129|108723008|SNOMEDCT_US|Respiratory syncytial virus immune globulin (substance)||S|PF|Y
C0388013|T116|120709004|SNOMEDCT_US|Respiratory syncytial virus immunoglobulin||S|PF|Y
C0388013|T121|120709004|SNOMEDCT_US|Respiratory syncytial virus immunoglobulin||S|PF|Y
C0388013|T129|120709004|SNOMEDCT_US|Respiratory syncytial virus immunoglobulin||S|PF|Y
C0593408|T121|77|CVX|tick-borne encephalitis||S|PF|N
C0593408|T129|77|CVX|tick-borne encephalitis||S|PF|N
C0593408|T116|77|CVX|tick-borne encephalitis||S|PF|N
C0593408|T121|77|CVX|tick-borne encephalitis vaccine||P|VC|Y
C0593408|T129|77|CVX|tick-borne encephalitis vaccine||P|VC|Y
C0593408|T116|77|CVX|tick-borne encephalitis vaccine||P|VC|Y
C0593408|T121|77|HL7V2.5|tick-borne encephalitis||S|PF|N
C0593408|T129|77|HL7V2.5|tick-borne encephalitis||S|PF|N
C0593408|T116|77|HL7V2.5|tick-borne encephalitis||S|PF|N
C0593408|T121|77|HL7V3.0|tick-borne encephalitis||S|PF|Y
C0593408|T129|77|HL7V3.0|tick-borne encephalitis||S|PF|Y
C0593408|T116|77|HL7V3.0|tick-borne encephalitis||S|PF|Y
C0593408|T121|NOCODE|MTH|Tick-borne encephalitis vaccine||P|PF|Y
C0593408|T129|NOCODE|MTH|Tick-borne encephalitis vaccine||P|PF|Y
C0593408|T116|NOCODE|MTH|Tick-borne encephalitis vaccine||P|PF|Y
C0593408|T121|333699008|SNOMEDCT_US|Tick-borne encephalitis vaccine||P|PF|N
C0593408|T129|333699008|SNOMEDCT_US|Tick-borne encephalitis vaccine||P|PF|N
C0593408|T116|333699008|SNOMEDCT_US|Tick-borne encephalitis vaccine||P|PF|N
C0593408|T121|333699008|SNOMEDCT_US|Tick-borne encephalitis vaccine (product)||S|PF|Y
C0593408|T129|333699008|SNOMEDCT_US|Tick-borne encephalitis vaccine (product)||S|PF|Y
C0593408|T116|333699008|SNOMEDCT_US|Tick-borne encephalitis vaccine (product)||S|PF|Y
C0593408|T121|333699008|SNOMEDCT_US|Tick-borne encephalitis vaccine (substance)||S|PF|N
C0593408|T129|333699008|SNOMEDCT_US|Tick-borne encephalitis vaccine (substance)||S|PF|N
C0593408|T116|333699008|SNOMEDCT_US|Tick-borne encephalitis vaccine (substance)||S|PF|N
C0593408|T121|398783009|SNOMEDCT_US|Tick-borne encephalitis vaccine||P|PF|N
C0593408|T129|398783009|SNOMEDCT_US|Tick-borne encephalitis vaccine||P|PF|N
C0593408|T116|398783009|SNOMEDCT_US|Tick-borne encephalitis vaccine||P|PF|N
C0593408|T121|398783009|SNOMEDCT_US|Tick-borne encephalitis vaccine (substance)||S|PF|Y
C0593408|T129|398783009|SNOMEDCT_US|Tick-borne encephalitis vaccine (substance)||S|PF|Y
C0593408|T116|398783009|SNOMEDCT_US|Tick-borne encephalitis vaccine (substance)||S|PF|Y
C0694727|T129|28|CVX|diphtheria and tetanus toxoids, adsorbed for pediatric use||P|PF|Y
C0694727|T121|28|CVX|diphtheria and tetanus toxoids, adsorbed for pediatric use||P|PF|Y
C0694727|T129|28|CVX|DT (pediatric)||S|PF|N
C0694727|T121|28|CVX|DT (pediatric)||S|PF|N
C0694727|T129|28|HL7V2.5|DT (pediatric)||S|PF|N
C0694727|T121|28|HL7V2.5|DT (pediatric)||S|PF|N
C0694727|T129|28|HL7V3.0|DT (pediatric)||S|PF|Y
C0694727|T121|28|HL7V3.0|DT (pediatric)||S|PF|Y
C0694730|T121|22|CVX|DTP-Haemophilus influenzae type b conjugate vaccine||P|PF|Y
C0694730|T129|22|CVX|DTP-Haemophilus influenzae type b conjugate vaccine||P|PF|Y
C0694730|T121|22|CVX|DTP-Hib||S|PF|N
C0694730|T129|22|CVX|DTP-Hib||S|PF|N
C0694730|T121|22|HL7V2.5|DTP-Hib||S|PF|N
C0694730|T129|22|HL7V2.5|DTP-Hib||S|PF|N
C0694730|T121|22|HL7V3.0|DTP-Hib||S|PF|Y
C0694730|T129|22|HL7V3.0|DTP-Hib||S|PF|Y
C0694731|T121|31|CVX|Hep A, pediatric, unspecified formulation||S|PF|Y
C0694731|T129|31|CVX|Hep A, pediatric, unspecified formulation||S|PF|Y
C0694731|T121|31|CVX|hepatitis A vaccine, pediatric dosage, unspecified formulation||P|PF|Y
C0694731|T129|31|CVX|hepatitis A vaccine, pediatric dosage, unspecified formulation||P|PF|Y
C0694731|T121|31|HL7V2.5|Hep A, pediatric, NOS||S|PF|N
C0694731|T129|31|HL7V2.5|Hep A, pediatric, NOS||S|PF|N
C0694731|T121|31|HL7V3.0|Hep A, pediatric, NOS||S|PF|Y
C0694731|T129|31|HL7V3.0|Hep A, pediatric, NOS||S|PF|Y
C0694733|T121|08|CVX|Hep B, adolescent or pediatric||S|PF|N
C0694733|T129|08|CVX|Hep B, adolescent or pediatric||S|PF|N
C0694733|T121|08|CVX|hepatitis B vaccine, pediatric or pediatric/adolescent dosage||P|PF|Y
C0694733|T129|08|CVX|hepatitis B vaccine, pediatric or pediatric/adolescent dosage||P|PF|Y
C0694733|T121|08|HL7V2.5|Hep B, adolescent or pediatric||S|PF|N
C0694733|T129|08|HL7V2.5|Hep B, adolescent or pediatric||S|PF|N
C0694733|T121|8|HL7V3.0|Hep B, adolescent or pediatric||S|PF|Y
C0694733|T129|8|HL7V3.0|Hep B, adolescent or pediatric||S|PF|Y
C0694736|T121|44|CVX|Hep B, dialysis||S|PF|N
C0694736|T129|44|CVX|Hep B, dialysis||S|PF|N
C0694736|T121|44|CVX|hepatitis B vaccine, dialysis patient dosage||P|PF|Y
C0694736|T129|44|CVX|hepatitis B vaccine, dialysis patient dosage||P|PF|Y
C0694736|T121|44|HL7V2.5|Hep B, dialysis||S|PF|N
C0694736|T129|44|HL7V2.5|Hep B, dialysis||S|PF|N
C0694736|T121|44|HL7V3.0|Hep B, dialysis||S|PF|Y
C0694736|T129|44|HL7V3.0|Hep B, dialysis||S|PF|Y
C0694739|T121|46|CVX|Haemophilus influenzae type b vaccine, PRP-D conjugate||P|PF|Y
C0694739|T129|46|CVX|Haemophilus influenzae type b vaccine, PRP-D conjugate||P|PF|Y
C0694739|T121|46|CVX|Hib (PRP-D)||S|PF|N
C0694739|T129|46|CVX|Hib (PRP-D)||S|PF|N
C0694739|T121|46|HL7V2.5|Hib (PRP-D)||S|PF|N
C0694739|T129|46|HL7V2.5|Hib (PRP-D)||S|PF|N
C0694739|T121|46|HL7V3.0|Hib (PRP-D)||S|PF|Y
C0694739|T129|46|HL7V3.0|Hib (PRP-D)||S|PF|Y
C0694740|T121|47|CVX|Haemophilus influenzae type b vaccine, HbOC conjugate||P|PF|Y
C0694740|T129|47|CVX|Haemophilus influenzae type b vaccine, HbOC conjugate||P|PF|Y
C0694740|T121|47|CVX|Hib (HbOC)||S|PF|N
C0694740|T129|47|CVX|Hib (HbOC)||S|PF|N
C0694740|T121|47|HL7V2.5|Hib (HbOC)||S|PF|N
C0694740|T129|47|HL7V2.5|Hib (HbOC)||S|PF|N
C0694740|T121|47|HL7V3.0|Hib (HbOC)||S|PF|Y
C0694740|T129|47|HL7V3.0|Hib (HbOC)||S|PF|Y
C0694741|T121|48|CVX|Haemophilus influenzae type b vaccine, PRP-T conjugate||P|PF|Y
C0694741|T129|48|CVX|Haemophilus influenzae type b vaccine, PRP-T conjugate||P|PF|Y
C0694741|T121|48|CVX|Hib (PRP-T)||S|PF|N
C0694741|T129|48|CVX|Hib (PRP-T)||S|PF|N
C0694741|T121|48|HL7V2.5|Hib (PRP-T)||S|PF|N
C0694741|T129|48|HL7V2.5|Hib (PRP-T)||S|PF|N
C0694741|T121|48|HL7V3.0|Hib (PRP-T)||S|PF|Y
C0694741|T129|48|HL7V3.0|Hib (PRP-T)||S|PF|Y
C0694742|T121|49|CVX|Haemophilus influenzae type b vaccine, PRP-OMP conjugate||P|PF|Y
C0694742|T129|49|CVX|Haemophilus influenzae type b vaccine, PRP-OMP conjugate||P|PF|Y
C0694742|T121|49|CVX|Hib (PRP-OMP)||S|PF|N
C0694742|T129|49|CVX|Hib (PRP-OMP)||S|PF|N
C0694742|T121|49|HL7V2.5|Hib (PRP-OMP)||S|PF|N
C0694742|T129|49|HL7V2.5|Hib (PRP-OMP)||S|PF|N
C0694742|T121|49|HL7V3.0|Hib (PRP-OMP)||S|PF|Y
C0694742|T129|49|HL7V3.0|Hib (PRP-OMP)||S|PF|Y
C0694743|T121|51|CVX|Haemophilus influenzae type b conjugate and Hepatitis B vaccine||P|PF|Y
C0694743|T129|51|CVX|Haemophilus influenzae type b conjugate and Hepatitis B vaccine||P|PF|Y
C0694743|T121|51|CVX|Hib-Hep B||S|PF|N
C0694743|T129|51|CVX|Hib-Hep B||S|PF|N
C0694743|T121|51|HL7V2.5|Hib-Hep B||S|PF|N
C0694743|T129|51|HL7V2.5|Hib-Hep B||S|PF|N
C0694743|T121|51|HL7V3.0|Hib-Hep B||S|PF|Y
C0694743|T129|51|HL7V3.0|Hib-Hep B||S|PF|Y
C0694744|T121|15|CVX|influenza virus vaccine, split virus (incl. purified surface antigen)-retired CODE||P|PF|Y
C0694744|T129|15|CVX|influenza virus vaccine, split virus (incl. purified surface antigen)-retired CODE||P|PF|Y
C0694744|T121|15|CVX|influenza, split (incl. purified surface antigen)||S|PF|N
C0694744|T129|15|CVX|influenza, split (incl. purified surface antigen)||S|PF|N
C0694744|T121|15|HL7V2.5|influenza, split (incl. purified surface antigen)||S|PF|N
C0694744|T129|15|HL7V2.5|influenza, split (incl. purified surface antigen)||S|PF|N
C0694744|T121|15|HL7V3.0|influenza, split (incl. purified surface antigen)||S|PF|Y
C0694744|T129|15|HL7V3.0|influenza, split (incl. purified surface antigen)||S|PF|Y
C0694745|T121|16|CVX|influenza virus vaccine, whole virus||P|PF|Y
C0694745|T129|16|CVX|influenza virus vaccine, whole virus||P|PF|Y
C0694745|T121|16|CVX|influenza, whole||S|PF|N
C0694745|T129|16|CVX|influenza, whole||S|PF|N
C0694745|T121|16|HL7V2.5|influenza, whole||S|PF|N
C0694745|T129|16|HL7V2.5|influenza, whole||S|PF|N
C0694745|T121|16|HL7V3.0|influenza, whole||S|PF|Y
C0694745|T129|16|HL7V3.0|influenza, whole||S|PF|Y
C0694746|T121|04|CVX|M/R||S|PF|N
C0694746|T129|04|CVX|M/R||S|PF|N
C0694746|T121|04|CVX|measles and rubella virus vaccine||S|VO|Y
C0694746|T129|04|CVX|measles and rubella virus vaccine||S|VO|Y
C0694746|T121|04|HL7V2.5|M/R||S|PF|N
C0694746|T129|04|HL7V2.5|M/R||S|PF|N
C0694746|T121|4|HL7V3.0|M/R||S|PF|Y
C0694746|T129|4|HL7V3.0|M/R||S|PF|Y
C0694746|T121|d03006|MMSL|measles-rubella virus vaccine||S|PF|Y
C0694746|T129|d03006|MMSL|measles-rubella virus vaccine||S|PF|Y
C0694746|T121|NOCODE|MTH|MR vaccine||P|PF|Y
C0694746|T129|NOCODE|MTH|MR vaccine||P|PF|Y
C0694749|T121|40|CVX|rabies vaccine, for intradermal injection||P|PF|Y
C0694749|T129|40|CVX|rabies vaccine, for intradermal injection||P|PF|Y
C0694749|T121|40|CVX|rabies, intradermal injection||S|PF|N
C0694749|T129|40|CVX|rabies, intradermal injection||S|PF|N
C0694749|T121|40|HL7V2.5|rabies, intradermal injection||S|PF|N
C0694749|T129|40|HL7V2.5|rabies, intradermal injection||S|PF|N
C0694749|T121|40|HL7V3.0|rabies, intradermal injection||S|PF|Y
C0694749|T129|40|HL7V3.0|rabies, intradermal injection||S|PF|Y
C0694750|T121|38|CVX|rubella and mumps virus vaccine||S|VO|Y
C0694750|T129|38|CVX|rubella and mumps virus vaccine||S|VO|Y
C0694750|T121|38|CVX|rubella/mumps||S|PF|N
C0694750|T129|38|CVX|rubella/mumps||S|PF|N
C0694750|T121|38|HL7V2.5|rubella/mumps||S|PF|N
C0694750|T129|38|HL7V2.5|rubella/mumps||S|PF|N
C0694750|T121|38|HL7V3.0|rubella/mumps||S|PF|Y
C0694750|T129|38|HL7V3.0|rubella/mumps||S|PF|Y
C0694750|T121|d03005|MMSL|mumps-rubella virus vaccine||S|PF|Y
C0694750|T129|d03005|MMSL|mumps-rubella virus vaccine||S|PF|Y
C0694750|T121|NOCODE|MTH|Rubella/Mumps vaccine||P|PF|Y
C0694750|T129|NOCODE|MTH|Rubella/Mumps vaccine||P|PF|Y
C0694750|T121|412300006|SNOMEDCT_US|Rubella and mumps vaccine||P|VO|Y
C0694750|T129|412300006|SNOMEDCT_US|Rubella and mumps vaccine||P|VO|Y
C0694750|T121|412300006|SNOMEDCT_US|Rubella and mumps vaccine (substance)||S|PF|Y
C0694750|T129|412300006|SNOMEDCT_US|Rubella and mumps vaccine (substance)||S|PF|Y
C0694751|T121|41|CVX|typhoid vaccine, parenteral, other than acetone-killed, dried||P|PF|Y
C0694751|T129|41|CVX|typhoid vaccine, parenteral, other than acetone-killed, dried||P|PF|Y
C0694751|T121|41|CVX|typhoid, parenteral||S|PF|N
C0694751|T129|41|CVX|typhoid, parenteral||S|PF|N
C0694751|T121|41|HL7V2.5|typhoid, parenteral||S|PF|N
C0694751|T129|41|HL7V2.5|typhoid, parenteral||S|PF|N
C0694751|T121|41|HL7V3.0|typhoid, parenteral||S|PF|Y
C0694751|T129|41|HL7V3.0|typhoid, parenteral||S|PF|Y
C0695129|T121|90476|CPT|ADENOVIRUS VACCINE TYPE 4||S|PF|Y
C0695129|T129|90476|CPT|ADENOVIRUS VACCINE TYPE 4||S|PF|Y
C0695129|T121|90476|CPT|ADENOVIRUS VACCINE TYPE 4 LIVE ORAL||S|PF|Y
C0695129|T129|90476|CPT|ADENOVIRUS VACCINE TYPE 4 LIVE ORAL||S|PF|Y
C0695129|T121|90476|CPT|Adenovirus vaccine, type 4, live, for oral use||S|PF|Y
C0695129|T129|90476|CPT|Adenovirus vaccine, type 4, live, for oral use||S|PF|Y
C0695129|T121|54|CVX|adenovirus vaccine, type 4, live, oral||S|VC|Y
C0695129|T129|54|CVX|adenovirus vaccine, type 4, live, oral||S|VC|Y
C0695129|T121|54|CVX|adenovirus, type 4||S|PF|N
C0695129|T129|54|CVX|adenovirus, type 4||S|PF|N
C0695129|T121|90476|HCPT|Adenovirus vaccine type 4||S|VC|Y
C0695129|T129|90476|HCPT|Adenovirus vaccine type 4||S|VC|Y
C0695129|T121|54|HL7V2.5|adenovirus, type 4||S|PF|N
C0695129|T129|54|HL7V2.5|adenovirus, type 4||S|PF|N
C0695129|T121|54|HL7V3.0|adenovirus, type 4||S|PF|Y
C0695129|T129|54|HL7V3.0|adenovirus, type 4||S|PF|Y
C0695129|T121|133325|MEDCIN|live adenovirus type 4 vaccine for oral use||S|VCW|Y
C0695129|T129|133325|MEDCIN|live adenovirus type 4 vaccine for oral use||S|VCW|Y
C0695129|T121|133325|MEDCIN|live adenovirus type 4 vaccine for oral use (medication)||S|PF|Y
C0695129|T129|133325|MEDCIN|live adenovirus type 4 vaccine for oral use (medication)||S|PF|Y
C0695129|T121|133325|MEDCIN|vaccines adenovirus type 4 live, for oral use||S|VO|Y
C0695129|T129|133325|MEDCIN|vaccines adenovirus type 4 live, for oral use||S|VO|Y
C0695129|T121|442560004|SNOMEDCT_US|Live adenovirus type 4 vaccine oral dosage form||P|PF|Y
C0695129|T129|442560004|SNOMEDCT_US|Live adenovirus type 4 vaccine oral dosage form||P|PF|Y
C0695129|T121|442560004|SNOMEDCT_US|Live adenovirus type 4 vaccine oral dosage form (product)||S|PF|Y
C0695129|T129|442560004|SNOMEDCT_US|Live adenovirus type 4 vaccine oral dosage form (product)||S|PF|Y
C0695130|T121|90477|CPT|ADENOVIRUS VACCINE TYPE 7||S|PF|Y
C0695130|T129|90477|CPT|ADENOVIRUS VACCINE TYPE 7||S|PF|Y
C0695130|T121|90477|CPT|ADENOVIRUS VACCINE TYPE 7 LIVE FOR ORAL||S|PF|Y
C0695130|T129|90477|CPT|ADENOVIRUS VACCINE TYPE 7 LIVE FOR ORAL||S|PF|Y
C0695130|T121|90477|CPT|Adenovirus vaccine, type 7, live, for oral use||S|PF|Y
C0695130|T129|90477|CPT|Adenovirus vaccine, type 7, live, for oral use||S|PF|Y
C0695130|T121|55|CVX|adenovirus vaccine, type 7, live, oral||S|VO|Y
C0695130|T129|55|CVX|adenovirus vaccine, type 7, live, oral||S|VO|Y
C0695130|T121|55|CVX|adenovirus, type 7||S|PF|N
C0695130|T129|55|CVX|adenovirus, type 7||S|PF|N
C0695130|T121|90477|HCPT|Adenovirus vaccine type 7||S|VC|Y
C0695130|T129|90477|HCPT|Adenovirus vaccine type 7||S|VC|Y
C0695130|T121|55|HL7V2.5|adenovirus, type 7||S|PF|N
C0695130|T129|55|HL7V2.5|adenovirus, type 7||S|PF|N
C0695130|T121|55|HL7V3.0|adenovirus, type 7||S|PF|Y
C0695130|T129|55|HL7V3.0|adenovirus, type 7||S|PF|Y
C0695130|T121|133326|MEDCIN|live adenovirus type 7 vaccine for oral use||S|VCW|Y
C0695130|T129|133326|MEDCIN|live adenovirus type 7 vaccine for oral use||S|VCW|Y
C0695130|T121|133326|MEDCIN|live adenovirus type 7 vaccine for oral use (medication)||S|PF|Y
C0695130|T129|133326|MEDCIN|live adenovirus type 7 vaccine for oral use (medication)||S|PF|Y
C0695130|T121|133326|MEDCIN|vaccines adenovirus type 7 live, for oral use||S|VO|Y
C0695130|T129|133326|MEDCIN|vaccines adenovirus type 7 live, for oral use||S|VO|Y
C0695130|T121|442561000|SNOMEDCT_US|Live adenovirus type 7 vaccine oral dosage form||P|PF|Y
C0695130|T129|442561000|SNOMEDCT_US|Live adenovirus type 7 vaccine oral dosage form||P|PF|Y
C0695130|T121|442561000|SNOMEDCT_US|Live adenovirus type 7 vaccine oral dosage form (product)||S|PF|Y
C0695130|T129|442561000|SNOMEDCT_US|Live adenovirus type 7 vaccine oral dosage form (product)||S|PF|Y
C0717360|T121|66|CVX|Lyme disease||S|PF|N
C0717360|T129|66|CVX|Lyme disease||S|PF|N
C0717360|T121|66|CVX|Lyme disease vaccine||P|VC|N
C0717360|T129|66|CVX|Lyme disease vaccine||P|VC|N
C0717360|T121|66|HL7V2.5|Lyme disease||S|PF|N
C0717360|T129|66|HL7V2.5|Lyme disease||S|PF|N
C0717360|T121|66|HL7V3.0|Lyme disease||S|PF|Y
C0717360|T129|66|HL7V3.0|Lyme disease||S|PF|Y
C0717360|T121|d04379|MMSL|Lyme disease vaccine||P|VC|N
C0717360|T129|d04379|MMSL|Lyme disease vaccine||P|VC|N
C0717360|T121|D022123|MSH|LYME DIS VACCINES||S|PF|Y
C0717360|T129|D022123|MSH|LYME DIS VACCINES||S|PF|Y
C0717360|T121|D022123|MSH|Lyme Disease Vaccines||P|VO|Y
C0717360|T129|D022123|MSH|Lyme Disease Vaccines||P|VO|Y
C0717360|T121|D022123|MSH|VACCINES LYME DIS||S|VW|Y
C0717360|T129|D022123|MSH|VACCINES LYME DIS||S|VW|Y
C0717360|T121|D022123|MSH|Vaccines, Lyme Disease||P|VO|Y
C0717360|T129|D022123|MSH|Vaccines, Lyme Disease||P|VO|Y
C0717360|T121|NOCODE|MTH|Lyme Disease Vaccine||P|PF|Y
C0717360|T129|NOCODE|MTH|Lyme Disease Vaccine||P|PF|Y
C0717360|T121|N0000148598|NDFRT|LYME DISEASE VACCINE||P|VC|N
C0717360|T129|N0000148598|NDFRT|LYME DISEASE VACCINE||P|VC|N
C0717360|T121|N0000170888|NDFRT|Lyme Disease Vaccines||P|VO|N
C0717360|T129|N0000170888|NDFRT|Lyme Disease Vaccines||P|VO|N
C0717360|T121|N0000170888|NDFRT|Lyme Disease Vaccines [Chemical/Ingredient]||S|PF|Y
C0717360|T129|N0000170888|NDFRT|Lyme Disease Vaccines [Chemical/Ingredient]||S|PF|Y
C0717360|T121|N0000170888|NDFRT|Vaccines, Lyme Disease||P|VO|N
C0717360|T129|N0000170888|NDFRT|Vaccines, Lyme Disease||P|VO|N
C0717360|T121|214177|RXNORM|Lyme Disease Vaccine||P|PF|N
C0717360|T129|214177|RXNORM|Lyme Disease Vaccine||P|PF|N
C0717360|T121|116083002|SNOMEDCT_US|Lyme disease vaccine||P|VC|Y
C0717360|T129|116083002|SNOMEDCT_US|Lyme disease vaccine||P|VC|Y
C0717360|T121|116083002|SNOMEDCT_US|Lyme disease vaccine (product)||S|PF|Y
C0717360|T129|116083002|SNOMEDCT_US|Lyme disease vaccine (product)||S|PF|Y
C0717360|T121|116083002|SNOMEDCT_US|Lyme disease vaccine (substance)||S|PF|N
C0717360|T129|116083002|SNOMEDCT_US|Lyme disease vaccine (substance)||S|PF|N
C0717360|T121|397236006|SNOMEDCT_US|Lyme disease vaccine||P|VC|N
C0717360|T129|397236006|SNOMEDCT_US|Lyme disease vaccine||P|VC|N
C0717360|T121|397236006|SNOMEDCT_US|Lyme disease vaccine (substance)||S|PF|Y
C0717360|T129|397236006|SNOMEDCT_US|Lyme disease vaccine (substance)||S|PF|Y
C0717360|T121|4021145|VANDF|LYME DISEASE VACCINE||P|VC|Y
C0717360|T129|4021145|VANDF|LYME DISEASE VACCINE||P|VC|Y
C0718003|T121|90713|CPT|Inactivated poliovirus vaccine||P|VCW|N
C0718003|T129|90713|CPT|Inactivated poliovirus vaccine||P|VCW|N
C0718003|T121|10|CVX|IPV||S|PF|N
C0718003|T129|10|CVX|IPV||S|PF|N
C0718003|T121|10|CVX|poliovirus vaccine, inactivated||P|VC|N
C0718003|T129|10|CVX|poliovirus vaccine, inactivated||P|VC|N
C0718003|T121|10|HL7V2.5|IPV||S|PF|N
C0718003|T129|10|HL7V2.5|IPV||S|PF|N
C0718003|T121|10|HL7V3.0|IPV||S|PF|N
C0718003|T129|10|HL7V3.0|IPV||S|PF|N
C0718003|T121|LP91385-2|LNC|Inactivated poliovirus vaccine||P|VCW|N
C0718003|T129|LP91385-2|LNC|Inactivated poliovirus vaccine||P|VCW|N
C0718003|T121|197498|MEDCIN|diphtheria + tetanus toxoid + inactivated polio vaccine (IPV)||S|PF|Y
C0718003|T129|197498|MEDCIN|diphtheria + tetanus toxoid + inactivated polio vaccine (IPV)||S|PF|Y
C0718003|T121|197498|MEDCIN|diphtheria + tetanus toxoid + inactivated polio vaccine (IPV) (medication)||S|PF|Y
C0718003|T129|197498|MEDCIN|diphtheria + tetanus toxoid + inactivated polio vaccine (IPV) (medication)||S|PF|Y
C0718003|T121|197498|MEDCIN|diphtheria + tetanus toxoid + poliovirus vaccine, IPV||S|PF|Y
C0718003|T129|197498|MEDCIN|diphtheria + tetanus toxoid + poliovirus vaccine, IPV||S|PF|Y
C0718003|T121|44452|MEDCIN|inactivated poliovirus vaccine, IPV||S|PF|Y
C0718003|T129|44452|MEDCIN|inactivated poliovirus vaccine, IPV||S|PF|Y
C0718003|T121|44452|MEDCIN|inactivated poliovirus vaccine, IPV (medication)||S|PF|Y
C0718003|T129|44452|MEDCIN|inactivated poliovirus vaccine, IPV (medication)||S|PF|Y
C0718003|T121|12383|MMSL|poliomyelitis vaccine (inactivated)||S|VCW|Y
C0718003|T129|12383|MMSL|poliomyelitis vaccine (inactivated)||S|VCW|Y
C0718003|T121|7423|MMSL|polio vaccine, inactivated (monkey kidney)||S|PF|Y
C0718003|T129|7423|MMSL|polio vaccine, inactivated (monkey kidney)||S|PF|Y
C0718003|T121|d01163|MMSL|poliovirus vaccine, inactivated||P|VC|Y
C0718003|T129|d01163|MMSL|poliovirus vaccine, inactivated||P|VC|Y
C0718003|T121|D011054|MSH|Inactivated Poliovirus Vaccine||P|VW|N
C0718003|T129|D011054|MSH|Inactivated Poliovirus Vaccine||P|VW|N
C0718003|T121|D011054|MSH|Poliovirus Vaccine, Inactivated||P|PF|N
C0718003|T129|D011054|MSH|Poliovirus Vaccine, Inactivated||P|PF|N
C0718003|T121|D011054|MSH|Vaccine, Inactivated Poliovirus||P|VW|Y
C0718003|T129|D011054|MSH|Vaccine, Inactivated Poliovirus||P|VW|Y
C0718003|T121|NOCODE|MTH|Poliovirus Vaccine, Inactivated||P|PF|Y
C0718003|T129|NOCODE|MTH|Poliovirus Vaccine, Inactivated||P|PF|Y
C0718003|T121|C91715|NCI|Inactivated Poliovirus Vaccine||P|VW|Y
C0718003|T129|C91715|NCI|Inactivated Poliovirus Vaccine||P|VW|Y
C0718003|T121|C91715|NCI|IPV||S|PF|N
C0718003|T129|C91715|NCI|IPV||S|PF|N
C0718003|T121|C91715|NCI_NICHD|Inactivated Poliovirus Vaccine||P|VW|N
C0718003|T129|C91715|NCI_NICHD|Inactivated Poliovirus Vaccine||P|VW|N
C0718003|T121|C91715|NCI_NICHD|IPV||S|PF|Y
C0718003|T129|C91715|NCI_NICHD|IPV||S|PF|Y
C0718003|T121|N0000148276|NDFRT|POLIOVIRUS VACCINE INACTIVATED||P|VC|N
C0718003|T129|N0000148276|NDFRT|POLIOVIRUS VACCINE INACTIVATED||P|VC|N
C0718003|T121|N0000170917|NDFRT|Poliovirus Vaccine, Inactivated||P|PF|N
C0718003|T129|N0000170917|NDFRT|Poliovirus Vaccine, Inactivated||P|PF|N
C0718003|T121|N0000170917|NDFRT|Poliovirus Vaccine, Inactivated [Chemical/Ingredient]||S|PF|Y
C0718003|T129|N0000170917|NDFRT|Poliovirus Vaccine, Inactivated [Chemical/Ingredient]||S|PF|Y
C0718003|T121|125688000|SNOMEDCT_US|Inactivated poliomyelitis vaccine||S|PF|Y
C0718003|T129|125688000|SNOMEDCT_US|Inactivated poliomyelitis vaccine||S|PF|Y
C0718003|T121|125688000|SNOMEDCT_US|Inactivated poliovirus vaccine||P|VCW|Y
C0718003|T129|125688000|SNOMEDCT_US|Inactivated poliovirus vaccine||P|VCW|Y
C0718003|T121|125688000|SNOMEDCT_US|Inactivated poliovirus vaccine (product)||S|PF|Y
C0718003|T129|125688000|SNOMEDCT_US|Inactivated poliovirus vaccine (product)||S|PF|Y
C0718003|T121|125688000|SNOMEDCT_US|Inactivated poliovirus vaccine (substance)||S|PF|N
C0718003|T129|125688000|SNOMEDCT_US|Inactivated poliovirus vaccine (substance)||S|PF|N
C0718003|T121|125688000|SNOMEDCT_US|Pol/Vac (inact)||S|PF|Y
C0718003|T129|125688000|SNOMEDCT_US|Pol/Vac (inact)||S|PF|Y
C0718003|T121|396435000|SNOMEDCT_US|Inactivated poliomyelitis vaccine||S|PF|N
C0718003|T129|396435000|SNOMEDCT_US|Inactivated poliomyelitis vaccine||S|PF|N
C0718003|T121|396435000|SNOMEDCT_US|Inactivated poliovirus vaccine||P|VCW|N
C0718003|T129|396435000|SNOMEDCT_US|Inactivated poliovirus vaccine||P|VCW|N
C0718003|T121|396435000|SNOMEDCT_US|Inactivated poliovirus vaccine (substance)||S|PF|Y
C0718003|T129|396435000|SNOMEDCT_US|Inactivated poliovirus vaccine (substance)||S|PF|Y
C0718003|T121|396435000|SNOMEDCT_US|Pol/Vac (inact)||S|PF|N
C0718003|T129|396435000|SNOMEDCT_US|Pol/Vac (inact)||S|PF|N
C0718003|T121|4020575|VANDF|POLIOVIRUS VACCINE INACTIVATED||P|VC|Y
C0718003|T129|4020575|VANDF|POLIOVIRUS VACCINE INACTIVATED||P|VC|Y
C0770715|T121|78|CVX|tularemia vaccine||P|PF|N
C0770715|T121|78|CVX|tularemia vaccine||P|PF|Y
C0770715|T109|78|CVX|tularemia vaccine||P|PF|N
C0770715|T109|78|CVX|tularemia vaccine||P|PF|Y
C0770715|T129|78|CVX|tularemia vaccine||P|PF|N
C0770715|T129|78|CVX|tularemia vaccine||P|PF|Y
C0770715|T121|78|HL7V2.5|tularemia vaccine||P|PF|N
C0770715|T109|78|HL7V2.5|tularemia vaccine||P|PF|N
C0770715|T129|78|HL7V2.5|tularemia vaccine||P|PF|N
C0770715|T121|78|HL7V3.0|tularemia vaccine||P|PF|N
C0770715|T109|78|HL7V3.0|tularemia vaccine||P|PF|N
C0770715|T129|78|HL7V3.0|tularemia vaccine||P|PF|N
C0770715|T121|133287|MEDCIN|tularemia vaccine||P|PF|N
C0770715|T109|133287|MEDCIN|tularemia vaccine||P|PF|N
C0770715|T129|133287|MEDCIN|tularemia vaccine||P|PF|N
C0770715|T121|133287|MEDCIN|tularemia vaccine (medication)||S|PF|Y
C0770715|T109|133287|MEDCIN|tularemia vaccine (medication)||S|PF|Y
C0770715|T129|133287|MEDCIN|tularemia vaccine (medication)||S|PF|Y
C0796561|T121|68|CVX|melanoma||S|PF|N
C0796561|T129|68|CVX|melanoma||S|PF|N
C0796561|T121|68|CVX|melanoma vaccine||P|VC|N
C0796561|T129|68|CVX|melanoma vaccine||P|VC|N
C0796561|T121|68|HL7V2.5|melanoma||S|PF|N
C0796561|T129|68|HL7V2.5|melanoma||S|PF|N
C0796561|T121|68|HL7V3.0|melanoma||S|PF|Y
C0796561|T129|68|HL7V3.0|melanoma||S|PF|Y
C0796561|T121|NOCODE|MTH|Melanoma vaccine||P|PF|Y
C0796561|T129|NOCODE|MTH|Melanoma vaccine||P|PF|Y
C0796561|T121|C2517|NCI|Melanoma Vaccine||P|VC|Y
C0796561|T129|C2517|NCI|Melanoma Vaccine||P|VC|Y
C0796561|T121|CDR0000046293|NCI_NCI-GLOSS|melanoma vaccine||P|VC|Y
C0796561|T129|CDR0000046293|NCI_NCI-GLOSS|melanoma vaccine||P|VC|Y
C0796561|T121|373869007|SNOMEDCT_US|Melanoma vaccine||P|PF|N
C0796561|T129|373869007|SNOMEDCT_US|Melanoma vaccine||P|PF|N
C0796561|T121|373869007|SNOMEDCT_US|Melanoma vaccine (product)||S|PF|Y
C0796561|T129|373869007|SNOMEDCT_US|Melanoma vaccine (product)||S|PF|Y
C0796561|T121|428026004|SNOMEDCT_US|Melanoma vaccine||P|PF|N
C0796561|T129|428026004|SNOMEDCT_US|Melanoma vaccine||P|PF|N
C0796561|T121|428026004|SNOMEDCT_US|Melanoma vaccine (substance)||S|PF|Y
C0796561|T129|428026004|SNOMEDCT_US|Melanoma vaccine (substance)||S|PF|Y
C0872996|T121|70|CVX|Q fever||S|PF|N
C0872996|T129|70|CVX|Q fever||S|PF|N
C0872996|T121|70|CVX|Q fever vaccine||P|PF|N
C0872996|T129|70|CVX|Q fever vaccine||P|PF|N
C0872996|T121|70|HL7V2.5|Q fever||S|PF|N
C0872996|T129|70|HL7V2.5|Q fever||S|PF|N
C0872996|T121|70|HL7V3.0|Q fever||S|PF|Y
C0872996|T129|70|HL7V3.0|Q fever||S|PF|Y
C0872996|T121|NOCODE|MTH|Q fever vaccine||P|PF|Y
C0872996|T129|NOCODE|MTH|Q fever vaccine||P|PF|Y
C0872996|T121|427533008|SNOMEDCT_US|Q fever vaccine||P|PF|N
C0872996|T129|427533008|SNOMEDCT_US|Q fever vaccine||P|PF|N
C0872996|T121|427533008|SNOMEDCT_US|Q fever vaccine (product)||S|PF|Y
C0872996|T129|427533008|SNOMEDCT_US|Q fever vaccine (product)||S|PF|Y
C0872996|T121|427674002|SNOMEDCT_US|Q fever vaccine||P|PF|N
C0872996|T129|427674002|SNOMEDCT_US|Q fever vaccine||P|PF|N
C0872996|T121|427674002|SNOMEDCT_US|Q fever vaccine (substance)||S|PF|Y
C0872996|T129|427674002|SNOMEDCT_US|Q fever vaccine (substance)||S|PF|Y
C0915344|T116|103|CVX|meningococcal C conjugate||S|PF|N
C0915344|T129|103|CVX|meningococcal C conjugate||S|PF|N
C0915344|T121|103|CVX|meningococcal C conjugate||S|PF|N
C0915344|T116|103|CVX|meningococcal C conjugate vaccine||S|VC|N
C0915344|T129|103|CVX|meningococcal C conjugate vaccine||S|VC|N
C0915344|T121|103|CVX|meningococcal C conjugate vaccine||S|VC|N
C0915344|T116|103|HL7V2.5|meningococcal C conjugate||S|PF|Y
C0915344|T129|103|HL7V2.5|meningococcal C conjugate||S|PF|Y
C0915344|T121|103|HL7V2.5|meningococcal C conjugate||S|PF|Y
C0915344|T116|257908|MEDCIN|meningococcal conjugate vaccine serogroup C||P|VW|Y
C0915344|T129|257908|MEDCIN|meningococcal conjugate vaccine serogroup C||P|VW|Y
C0915344|T121|257908|MEDCIN|meningococcal conjugate vaccine serogroup C||P|VW|Y
C0915344|T116|257908|MEDCIN|meningococcal conjugate vaccine serogroup C (medication)||S|PF|Y
C0915344|T129|257908|MEDCIN|meningococcal conjugate vaccine serogroup C (medication)||S|PF|Y
C0915344|T121|257908|MEDCIN|meningococcal conjugate vaccine serogroup C (medication)||S|PF|Y
C0915344|T116|C410218|MSH|CMC vaccine||S|PF|Y
C0915344|T129|C410218|MSH|CMC vaccine||S|PF|Y
C0915344|T121|C410218|MSH|CMC vaccine||S|PF|Y
C0915344|T116|C410218|MSH|meningococcal C conjugate vaccine||S|VC|Y
C0915344|T129|C410218|MSH|meningococcal C conjugate vaccine||S|VC|Y
C0915344|T121|C410218|MSH|meningococcal C conjugate vaccine||S|VC|Y
C0915344|T116|C410218|MSH|meningococcal type C conjugate vaccine||S|PF|Y
C0915344|T129|C410218|MSH|meningococcal type C conjugate vaccine||S|PF|Y
C0915344|T121|C410218|MSH|meningococcal type C conjugate vaccine||S|PF|Y
C0915344|T116|C410218|MSH|serogroup C meningococcal conjugate vaccine||P|PF|Y
C0915344|T129|C410218|MSH|serogroup C meningococcal conjugate vaccine||P|PF|Y
C0915344|T121|C410218|MSH|serogroup C meningococcal conjugate vaccine||P|PF|Y
C0915344|T116|359068008|SNOMEDCT_US|Meningococcal C conjugate vaccine||S|PF|Y
C0915344|T129|359068008|SNOMEDCT_US|Meningococcal C conjugate vaccine||S|PF|Y
C0915344|T121|359068008|SNOMEDCT_US|Meningococcal C conjugate vaccine||S|PF|Y
C0915344|T116|359068008|SNOMEDCT_US|Meningococcal C conjugate vaccine (product)||S|PF|Y
C0915344|T129|359068008|SNOMEDCT_US|Meningococcal C conjugate vaccine (product)||S|PF|Y
C0915344|T121|359068008|SNOMEDCT_US|Meningococcal C conjugate vaccine (product)||S|PF|Y
C0915344|T116|359068008|SNOMEDCT_US|Meningococcal C conjugate vaccine (substance)||S|PF|Y
C0915344|T129|359068008|SNOMEDCT_US|Meningococcal C conjugate vaccine (substance)||S|PF|Y
C0915344|T121|359068008|SNOMEDCT_US|Meningococcal C conjugate vaccine (substance)||S|PF|Y
C0961101|T121|90732|CPT|Pneumococcal polysaccharide vaccine, 23-valent||S|PF|Y
C0961101|T129|90732|CPT|Pneumococcal polysaccharide vaccine, 23-valent||S|PF|Y
C0961101|T121|33|CVX|pneumococcal polysaccharide PPV23||S|PF|Y
C0961101|T129|33|CVX|pneumococcal polysaccharide PPV23||S|PF|Y
C0961101|T121|33|CVX|pneumococcal polysaccharide vaccine, 23 valent||S|VC|Y
C0961101|T129|33|CVX|pneumococcal polysaccharide vaccine, 23 valent||S|VC|Y
C0961101|T121|C414006|MSH|23-valent pneumococcal capsular polysaccharide vaccine||P|PF|N
C0961101|T129|C414006|MSH|23-valent pneumococcal capsular polysaccharide vaccine||P|PF|N
C0961101|T121|C414006|MSH|23-valent vaccine||S|PF|Y
C0961101|T129|C414006|MSH|23-valent vaccine||S|PF|Y
C0961101|T121|NOCODE|MTH|23-valent pneumococcal capsular polysaccharide vaccine||P|PF|Y
C0961101|T129|NOCODE|MTH|23-valent pneumococcal capsular polysaccharide vaccine||P|PF|Y
C0961101|T121|C1643|NCI_NICHD|PCV 23||S|PF|Y
C0961101|T129|C1643|NCI_NICHD|PCV 23||S|PF|Y
C0961101|T121|C1643|NCI_NICHD|Pneumococcal 23-valent Polysaccharide Vaccine||S|VCW|Y
C0961101|T129|C1643|NCI_NICHD|Pneumococcal 23-valent Polysaccharide Vaccine||S|VCW|Y
C0979582|T121|100|CVX|pneumococcal conjugate PCV 7||S|PF|Y
C0979582|T129|100|CVX|pneumococcal conjugate PCV 7||S|PF|Y
C0979582|T121|100|CVX|pneumococcal conjugate vaccine, 7 valent||P|VCW|Y
C0979582|T129|100|CVX|pneumococcal conjugate vaccine, 7 valent||P|VCW|Y
C0979582|T121|d04920|MMSL|pneumococcal 7-valent conjugate vaccine||P|VC|Y
C0979582|T129|d04920|MMSL|pneumococcal 7-valent conjugate vaccine||P|VC|Y
C0979582|T121|C38141|NCI|Pneumococcal 7-Valent Conjugate Vaccine||P|VC|Y
C0979582|T129|C38141|NCI|Pneumococcal 7-Valent Conjugate Vaccine||P|VC|Y
C0979582|T121|C38141|NCI|Pneumococcal 7-valent Conjugate Vaccine (Diphtheria CRM197 Protein)||S|PF|Y
C0979582|T129|C38141|NCI|Pneumococcal 7-valent Conjugate Vaccine (Diphtheria CRM197 Protein)||S|PF|Y
C0979582|T121|C38141|NCI_NICHD|PCV 7||S|PF|Y
C0979582|T129|C38141|NCI_NICHD|PCV 7||S|PF|Y
C0979582|T121|C38141|NCI_NICHD|Pneumococcal 7-Valent Conjugate Vaccine||P|VC|N
C0979582|T129|C38141|NCI_NICHD|Pneumococcal 7-Valent Conjugate Vaccine||P|VC|N
C0979582|T121|N0000162690|NDFRT|PNEUMOCOCCAL 7-VALENT CONJUGATE VACCINE||P|VC|N
C0979582|T129|N0000162690|NDFRT|PNEUMOCOCCAL 7-VALENT CONJUGATE VACCINE||P|VC|N
C0979582|T121|N0000162690|NDFRT|PNEUMOCOCCAL 7-VALENT CONJUGATE VACCINE [VA Product]||S|PF|Y
C0979582|T129|N0000162690|NDFRT|PNEUMOCOCCAL 7-VALENT CONJUGATE VACCINE [VA Product]||S|PF|Y
C0979582|T121|125714002|SNOMEDCT_US|Pneumococcal 7-valent conjugate vaccine||P|PF|Y
C0979582|T129|125714002|SNOMEDCT_US|Pneumococcal 7-valent conjugate vaccine||P|PF|Y
C0979582|T121|125714002|SNOMEDCT_US|Pneumococcal 7-valent conjugate vaccine (product)||S|PF|Y
C0979582|T129|125714002|SNOMEDCT_US|Pneumococcal 7-valent conjugate vaccine (product)||S|PF|Y
C0979582|T121|125714002|SNOMEDCT_US|Pneumococcal 7-valent conjugate vaccine (substance)||S|PF|Y
C0979582|T129|125714002|SNOMEDCT_US|Pneumococcal 7-valent conjugate vaccine (substance)||S|PF|Y
C0979582|T121|4014972|VANDF|PNEUMOCOCCAL 7-VALENT CONJUGATE VACCINE||P|VC|N
C0979582|T121|4014972|VANDF|PNEUMOCOCCAL 7-VALENT CONJUGATE VACCINE||P|VC|Y
C0979582|T129|4014972|VANDF|PNEUMOCOCCAL 7-VALENT CONJUGATE VACCINE||P|VC|N
C0979582|T129|4014972|VANDF|PNEUMOCOCCAL 7-VALENT CONJUGATE VACCINE||P|VC|Y
C1170008|T121|90636|CPT|Hepatitis A and hepatitis B vaccine||P|VO|Y
C1170008|T129|90636|CPT|Hepatitis A and hepatitis B vaccine||P|VO|Y
C1170008|T121|104|CVX|Hep A-Hep B||S|PF|N
C1170008|T129|104|CVX|Hep A-Hep B||S|PF|N
C1170008|T121|104|CVX|hepatitis A and hepatitis B vaccine||P|VO|Y
C1170008|T129|104|CVX|hepatitis A and hepatitis B vaccine||P|VO|Y
C1170008|T121|104|HL7V2.5|Hep A-Hep B||S|PF|Y
C1170008|T129|104|HL7V2.5|Hep A-Hep B||S|PF|Y
C1170008|T121|d04685|MMSL|hepatitis A-hepatitis B vaccine||P|PF|Y
C1170008|T129|d04685|MMSL|hepatitis A-hepatitis B vaccine||P|PF|Y
C1249366|T121|18|CVX|rabies vaccine, for intramuscular injection||P|PF|Y
C1249366|T129|18|CVX|rabies vaccine, for intramuscular injection||P|PF|Y
C1249366|T121|18|CVX|rabies, intramuscular injection||S|PF|N
C1249366|T129|18|CVX|rabies, intramuscular injection||S|PF|N
C1249366|T121|18|HL7V2.5|rabies, intramuscular injection||S|PF|N
C1249366|T129|18|HL7V2.5|rabies, intramuscular injection||S|PF|N
C1249366|T121|18|HL7V3.0|rabies, intramuscular injection||S|PF|Y
C1249366|T129|18|HL7V3.0|rabies, intramuscular injection||S|PF|Y
C1548467|T129|102|CVX|DTaP/DTP-Hib-Hep B||S|PF|Y
C1548467|T121|102|CVX|DTaP/DTP-Hib-Hep B||S|PF|Y
C1548467|T129|102|CVX|DTP- Haemophilus influenzae type b conjugate and hepatitis b vaccine||P|PF|Y
C1548467|T121|102|CVX|DTP- Haemophilus influenzae type b conjugate and hepatitis b vaccine||P|PF|Y
C1548467|T129|102|HL7V2.5|DTP-Hib-Hep B||S|PF|Y
C1548467|T121|102|HL7V2.5|DTP-Hib-Hep B||S|PF|Y
C1548470|T129|105|CVX|vaccinia (smallpox) diluted||S|PF|Y
C1548470|T121|105|CVX|vaccinia (smallpox) diluted||S|PF|Y
C1548470|T129|105|CVX|vaccinia (smallpox) vaccine, diluted||P|PF|Y
C1548470|T121|105|CVX|vaccinia (smallpox) vaccine, diluted||P|PF|Y
C1548470|T129|105|HL7V2.5|smallpox, diluted||S|PF|Y
C1548470|T121|105|HL7V2.5|smallpox, diluted||S|PF|Y
C1548471|T129|106|CVX|diphtheria, tetanus toxoids and acellular pertussis vaccine, 5 pertussis antigens||P|PF|Y
C1548471|T121|106|CVX|diphtheria, tetanus toxoids and acellular pertussis vaccine, 5 pertussis antigens||P|PF|Y
C1548471|T129|106|CVX|DTaP, 5 pertussis antigens||S|PF|N
C1548471|T121|106|CVX|DTaP, 5 pertussis antigens||S|PF|N
C1548471|T129|106|HL7V2.5|DTaP, 5 pertussis antigens||S|PF|Y
C1548471|T121|106|HL7V2.5|DTaP, 5 pertussis antigens||S|PF|Y
C1548473|T121|34|CVX|rabies immune globulin||P|PF|N
C1548473|T129|34|CVX|rabies immune globulin||P|PF|N
C1548473|T116|34|CVX|rabies immune globulin||P|PF|N
C1548473|T121|34|CVX|RIG||S|PF|N
C1548473|T129|34|CVX|RIG||S|PF|N
C1548473|T116|34|CVX|RIG||S|PF|N
C1548473|T121|34|HL7V2.5|RIG||S|PF|N
C1548473|T129|34|HL7V2.5|RIG||S|PF|N
C1548473|T116|34|HL7V2.5|RIG||S|PF|N
C1548473|T121|34|HL7V3.0|RIG||S|PF|Y
C1548473|T129|34|HL7V3.0|RIG||S|PF|Y
C1548473|T116|34|HL7V3.0|RIG||S|PF|Y
C1548473|T121|133256|MEDCIN|human rabies immune globulin for intramuscular use||S|PF|Y
C1548473|T129|133256|MEDCIN|human rabies immune globulin for intramuscular use||S|PF|Y
C1548473|T116|133256|MEDCIN|human rabies immune globulin for intramuscular use||S|PF|Y
C1548473|T121|133256|MEDCIN|human rabies immune globulin for intramuscular use (medication)||S|PF|Y
C1548473|T129|133256|MEDCIN|human rabies immune globulin for intramuscular use (medication)||S|PF|Y
C1548473|T116|133256|MEDCIN|human rabies immune globulin for intramuscular use (medication)||S|PF|Y
C1548473|T121|133257|MEDCIN|human rabies immune globulin for subcutaneous use||S|PF|Y
C1548473|T129|133257|MEDCIN|human rabies immune globulin for subcutaneous use||S|PF|Y
C1548473|T116|133257|MEDCIN|human rabies immune globulin for subcutaneous use||S|PF|Y
C1548473|T121|133257|MEDCIN|human rabies immune globulin for subcutaneous use (medication)||S|PF|Y
C1548473|T129|133257|MEDCIN|human rabies immune globulin for subcutaneous use (medication)||S|PF|Y
C1548473|T116|133257|MEDCIN|human rabies immune globulin for subcutaneous use (medication)||S|PF|Y
C1548473|T121|NOCODE|MTH|rabies immune globulin||P|PF|Y
C1548473|T129|NOCODE|MTH|rabies immune globulin||P|PF|Y
C1548473|T116|NOCODE|MTH|rabies immune globulin||P|PF|Y
C1548476|T129|53|CVX|typhoid vaccine, parenteral, acetone-killed, dried (U.S. military)||P|PF|Y
C1548476|T121|53|CVX|typhoid vaccine, parenteral, acetone-killed, dried (U.S. military)||P|PF|Y
C1548476|T129|53|CVX|typhoid, parenteral, AKD (U.S. military)||S|PF|N
C1548476|T121|53|CVX|typhoid, parenteral, AKD (U.S. military)||S|PF|N
C1548476|T129|53|HL7V2.5|typhoid, parenteral, AKD (U.S. military)||S|PF|N
C1548476|T121|53|HL7V2.5|typhoid, parenteral, AKD (U.S. military)||S|PF|N
C1548476|T129|53|HL7V3.0|typhoid, parenteral, AKD (U.S. military)||S|PF|Y
C1548476|T121|53|HL7V3.0|typhoid, parenteral, AKD (U.S. military)||S|PF|Y
C1548477|T129|56|CVX|dengue fever||S|PF|N
C1548477|T121|56|CVX|dengue fever||S|PF|N
C1548477|T129|56|CVX|dengue fever vaccine||P|VC|Y
C1548477|T121|56|CVX|dengue fever vaccine||P|VC|Y
C1548477|T129|56|HL7V2.5|dengue fever||S|PF|N
C1548477|T121|56|HL7V2.5|dengue fever||S|PF|N
C1548477|T129|56|HL7V3.0|dengue fever||S|PF|Y
C1548477|T121|56|HL7V3.0|dengue fever||S|PF|Y
C1548477|T129|D053059|MSH|Dengue Vaccines||S|PF|Y
C1548477|T121|D053059|MSH|Dengue Vaccines||S|PF|Y
C1548477|T129|D053059|MSH|Vaccines, Dengue||S|VW|Y
C1548477|T121|D053059|MSH|Vaccines, Dengue||S|VW|Y
C1548477|T129|NOCODE|MTH|Dengue fever vaccine||P|PF|Y
C1548477|T121|NOCODE|MTH|Dengue fever vaccine||P|PF|Y
C1548477|T129|N0000175338|NDFRT|Dengue Vaccines||S|PF|N
C1548477|T121|N0000175338|NDFRT|Dengue Vaccines||S|PF|N
C1548477|T129|N0000175338|NDFRT|Dengue Vaccines [Chemical/Ingredient]||S|PF|Y
C1548477|T121|N0000175338|NDFRT|Dengue Vaccines [Chemical/Ingredient]||S|PF|Y
C1548478|T129|57|CVX|hantavirus||S|VC|N
C1548478|T121|57|CVX|hantavirus||S|VC|N
C1548478|T129|57|CVX|hantavirus vaccine||P|PF|N
C1548478|T121|57|CVX|hantavirus vaccine||P|PF|N
C1548478|T129|57|HL7V2.5|hantavirus||S|VC|Y
C1548478|T121|57|HL7V2.5|hantavirus||S|VC|Y
C1548478|T129|57|HL7V3.0|Hantavirus||S|PF|Y
C1548478|T121|57|HL7V3.0|Hantavirus||S|PF|Y
C1548478|T129|NOCODE|MTH|hantavirus vaccine||P|PF|Y
C1548478|T121|NOCODE|MTH|hantavirus vaccine||P|PF|Y
C1548480|T129|59|CVX|Hep E||P|PF|N
C1548480|T121|59|CVX|Hep E||P|PF|N
C1548480|T129|59|CVX|hepatitis E vaccine||S|PF|Y
C1548480|T121|59|CVX|hepatitis E vaccine||S|PF|Y
C1548480|T129|59|HL7V2.5|Hep E||P|PF|N
C1548480|T121|59|HL7V2.5|Hep E||P|PF|N
C1548480|T129|59|HL7V3.0|Hep E||P|PF|Y
C1548480|T121|59|HL7V3.0|Hep E||P|PF|Y
C1548481|T129|60|CVX|herpes simplex 2||S|PF|N
C1548481|T121|60|CVX|herpes simplex 2||S|PF|N
C1548481|T129|60|CVX|herpes simplex virus, type 2 vaccine||P|PF|N
C1548481|T121|60|CVX|herpes simplex virus, type 2 vaccine||P|PF|N
C1548481|T129|60|HL7V2.5|herpes simplex 2||S|PF|N
C1548481|T121|60|HL7V2.5|herpes simplex 2||S|PF|N
C1548481|T129|60|HL7V3.0|herpes simplex 2||S|PF|Y
C1548481|T121|60|HL7V3.0|herpes simplex 2||S|PF|Y
C1548481|T129|NOCODE|MTH|herpes simplex virus, type 2 vaccine||P|PF|Y
C1548481|T121|NOCODE|MTH|herpes simplex virus, type 2 vaccine||P|PF|Y
C1548482|T129|63|CVX|Junin virus||S|PF|N
C1548482|T121|63|CVX|Junin virus||S|PF|N
C1548482|T129|63|CVX|Junin virus vaccine||P|PF|N
C1548482|T121|63|CVX|Junin virus vaccine||P|PF|N
C1548482|T129|63|HL7V2.5|Junin virus||S|PF|N
C1548482|T121|63|HL7V2.5|Junin virus||S|PF|N
C1548482|T129|63|HL7V3.0|Junin virus||S|PF|Y
C1548482|T121|63|HL7V3.0|Junin virus||S|PF|Y
C1548482|T129|NOCODE|MTH|Junin virus vaccine||P|PF|Y
C1548482|T121|NOCODE|MTH|Junin virus vaccine||P|PF|Y
C1548483|T129|64|CVX|leishmaniasis||S|PF|N
C1548483|T121|64|CVX|leishmaniasis||S|PF|N
C1548483|T129|64|CVX|leishmaniasis vaccine||P|VC|Y
C1548483|T121|64|CVX|leishmaniasis vaccine||P|VC|Y
C1548483|T129|64|HL7V2.5|leishmaniasis||S|PF|N
C1548483|T121|64|HL7V2.5|leishmaniasis||S|PF|N
C1548483|T129|64|HL7V3.0|leishmaniasis||S|PF|Y
C1548483|T121|64|HL7V3.0|leishmaniasis||S|PF|Y
C1548483|T129|D054332|MSH|Leishmania Vaccines||S|PF|Y
C1548483|T121|D054332|MSH|Leishmania Vaccines||S|PF|Y
C1548483|T129|D054332|MSH|Leishmaniasis Vaccines||P|VO|Y
C1548483|T121|D054332|MSH|Leishmaniasis Vaccines||P|VO|Y
C1548483|T129|D054332|MSH|Vaccines, Leishmania||S|VW|Y
C1548483|T121|D054332|MSH|Vaccines, Leishmania||S|VW|Y
C1548483|T129|D054332|MSH|Vaccines, Leishmaniasis||P|VO|Y
C1548483|T121|D054332|MSH|Vaccines, Leishmaniasis||P|VO|Y
C1548483|T129|NOCODE|MTH|Leishmaniasis Vaccine||P|PF|Y
C1548483|T121|NOCODE|MTH|Leishmaniasis Vaccine||P|PF|Y
C1548483|T129|N0000178730|NDFRT|Leishmania Vaccines||S|PF|N
C1548483|T121|N0000178730|NDFRT|Leishmania Vaccines||S|PF|N
C1548483|T129|N0000178730|NDFRT|Leishmaniasis Vaccines||P|VO|N
C1548483|T121|N0000178730|NDFRT|Leishmaniasis Vaccines||P|VO|N
C1548483|T129|N0000178730|NDFRT|Leishmaniasis Vaccines [Chemical/Ingredient]||S|PF|Y
C1548483|T121|N0000178730|NDFRT|Leishmaniasis Vaccines [Chemical/Ingredient]||S|PF|Y
C1548484|T129|72|CVX|rheumatic fever||S|PF|N
C1548484|T121|72|CVX|rheumatic fever||S|PF|N
C1548484|T129|72|CVX|rheumatic fever vaccine||P|PF|N
C1548484|T121|72|CVX|rheumatic fever vaccine||P|PF|N
C1548484|T129|72|HL7V2.5|rheumatic fever||S|PF|N
C1548484|T121|72|HL7V2.5|rheumatic fever||S|PF|N
C1548484|T129|72|HL7V3.0|rheumatic fever||S|PF|Y
C1548484|T121|72|HL7V3.0|rheumatic fever||S|PF|Y
C1548484|T129|NOCODE|MTH|rheumatic fever vaccine||P|PF|Y
C1548484|T121|NOCODE|MTH|rheumatic fever vaccine||P|PF|Y
C1548485|T129|73|CVX|Rift Valley fever||S|PF|N
C1548485|T121|73|CVX|Rift Valley fever||S|PF|N
C1548485|T129|73|CVX|Rift Valley fever vaccine||P|PF|N
C1548485|T121|73|CVX|Rift Valley fever vaccine||P|PF|N
C1548485|T129|73|HL7V2.5|Rift Valley fever||S|PF|N
C1548485|T121|73|HL7V2.5|Rift Valley fever||S|PF|N
C1548485|T129|73|HL7V3.0|Rift Valley fever||S|PF|Y
C1548485|T121|73|HL7V3.0|Rift Valley fever||S|PF|Y
C1548485|T129|NOCODE|MTH|Rift Valley fever vaccine||P|PF|Y
C1548485|T121|NOCODE|MTH|Rift Valley fever vaccine||P|PF|Y
C1548486|T129|76|CVX|Staphylococcus bacterio lysate||S|PF|N
C1548486|T121|76|CVX|Staphylococcus bacterio lysate||S|PF|N
C1548486|T129|76|CVX|Staphylococcus bacteriophage lysate||P|PF|Y
C1548486|T121|76|CVX|Staphylococcus bacteriophage lysate||P|PF|Y
C1548486|T129|76|HL7V2.5|Staphylococcus bacterio lysate||S|PF|N
C1548486|T121|76|HL7V2.5|Staphylococcus bacterio lysate||S|PF|N
C1548486|T129|76|HL7V3.0|Staphylococcus bacterio lysate||S|PF|Y
C1548486|T121|76|HL7V3.0|Staphylococcus bacterio lysate||S|PF|Y
C1548487|T129|79|CVX|vaccinia immune globulin||P|PF|N
C1548487|T121|79|CVX|vaccinia immune globulin||P|PF|N
C1548487|T109|79|CVX|vaccinia immune globulin||P|PF|N
C1548487|T129|79|HL7V2.5|vaccinia immune globulin||P|PF|N
C1548487|T121|79|HL7V2.5|vaccinia immune globulin||P|PF|N
C1548487|T109|79|HL7V2.5|vaccinia immune globulin||P|PF|N
C1548487|T129|79|HL7V3.0|vaccinia immune globulin||P|PF|N
C1548487|T121|79|HL7V3.0|vaccinia immune globulin||P|PF|N
C1548487|T109|79|HL7V3.0|vaccinia immune globulin||P|PF|N
C1548487|T129|d05490|MMSL|vaccinia immune globulin||P|PF|Y
C1548487|T121|d05490|MMSL|vaccinia immune globulin||P|PF|Y
C1548487|T109|d05490|MMSL|vaccinia immune globulin||P|PF|Y
C1548488|T129|80|CVX|VEE, live||S|PF|N
C1548488|T121|80|CVX|VEE, live||S|PF|N
C1548488|T129|80|CVX|Venezuelan equine encephalitis, live, attenuated||P|PF|Y
C1548488|T121|80|CVX|Venezuelan equine encephalitis, live, attenuated||P|PF|Y
C1548488|T129|80|HL7V2.5|VEE, live||S|PF|N
C1548488|T121|80|HL7V2.5|VEE, live||S|PF|N
C1548488|T129|80|HL7V3.0|VEE, live||S|PF|Y
C1548488|T121|80|HL7V3.0|VEE, live||S|PF|Y
C1548489|T129|81|CVX|VEE, inactivated||S|PF|N
C1548489|T121|81|CVX|VEE, inactivated||S|PF|N
C1548489|T129|81|CVX|Venezuelan equine encephalitis, inactivated||P|PF|Y
C1548489|T121|81|CVX|Venezuelan equine encephalitis, inactivated||P|PF|Y
C1548489|T129|81|HL7V2.5|VEE, inactivated||S|PF|N
C1548489|T121|81|HL7V2.5|VEE, inactivated||S|PF|N
C1548489|T129|81|HL7V3.0|VEE, inactivated||S|PF|Y
C1548489|T121|81|HL7V3.0|VEE, inactivated||S|PF|Y
C1548490|T129|82|CVX|adenovirus vaccine, unspecified formulation||P|PF|Y
C1548490|T121|82|CVX|adenovirus vaccine, unspecified formulation||P|PF|Y
C1548490|T129|82|CVX|adenovirus, unspecified formulation||S|PF|Y
C1548490|T121|82|CVX|adenovirus, unspecified formulation||S|PF|Y
C1548490|T129|82|HL7V2.5|adenovirus, NOS1||S|PF|Y
C1548490|T121|82|HL7V2.5|adenovirus, NOS1||S|PF|Y
C1548491|T129|83|CVX|Hep A, ped/adol, 2 dose||S|PF|N
C1548491|T121|83|CVX|Hep A, ped/adol, 2 dose||S|PF|N
C1548491|T129|83|CVX|hepatitis A vaccine, pediatric/adolescent dosage, 2 dose schedule||P|PF|Y
C1548491|T121|83|CVX|hepatitis A vaccine, pediatric/adolescent dosage, 2 dose schedule||P|PF|Y
C1548491|T129|83|HL7V2.5|Hep A, ped/adol, 2 dose||S|PF|N
C1548491|T121|83|HL7V2.5|Hep A, ped/adol, 2 dose||S|PF|N
C1548491|T129|83|HL7V3.0|Hep A, ped/adol, 2 dose||S|PF|Y
C1548491|T121|83|HL7V3.0|Hep A, ped/adol, 2 dose||S|PF|Y
C1548492|T129|84|CVX|Hep A, ped/adol, 3 dose||S|PF|N
C1548492|T121|84|CVX|Hep A, ped/adol, 3 dose||S|PF|N
C1548492|T129|84|CVX|hepatitis A vaccine, pediatric/adolescent dosage, 3 dose schedule||P|PF|Y
C1548492|T121|84|CVX|hepatitis A vaccine, pediatric/adolescent dosage, 3 dose schedule||P|PF|Y
C1548492|T129|84|HL7V2.5|Hep A, ped/adol, 3 dose||S|PF|N
C1548492|T121|84|HL7V2.5|Hep A, ped/adol, 3 dose||S|PF|N
C1548492|T129|84|HL7V3.0|Hep A, ped/adol, 3 dose||S|PF|Y
C1548492|T121|84|HL7V3.0|Hep A, ped/adol, 3 dose||S|PF|Y
C1548495|T129|93|CVX|respiratory syncytial virus monoclonal antibody (palivizumab), intramuscular||P|PF|Y
C1548495|T121|93|CVX|respiratory syncytial virus monoclonal antibody (palivizumab), intramuscular||P|PF|Y
C1548495|T129|93|CVX|RSV-MAb||S|VC|N
C1548495|T121|93|CVX|RSV-MAb||S|VC|N
C1548495|T129|93|HL7V2.5|RSV-MAb||S|VC|Y
C1548495|T121|93|HL7V2.5|RSV-MAb||S|VC|Y
C1548495|T129|93|HL7V3.0|RSV-Mab||S|PF|Y
C1548495|T121|93|HL7V3.0|RSV-Mab||S|PF|Y
C1548496|T074|95|CVX|TST-OT tine test||S|PF|N
C1548496|T074|95|CVX|tuberculin skin test; old tuberculin, multipuncture device||P|PF|Y
C1548496|T074|95|HL7V2.5|TST-OT tine test||S|PF|N
C1548496|T074|95|HL7V3.0|TST-OT tine test||S|PF|Y
C1548497|T121|96|CVX|TST-PPD intradermal||S|PF|N
C1548497|T129|96|CVX|TST-PPD intradermal||S|PF|N
C1548497|T121|96|CVX|tuberculin skin test; purified protein derivative solution, intradermal||P|PF|Y
C1548497|T129|96|CVX|tuberculin skin test; purified protein derivative solution, intradermal||P|PF|Y
C1548497|T121|96|HL7V2.5|TST-PPD intradermal||S|PF|N
C1548497|T129|96|HL7V2.5|TST-PPD intradermal||S|PF|N
C1548497|T121|96|HL7V3.0|TST-PPD intradermal||S|PF|Y
C1548497|T129|96|HL7V3.0|TST-PPD intradermal||S|PF|Y
C1548498|T074|97|CVX|TST-PPD tine test||S|PF|N
C1548498|T074|97|CVX|tuberculin skin test; purified protein derivative, multipuncture device||P|PF|Y
C1548498|T074|97|HL7V2.5|TST-PPD tine test||S|PF|N
C1548498|T074|97|HL7V3.0|TST-PPD tine test||S|PF|Y
C1548500|T077|99|CVX|RESERVED - do not use||P|VO|Y
C1548500|T077|99|CVX|RESERVED - do not use||P|VO|N
C1548500|T077|99|HL7V2.5|RESERVED _ do not use||P|PF|Y
C1548501|T078|998|CVX|no vaccine administered||P|PF|N
C1548501|T078|998|CVX|no vaccine administered||P|PF|Y
C1548501|T078|998|HL7V2.5|no vaccine administered||P|PF|N
C1552908|T129|42|CVX|Hep B, adolescent/high risk infant||S|PF|N
C1552908|T121|42|CVX|Hep B, adolescent/high risk infant||S|PF|N
C1552908|T129|42|CVX|hepatitis B vaccine, adolescent/high risk infant dosage||P|PF|Y
C1552908|T121|42|CVX|hepatitis B vaccine, adolescent/high risk infant dosage||P|PF|Y
C1552908|T129|42|HL7V3.0|Hep B, adolescent/high risk infant||S|PF|Y
C1552908|T121|42|HL7V3.0|Hep B, adolescent/high risk infant||S|PF|Y
C1552909|T129|43|CVX|Hep B, adult||S|PF|N
C1552909|T121|43|CVX|Hep B, adult||S|PF|N
C1552909|T129|43|CVX|hepatitis B vaccine, adult dosage||P|PF|Y
C1552909|T121|43|CVX|hepatitis B vaccine, adult dosage||P|PF|Y
C1552909|T129|43|HL7V3.0|Hep B, adult||S|PF|Y
C1552909|T121|43|HL7V3.0|Hep B, adult||S|PF|Y
C1720918|T129|121|CVX|zoster||S|PF|Y
C1720918|T121|121|CVX|zoster||S|PF|Y
C1720918|T129|121|CVX|zoster vaccine, live||S|VO|Y
C1720918|T121|121|CVX|zoster vaccine, live||S|VO|Y
C1720918|T129|302157|MEDCIN|live herpes zoster vaccine||S|PF|Y
C1720918|T121|302157|MEDCIN|live herpes zoster vaccine||S|PF|Y
C1720918|T129|302157|MEDCIN|live herpes zoster vaccine (medication)||S|PF|Y
C1720918|T121|302157|MEDCIN|live herpes zoster vaccine (medication)||S|PF|Y
C1720918|T129|302157|MEDCIN|zoster vaccine, live||S|VO|N
C1720918|T121|302157|MEDCIN|zoster vaccine, live||S|VO|N
C1720918|T129|21429|MMSL|zoster vaccine live||S|PF|N
C1720918|T121|21429|MMSL|zoster vaccine live||S|PF|N
C1720918|T129|d05813|MMSL|zoster vaccine live||S|PF|Y
C1720918|T121|d05813|MMSL|zoster vaccine live||S|PF|Y
C1720918|T129|D053061|MSH|Herpes Zoster Vaccine||P|PF|N
C1720918|T121|D053061|MSH|Herpes Zoster Vaccine||P|PF|N
C1720918|T129|D053061|MSH|Shingles Vaccine||S|PF|Y
C1720918|T121|D053061|MSH|Shingles Vaccine||S|PF|Y
C1720918|T129|D053061|MSH|Vaccine, Herpes Zoster||P|VW|Y
C1720918|T121|D053061|MSH|Vaccine, Herpes Zoster||P|VW|Y
C1720918|T129|D053061|MSH|Vaccine, Shingles||S|VW|Y
C1720918|T121|D053061|MSH|Vaccine, Shingles||S|VW|Y
C1720918|T129|D053061|MSH|Vaccine, Zoster||S|VW|Y
C1720918|T121|D053061|MSH|Vaccine, Zoster||S|VW|Y
C1720918|T129|D053061|MSH|Zoster Vaccine||S|PF|Y
C1720918|T121|D053061|MSH|Zoster Vaccine||S|PF|Y
C1720918|T129|NOCODE|MTH|Herpes Zoster Vaccine||P|PF|Y
C1720918|T121|NOCODE|MTH|Herpes Zoster Vaccine||P|PF|Y
C1720918|T129|N0000175337|NDFRT|Herpes Zoster Vaccine||P|PF|N
C1720918|T121|N0000175337|NDFRT|Herpes Zoster Vaccine||P|PF|N
C1720918|T129|N0000175337|NDFRT|Herpes Zoster Vaccine [Chemical/Ingredient]||S|PF|Y
C1720918|T121|N0000175337|NDFRT|Herpes Zoster Vaccine [Chemical/Ingredient]||S|PF|Y
C1720918|T129|N0000175337|NDFRT|Shingles Vaccine||S|PF|N
C1720918|T121|N0000175337|NDFRT|Shingles Vaccine||S|PF|N
C1720918|T129|N0000175337|NDFRT|Zoster Vaccine||S|PF|N
C1720918|T121|N0000175337|NDFRT|Zoster Vaccine||S|PF|N
C1720918|T129|N0000176171|NDFRT|ZOSTER VACCINE||S|VC|N
C1720918|T121|N0000176171|NDFRT|ZOSTER VACCINE||S|VC|N
C1720918|T129|4025495|VANDF|ZOSTER VACCINE||S|VC|Y
C1720918|T121|4025495|VANDF|ZOSTER VACCINE||S|VC|Y
C2047258|T129|62|CVX|HPV, quadrivalent||S|PF|Y
C2047258|T121|62|CVX|HPV, quadrivalent||S|PF|Y
C2047258|T129|62|CVX|human papilloma virus vaccine, quadrivalent||P|PF|Y
C2047258|T121|62|CVX|human papilloma virus vaccine, quadrivalent||P|PF|Y
C2047258|T129|302156|MEDCIN|human papilloma virus vaccine, quadrivalent||P|PF|N
C2047258|T121|302156|MEDCIN|human papilloma virus vaccine, quadrivalent||P|PF|N
C2047258|T129|302156|MEDCIN|human papilloma virus vaccine, quadrivalent (medication)||S|PF|Y
C2047258|T121|302156|MEDCIN|human papilloma virus vaccine, quadrivalent (medication)||S|PF|Y
C2094631|T129|50|CVX|DTaP-Haemophilus influenzae type b conjugate vaccine||P|PF|Y
C2094631|T121|50|CVX|DTaP-Haemophilus influenzae type b conjugate vaccine||P|PF|Y
C2094631|T129|50|CVX|DTaP-Hib||S|PF|N
C2094631|T121|50|CVX|DTaP-Hib||S|PF|N
C2094631|T129|50|HL7V2.5|DTaP-Hib||S|PF|Y
C2094631|T121|50|HL7V2.5|DTaP-Hib||S|PF|Y
C2094631|T129|50|HL7V3.0|DTaPHib||S|PF|Y
C2094631|T121|50|HL7V3.0|DTaPHib||S|PF|Y
C2094631|T129|76711|MEDCIN|diphtheria, tetanus, and acellular pertussis (DTaP) vaccine + active Haemophilus influenzae type B (HIB) vaccine||S|PF|Y
C2094631|T121|76711|MEDCIN|diphtheria, tetanus, and acellular pertussis (DTaP) vaccine + active Haemophilus influenzae type B (HIB) vaccine||S|PF|Y
C2094631|T129|76711|MEDCIN|diphtheria, tetanus, and acellular pertussis (DTaP) vaccine + active Haemophilus influenzae type B (HIB) vaccine (medication)||S|PF|Y
C2094631|T121|76711|MEDCIN|diphtheria, tetanus, and acellular pertussis (DTaP) vaccine + active Haemophilus influenzae type B (HIB) vaccine (medication)||S|PF|Y
C2148557|T129|58|CVX|Hep C||S|PF|N
C2148557|T121|58|CVX|Hep C||S|PF|N
C2148557|T129|58|CVX|hepatitis C vaccine||P|PF|N
C2148557|T121|58|CVX|hepatitis C vaccine||P|PF|N
C2148557|T129|58|HL7V2.5|Hep C||S|PF|N
C2148557|T121|58|HL7V2.5|Hep C||S|PF|N
C2148557|T129|58|HL7V3.0|Hep C||S|PF|Y
C2148557|T121|58|HL7V3.0|Hep C||S|PF|Y
C2148557|T129|133272|MEDCIN|hepatitis C vaccine||P|PF|Y
C2148557|T121|133272|MEDCIN|hepatitis C vaccine||P|PF|Y
C2148557|T129|133272|MEDCIN|hepatitis C vaccine (medication)||S|PF|Y
C2148557|T121|133272|MEDCIN|hepatitis C vaccine (medication)||S|PF|Y
C2342811|T200|119|CVX|rotavirus, live, monovalent vaccine||P|VW|Y
C2342811|T200|119|CVX|rotavirus, monovalent||S|PF|Y
C2342811|T200|21736|MMSL|rotavirus vaccine, live, monovalent||P|PF|Y
C2367757|T129|118|CVX|HPV, bivalent||S|PF|Y
C2367757|T121|118|CVX|HPV, bivalent||S|PF|Y
C2367757|T129|118|CVX|human papilloma virus vaccine, bivalent||P|PF|Y
C2367757|T121|118|CVX|human papilloma virus vaccine, bivalent||P|PF|Y
C2367757|T129|304017|MEDCIN|bivalent HPV vaccine||S|PF|Y
C2367757|T121|304017|MEDCIN|bivalent HPV vaccine||S|PF|Y
C2367757|T129|304017|MEDCIN|bivalent human papilloma virus vaccine||P|VW|Y
C2367757|T121|304017|MEDCIN|bivalent human papilloma virus vaccine||P|VW|Y
C2367757|T129|304017|MEDCIN|bivalent human papilloma virus vaccine (medication)||S|PF|Y
C2367757|T121|304017|MEDCIN|bivalent human papilloma virus vaccine (medication)||S|PF|Y
C2367757|T129|304017|MEDCIN|human papilloma virus vaccine, bivalent||P|PF|N
C2367757|T121|304017|MEDCIN|human papilloma virus vaccine, bivalent||P|PF|N
C2716396|T129|120|CVX|diphtheria, tetanus toxoids and acellular pertussis vaccine, Haemophilus influenzae type b conjugate, and poliovirus vaccine, inactivated (DTaP-Hib-IPV)||S|PF|Y
C2716396|T121|120|CVX|diphtheria, tetanus toxoids and acellular pertussis vaccine, Haemophilus influenzae type b conjugate, and poliovirus vaccine, inactivated (DTaP-Hib-IPV)||S|PF|Y
C2716396|T129|120|CVX|DTaP-Hib-IPV||S|VW|Y
C2716396|T121|120|CVX|DTaP-Hib-IPV||S|VW|Y
C2716396|T129|C541234|MSH|diphtheria-tetanus-five component acellular pertussis-inactivated poliomyelitis -Haemophilus influenzae type b conjugate vaccine||P|PF|Y
C2716396|T121|C541234|MSH|diphtheria-tetanus-five component acellular pertussis-inactivated poliomyelitis -Haemophilus influenzae type b conjugate vaccine||P|PF|Y
C2716396|T129|C541234|MSH|DTaP-IPV-Hib conjugate vaccine||S|PF|Y
C2716396|T121|C541234|MSH|DTaP-IPV-Hib conjugate vaccine||S|PF|Y
C2716396|T129|C122399|NCI|Diphtheria-Tetanus-Acellular Pertussis-Inactivated Poliomyelitis-Haemophilus influenzae Type B Vaccine||S|PF|Y
C2716396|T121|C122399|NCI|Diphtheria-Tetanus-Acellular Pertussis-Inactivated Poliomyelitis-Haemophilus influenzae Type B Vaccine||S|PF|Y
C2716396|T129|C122399|NCI|DTaP-IPV-Hib||S|PF|Y
C2716396|T121|C122399|NCI|DTaP-IPV-Hib||S|PF|Y
C2716396|T129|C122399|NCI|DTaP(5)-IPV-Hib||S|PF|Y
C2716396|T121|C122399|NCI|DTaP(5)-IPV-Hib||S|PF|Y
C2716397|T129|146|CVX|Diphtheria and Tetanus Toxoids and Acellular Pertussis Adsorbed, Inactivated Poliovirus, Haemophilus b Conjugate (Meningococcal Protein Conjugate), and Hepatitis B (Recombinant) Vaccine.||S|PF|Y
C2716397|T121|146|CVX|Diphtheria and Tetanus Toxoids and Acellular Pertussis Adsorbed, Inactivated Poliovirus, Haemophilus b Conjugate (Meningococcal Protein Conjugate), and Hepatitis B (Recombinant) Vaccine.||S|PF|Y
C2716397|T129|146|CVX|DTaP,IPV,Hib,HepB||S|VC|Y
C2716397|T121|146|CVX|DTaP,IPV,Hib,HepB||S|VC|Y
C2716397|T129|306116|MEDCIN|dtap-ipv-hib-hepb||S|PF|Y
C2716397|T121|306116|MEDCIN|dtap-ipv-hib-hepb||S|PF|Y
C2716397|T129|306116|MEDCIN|dtap-ipv-hib-hepb (medication)||S|PF|Y
C2716397|T121|306116|MEDCIN|dtap-ipv-hib-hepb (medication)||S|PF|Y
C2716397|T129|C541235|MSH|diphtheria-tetanus-acellular pertussis-inactivated poliovirus-Haemophilus influenzae b conjugate-hepatitis B vaccine||P|PF|Y
C2716397|T121|C541235|MSH|diphtheria-tetanus-acellular pertussis-inactivated poliovirus-Haemophilus influenzae b conjugate-hepatitis B vaccine||P|PF|Y
C2716397|T129|C541235|MSH|DTaP-IPV-Hib-HBV conjugate vaccine||S|PF|Y
C2716397|T121|C541235|MSH|DTaP-IPV-Hib-HBV conjugate vaccine||S|PF|Y
C2716397|T129|C541235|MSH|DTaP-IPV-Hib-HBV vaccine||S|PF|Y
C2716397|T121|C541235|MSH|DTaP-IPV-Hib-HBV vaccine||S|PF|Y
C2719522|T129|90680|CPT|Live rotavirus vaccine, pentavalent||P|VCW|Y
C2719522|T121|90680|CPT|Live rotavirus vaccine, pentavalent||P|VCW|Y
C2719522|T129|116|CVX|rotavirus, live, pentavalent vaccine||P|VW|Y
C2719522|T121|116|CVX|rotavirus, live, pentavalent vaccine||P|VW|Y
C2719522|T129|116|CVX|rotavirus, pentavalent||S|PF|Y
C2719522|T121|116|CVX|rotavirus, pentavalent||S|PF|Y
C2719522|T129|26561|MMSL|rotavirus vaccine, live, pentavalent||P|PF|Y
C2719522|T121|26561|MMSL|rotavirus vaccine, live, pentavalent||P|PF|Y
C3152625|T129|90670|CPT|Pneumococcal conjugate vaccine, 13 valent||P|VW|Y
C3152625|T121|90670|CPT|Pneumococcal conjugate vaccine, 13 valent||P|VW|Y
C3152625|T129|133|CVX|Pneumococcal conjugate PCV 13||S|PF|Y
C3152625|T121|133|CVX|Pneumococcal conjugate PCV 13||S|PF|Y
C3152625|T129|133|CVX|pneumococcal conjugate vaccine, 13 valent||P|VCW|Y
C3152625|T121|133|CVX|pneumococcal conjugate vaccine, 13 valent||P|VCW|Y
C3152625|T129|d07586|MMSL|pneumococcal 13-valent conjugate vaccine||P|VC|Y
C3152625|T121|d07586|MMSL|pneumococcal 13-valent conjugate vaccine||P|VC|Y
C3152625|T129|C568598|MSH|PCV13 vaccine||S|PF|Y
C3152625|T121|C568598|MSH|PCV13 vaccine||S|PF|Y
C3152625|T129|C97121|NCI|PCV 13||S|PF|N
C3152625|T121|C97121|NCI|PCV 13||S|PF|N
C3152625|T129|C97121|NCI|PCV13 Vaccine||S|VC|Y
C3152625|T121|C97121|NCI|PCV13 Vaccine||S|VC|Y
C3152625|T129|C97121|NCI|Pneumococcal 13-valent Conjugate Vaccine||P|VC|Y
C3152625|T121|C97121|NCI|Pneumococcal 13-valent Conjugate Vaccine||P|VC|Y
C3152625|T129|C97121|NCI_NICHD|PCV 13||S|PF|Y
C3152625|T121|C97121|NCI_NICHD|PCV 13||S|PF|Y
C3152625|T129|C97121|NCI_NICHD|Pneumococcal 13-valent Conjugate Vaccine||P|VC|N
C3152625|T121|C97121|NCI_NICHD|Pneumococcal 13-valent Conjugate Vaccine||P|VC|N
C3152625|T129|N0000183831|NDFRT|PNEUMOCOCCAL 13-VALENT CONJUGATE VACCINE||P|VC|N
C3152625|T121|N0000183831|NDFRT|PNEUMOCOCCAL 13-VALENT CONJUGATE VACCINE||P|VC|N
C3152625|T129|N0000183831|NDFRT|PNEUMOCOCCAL 13-VALENT CONJUGATE VACCINE [VA Product]||S|PF|Y
C3152625|T121|N0000183831|NDFRT|PNEUMOCOCCAL 13-VALENT CONJUGATE VACCINE [VA Product]||S|PF|Y
C3152625|T129|448964007|SNOMEDCT_US|Pneumococcal 13-valent conjugate vaccine||P|PF|Y
C3152625|T121|448964007|SNOMEDCT_US|Pneumococcal 13-valent conjugate vaccine||P|PF|Y
C3152625|T129|448964007|SNOMEDCT_US|Pneumococcal 13-valent conjugate vaccine (product)||S|PF|Y
C3152625|T121|448964007|SNOMEDCT_US|Pneumococcal 13-valent conjugate vaccine (product)||S|PF|Y
C3152625|T129|4031027|VANDF|PNEUMOCOCCAL 13-VALENT CONJUGATE VACCINE||P|VC|Y
C3152625|T129|4031027|VANDF|PNEUMOCOCCAL 13-VALENT CONJUGATE VACCINE||P|VC|N
C3152625|T121|4031027|VANDF|PNEUMOCOCCAL 13-VALENT CONJUGATE VACCINE||P|VC|Y
C3152625|T121|4031027|VANDF|PNEUMOCOCCAL 13-VALENT CONJUGATE VACCINE||P|VC|N
C3161510|T129|142|CVX|tetanus toxoid, not adsorbed||P|PF|N
C3161510|T129|142|CVX|tetanus toxoid, not adsorbed||P|PF|Y
C3161510|T121|142|CVX|tetanus toxoid, not adsorbed||P|PF|N
C3161510|T121|142|CVX|tetanus toxoid, not adsorbed||P|PF|Y
C3161510|T129|307941|MEDCIN|tetanus toxoid, not adsorbed||P|PF|N
C3161510|T121|307941|MEDCIN|tetanus toxoid, not adsorbed||P|PF|N
C3161510|T129|307941|MEDCIN|tetanus toxoid, not adsorbed (medication)||S|PF|Y
C3161510|T121|307941|MEDCIN|tetanus toxoid, not adsorbed (medication)||S|PF|Y
C3272840|T129|32|CVX|meningococcal MPSV4||S|PF|Y
C3272840|T121|32|CVX|meningococcal MPSV4||S|PF|Y
C3272840|T129|32|CVX|meningococcal polysaccharide vaccine (MPSV4)||P|PF|N
C3272840|T121|32|CVX|meningococcal polysaccharide vaccine (MPSV4)||P|PF|N
C3272840|T129|32|HL7V2.5|meningococcal||S|PF|N
C3272840|T121|32|HL7V2.5|meningococcal||S|PF|N
C3272840|T129|32|HL7V3.0|meningococcal||S|PF|Y
C3272840|T121|32|HL7V3.0|meningococcal||S|PF|Y
C3272840|T129|NOCODE|MTH|meningococcal polysaccharide vaccine (MPSV4)||P|PF|Y
C3272840|T121|NOCODE|MTH|meningococcal polysaccharide vaccine (MPSV4)||P|PF|Y
C3272840|T129|C96519|NCI|Meningococcal Polysaccharide Vaccine MPS-4||S|PF|Y
C3272840|T121|C96519|NCI|Meningococcal Polysaccharide Vaccine MPS-4||S|PF|Y
C3272840|T129|C96519|NCI|Meningococcal Polysaccharide Vaccine MPSV4||P|VC|Y
C3272840|T121|C96519|NCI|Meningococcal Polysaccharide Vaccine MPSV4||P|VC|Y
C3272840|T129|C96519|NCI|Meningococcal Polysaccharide Vaccine, Groups A, C, Y and W-135 Combination||S|PF|Y
C3272840|T121|C96519|NCI|Meningococcal Polysaccharide Vaccine, Groups A, C, Y and W-135 Combination||S|PF|Y
C3272840|T129|C96519|NCI_NICHD|Meningococcal Polysaccharide Vaccine MPSV-4||S|PF|Y
C3272840|T121|C96519|NCI_NICHD|Meningococcal Polysaccharide Vaccine MPSV-4||S|PF|Y
C3272840|T129|C96519|NCI_NICHD|Meningococcal Polysaccharide Vaccine MPSV4||P|VC|N
C3272840|T121|C96519|NCI_NICHD|Meningococcal Polysaccharide Vaccine MPSV4||P|VC|N
C3273244|T129|90691|CPT|Typhoid vaccine, Vi capsular polysaccharide||P|VCW|Y
C3273244|T121|90691|CPT|Typhoid vaccine, Vi capsular polysaccharide||P|VCW|Y
C3273244|T129|101|CVX|typhoid Vi capsular polysaccharide vaccine||P|VCW|Y
C3273244|T121|101|CVX|typhoid Vi capsular polysaccharide vaccine||P|VCW|Y
C3273244|T129|101|CVX|typhoid, ViCPs||S|PF|N
C3273244|T121|101|CVX|typhoid, ViCPs||S|PF|N
C3273244|T129|101|HL7V2.5|typhoid, ViCPs||S|PF|N
C3273244|T121|101|HL7V2.5|typhoid, ViCPs||S|PF|N
C3273244|T129|101|HL7V3.0|typhoid, ViCPs||S|PF|Y
C3273244|T121|101|HL7V3.0|typhoid, ViCPs||S|PF|Y
C3273244|T129|NOCODE|MTH|Vi Capsular Polysaccharide Typhoid Vaccine||P|PF|Y
C3273244|T121|NOCODE|MTH|Vi Capsular Polysaccharide Typhoid Vaccine||P|PF|Y
C3273244|T129|C97127|NCI|Vi Capsular Polysaccharide Typhoid Vaccine||P|PF|N
C3273244|T121|C97127|NCI|Vi Capsular Polysaccharide Typhoid Vaccine||P|PF|N
C3273244|T129|C97127|NCI_NICHD|Vi||S|PF|Y
C3273244|T121|C97127|NCI_NICHD|Vi||S|PF|Y
C3273244|T129|C97127|NCI_NICHD|Vi Capsular Polysaccharide Typhoid Vaccine||P|PF|N
C3273244|T121|C97127|NCI_NICHD|Vi Capsular Polysaccharide Typhoid Vaccine||P|PF|N
C3273244|T129|C97127|NCI_NICHD|ViCPS||S|PF|Y
C3273244|T121|C97127|NCI_NICHD|ViCPS||S|PF|Y
C3494357|T129|143|CVX|Adenovirus types 4 and 7||S|PF|Y
C3494357|T121|143|CVX|Adenovirus types 4 and 7||S|PF|Y
C3494357|T129|143|CVX|Adenovirus, type 4 and type 7, live, oral||S|PF|Y
C3494357|T121|143|CVX|Adenovirus, type 4 and type 7, live, oral||S|PF|Y
C3494357|T129|D062705|MSH|Adenovirus Type 4 and Type 7 Vaccine, Live, Oral||P|PF|Y
C3494357|T121|D062705|MSH|Adenovirus Type 4 and Type 7 Vaccine, Live, Oral||P|PF|Y
C3494357|T129|D062705|MSH|Adenovirus Type 4 and Type 7 Vaccines, Live, Oral||P|VO|Y
C3494357|T121|D062705|MSH|Adenovirus Type 4 and Type 7 Vaccines, Live, Oral||P|VO|Y
C3511581|T121|149|CVX|influenza, live, intranasal, quadrivalent||P|PF|N
C3511581|T121|149|CVX|influenza, live, intranasal, quadrivalent||P|PF|Y
C3511581|T129|149|CVX|influenza, live, intranasal, quadrivalent||P|PF|N
C3511581|T129|149|CVX|influenza, live, intranasal, quadrivalent||P|PF|Y
C3511581|T121|309648|MEDCIN|influenza virus vaccine live intranasal quadrivalent||S|PF|Y
C3511581|T129|309648|MEDCIN|influenza virus vaccine live intranasal quadrivalent||S|PF|Y
C3511581|T121|309648|MEDCIN|influenza virus vaccine live intranasal quadrivalent (medication)||S|PF|Y
C3511581|T129|309648|MEDCIN|influenza virus vaccine live intranasal quadrivalent (medication)||S|PF|Y
C3526526|T129|90632|CPT|Hepatitis A vaccine, adult dosage||P|PF|Y
C3526526|T121|90632|CPT|Hepatitis A vaccine, adult dosage||P|PF|Y
C3526526|T129|52|CVX|Hep A, adult||S|PF|N
C3526526|T121|52|CVX|Hep A, adult||S|PF|N
C3526526|T129|52|CVX|hepatitis A vaccine, adult dosage||P|VC|Y
C3526526|T121|52|CVX|hepatitis A vaccine, adult dosage||P|VC|Y
C3526526|T129|52|HL7V2.5|Hep A, adult||S|PF|N
C3526526|T121|52|HL7V2.5|Hep A, adult||S|PF|N
C3526526|T129|52|HL7V3.0|Hep A, adult||S|PF|Y
C3526526|T121|52|HL7V3.0|Hep A, adult||S|PF|Y
C3526551|T121|90696|CPT|Diphtheria, tetanus toxoids, acellular pertussis vaccine and poliovirus vaccine, inactivated||P|PF|Y
C3526551|T129|90696|CPT|Diphtheria, tetanus toxoids, acellular pertussis vaccine and poliovirus vaccine, inactivated||P|PF|Y
C3526551|T121|130|CVX|Diphtheria, tetanus toxoids and acellular pertussis vaccine, and poliovirus vaccine, inactivated||P|VO|Y
C3526551|T129|130|CVX|Diphtheria, tetanus toxoids and acellular pertussis vaccine, and poliovirus vaccine, inactivated||P|VO|Y
C3526551|T121|130|CVX|DTaP-IPV||S|PF|N
C3526551|T129|130|CVX|DTaP-IPV||S|PF|N
C3526551|T121|303949|MEDCIN|DTaP-IPV||S|PF|Y
C3526551|T129|303949|MEDCIN|DTaP-IPV||S|PF|Y
C3526551|T121|303949|MEDCIN|DTaP-IPV (medication)||S|PF|Y
C3526551|T129|303949|MEDCIN|DTaP-IPV (medication)||S|PF|Y
C3526553|T129|90700|CPT|Diphtheria, tetanus toxoids, and acellular pertussis vaccine||P|PF|N
C3526553|T121|90700|CPT|Diphtheria, tetanus toxoids, and acellular pertussis vaccine||P|PF|N
C3526553|T129|20|CVX|diphtheria, tetanus toxoids and acellular pertussis vaccine||P|VC|Y
C3526553|T121|20|CVX|diphtheria, tetanus toxoids and acellular pertussis vaccine||P|VC|Y
C3526553|T129|20|CVX|DTaP||S|PF|Y
C3526553|T121|20|CVX|DTaP||S|PF|Y
C3526553|T129|NOCODE|MTH|Diphtheria, tetanus toxoids, and acellular pertussis vaccine||P|PF|Y
C3526553|T121|NOCODE|MTH|Diphtheria, tetanus toxoids, and acellular pertussis vaccine||P|PF|Y
C3536784|T129|29|CVX|CMVIG||S|PF|N
C3536784|T121|29|CVX|CMVIG||S|PF|N
C3536784|T129|29|CVX|cytomegalovirus immune globulin, intravenous||P|PF|N
C3536784|T121|29|CVX|cytomegalovirus immune globulin, intravenous||P|PF|N
C3536784|T129|29|HL7V2.5|CMVIG||S|PF|N
C3536784|T121|29|HL7V2.5|CMVIG||S|PF|N
C3536784|T129|29|HL7V3.0|CMVIG||S|PF|Y
C3536784|T121|29|HL7V3.0|CMVIG||S|PF|Y
C3536784|T129|NOCODE|MTH|cytomegalovirus immune globulin, intravenous||P|PF|Y
C3536784|T121|NOCODE|MTH|cytomegalovirus immune globulin, intravenous||P|PF|Y
C3536964|T129|74|CVX|rotavirus, live, tetravalent vaccine||P|PF|N
C3536964|T121|74|CVX|rotavirus, live, tetravalent vaccine||P|PF|N
C3536964|T129|74|CVX|rotavirus, tetravalent||S|PF|Y
C3536964|T121|74|CVX|rotavirus, tetravalent||S|PF|Y
C3536964|T129|74|HL7V2.5|rotavirus||S|PF|N
C3536964|T121|74|HL7V2.5|rotavirus||S|PF|N
C3536964|T129|74|HL7V3.0|rotavirus||S|PF|Y
C3536964|T121|74|HL7V3.0|rotavirus||S|PF|Y
C3536964|T129|NOCODE|MTH|rotavirus, live, tetravalent vaccine||P|PF|Y
C3536964|T121|NOCODE|MTH|rotavirus, live, tetravalent vaccine||P|PF|Y
C3536988|T129|39|CVX|Japanese encephalitis SC||S|PF|Y
C3536988|T121|39|CVX|Japanese encephalitis SC||S|PF|Y
C3536988|T129|39|CVX|Japanese Encephalitis Vaccine SC||P|PF|Y
C3536988|T121|39|CVX|Japanese Encephalitis Vaccine SC||P|PF|Y
C3536988|T129|44436|MEDCIN|inactivated Japanese encephalitis vaccine for subcutaneous use||S|PF|Y
C3536988|T121|44436|MEDCIN|inactivated Japanese encephalitis vaccine for subcutaneous use||S|PF|Y
C3536988|T129|44436|MEDCIN|inactivated Japanese encephalitis vaccine for subcutaneous use (medication)||S|PF|Y
C3536988|T121|44436|MEDCIN|inactivated Japanese encephalitis vaccine for subcutaneous use (medication)||S|PF|Y
C3536988|T129|44436|MEDCIN|vaccines viral Japanese encephalitis||S|PF|Y
C3536988|T121|44436|MEDCIN|vaccines viral Japanese encephalitis||S|PF|Y
C3539056|T129|138|CVX|Td (adult)||S|PF|Y
C3539056|T121|138|CVX|Td (adult)||S|PF|Y
C3539056|T129|138|CVX|tetanus and diphtheria toxoids, not adsorbed, for adult use||P|PF|N
C3539056|T121|138|CVX|tetanus and diphtheria toxoids, not adsorbed, for adult use||P|PF|N
C3539056|T129|NOCODE|MTH|tetanus and diphtheria toxoids, not adsorbed, for adult use||P|PF|Y
C3539056|T121|NOCODE|MTH|tetanus and diphtheria toxoids, not adsorbed, for adult use||P|PF|Y
C3541433|T121|999|CVX|unknown||S|PF|Y
C3541433|T129|999|CVX|unknown||S|PF|Y
C3541433|T121|999|CVX|unknown vaccine or immune globulin||P|PF|N
C3541433|T129|999|CVX|unknown vaccine or immune globulin||P|PF|N
C3541433|T121|NOCODE|MTH|unknown vaccine or immune globulin||P|PF|Y
C3541433|T129|NOCODE|MTH|unknown vaccine or immune globulin||P|PF|Y
C3644154|T129|107|CVX|diphtheria, tetanus toxoids and acellular pertussis vaccine, unspecified formulation||P|PF|Y
C3644154|T121|107|CVX|diphtheria, tetanus toxoids and acellular pertussis vaccine, unspecified formulation||P|PF|Y
C3644154|T129|107|CVX|DTaP, unspecified formulation||S|PF|Y
C3644154|T121|107|CVX|DTaP, unspecified formulation||S|PF|Y
C3644155|T121|110|CVX|DTaP-Hep B-IPV||S|PF|Y
C3644155|T129|110|CVX|DTaP-Hep B-IPV||S|PF|Y
C3644155|T121|110|CVX|DTaP-hepatitis B and poliovirus vaccine||P|PF|Y
C3644155|T129|110|CVX|DTaP-hepatitis B and poliovirus vaccine||P|PF|Y
C3644157|T121|85|CVX|Hep A, unspecified formulation||S|PF|Y
C3644157|T129|85|CVX|Hep A, unspecified formulation||S|PF|Y
C3644157|T121|85|CVX|hepatitis A vaccine, unspecified formulation||P|PF|Y
C3644157|T129|85|CVX|hepatitis A vaccine, unspecified formulation||P|PF|Y
C3644158|T121|45|CVX|Hep B, unspecified formulation||S|PF|Y
C3644158|T129|45|CVX|Hep B, unspecified formulation||S|PF|Y
C3644158|T121|45|CVX|hepatitis B vaccine, unspecified formulation||P|PF|Y
C3644158|T129|45|CVX|hepatitis B vaccine, unspecified formulation||P|PF|Y
C3644159|T121|17|CVX|Haemophilus influenzae type b vaccine, conjugate unspecified formulation||P|PF|Y
C3644159|T129|17|CVX|Haemophilus influenzae type b vaccine, conjugate unspecified formulation||P|PF|Y
C3644159|T121|17|CVX|Hib, unspecified formulation||S|PF|Y
C3644159|T129|17|CVX|Hib, unspecified formulation||S|PF|Y
C3644160|T121|14|CVX|IG, unspecified formulation||S|PF|Y
C3644160|T129|14|CVX|IG, unspecified formulation||S|PF|Y
C3644160|T121|14|CVX|immune globulin, unspecified formulation||P|PF|Y
C3644160|T129|14|CVX|immune globulin, unspecified formulation||P|PF|Y
C3644161|T121|111|CVX|influenza virus vaccine, live, attenuated, for intranasal use||P|PF|Y
C3644161|T129|111|CVX|influenza virus vaccine, live, attenuated, for intranasal use||P|PF|Y
C3644161|T121|111|CVX|influenza, live, intranasal||S|PF|Y
C3644161|T129|111|CVX|influenza, live, intranasal||S|PF|Y
C3644162|T129|88|CVX|influenza virus vaccine, unspecified formulation||P|PF|Y
C3644162|T121|88|CVX|influenza virus vaccine, unspecified formulation||P|PF|Y
C3644162|T129|88|CVX|influenza, unspecified formulation||S|PF|Y
C3644162|T121|88|CVX|influenza, unspecified formulation||S|PF|Y
C3644163|T121|123|CVX|influenza virus vaccine, H5N1, A/Vietnam/1203/2004 (national stockpile)||P|PF|Y
C3644163|T129|123|CVX|influenza virus vaccine, H5N1, A/Vietnam/1203/2004 (national stockpile)||P|PF|Y
C3644163|T121|123|CVX|influenza, H5N1-1203||S|PF|Y
C3644163|T129|123|CVX|influenza, H5N1-1203||S|PF|Y
C3644164|T121|89|CVX|polio, unspecified formulation||S|PF|Y
C3644164|T129|89|CVX|polio, unspecified formulation||S|PF|Y
C3644164|T121|89|CVX|poliovirus vaccine, unspecified formulation||P|PF|Y
C3644164|T129|89|CVX|poliovirus vaccine, unspecified formulation||P|PF|Y
C3644165|T129|114|CVX|meningococcal MCV4P||S|PF|Y
C3644165|T121|114|CVX|meningococcal MCV4P||S|PF|Y
C3644165|T129|114|CVX|meningococcal polysaccharide (groups A, C, Y and W-135) diphtheria toxoid conjugate vaccine (MCV4P)||P|PF|Y
C3644165|T121|114|CVX|meningococcal polysaccharide (groups A, C, Y and W-135) diphtheria toxoid conjugate vaccine (MCV4P)||P|PF|Y
C3644167|T121|109|CVX|pneumococcal vaccine, unspecified formulation||P|PF|Y
C3644167|T129|109|CVX|pneumococcal vaccine, unspecified formulation||P|PF|Y
C3644167|T121|109|CVX|pneumococcal, unspecified formulation||S|PF|Y
C3644167|T129|109|CVX|pneumococcal, unspecified formulation||S|PF|Y
C3644168|T129|90|CVX|rabies vaccine, unspecified formulation||P|PF|Y
C3644168|T121|90|CVX|rabies vaccine, unspecified formulation||P|PF|Y
C3644168|T129|90|CVX|rabies, unspecified formulation||S|PF|Y
C3644168|T121|90|CVX|rabies, unspecified formulation||S|PF|Y
C3644169|T129|122|CVX|rotavirus vaccine, unspecified formulation||P|PF|Y
C3644169|T121|122|CVX|rotavirus vaccine, unspecified formulation||P|PF|Y
C3644169|T129|122|CVX|rotavirus, unspecified formulation||S|PF|Y
C3644169|T121|122|CVX|rotavirus, unspecified formulation||S|PF|Y
C3644170|T129|113|CVX|Td (adult) preservative free||S|PF|Y
C3644170|T121|113|CVX|Td (adult) preservative free||S|PF|Y
C3644170|T129|113|CVX|tetanus and diphtheria toxoids, adsorbed, preservative free, for adult use||P|PF|Y
C3644170|T121|113|CVX|tetanus and diphtheria toxoids, adsorbed, preservative free, for adult use||P|PF|Y
C3644171|T121|115|CVX|Tdap||S|PF|Y
C3644171|T129|115|CVX|Tdap||S|PF|Y
C3644171|T121|115|CVX|tetanus toxoid, reduced diphtheria toxoid, and acellular pertussis vaccine, adsorbed||P|PF|Y
C3644171|T129|115|CVX|tetanus toxoid, reduced diphtheria toxoid, and acellular pertussis vaccine, adsorbed||P|PF|Y
C3644172|T121|112|CVX|tetanus toxoid, unspecified formulation||P|PF|N
C3644172|T121|112|CVX|tetanus toxoid, unspecified formulation||P|PF|Y
C3644172|T129|112|CVX|tetanus toxoid, unspecified formulation||P|PF|N
C3644172|T129|112|CVX|tetanus toxoid, unspecified formulation||P|PF|Y
C3644173|T130|98|CVX|TST, unspecified formulation||S|PF|Y
C3644173|T129|98|CVX|TST, unspecified formulation||S|PF|Y
C3644173|T130|98|CVX|tuberculin skin test; unspecified formulation||P|PF|Y
C3644173|T129|98|CVX|tuberculin skin test; unspecified formulation||P|PF|Y
C3644174|T129|91|CVX|typhoid vaccine, unspecified formulation||P|PF|Y
C3644174|T121|91|CVX|typhoid vaccine, unspecified formulation||P|PF|Y
C3644174|T129|91|CVX|typhoid, unspecified formulation||S|PF|Y
C3644174|T121|91|CVX|typhoid, unspecified formulation||S|PF|Y
C3644175|T129|92|CVX|VEE, unspecified formulation||S|PF|Y
C3644175|T121|92|CVX|VEE, unspecified formulation||S|PF|Y
C3644175|T129|92|CVX|Venezuelan equine encephalitis vaccine, unspecified formulation||P|PF|Y
C3644175|T121|92|CVX|Venezuelan equine encephalitis vaccine, unspecified formulation||P|PF|Y
C3644176|T129|117|CVX|varicella zoster immune globulin (Investigational New Drug)||P|PF|Y
C3644176|T121|117|CVX|varicella zoster immune globulin (Investigational New Drug)||P|PF|Y
C3644176|T129|117|CVX|VZIG (IND)||S|PF|Y
C3644176|T121|117|CVX|VZIG (IND)||S|PF|Y
C3644177|T129|134|CVX|Japanese Encephalitis IM||S|PF|Y
C3644177|T121|134|CVX|Japanese Encephalitis IM||S|PF|Y
C3644177|T129|134|CVX|Japanese Encephalitis vaccine for intramuscular administration||P|PF|Y
C3644177|T121|134|CVX|Japanese Encephalitis vaccine for intramuscular administration||P|PF|Y
C3644178|T129|137|CVX|HPV, unspecified formulation||P|PF|Y
C3644178|T129|137|CVX|HPV, unspecified formulation||P|PF|N
C3644178|T121|137|CVX|HPV, unspecified formulation||P|PF|Y
C3644178|T121|137|CVX|HPV, unspecified formulation||P|PF|N
C3644179|T121|136|CVX|Meningococcal MCV4O||S|PF|Y
C3644179|T129|136|CVX|Meningococcal MCV4O||S|PF|Y
C3644179|T121|136|CVX|meningococcal oligosaccharide (groups A, C, Y and W-135) diphtheria toxoid conjugate vaccine (MCV4O)||P|PF|Y
C3644179|T129|136|CVX|meningococcal oligosaccharide (groups A, C, Y and W-135) diphtheria toxoid conjugate vaccine (MCV4O)||P|PF|Y
C3644180|T129|135|CVX|Influenza, high dose seasonal||S|PF|Y
C3644180|T121|135|CVX|Influenza, high dose seasonal||S|PF|Y
C3644180|T129|135|CVX|influenza, high dose seasonal, preservative-free||P|PF|Y
C3644180|T121|135|CVX|influenza, high dose seasonal, preservative-free||P|PF|Y
C3644181|T033|131|CVX|Historical record of a typhus vaccination||P|PF|Y
C3644181|T033|131|CVX|typhus, historical||S|PF|Y
C3644182|T033|132|CVX|DTaP-IPV-HIB-HEP B, historical||S|PF|Y
C3644182|T033|132|CVX|Historical record of vaccine containing * diphtheria, tetanus toxoids and acellular pertussis, * poliovirus, inactivated, * Haemophilus influenzae type b conjugate, * Hepatitis B||P|PF|Y
C3644183|T121|128|CVX|Novel influenza-H1N1-09, all formulations||P|PF|Y
C3644183|T121|128|CVX|Novel Influenza-H1N1-09, all formulations||P|VC|Y
C3644183|T129|128|CVX|Novel influenza-H1N1-09, all formulations||P|PF|Y
C3644183|T129|128|CVX|Novel Influenza-H1N1-09, all formulations||P|VC|Y
C3644184|T121|125|CVX|Novel Influenza-H1N1-09, live virus for nasal administration||P|PF|Y
C3644184|T129|125|CVX|Novel Influenza-H1N1-09, live virus for nasal administration||P|PF|Y
C3644184|T121|125|CVX|Novel Influenza-H1N1-09, nasal||S|PF|Y
C3644184|T129|125|CVX|Novel Influenza-H1N1-09, nasal||S|PF|Y
C3644185|T121|126|CVX|Novel influenza-H1N1-09, preservative-free||S|PF|Y
C3644185|T129|126|CVX|Novel influenza-H1N1-09, preservative-free||S|PF|Y
C3644185|T121|126|CVX|Novel influenza-H1N1-09, preservative-free, injectable||P|PF|Y
C3644185|T129|126|CVX|Novel influenza-H1N1-09, preservative-free, injectable||P|PF|Y
C3644186|T121|127|CVX|Novel influenza-H1N1-09||S|PF|Y
C3644186|T129|127|CVX|Novel influenza-H1N1-09||S|PF|Y
C3644186|T121|127|CVX|Novel influenza-H1N1-09, injectable||P|PF|Y
C3644186|T129|127|CVX|Novel influenza-H1N1-09, injectable||P|PF|Y
C3644187|T129|139|CVX|Td(adult) unspecified formulation||P|PF|Y
C3644187|T129|139|CVX|Td(adult) unspecified formulation||P|PF|N
C3644187|T121|139|CVX|Td(adult) unspecified formulation||P|PF|Y
C3644187|T121|139|CVX|Td(adult) unspecified formulation||P|PF|N
C3644188|T121|140|CVX|Influenza, seasonal, injectable, preservative free||P|PF|Y
C3644188|T121|140|CVX|Influenza, seasonal, injectable, preservative free||P|PF|N
C3644188|T129|140|CVX|Influenza, seasonal, injectable, preservative free||P|PF|Y
C3644188|T129|140|CVX|Influenza, seasonal, injectable, preservative free||P|PF|N
C3644189|T129|129|CVX|Japanese Encephalitis vaccine, unspecified formulation||P|PF|Y
C3644189|T121|129|CVX|Japanese Encephalitis vaccine, unspecified formulation||P|PF|Y
C3644189|T129|129|CVX|Japanese Encephalitis, unspecified formulation||S|PF|Y
C3644189|T121|129|CVX|Japanese Encephalitis, unspecified formulation||S|PF|Y
C3644190|T121|141|CVX|Influenza, seasonal, injectable||P|PF|N
C3644190|T121|141|CVX|Influenza, seasonal, injectable||P|PF|Y
C3644190|T129|141|CVX|Influenza, seasonal, injectable||P|PF|N
C3644190|T129|141|CVX|Influenza, seasonal, injectable||P|PF|Y
C3644191|T121|144|CVX|influenza, seasonal, intradermal, preservative free||P|VW|Y
C3644191|T129|144|CVX|influenza, seasonal, intradermal, preservative free||P|VW|Y
C3644191|T121|144|CVX|seasonal influenza, intradermal, preservative free||P|PF|Y
C3644191|T129|144|CVX|seasonal influenza, intradermal, preservative free||P|PF|Y
C3644192|T121|145|CVX|respiratory syncytial virus monoclonal antibody (motavizumab), intramuscular||P|PF|Y
C3644192|T129|145|CVX|respiratory syncytial virus monoclonal antibody (motavizumab), intramuscular||P|PF|Y
C3644192|T121|145|CVX|RSV-MAb (new)||S|PF|Y
C3644192|T129|145|CVX|RSV-MAb (new)||S|PF|Y
C3644194|T121|147|CVX|meningococcal MCV4, unspecified formulation||S|PF|Y
C3644194|T129|147|CVX|meningococcal MCV4, unspecified formulation||S|PF|Y
C3644194|T121|147|CVX|Meningococcal, MCV4, unspecified conjugate formulation(groups A, C, Y and W-135)||P|PF|Y
C3644194|T129|147|CVX|Meningococcal, MCV4, unspecified conjugate formulation(groups A, C, Y and W-135)||P|PF|Y
C3644195|T121|148|CVX|Meningococcal C/Y-HIB PRP||S|PF|Y
C3644195|T129|148|CVX|Meningococcal C/Y-HIB PRP||S|PF|Y
C3644195|T121|148|CVX|Meningococcal Groups C and Y and Haemophilus b Tetanus Toxoid Conjugate Vaccine||P|PF|Y
C3644195|T129|148|CVX|Meningococcal Groups C and Y and Haemophilus b Tetanus Toxoid Conjugate Vaccine||P|PF|Y
C3644196|T121|150|CVX|Influenza, injectable, quadrivalent, preservative free||P|PF|Y
C3644196|T121|150|CVX|influenza, injectable, quadrivalent, preservative free||P|VC|Y
C3644196|T129|150|CVX|Influenza, injectable, quadrivalent, preservative free||P|PF|Y
C3644196|T129|150|CVX|influenza, injectable, quadrivalent, preservative free||P|VC|Y
C3644197|T121|151|CVX|influenza nasal, unspecified formulation||P|PF|Y
C3644197|T121|151|CVX|influenza nasal, unspecified formulation||P|PF|N
C3644197|T129|151|CVX|influenza nasal, unspecified formulation||P|PF|Y
C3644197|T129|151|CVX|influenza nasal, unspecified formulation||P|PF|N
C3644198|T129|152|CVX|Pneumococcal Conjugate, unspecified formulation||P|PF|Y
C3644198|T129|152|CVX|Pneumococcal Conjugate, unspecified formulation||P|PF|N
C3644198|T121|152|CVX|Pneumococcal Conjugate, unspecified formulation||P|PF|Y
C3644198|T121|152|CVX|Pneumococcal Conjugate, unspecified formulation||P|PF|N
C3644199|T121|153|CVX|Influenza, injectable, Madin Darby Canine Kidney, preservative free||P|PF|Y
C3644199|T129|153|CVX|Influenza, injectable, Madin Darby Canine Kidney, preservative free||P|PF|Y
C3644199|T121|153|CVX|Influenza, injectable, MDCK, preservative free||S|PF|Y
C3644199|T129|153|CVX|Influenza, injectable, MDCK, preservative free||S|PF|Y
C3644200|T121|154|CVX|Hep A, IG||S|PF|Y
C3644200|T129|154|CVX|Hep A, IG||S|PF|Y
C3644200|T121|154|CVX|Hepatitis A immune globulin||P|PF|Y
C3644200|T129|154|CVX|Hepatitis A immune globulin||P|PF|Y
C3644201|T129|155|CVX|influenza, recombinant, injectable, preservative free||S|PF|Y
C3644201|T121|155|CVX|influenza, recombinant, injectable, preservative free||S|PF|Y
C3644201|T129|155|CVX|Seasonal, trivalent, recombinant, injectable influenza vaccine, preservative free||P|PF|Y
C3644201|T121|155|CVX|Seasonal, trivalent, recombinant, injectable influenza vaccine, preservative free||P|PF|Y
C3833494|T121|156|CVX|Rho(D) Immune globulin- IV or IM||P|PF|Y
C3833494|T129|156|CVX|Rho(D) Immune globulin- IV or IM||P|PF|Y
C3833494|T121|156|CVX|Rho(D)-IG||S|PF|Y
C3833494|T129|156|CVX|Rho(D)-IG||S|PF|Y
C3833495|T121|157|CVX|Rho(D) -IG IM||S|PF|Y
C3833495|T129|157|CVX|Rho(D) -IG IM||S|PF|Y
C3833495|T121|157|CVX|Rho(D) Immune globulin - IM||P|PF|Y
C3833495|T129|157|CVX|Rho(D) Immune globulin - IM||P|PF|Y
C3833496|T121|158|CVX|influenza, injectable, quadrivalent||S|PF|Y
C3833496|T129|158|CVX|influenza, injectable, quadrivalent||S|PF|Y
C3833496|T121|158|CVX|influenza, injectable, quadrivalent, contains preservative||P|PF|Y
C3833496|T129|158|CVX|influenza, injectable, quadrivalent, contains preservative||P|PF|Y
C3833497|T121|159|CVX|Rho(D) - Unspecified formulation||P|VO|Y
C3833497|T129|159|CVX|Rho(D) - Unspecified formulation||P|VO|Y
C3833497|T121|159|CVX|Rho(D) Unspecified formulation||P|PF|Y
C3833497|T129|159|CVX|Rho(D) Unspecified formulation||P|PF|Y
C3833498|T121|160|CVX|Influenza A monovalent (H5N1), ADJUVANTED-2013||S|PF|Y
C3833498|T129|160|CVX|Influenza A monovalent (H5N1), ADJUVANTED-2013||S|PF|Y
C3833498|T121|160|CVX|Influenza A monovalent (H5N1), adjuvanted, National stockpile 2013||P|PF|Y
C3833498|T129|160|CVX|Influenza A monovalent (H5N1), adjuvanted, National stockpile 2013||P|PF|Y
C3833499|T121|801|CVX|AS03 Adjuvant||P|PF|N
C3833499|T121|801|CVX|AS03 Adjuvant||P|PF|Y
C3833499|T129|801|CVX|AS03 Adjuvant||P|PF|N
C3833499|T129|801|CVX|AS03 Adjuvant||P|PF|Y
C3864305|T129|161|CVX|Influenza, injectable,quadrivalent, preservative free, pediatric||P|PF|N
C3864305|T129|161|CVX|Influenza, injectable,quadrivalent, preservative free, pediatric||P|PF|Y
C3864305|T121|161|CVX|Influenza, injectable,quadrivalent, preservative free, pediatric||P|PF|N
C3864305|T121|161|CVX|Influenza, injectable,quadrivalent, preservative free, pediatric||P|PF|Y
C3864306|T121|162|CVX|meningococcal B vaccine, fully recombinant||P|PF|Y
C3864306|T129|162|CVX|meningococcal B vaccine, fully recombinant||P|PF|Y
C3864306|T121|162|CVX|meningococcal B, recombinant||S|PF|Y
C3864306|T129|162|CVX|meningococcal B, recombinant||S|PF|Y
C3864307|T121|163|CVX|meningococcal B vaccine, recombinant, OMV, adjuvanted||P|PF|Y
C3864307|T129|163|CVX|meningococcal B vaccine, recombinant, OMV, adjuvanted||P|PF|Y
C3864307|T121|163|CVX|meningococcal B, OMV||S|PF|Y
C3864307|T129|163|CVX|meningococcal B, OMV||S|PF|Y
C3864308|T121|164|CVX|meningococcal B, unspecified||S|PF|Y
C3864308|T129|164|CVX|meningococcal B, unspecified||S|PF|Y
C3864308|T121|164|CVX|meningococcal B, unspecified formulation||P|PF|Y
C3864308|T129|164|CVX|meningococcal B, unspecified formulation||P|PF|Y
C3864309|T129|165|CVX|HPV9||S|PF|Y
C3864309|T121|165|CVX|HPV9||S|PF|Y
C3864309|T129|165|CVX|Human Papillomavirus 9-valent vaccine||P|VCW|Y
C3864309|T121|165|CVX|Human Papillomavirus 9-valent vaccine||P|VCW|Y
C3864309|T129|N0000191285|NDFRT|PAPILLOMAVIRUS HUMAN 9-VALENT VACCINE||P|PF|N
C3864309|T121|N0000191285|NDFRT|PAPILLOMAVIRUS HUMAN 9-VALENT VACCINE||P|PF|N
C3864309|T129|4033963|VANDF|PAPILLOMAVIRUS HUMAN 9-VALENT VACCINE||P|PF|Y
C3864309|T121|4033963|VANDF|PAPILLOMAVIRUS HUMAN 9-VALENT VACCINE||P|PF|Y
C3864310|T129|166|CVX|influenza, intradermal, quadrivalent, preservative free||S|PF|Y
C3864310|T121|166|CVX|influenza, intradermal, quadrivalent, preservative free||S|PF|Y
C3864310|T129|166|CVX|influenza, intradermal, quadrivalent, preservative free, injectable||P|PF|Y
C3864310|T121|166|CVX|influenza, intradermal, quadrivalent, preservative free, injectable||P|PF|Y
C4048265|T129|13|CVX|tetanus immune globulin||P|VC|N
C4048265|T116|13|CVX|tetanus immune globulin||P|VC|N
C4048265|T121|13|CVX|tetanus immune globulin||P|VC|N
C4048265|T129|13|CVX|TIG||S|PF|N
C4048265|T116|13|CVX|TIG||S|PF|N
C4048265|T121|13|CVX|TIG||S|PF|N
C4048265|T129|13|HL7V2.5|TIG||S|PF|N
C4048265|T116|13|HL7V2.5|TIG||S|PF|N
C4048265|T121|13|HL7V2.5|TIG||S|PF|N
C4048265|T129|13|HL7V3.0|TIG||S|PF|Y
C4048265|T116|13|HL7V3.0|TIG||S|PF|Y
C4048265|T121|13|HL7V3.0|TIG||S|PF|Y
C4048265|T129|5557|MMSL|tetanus immune globulin||P|VC|N
C4048265|T116|5557|MMSL|tetanus immune globulin||P|VC|N
C4048265|T121|5557|MMSL|tetanus immune globulin||P|VC|N
C4048265|T129|d01137|MMSL|tetanus immune globulin||P|VC|Y
C4048265|T116|d01137|MMSL|tetanus immune globulin||P|VC|Y
C4048265|T121|d01137|MMSL|tetanus immune globulin||P|VC|Y
C4048265|T129|NOCODE|MTH|Tetanus immune globulin||P|PF|Y
C4048265|T116|NOCODE|MTH|Tetanus immune globulin||P|PF|Y
C4048265|T121|NOCODE|MTH|Tetanus immune globulin||P|PF|Y
C4048265|T129|N0000020185|NDFRT|TETANUS IMMUNE GLOBULIN||P|VC|N
C4048265|T116|N0000020185|NDFRT|TETANUS IMMUNE GLOBULIN||P|VC|N
C4048265|T121|N0000020185|NDFRT|TETANUS IMMUNE GLOBULIN||P|VC|N
C4048265|T129|1727875|RXNORM|Tetanus immune globulin||P|PF|N
C4048265|T116|1727875|RXNORM|Tetanus immune globulin||P|PF|N
C4048265|T121|1727875|RXNORM|Tetanus immune globulin||P|PF|N
C4048265|T129|170458003|SNOMEDCT_US|Anti-Tetanus immunoglobulin||S|PF|Y
C4048265|T116|170458003|SNOMEDCT_US|Anti-Tetanus immunoglobulin||S|PF|Y
C4048265|T121|170458003|SNOMEDCT_US|Anti-Tetanus immunoglobulin||S|PF|Y
C4048265|T129|412313000|SNOMEDCT_US|Tetanus immunoglobulin||S|PF|N
C4048265|T116|412313000|SNOMEDCT_US|Tetanus immunoglobulin||S|PF|N
C4048265|T121|412313000|SNOMEDCT_US|Tetanus immunoglobulin||S|PF|N
C4048265|T129|425682001|SNOMEDCT_US|Tetanus immunoglobulin||S|PF|Y
C4048265|T116|425682001|SNOMEDCT_US|Tetanus immunoglobulin||S|PF|Y
C4048265|T121|425682001|SNOMEDCT_US|Tetanus immunoglobulin||S|PF|Y
C4048265|T129|425682001|SNOMEDCT_US|Tetanus immunoglobulin (substance)||S|PF|Y
C4048265|T116|425682001|SNOMEDCT_US|Tetanus immunoglobulin (substance)||S|PF|Y
C4048265|T121|425682001|SNOMEDCT_US|Tetanus immunoglobulin (substance)||S|PF|Y
C4048265|T129|4022179|VANDF|TETANUS IMMUNE GLOBULIN||P|VC|Y
C4048265|T116|4022179|VANDF|TETANUS IMMUNE GLOBULIN||P|VC|Y
C4048265|T121|4022179|VANDF|TETANUS IMMUNE GLOBULIN||P|VC|Y
C4067702|T121|108|CVX|meningococcal ACWY vaccine, unspecified formulation||P|PF|Y
C4067702|T129|108|CVX|meningococcal ACWY vaccine, unspecified formulation||P|PF|Y
C4067702|T121|108|CVX|meningococcal ACWY, unspecified formulation||S|PF|Y
C4067702|T129|108|CVX|meningococcal ACWY, unspecified formulation||S|PF|Y
C4067703|T129|167|CVX|meningococcal vaccine of unknown formulation and unknown serogroups||P|PF|Y
C4067703|T121|167|CVX|meningococcal vaccine of unknown formulation and unknown serogroups||P|PF|Y
C4067703|T129|167|CVX|meningococcal, unknown serogroups||S|PF|Y
C4067703|T121|167|CVX|meningococcal, unknown serogroups||S|PF|Y
C4067704|T121|168|CVX|influenza, trivalent, adjuvanted||S|PF|Y
C4067704|T129|168|CVX|influenza, trivalent, adjuvanted||S|PF|Y
C4067704|T121|168|CVX|Seasonal trivalent influenza vaccine, adjuvanted, preservative free||P|PF|Y
C4067704|T129|168|CVX|Seasonal trivalent influenza vaccine, adjuvanted, preservative free||P|PF|Y