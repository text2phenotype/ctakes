// CUI|TUI|CODE|VOCAB|TXT|PREF TEXT
C000001|T034|6|CUSTOM|Sodium|Sodium