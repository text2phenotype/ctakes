C0419735|T129||CVX|PATIENT IMMUNE TO HEPATITIS A
C0419735|T129||CVX|PATIENT IMMUNE TO HEP A
C0419735|T129||CVX|PATIENT VACCINATED FOR HEP A
C1170008|T129||CVX|HEPATITIS A AND HEPATITIS B VACCINE
C0419735|T129||CVX|HEPATITIS A IMMUNIZATION (SNOMED:243789007)
C3526526|T129||CVX|HEPATITIS A VACCINE, ADULT DOSAGE
C0694731|T129||CVX|HEPATITIS A VACCINE, PEDIATRIC DOSAGE, UNSPECIFIED FORMULATION
C1548491|T129|83|CVX|HEPATITIS A VACCINE, PEDIATRIC/ADOLESCENT DOSAGE, 2 DOSE SCHEDULE|HEP A, PED/ADOL, 2 DOSE
C1548492|T129|84|CVX|HEPATITIS A VACCINE, PEDIATRIC/ADOLESCENT DOSAGE, 3 DOSE SCHEDULE|HEP A, PED/ADOL, 3 DOSE
C3644157|T129||CVX|HEPATITIS A VACCINE, UNSPECIFIED FORMULATION
C1548491|T129|83|CVX|HEP A, PED/ADOL, 2 DOSE|HEP A, PED/ADOL, 2 DOSE
C1548492|T129|84|CVX|HEP A, PED/ADOL, 3 DOSE|HEP A, PED/ADOL, 3 DOSE
C0694731|T129||CVX|HEP A, PEDIATRIC, UNSPECIFIED FORMULATION
C3644157|T129||CVX|HEP A, UNSPECIFIED FORMULATION
C1170008|T129||CVX|HEP A-HEP B
C0730242|T129||CVX|COMBINED HEPATITIS A & HEPATITIS B VACCINATION
C0730242|T129||CVX|COMBINED HEPATITIS A AND HEPATITIS B VACCINATION 
C0730242|T129||CVX|COMBINED HEPATITIS A AND HEPATITIS B VACCINATION
C0730242|T129||CVX|COMBINED HEPATITIS A AND B VACCINATION
C0730242|T129||CVX|COMBINED HEPATITIS A AND B VACCINATION 
C1281986|T129||CVX|HEPATITIS A AND TYPHOID VACCINATION 
C1281986|T129||CVX|HEPATITIS A AND TYPHOID VACCINATION
C0419735|T129||CVX|IMMUNISATION;HEPATITIS A
C0419735|T129||CVX|HEPATITIS A IMMUNIZATION
C0419735|T129||CVX|HEPATITIS A IMMUNISATION
C0419735|T129||CVX|HEPATITIS A IMMUNISATION 
C0419735|T129||CVX|HEPATITIS A VACCINE ADMINISTRATION 
C0419735|T129||CVX|HEPATITIS A VACCINE ADMINISTRATION
C0419735|T129||CVX|HEPATITIS A VACCINATION
C0419735|T129||CVX|HEPATITIS A VACCINATION, UNSPECIFIED
C0419735|T129||CVX|HEPATITIS A IMMUNIZATION 
C0419735|T129||CVX|IMMUNIZATION;HEPATITIS A
C0419736|T129||CVX|FIRST HEPATITIS A VACCINATION 
C0419736|T129||CVX|FIRST HEPATITIS A VACCINATION
C0419736|T129||CVX|FIRST HEPATITIS A VACCINATION 
C0419736|T129||CVX|HEPATITIS A VACCINES FIRST VACCINATION
C0419736|T129||CVX|1ST HEPATITIS A VACCINATION
C0419737|T129||CVX|SECOND HEPATITIS A VACCINATION
C0419737|T129||CVX|SECOND HEPATITIS A VACCINATION 
C0419737|T129||CVX|SECOND HEPATITIS A VACCINATION 
C0419737|T129||CVX|HEPATITIS A VACCINES SECOND VACCINATION
C0419737|T129||CVX|2ND HEPATITIS A VACCINATION
C0419739|T129||CVX|BOOSTER HEPATITIS A VACCINATION
C0419739|T129||CVX|BOOSTER HEPATITIS A VACCINATION 
C0419738|T129||CVX|THIRD HEPATITIS A VACCINATION
C0419738|T129||CVX|THIRD HEPATITIS A VACCINATION 
C0419738|T129||CVX|3RD HEPATITIS A VACCINATION
C1170689|T129||CVX|TWINRIX JUNIOR
C1170008|T129||CVX|HEPATITIS A AND HEPATITIS B VACCINE
C1170008|T129||CVX|HEP A-HEP B
C1170008|T129||CVX|HEPATITIS A-HEPATITIS B VACCINE
C3526526|T129||CVX|HEPATITIS A VACCINE, ADULT DOSAGE
C3526526|T129||CVX|HEP A, ADULT
C0694731|T129||CVX|HEP A, PEDIATRIC, UNSPECIFIED FORMULATION
C0694731|T129||CVX|HEPATITIS A VACCINE, PEDIATRIC DOSAGE, UNSPECIFIED FORMULATION
C0694731|T129||CVX|HEP A, PEDIATRIC, NOS
C1548491|T129|83|CVX|HEP A, PED/ADOL, 2 DOSE|HEP A, PED/ADOL, 2 DOSE
C1548491|T129|83|CVX|HEPATITIS A VACCINE, PEDIATRIC/ADOLESCENT DOSAGE, 2 DOSE SCHEDULE|HEP A, PED/ADOL, 2 DOSE
C1548492|T129|84|CVX|HEPATITIS A VACCINE, PEDIATRIC/ADOLESCENT DOSAGE, 3 DOSE SCHEDULE|HEP A, PED/ADOL, 3 DOSE
C1548492|T129|84|CVX|HEP A, PED/ADOL, 3 DOSE|HEP A, PED/ADOL, 3 DOSE
C3644157|T129||CVX|HEP A, UNSPECIFIED FORMULATION
C3644157|T129||CVX|HEPATITIS A VACCINE, UNSPECIFIED FORMULATION
