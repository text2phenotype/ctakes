C3871344|T033||HCPCS|CURRENT OR FORMER INJECTION DRUG USER (EVEN ONCE)
C3871344|T033||HCPCS|CURRENT OR FORMER INJECTION DRUG USER
C3871344|T033||HCPCS|CURRENT OR FORMER IV DRUG USER
C3871344|T033||HCPCS|CURRENT OR FORMER IV USER
C3871344|T033||HCPCS|CURRENT IV USER
C3871344|T033||HCPCS|FORMER IV USER
C3871344|T033||HCPCS|FORMER IV DRUG USER
C3871344|T033||HCPCS|HISTORY OF INJECTION DRUG USE
C3871344|T033||HCPCS|HISTORY OF IV DRUG USE
C3871344|T033||HCPCS|HISTORY OF IV USE
C3871344|T033||HCPCS|HX INJEC DRUG USE
C3871344|T033||HCPCS|HX IV USE
C3871344|T033||HCPCS|HISTORY IV USE
C3871344|T033||HCPCS|USES IV NEEDLES
C3871344|T033||HCPCS|IV DRUG USER
C3871344|T033||HCPCS|HISTORY OF INJECTION DRUG USE
C3871344|T033||HCPCS|HX INJEC DRUG USE
