C0004096|T047|195979001|SNOMEDCT_US|ASTHMA|ASTHMA UNSPECIFIED (DISORDER)
C0340067|T047|93432008|SNOMEDCT_US|DRUG-INDUCED ASTHMA |DRUG-INDUCED ASTHMA (DISORDER)
C0340067|T047|93432008|SNOMEDCT_US|ASTHMA DRUG-INDUCED|DRUG-INDUCED ASTHMA (DISORDER)
C0340067|T047|93432008|SNOMEDCT_US|DRUG-INDUCED ASTHMA|DRUG-INDUCED ASTHMA (DISORDER)
C0340067|T047|93432008|SNOMEDCT_US|DRUG-INDUCED ASTHMA |DRUG-INDUCED ASTHMA (DISORDER)
C0340067|T047|93432008|SNOMEDCT_US|DRUG-INDUCED ASTHMA, NOS|DRUG-INDUCED ASTHMA (DISORDER)
C0348819|T047|195977004|SNOMEDCT_US|MIXED ASTHMA|MIXED ASTHMA (DISORDER)
C0348819|T047|195977004|SNOMEDCT_US|ASTHMA MIXED|MIXED ASTHMA (DISORDER)
C0348819|T047|195977004|SNOMEDCT_US|MIXED ASTHMA |MIXED ASTHMA (DISORDER)
C0348819|T047|195977004|SNOMEDCT_US|MIXED ASTHMA |MIXED ASTHMA (DISORDER)
C0348819|T047|195977004|SNOMEDCT_US|ASTHMA; MIXED|MIXED ASTHMA (DISORDER)
C0348819|T047|195977004|SNOMEDCT_US|MIXED; ASTHMA|MIXED ASTHMA (DISORDER)
C0858626|T047||SNOMEDCT_US|ASTHMATIC ATTACK INDUCED
C0856716|T047||SNOMEDCT_US|ASPIRIN-SENSITIVE ASTHMA
C0856716|T047||SNOMEDCT_US|ASPIRIN ASTHMA
C0856716|T047||SNOMEDCT_US|ASTHMA ASPIRIN-SENSITIVE
C0859194|T047||SNOMEDCT_US|CHRONIC OBSTRUCTIVE ASTHMA (WITH OBSTRUCTIVE PULMONARY DISEASE), W/O-MENT OF STATUS ASTHMATICUS
C0859194|T047||SNOMEDCT_US|CHRONIC OBSTRUCTIVE ASTHMA (WITH OBSTRUCTIVE PULMONARY DISEASE), W/O MENT OF STATUS ASTHMATICUS
C0494660|T047||SNOMEDCT_US|PREDOMINANTLY ALLERGIC ASTHMA
C0494660|T047||SNOMEDCT_US|ALLERGIC (PREDOMINANTLY) ASTHMA
C0494660|T047||SNOMEDCT_US|ASTHMA; PREDOMINANTLY ALLERGIC
C0494660|T047||SNOMEDCT_US|PREDOMINANTLY ALLERGIC; ASTHMA
C0155883|T047||SNOMEDCT_US|CHRONIC OBSTRUCTIVE ASTHMA
C0155883|T047||SNOMEDCT_US|CHRONIC OBSTRUCTIVE ASTHMA 
C0155883|T047||SNOMEDCT_US|CHRONIC OBSTRUCTIVE ASTHMA (WITH OBSTRUCTIVE PULMONARY DISEASE)
C0948683|T047||SNOMEDCT_US|ASTHMATIC ATTACK ATOPIC
C0155879|T047|266360009|SNOMEDCT_US|EXTRINSIC ASTHMA WITH STATUS ASTHMATICUS|EXTRINSIC ASTHMA WITH STATUS ASTHMATICUS (DISORDER)
C0155879|T047|266360009|SNOMEDCT_US|EXTRINSIC ASTHMA WITH STATUS ASTHMATICUS |EXTRINSIC ASTHMA WITH STATUS ASTHMATICUS (DISORDER)
C0155879|T047|266360009|SNOMEDCT_US|EXT ASTHMA W STATUS ASTH|EXTRINSIC ASTHMA WITH STATUS ASTHMATICUS (DISORDER)
C0155879|T047|266360009|SNOMEDCT_US|EXTRINSIC ASTHMA WITH STATUS ASTHMATICUS |EXTRINSIC ASTHMA WITH STATUS ASTHMATICUS (DISORDER)
C0155880|T047|195976008|SNOMEDCT_US|NONALLERGIC ASTHMA|INTRINSIC ASTHMA NOS (DISORDER)
C0155880|T047|195976008|SNOMEDCT_US|INTRINSIC ASTHMA|INTRINSIC ASTHMA NOS (DISORDER)
C0155880|T047|195976008|SNOMEDCT_US|INTRINSIC ASTHMA |INTRINSIC ASTHMA NOS (DISORDER)
C0155880|T047|195976008|SNOMEDCT_US|INTRINSIC NONALLERGIC ASTHMA|INTRINSIC ASTHMA NOS (DISORDER)
C0155880|T047|195976008|SNOMEDCT_US|INTRINSIC ASTHMA |INTRINSIC ASTHMA NOS (DISORDER)
C0155880|T047|195976008|SNOMEDCT_US|INTRINSIC ASTHMA NOS|INTRINSIC ASTHMA NOS (DISORDER)
C0155880|T047|195976008|SNOMEDCT_US|INTRINSIC ASTHMA NOS |INTRINSIC ASTHMA NOS (DISORDER)
C0155880|T047|195976008|SNOMEDCT_US|NON-ALLERGIC ASTHMA|INTRINSIC ASTHMA NOS (DISORDER)
C0155880|T047|195976008|SNOMEDCT_US|NON-ALLERGIC ASTHMA |INTRINSIC ASTHMA NOS (DISORDER)
C0155880|T047|195976008|SNOMEDCT_US|ASTHMA NON-ALLERGIC|INTRINSIC ASTHMA NOS (DISORDER)
C0155880|T047|195976008|SNOMEDCT_US|ASTHMA DUE TO INTERNAL IMMUNOLOGICAL PROCESS|INTRINSIC ASTHMA NOS (DISORDER)
C0155880|T047|195976008|SNOMEDCT_US|NON-ALLERGIC ASTHMA |INTRINSIC ASTHMA NOS (DISORDER)
C0155880|T047|195976008|SNOMEDCT_US|ASTHMA; INTRINSIC, NONALLERGIC|INTRINSIC ASTHMA NOS (DISORDER)
C0155880|T047|195976008|SNOMEDCT_US|ASTHMA; INTRINSIC|INTRINSIC ASTHMA NOS (DISORDER)
C0155880|T047|195976008|SNOMEDCT_US|ASTHMA; NONALLERGIC|INTRINSIC ASTHMA NOS (DISORDER)
C0155880|T047|195976008|SNOMEDCT_US|INTRINSIC; ASTHMA, NONALLERGIC|INTRINSIC ASTHMA NOS (DISORDER)
C0155880|T047|195976008|SNOMEDCT_US|INTRINSIC; ASTHMA|INTRINSIC ASTHMA NOS (DISORDER)
C0155880|T047|195976008|SNOMEDCT_US|NONALLERGIC; ASTHMA|INTRINSIC ASTHMA NOS (DISORDER)
C0155880|T047|195976008|SNOMEDCT_US|INTRINSIC ASTHMA  [AMBIGUOUS]|INTRINSIC ASTHMA NOS (DISORDER)
C0155882|T047|266362001|SNOMEDCT_US|INTRINSIC ASTHMA WITH STATUS ASTHMATICUS |INTRINSIC ASTHMA WITH STATUS ASTHMATICUS (DISORDER)
C0155882|T047|266362001|SNOMEDCT_US|INTRINSIC ASTHMA WITH STATUS ASTHMATICUS|INTRINSIC ASTHMA WITH STATUS ASTHMATICUS (DISORDER)
C0155882|T047|266362001|SNOMEDCT_US|INT ASTHMA W STATUS ASTH|INTRINSIC ASTHMA WITH STATUS ASTHMATICUS (DISORDER)
C0155882|T047|266362001|SNOMEDCT_US|INTRINSIC ASTHMA WITH STATUS ASTHMATICUS |INTRINSIC ASTHMA WITH STATUS ASTHMATICUS (DISORDER)
C0155878|T047||SNOMEDCT_US|EXTRINSIC ASTHMA WITHOUT MENTION OF STATUS ASTHMATICUS
C0155878|T047||SNOMEDCT_US|EXTRINSIC ASTHMA NOS
C0155878|T047||SNOMEDCT_US|EXTRINSIC ASTHMA, UNSPECIFIED
C0155881|T047||SNOMEDCT_US|INTRINSIC ASTHMA WITHOUT MENTION OF STATUS ASTHMATICUS
C0155881|T047||SNOMEDCT_US|INTRINSIC ASTHMA NOS
C0155881|T047||SNOMEDCT_US|INTRINSIC ASTHMA, UNSPECIFIED
C0155886|T047||SNOMEDCT_US|ASTHMA, UNSPECIFIED TYPE, WITHOUT MENTION OF STATUS ASTHMATICUS
C0155886|T047||SNOMEDCT_US|ASTHMA NOS
C0155886|T047||SNOMEDCT_US|ASTHMA, UNSPECIFIED TYPE, UNSPECIFIED
C0549336|T047||SNOMEDCT_US|ASTHMA AGGRAVATED
C0347950|T047|266364000|SNOMEDCT_US|ASTHMA ATTACK|ASTHMA ATTACK (DISORDER)
C0347950|T047|266364000|SNOMEDCT_US|ASTHMA ATTACK NOS |ASTHMA ATTACK (DISORDER)
C0347950|T047|266364000|SNOMEDCT_US|ASTHMA ATTACK (& NOS) |ASTHMA ATTACK (DISORDER)
C0347950|T047|266364000|SNOMEDCT_US|ASTHMA ATTACK (& NOS)|ASTHMA ATTACK (DISORDER)
C0347950|T047|266364000|SNOMEDCT_US|ASTHMA ATTACK NOS|ASTHMA ATTACK (DISORDER)
C0347950|T047|266364000|SNOMEDCT_US|ASTHMA ATTACK |ASTHMA ATTACK (DISORDER)
C0347950|T047|266364000|SNOMEDCT_US|ASTHMA ATTACK |ASTHMA ATTACK (DISORDER)
C0347950|T047|266364000|SNOMEDCT_US|ACUTE EXACERBATION OF ASTHMA|ASTHMA ATTACK (DISORDER)
C0347950|T047|266364000|SNOMEDCT_US|ACUTE EXACERBATION OF ASTHMA |ASTHMA ATTACK (DISORDER)
C0347950|T047|266364000|SNOMEDCT_US|ASTHMATIC ATTACK|ASTHMA ATTACK (DISORDER)
C0810292|T047||SNOMEDCT_US|OTHER AND UNSPECIFIED ASTHMA
C0004096|T047|195979001|SNOMEDCT_US|ASTHMA|ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|ASTHMAS|ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|ASTHMA, UNSPECIFIED|ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|BRONCHIAL ASTHMA|ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|ASTHMA |ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|BR. ASTHMA|ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|ASTHMA NOS|ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|UNSPECIFIED ASTHMA|ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|ASTHMA [DISEASE/FINDING]|ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|ASTHMA, BRONCHIAL|ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|ASTHMA |ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|ASTHMA UNSPECIFIED |ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|ASTHMA NOS |ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|ASTHMA UNSPECIFIED|ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|-- ASTHMA|ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|ASTHMATIC|ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|ASTHMA BRONCHIAL|ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|BRONCHITIC ASTHMA|ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|CARDIO/PULM: ASTHMA|ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|AIRWAY HYPERREACTIVITY|ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|ASTHMA, NOS|ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|BRONCHIAL ASTHMA, NOS|ASTHMA UNSPECIFIED (DISORDER)
C0004096|T047|195979001|SNOMEDCT_US|ASTHMA  [AMBIGUOUS]|ASTHMA UNSPECIFIED (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|ASTHMATIC CRISES|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|ASTHMATIC SHOCKS|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|ASTHMATICUS, STATUS|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|CRISES, ASTHMATIC|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|CRISIS, ASTHMATIC|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|SHOCK, ASTHMATIC|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|SHOCKS, ASTHMATIC|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|STATUS ASTHMATICUS|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|STATUS ASTHMATICUS -RETIRED-|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|ASTHMA W STATUS ASTHMAT|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|ASTHMATIC SHOCK|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|STATUS ASTHMATICUS [DISEASE/FINDING]|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|ASTHMATIC CRISIS|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|STATUS ASTHMATICUS NOS|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS)|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|STATUS ASTHMATICUS NOS |(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|STATUS ASTHMATICUS |(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|SEVERE ASTHMA ATTACK|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) |(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|ACUTE SEVERE ASTHMA|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|ASTHMA WITH STATUS ASTHMATICUS|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|ACUTE SEVERE EXACERBATION OF ASTHMA|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|ASTHMA WITH STATUS ASTHMATICUS |(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|ACUTE SEVERE EXACERBATION OF ASTHMA |(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|ASTHMA, UNSPECIFIED TYPE, WITH STATUS ASTHMATICUS|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|ASTHMA WITH STATUS ASTHMATICUS |(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|ASTHMATICUS; STATUS|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0038218|T047|195980003|SNOMEDCT_US|STATUS; ASTHMATICUS|(SEVERE ASTHMA ATTACK) OR (STATUS ASTHMATICUS NOS) (DISORDER)
C0004099|T047|139202009|SNOMEDCT_US|ASTHMA, EXERCISE INDUCED|EXERCISE-INDUCED ASTHMA (FINDING)
C0004099|T047|139202009|SNOMEDCT_US|ASTHMA, EXERCISE-INDUCED|EXERCISE-INDUCED ASTHMA (FINDING)
C0004099|T047|139202009|SNOMEDCT_US|ASTHMAS, EXERCISE-INDUCED|EXERCISE-INDUCED ASTHMA (FINDING)
C0004099|T047|139202009|SNOMEDCT_US|EXERCISE INDUCED ASTHMA|EXERCISE-INDUCED ASTHMA (FINDING)
C0004099|T047|139202009|SNOMEDCT_US|EXERCISE-INDUCED ASTHMAS|EXERCISE-INDUCED ASTHMA (FINDING)
C0004099|T047|139202009|SNOMEDCT_US|EXERCISE IND ASTHMA|EXERCISE-INDUCED ASTHMA (FINDING)
C0004099|T047|139202009|SNOMEDCT_US|ASTHMA EXERCISE IND|EXERCISE-INDUCED ASTHMA (FINDING)
C0004099|T047|139202009|SNOMEDCT_US|EXERCISE-INDUCED ASTHMA|EXERCISE-INDUCED ASTHMA (FINDING)
C0004099|T047|139202009|SNOMEDCT_US|EXERCISE-INDUCED ASTHMA |EXERCISE-INDUCED ASTHMA (FINDING)
C0004099|T047|139202009|SNOMEDCT_US|EIA (EXERCISE-INDUCED ASTHMA)|EXERCISE-INDUCED ASTHMA (FINDING)
C0004099|T047|139202009|SNOMEDCT_US|ASTHMA EXERCISE INDUCED|EXERCISE-INDUCED ASTHMA (FINDING)
C0004099|T047|139202009|SNOMEDCT_US|ASTHMA, EXERCISE-INDUCED [DISEASE/FINDING]|EXERCISE-INDUCED ASTHMA (FINDING)
C0004099|T047|139202009|SNOMEDCT_US|EXERCISE-INDUCED ASTHMA |EXERCISE-INDUCED ASTHMA (FINDING)
C0004099|T047|139202009|SNOMEDCT_US|EIA - EXERCISE-INDUCED ASTHMA|EXERCISE-INDUCED ASTHMA (FINDING)
C0004099|T047|139202009|SNOMEDCT_US|EXERCISE-INDUCED ASTHMA |EXERCISE-INDUCED ASTHMA (FINDING)
C1319853|T047|407674008|SNOMEDCT_US|ASPIRIN INDUCED ASTHMAS|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|ASPIRIN-INDUCED ASTHMAS|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|NSAID-INDUCED ASTHMAS|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|ASPIRIN-INDUCED ASTHMA SYNDROMES|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|ASTHMA SYNDROME, ASPIRIN-INDUCED|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|ASTHMA, NSAID INDUCED|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|SYNDROME, ASPIRIN-INDUCED ASTHMA|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|SYNDROMES, ASPIRIN-INDUCED ASTHMA|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|ASTHMAS, ASPIRIN-INDUCED|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|ASTHMA, ASPIRIN INDUCED|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|ASTHMA SYNDROMES, ASPIRIN-INDUCED|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|ASTHMAS, ASPIRIN INDUCED|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|INDUCED ASTHMAS, ASPIRIN|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|ASTHMA, ASPIRIN-INDUCED|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|ASTHMAS, NSAID-INDUCED|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|NSAID-INDUCED ASTHMA|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|ASPIRIN INDUCED ASTHMA SYNDROME|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|INDUCED ASTHMA, ASPIRIN|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|ASTHMA, NSAID-INDUCED|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|ASTHMA, ASPIRIN-INDUCED [DISEASE/FINDING]|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|ASPIRIN INDUCED ASTHMA|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|ASPIRIN-INDUCED ASTHMA|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|ASPIRIN-INDUCED ASTHMA SYNDROME|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|ASPIRIN-INDUCED ASTHMA |ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|ASTHMA DRUG-INDUCED ASPIRIN|ASPIRIN-INDUCED ASTHMA (DISORDER)
C1319853|T047|407674008|SNOMEDCT_US|ASPIRIN-INDUCED ASTHMA |ASPIRIN-INDUCED ASTHMA (DISORDER)
C1960045|T047|427679007|SNOMEDCT_US|MILD INTERMITTENT ASTHMA|MILD INTERMITTENT ASTHMA (DISORDER)
C1960045|T047|427679007|SNOMEDCT_US|MILD INTERMITTENT ASTHMA |MILD INTERMITTENT ASTHMA (DISORDER)
C1960045|T047|427679007|SNOMEDCT_US|MILD INTERMITTENT ASTHMA |MILD INTERMITTENT ASTHMA (DISORDER)
C1960045|T047|427679007|SNOMEDCT_US|MILD INTERMITTENT ASTHMA NOS|MILD INTERMITTENT ASTHMA (DISORDER)
C1960046|T047|426979002|SNOMEDCT_US|MILD PERSISTENT ASTHMA |MILD PERSISTENT ASTHMA (DISORDER)
C1960046|T047|426979002|SNOMEDCT_US|MILD PERSISTENT ASTHMA|MILD PERSISTENT ASTHMA (DISORDER)
C1960046|T047|426979002|SNOMEDCT_US|MILD PERSISTENT ASTHMA |MILD PERSISTENT ASTHMA (DISORDER)
C1960046|T047|426979002|SNOMEDCT_US|MILD PERSISTENT ASTHMA NOS|MILD PERSISTENT ASTHMA (DISORDER)
C1960047|T047|427295004|SNOMEDCT_US|MODERATE PERSISTENT ASTHMA|MODERATE PERSISTENT ASTHMA (DISORDER)
C1960047|T047|427295004|SNOMEDCT_US|MODERATE PERSISTENT ASTHMA |MODERATE PERSISTENT ASTHMA (DISORDER)
C1960047|T047|427295004|SNOMEDCT_US|MODERATE PERSISTENT ASTHMA |MODERATE PERSISTENT ASTHMA (DISORDER)
C1960047|T047|427295004|SNOMEDCT_US|MODERATE PERSISTENT ASTHMA NOS|MODERATE PERSISTENT ASTHMA (DISORDER)
C1960048|T047|426656000|SNOMEDCT_US|SEVERE PERSISTENT ASTHMA |SEVERE PERSISTENT ASTHMA (DISORDER)
C1960048|T047|426656000|SNOMEDCT_US|SEVERE PERSISTENT ASTHMA|SEVERE PERSISTENT ASTHMA (DISORDER)
C1960048|T047|426656000|SNOMEDCT_US|SEVERE PERSISTENT ASTHMA |SEVERE PERSISTENT ASTHMA (DISORDER)
C1960048|T047|426656000|SNOMEDCT_US|SEVERE PERSISTENT ASTHMA NOS|SEVERE PERSISTENT ASTHMA (DISORDER)
C2887463|T047||SNOMEDCT_US|UNSPECIFIED ASTHMA WITH (ACUTE) EXACERBATION
C2887464|T047||SNOMEDCT_US|UNSPECIFIED ASTHMA WITH STATUS ASTHMATICUS
C2887465|T047||SNOMEDCT_US|UNSPECIFIED ASTHMA, UNCOMPLICATED
C2919352|T047|445427006|SNOMEDCT_US|SEASONAL ASTHMA |SEASONAL ASTHMA (DISORDER)
C2919352|T047|445427006|SNOMEDCT_US|SEASONAL ASTHMA|SEASONAL ASTHMA (DISORDER)
C2919352|T047|445427006|SNOMEDCT_US|SEASONAL ASTHMA |SEASONAL ASTHMA (DISORDER)
C2919352|T047|445427006|SNOMEDCT_US|ASTHMA SEASONAL|SEASONAL ASTHMA (DISORDER)
C0349790|T047|281239006|SNOMEDCT_US|ASTHMA WITH ACUTE EXACERBATION|EXACERBATION OF ASTHMA (DISORDER)
C0349790|T047|281239006|SNOMEDCT_US|ASTHMA WITH ACUTE EXACERBATION |EXACERBATION OF ASTHMA (DISORDER)
C0349790|T047|281239006|SNOMEDCT_US|EXACERBATION OF ASTHMA |EXACERBATION OF ASTHMA (DISORDER)
C0349790|T047|281239006|SNOMEDCT_US|EXACERBATION OF ASTHMA|EXACERBATION OF ASTHMA (DISORDER)
C0349790|T047|281239006|SNOMEDCT_US|ACUTE EXACERBATION OF ASTHMA|EXACERBATION OF ASTHMA (DISORDER)
C0694548|T047|409663006|SNOMEDCT_US|COUGH VARIANT ASTHMA|COUGH VARIANT ASTHMA (DISORDER)
C0694548|T047|409663006|SNOMEDCT_US|COUGH VARIANT ASTHMA |COUGH VARIANT ASTHMA (DISORDER)
C0694548|T047|409663006|SNOMEDCT_US|COUGH VARIANT ASTHMA |COUGH VARIANT ASTHMA (DISORDER)
C0264408|T047|233678006|SNOMEDCT_US|CHILDHOOD ASTHMA |CHILDHOOD ASTHMA (DISORDER)
C0264408|T047|233678006|SNOMEDCT_US|CHILDHOOD ASTHMA|CHILDHOOD ASTHMA (DISORDER)
C0264408|T047|233678006|SNOMEDCT_US|CHILDHOOD ASTHMA NOS|CHILDHOOD ASTHMA (DISORDER)
C0264408|T047|233678006|SNOMEDCT_US|ASTHMA IN CHILDREN|CHILDHOOD ASTHMA (DISORDER)
C0264408|T047|233678006|SNOMEDCT_US|CHILDHOOD ASTHMA |CHILDHOOD ASTHMA (DISORDER)
C0264408|T047|233678006|SNOMEDCT_US|ASTHMA; CHILDHOOD|CHILDHOOD ASTHMA (DISORDER)
C0264408|T047|233678006|SNOMEDCT_US|CHILDHOOD; ASTHMA|CHILDHOOD ASTHMA (DISORDER)
C0264408|T047|233678006|SNOMEDCT_US|ASTHMA, CHILDHOOD|CHILDHOOD ASTHMA (DISORDER)
C1740754|T047|427603009|SNOMEDCT_US|INTERMITTENT ASTHMA|INTERMITTENT ASTHMA (DISORDER)
C1740754|T047|427603009|SNOMEDCT_US|INTERMITTENT ASTHMA (ASTHMA)|INTERMITTENT ASTHMA (DISORDER)
C1740754|T047|427603009|SNOMEDCT_US|INTERMITTENT ASTHMA |INTERMITTENT ASTHMA (DISORDER)
C1740754|T047|427603009|SNOMEDCT_US|INTERMITTENT ASTHMA |INTERMITTENT ASTHMA (DISORDER)
C0264423|T047|57607007|SNOMEDCT_US|OCCUPATIONAL ASTHMA |OCCUPATIONAL ASTHMA (DISORDER)
C0264423|T047|57607007|SNOMEDCT_US|OCCUPATIONAL ASTHMA|OCCUPATIONAL ASTHMA (DISORDER)
C0264423|T047|57607007|SNOMEDCT_US|ASTHMAS, OCCUPATIONAL|OCCUPATIONAL ASTHMA (DISORDER)
C0264423|T047|57607007|SNOMEDCT_US|ASTHMA, OCCUPATIONAL|OCCUPATIONAL ASTHMA (DISORDER)
C0264423|T047|57607007|SNOMEDCT_US|OCCUPATIONAL ASTHMAS|OCCUPATIONAL ASTHMA (DISORDER)
C0264423|T047|57607007|SNOMEDCT_US|ASTHMA, OCCUPATIONAL [DISEASE/FINDING]|OCCUPATIONAL ASTHMA (DISORDER)
C0264423|T047|57607007|SNOMEDCT_US|INDUSTRIAL ASTHMA|OCCUPATIONAL ASTHMA (DISORDER)
C0264423|T047|57607007|SNOMEDCT_US|OCCUPATIONAL ASTHMA |OCCUPATIONAL ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|ALLERGIC ASTHMA|ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|EXTRINSIC ASTHMA|ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|EXTRINSIC ASTHMA |ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|ATOPIC ASTHMA|ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|EXTRINSIC ALLERGIC ASTHMA|ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|EXTRINSIC ASTHMA |ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|EXTRINSIC ASTHMA NOS |ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|ALLERGIC ATOPIC ASTHMA |ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|ALLERGIC ATOPIC ASTHMA|ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|EXTRINSIC ASTHMA NOS|ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|ALLERGIC ASTHMA |ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|ASTHMA ALLERGIC|ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|ALLERGIC ASTHMA |ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|ASTHMA, ATOPIC|ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|ASTHMA EXTRINSIC|ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|ASTHMA; ALLERGIC EXTRINSIC|ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|ASTHMA; ATOPIC|ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|ASTHMA; EXTRINSIC|ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|ATOPIC; ASTHMA|ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|EXTRINSIC; ASTHMA|ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|ALLERGIC; ASTHMA, EXTRINSIC|ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|ALLERGIC; EXTRINSIC ASTHMA|ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|EXTRINSIC ASTHMA [AMBIGUOUS] |ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|ALLERGIC ATOPIC ASTHMA [AMBIGUOUS]|ALLERGIC ATOPIC ASTHMA (DISORDER)
C0155877|T047|266358007|SNOMEDCT_US|ASTHMA, ALLERGIC NOS|ALLERGIC ATOPIC ASTHMA (DISORDER)
C0264413|T047|155576005|SNOMEDCT_US|ASTHMA LATE ONSET|LATE-ONSET ASTHMA (LOA)
C0264413|T047|155576005|SNOMEDCT_US|LATE ONSET ASTHMA|LATE-ONSET ASTHMA (LOA)
C0264413|T047|155576005|SNOMEDCT_US|LOA - LATE ONSET ASTHMA|LATE-ONSET ASTHMA (LOA)
C0264413|T047|155576005|SNOMEDCT_US|LATE ONSET ASTHMA |LATE-ONSET ASTHMA (LOA)
C0264413|T047|155576005|SNOMEDCT_US|LATE-ONSET ASTHMA|LATE-ONSET ASTHMA (LOA)
C0264413|T047|155576005|SNOMEDCT_US|LATE-ONSET ASTHMA (LOA)|LATE-ONSET ASTHMA (LOA)
C0264413|T047|155576005|SNOMEDCT_US|ASTHMA LATE-ONSET|LATE-ONSET ASTHMA (LOA)
C0264413|T047|155576005|SNOMEDCT_US|LATE-ONSET ASTHMA |LATE-ONSET ASTHMA (LOA)
C0264413|T047|155576005|SNOMEDCT_US|ASTHMA; LATE ONSET|LATE-ONSET ASTHMA (LOA)
C0264413|T047|155576005|SNOMEDCT_US|LATE ONSET; ASTHMA|LATE-ONSET ASTHMA (LOA)
C0729337|T047|225057002|SNOMEDCT_US|ASTHMA BRITTLE|BRITTLE ASTHMA (DISORDER)
C0729337|T047|225057002|SNOMEDCT_US|ASTHMA BRITTLE |BRITTLE ASTHMA (DISORDER)
C0729337|T047|225057002|SNOMEDCT_US|BRITTLE ASTHMA|BRITTLE ASTHMA (DISORDER)
C0729337|T047|225057002|SNOMEDCT_US|BRITTLE ASTHMA |BRITTLE ASTHMA (DISORDER)
C3508931|T047|707444001|SNOMEDCT_US|ASTHMA UNCOMPLICATED|UNCOMPLICATED ASTHMA (DISORDER)
C3508931|T047|707444001|SNOMEDCT_US|ASTHMA UNCOMPLICATED |UNCOMPLICATED ASTHMA (DISORDER)
C3508931|T047|707444001|SNOMEDCT_US|UNCOMPLICATED ASTHMA |UNCOMPLICATED ASTHMA (DISORDER)
C3508931|T047|707444001|SNOMEDCT_US|UNCOMPLICATED ASTHMA|UNCOMPLICATED ASTHMA (DISORDER)
C0264508|T047|41997000|SNOMEDCT_US|ASTHMATIC PULMONARY ALVEOLITIS|ASTHMATIC PULMONARY ALVEOLITIS (DISORDER)
C0264508|T047|41997000|SNOMEDCT_US|ASTHMATIC PULMONARY ALVEOLITIS |ASTHMATIC PULMONARY ALVEOLITIS (DISORDER)
C0264411|T047|67415000|SNOMEDCT_US|HAY FEVER WITH ASTHMA|HAY ASTHMA (DISORDER)
C0264411|T047|67415000|SNOMEDCT_US|EXTRINSIC ASTHMA - ATOPY|HAY ASTHMA (DISORDER)
C0264411|T047|67415000|SNOMEDCT_US|HAY ASTHMA |HAY ASTHMA (DISORDER)
C0264411|T047|67415000|SNOMEDCT_US|POLLEN ASTHMA|HAY ASTHMA (DISORDER)
C0264411|T047|67415000|SNOMEDCT_US|EXTRINSIC (ATOPIC) ASTHMA|HAY ASTHMA (DISORDER)
C0264411|T047|67415000|SNOMEDCT_US|HAY ASTHMA|HAY ASTHMA (DISORDER)
C0264411|T047|67415000|SNOMEDCT_US|HAY FEVER WITH ASTHMA |HAY ASTHMA (DISORDER)
C0264411|T047|67415000|SNOMEDCT_US|HAY FEVER WITH ASTHMA |HAY ASTHMA (DISORDER)
C0264411|T047|67415000|SNOMEDCT_US|ASTHMA; HAY FEVER|HAY ASTHMA (DISORDER)
C0264411|T047|67415000|SNOMEDCT_US|HAY FEVER; ASTHMA|HAY ASTHMA (DISORDER)
C0264411|T047|67415000|SNOMEDCT_US|ASTHMA, HAY|HAY ASTHMA (DISORDER)
C0684913|T047|92807009|SNOMEDCT_US|CHEMICAL-INDUCED ASTHMA|CHEMICAL-INDUCED ASTHMA (DISORDER)
C0684913|T047|92807009|SNOMEDCT_US|ASTHMA CHEMICAL-INDUCED|CHEMICAL-INDUCED ASTHMA (DISORDER)
C0684913|T047|92807009|SNOMEDCT_US|CHEMICAL-INDUCED ASTHMA |CHEMICAL-INDUCED ASTHMA (DISORDER)
C0684913|T047|92807009|SNOMEDCT_US|CHEMICAL-INDUCED ASTHMA |CHEMICAL-INDUCED ASTHMA (DISORDER)
C0684913|T047|92807009|SNOMEDCT_US|CHEMICAL-INDUCED ASTHMA, NOS|CHEMICAL-INDUCED ASTHMA (DISORDER)
C1956414|T047|71892000|SNOMEDCT_US|CARDIAC ASTHMA|CARDIAC ASTHMA (DISORDER)
C1956414|T047|71892000|SNOMEDCT_US|ASTHMA, CARDIAC|CARDIAC ASTHMA (DISORDER)
C1956414|T047|71892000|SNOMEDCT_US|ASTHMA - CARDIAC|CARDIAC ASTHMA (DISORDER)
C1956414|T047|71892000|SNOMEDCT_US|ASTHMA CARDIAC|CARDIAC ASTHMA (DISORDER)
C1956414|T047|71892000|SNOMEDCT_US|CARDIAC ASTHMA |CARDIAC ASTHMA (DISORDER)
C1956414|T047|71892000|SNOMEDCT_US|ASTHMA; CARDIAC|CARDIAC ASTHMA (DISORDER)
C1956414|T047|71892000|SNOMEDCT_US|CARDIAC; ASTHMA|CARDIAC ASTHMA (DISORDER)
C0264404|T047|89099002|SNOMEDCT_US|CHRONIC ALLERGIC BRONCHITIS |CHRONIC ALLERGIC BRONCHITIS (DISORDER)
C0264404|T047|89099002|SNOMEDCT_US|CHRONIC ALLERGIC BRONCHITIS|CHRONIC ALLERGIC BRONCHITIS (DISORDER)
C0264404|T047|89099002|SNOMEDCT_US|ALLERGIC BRONCHITIS CHRONIC|CHRONIC ALLERGIC BRONCHITIS (DISORDER)
C0264404|T047|89099002|SNOMEDCT_US|CHRONIC ALLERGIC BRONCHITIS |CHRONIC ALLERGIC BRONCHITIS (DISORDER)
C0340070|T047|11641008|SNOMEDCT_US|MILLERS' ASTHMA|MILLERS' ASTHMA (DISORDER)
C0340070|T047|11641008|SNOMEDCT_US|MILLERS' ASTHMA |MILLERS' ASTHMA (DISORDER)
C0340070|T047|11641008|SNOMEDCT_US|ASTHMA MILLERS'|MILLERS' ASTHMA (DISORDER)
C0340070|T047|11641008|SNOMEDCT_US|MILL-WORKERS' ASTHMA|MILLERS' ASTHMA (DISORDER)
C0340070|T047|11641008|SNOMEDCT_US|GRAIN WORKER'S ASTHMA|MILLERS' ASTHMA (DISORDER)
C0340070|T047|11641008|SNOMEDCT_US|MILLERS' ASTHMA |MILLERS' ASTHMA (DISORDER)
C0006542|T047|233689004|SNOMEDCT_US|BYSSINOSES|MILL FEVER (DISORDER)
C0006542|T047|233689004|SNOMEDCT_US|BYSSINOSIS|MILL FEVER (DISORDER)
C0006542|T047|233689004|SNOMEDCT_US|MILL FEVER|MILL FEVER (DISORDER)
C0006542|T047|233689004|SNOMEDCT_US|COTTON DUST ASTHMA|MILL FEVER (DISORDER)
C0006542|T047|233689004|SNOMEDCT_US|BROWN LUNG|MILL FEVER (DISORDER)
C0006542|T047|233689004|SNOMEDCT_US|COTTON MILL FEVER|MILL FEVER (DISORDER)
C0006542|T047|233689004|SNOMEDCT_US|BYSSINOSIS |MILL FEVER (DISORDER)
C0006542|T047|233689004|SNOMEDCT_US|OCCUPATIONAL ASTHMA (BYSSINOSIS)|MILL FEVER (DISORDER)
C0006542|T047|233689004|SNOMEDCT_US|BROWN LUNGS|MILL FEVER (DISORDER)
C0006542|T047|233689004|SNOMEDCT_US|BROWN LUNG DISEASES|MILL FEVER (DISORDER)
C0006542|T047|233689004|SNOMEDCT_US|BYSSINOSIS [DISEASE/FINDING]|MILL FEVER (DISORDER)
C0006542|T047|233689004|SNOMEDCT_US|BROWN LUNG DISEASE|MILL FEVER (DISORDER)
C0006542|T047|233689004|SNOMEDCT_US|MILL FEVER |MILL FEVER (DISORDER)
C0006542|T047|233689004|SNOMEDCT_US|COTTON WORKERS' LUNG DISEASE|MILL FEVER (DISORDER)
C0006542|T047|233689004|SNOMEDCT_US|COTTON-DUST ASTHMA|MILL FEVER (DISORDER)
C0006542|T047|233689004|SNOMEDCT_US|BYSSINOSIS |MILL FEVER (DISORDER)
C0006542|T047|233689004|SNOMEDCT_US|DISEASE (OR DISORDER); RESPIRATORY TRACT, DUE TO COTTON DUST|MILL FEVER (DISORDER)
C0006542|T047|233689004|SNOMEDCT_US|FIBROSIS; LUNG, WITH BYSSINOSIS|MILL FEVER (DISORDER)
C0006542|T047|233689004|SNOMEDCT_US|LUNG; FIBROSIS, WITH BYSSINOSIS|MILL FEVER (DISORDER)
C1563057|T047|416601004|SNOMEDCT_US|WORK AGGRAVATED ASTHMA|WORK AGGRAVATED ASTHMA (DISORDER)
C1563057|T047|416601004|SNOMEDCT_US|WORK AGGRAVATED ASTHMA |WORK AGGRAVATED ASTHMA (DISORDER)
C1260881|T047|405720007|SNOMEDCT_US|FELINE ASTHMA|ALLERGIC BRONCHITIS (DISORDER)
C1319018|T047|405944004|SNOMEDCT_US|ASTHMATIC BRONCHITIS|ASTHMATIC BRONCHITIS (DISORDER)
C1319018|T047|405944004|SNOMEDCT_US|ASTHMATIC BRONCHITIS |ASTHMATIC BRONCHITIS (DISORDER)
C1319018|T047|405944004|SNOMEDCT_US|ASTHMA/BRONCHITIS|ASTHMATIC BRONCHITIS (DISORDER)
C1319018|T047|405944004|SNOMEDCT_US|ASTHMATIC BRONCHITIS NOS|ASTHMATIC BRONCHITIS (DISORDER)
C1319018|T047|405944004|SNOMEDCT_US|BRONCHITIS;ASTHMATIC|ASTHMATIC BRONCHITIS (DISORDER)
C1319018|T047|405944004|SNOMEDCT_US|BRONCHITIS;WHEEZY|ASTHMATIC BRONCHITIS (DISORDER)
C1319018|T047|405944004|SNOMEDCT_US|ASTHMATIC BRONCHITIS |ASTHMATIC BRONCHITIS (DISORDER)
C1319018|T047|405944004|SNOMEDCT_US|WHEEZY BRONCHITIS|ASTHMATIC BRONCHITIS (DISORDER)
C1319018|T047|405944004|SNOMEDCT_US|BRONCHITIS ASTHMATIC|ASTHMATIC BRONCHITIS (DISORDER)
C1319018|T047|405944004|SNOMEDCT_US|ASTHMATIC BRONCHITIS, NOS|ASTHMATIC BRONCHITIS (DISORDER)
C1319018|T047|405944004|SNOMEDCT_US|BRONCHITIS, ASTHMATIC|ASTHMATIC BRONCHITIS (DISORDER)
C3266628|T047|5281000124103|SNOMEDCT_US|PERSISTENT ASTHMA|PERSISTENT ASTHMA (DISORDER)
C3266628|T047|5281000124103|SNOMEDCT_US|PERSISTENT ASTHMA |PERSISTENT ASTHMA (DISORDER)
C3266628|T047|5281000124103|SNOMEDCT_US|PERSISTENT ASTHMA |PERSISTENT ASTHMA (DISORDER)
C3266628|T047|5281000124103|SNOMEDCT_US|ASTHMA PERSISTENT|PERSISTENT ASTHMA (DISORDER)
C3662842|T047|1761000119103|SNOMEDCT_US|CHRONIC OBSTRUCTIVE AIRWAY DISEASE WITH ASTHMA |CHRONIC OBSTRUCTIVE AIRWAY DISEASE WITH ASTHMA (DISORDER)
C3662842|T047|1761000119103|SNOMEDCT_US|CHRONIC OBSTRUCTIVE AIRWAY DISEASE WITH ASTHMA|CHRONIC OBSTRUCTIVE AIRWAY DISEASE WITH ASTHMA (DISORDER)
C3661951|T047|401000119107|SNOMEDCT_US|ASTHMA WITH IRREVERSIBLE AIRWAY OBSTRUCTION|ASTHMA WITH IRREVERSIBLE AIRWAY OBSTRUCTION (DISORDER)
C3661951|T047|401000119107|SNOMEDCT_US|ASTHMA WITH IRREVERSIBLE AIRWAY OBSTRUCTION |ASTHMA WITH IRREVERSIBLE AIRWAY OBSTRUCTION (DISORDER)
C0582415|T047|304527002|SNOMEDCT_US|ASTHMA ACUTE|ACUTE ASTHMA (DISORDER)
C0582415|T047|304527002|SNOMEDCT_US|ACUTE ASTHMA|ACUTE ASTHMA (DISORDER)
C0582415|T047|304527002|SNOMEDCT_US|ACUTE ASTHMA |ACUTE ASTHMA (DISORDER)
C0582415|T047|304527002|SNOMEDCT_US|ACUTE ASTHMA |ACUTE ASTHMA (DISORDER)
C0582415|T047|304527002|SNOMEDCT_US|ASTHMA; ACUTE|ACUTE ASTHMA (DISORDER)
C0582415|T047|304527002|SNOMEDCT_US|ACUTE; ASTHMA|ACUTE ASTHMA (DISORDER)
C1828277|T047|424199006|SNOMEDCT_US|SUBSTANCE INDUCED ASTHMA|SUBSTANCE INDUCED ASTHMA (DISORDER)
C1828277|T047|424199006|SNOMEDCT_US|SUBSTANCE INDUCED ASTHMA |SUBSTANCE INDUCED ASTHMA (DISORDER)
C1828277|T047|424199006|SNOMEDCT_US|SUBSTANCE-INDUCED ASTHMA|SUBSTANCE INDUCED ASTHMA (DISORDER)
C1828277|T047|424199006|SNOMEDCT_US|ASTHMA SUBSTANCE-INDUCED|SUBSTANCE INDUCED ASTHMA (DISORDER)
C1828277|T047|424199006|SNOMEDCT_US|SUBSTANCE-INDUCED ASTHMA |SUBSTANCE INDUCED ASTHMA (DISORDER)
C0581124|T047|370218001|SNOMEDCT_US|MILD ASTHMA |MILD ASTHMA (DISORDER)
C0581124|T047|370218001|SNOMEDCT_US|MILD ASTHMA |MILD ASTHMA (DISORDER)
C0581124|T047|370218001|SNOMEDCT_US|MILD ASTHMA|MILD ASTHMA (DISORDER)
C0581124|T047|370218001|SNOMEDCT_US|MILD ASTHMA |MILD ASTHMA (DISORDER)
C0581124|T047|370218001|SNOMEDCT_US|ASTHMA MILD|MILD ASTHMA (DISORDER)
C0581124|T047|370218001|SNOMEDCT_US|MILD ASTHMA |MILD ASTHMA (DISORDER)
C0581123|T047|370220003|SNOMEDCT_US|OCCASIONAL ASTHMA |OCCASIONAL ASTHMA (DISORDER)
C0581123|T047|370220003|SNOMEDCT_US|OCCASIONAL ASTHMA |OCCASIONAL ASTHMA (DISORDER)
C0581123|T047|370220003|SNOMEDCT_US|OCCASIONAL ASTHMA|OCCASIONAL ASTHMA (DISORDER)
C0581123|T047|370220003|SNOMEDCT_US|OCCASIONAL ASTHMA |OCCASIONAL ASTHMA (DISORDER)
C0581123|T047|370220003|SNOMEDCT_US|ASTHMA OCCASIONAL|OCCASIONAL ASTHMA (DISORDER)
C0581123|T047|370220003|SNOMEDCT_US|OCCASIONAL ASTHMA |OCCASIONAL ASTHMA (DISORDER)
C0264405|T047|55570000|SNOMEDCT_US|ASTHMA WITHOUT STATUS ASTHMATICUS |ASTHMA WITHOUT STATUS ASTHMATICUS (DISORDER)
C0264405|T047|55570000|SNOMEDCT_US|ASTHMA WITHOUT STATUS ASTHMATICUS|ASTHMA WITHOUT STATUS ASTHMATICUS (DISORDER)
C0264405|T047|55570000|SNOMEDCT_US|ASTHMA WITHOUT STATUS ASTHMATICUS |ASTHMA WITHOUT STATUS ASTHMATICUS (DISORDER)
C0581125|T047|370219009|SNOMEDCT_US|MODERATE ASTHMA |MODERATE ASTHMA (DISORDER)
C0581125|T047|370219009|SNOMEDCT_US|MODERATE ASTHMA |MODERATE ASTHMA (DISORDER)
C0581125|T047|370219009|SNOMEDCT_US|MODERATE ASTHMA|MODERATE ASTHMA (DISORDER)
C0581125|T047|370219009|SNOMEDCT_US|MODERATE ASTHMA |MODERATE ASTHMA (DISORDER)
C0581125|T047|370219009|SNOMEDCT_US|ASTHMA MODERATE|MODERATE ASTHMA (DISORDER)
C0581125|T047|370219009|SNOMEDCT_US|MODERATE ASTHMA |MODERATE ASTHMA (DISORDER)
C0340073|T047|233690008|SNOMEDCT_US|FACTITIOUS ASTHMA|FACTITIOUS ASTHMA (DISORDER)
C0340073|T047|233690008|SNOMEDCT_US|ASTHMA FACTITIOUS|FACTITIOUS ASTHMA (DISORDER)
C0340073|T047|233690008|SNOMEDCT_US|FACTITIOUS ASTHMA |FACTITIOUS ASTHMA (DISORDER)
C0340073|T047|233690008|SNOMEDCT_US|EMOTIONAL LARYNGEAL WHEEZING|FACTITIOUS ASTHMA (DISORDER)
C0340073|T047|233690008|SNOMEDCT_US|FUNCTIONAL LARYNGEAL STRIDOR|FACTITIOUS ASTHMA (DISORDER)
C0340073|T047|233690008|SNOMEDCT_US|FACTITIOUS ASTHMA |FACTITIOUS ASTHMA (DISORDER)
C0581126|T047|370221004|SNOMEDCT_US|SEVERE ASTHMA |SEVERE ASTHMA (DISORDER)
C0581126|T047|370221004|SNOMEDCT_US|SEVERE ASTHMA |SEVERE ASTHMA (DISORDER)
C0581126|T047|370221004|SNOMEDCT_US|SEVERE ASTHMA |SEVERE ASTHMA (DISORDER)
C0581126|T047|370221004|SNOMEDCT_US|SEVERE ASTHMA|SEVERE ASTHMA (DISORDER)
C0581126|T047|370221004|SNOMEDCT_US|ASTHMA SEVERE|SEVERE ASTHMA (DISORDER)
C0581126|T047|370221004|SNOMEDCT_US|SEVERE ASTHMA |SEVERE ASTHMA (DISORDER)
C0581126|T047|370221004|SNOMEDCT_US|ASTHMA; SEVERE|SEVERE ASTHMA (DISORDER)
C0581126|T047|370221004|SNOMEDCT_US|SEVERE; ASTHMA|SEVERE ASTHMA (DISORDER)
C1859647|T047||SNOMEDCT_US|ASTHMA, SHORT STATURE, AND ELEVATED IGA
C1853964|T047||SNOMEDCT_US|DERMATITIS, ATOPIC, WITH ASTHMA
C3280315|T047||SNOMEDCT_US| ASSOCIATED WITH SEVERE ASTHMA
C1858067|T047||SNOMEDCT_US|ASTHMA AND NASAL POLYPS
C1869116|T047||SNOMEDCT_US|ASTHMA, SUSCEPTIBILITY TO
C1869116|T047||SNOMEDCT_US|ASTHMA, SUSCEPTIBILITY TO 
C1869116|T047||SNOMEDCT_US|ASTHMA SUSCEPTIBILITY
C1869116|T047||SNOMEDCT_US|ASTHMA SUSCEPTIBILITY 
C1869116|T047||SNOMEDCT_US|ASTHMA-RELATED TRAITS, SUSCEPTIBILITY TO
C1869116|T047||SNOMEDCT_US|ASTHMA, BRONCHIAL
C3838502|T047||SNOMEDCT_US|ASTHMA PROTECTION 
C3838502|T047||SNOMEDCT_US|ASTHMA PROTECTION
C3838894|T047|10742121000119104|SNOMEDCT_US|ASTHMA IN MOTHER COMPLICATING CHILDBIRTH |ASTHMA IN CHILDBIRTH
C3838894|T047|10742121000119104|SNOMEDCT_US|ASTHMA IN CHILDBIRTH|ASTHMA IN CHILDBIRTH
C3838894|T047|10742121000119104|SNOMEDCT_US|ASTHMA IN MOTHER COMPLICATING CHILDBIRTH|ASTHMA IN CHILDBIRTH
C4038730|T047|10692761000119107|SNOMEDCT_US|ASTHMA-CHRONIC OBSTRUCTIVE PULMONARY DISEASE OVERLAP SYNDROME|ASTHMA-CHRONIC OBSTRUCTIVE PULMONARY DISEASE OVERLAP SYNDROME (DISORDER)
C4038730|T047|10692761000119107|SNOMEDCT_US|ASTHMA-CHRONIC OBSTRUCTIVE PULMONARY DISEASE OVERLAP SYNDROME |ASTHMA-CHRONIC OBSTRUCTIVE PULMONARY DISEASE OVERLAP SYNDROME (DISORDER)
C4038730|T047|10692761000119107|SNOMEDCT_US|ASTHMA-COPD OVERLAP SYNDROME (ACOS)|ASTHMA-CHRONIC OBSTRUCTIVE PULMONARY DISEASE OVERLAP SYNDROME (DISORDER)
C4038730|T047|10692761000119107|SNOMEDCT_US|ASTHMA-COPD OVERLAP SYNDROME|ASTHMA-CHRONIC OBSTRUCTIVE PULMONARY DISEASE OVERLAP SYNDROME (DISORDER)
C0741267|T047|2360001000004109|SNOMEDCT_US|STEROID DEPENDENT ASTHMA|STEROID DEPENDENT ASTHMA (DISORDER)
C0741267|T047|2360001000004109|SNOMEDCT_US|STEROID DEPENDENT ASTHMA |STEROID DEPENDENT ASTHMA (DISORDER)
C1388871|T047||SNOMEDCT_US|ASTHMA; CROUP
C1388871|T047||SNOMEDCT_US|CROUP; ASTHMA
C1388880|T047||SNOMEDCT_US|ASTHMATIC; DYSPNEA
C1388880|T047||SNOMEDCT_US|DYSPNEA; ASTHMATIC
C1388882|T047||SNOMEDCT_US|ASTHMATIC; DYSPNEA, WITH BRONCHITIS
C1388882|T047||SNOMEDCT_US|DYSPNEA; ASTHMATIC, WITH BRONCHITIS
C1403212|T047||SNOMEDCT_US|OBSTRUCTION; AIRWAY, WITH ASTHMA
C1403212|T047||SNOMEDCT_US|AIRWAY; OBSTRUCTION, WITH ASTHMA
C1260416|T047||SNOMEDCT_US|OTHER FORMS OF ASTHMA
C1176342|T047||SNOMEDCT_US|ASTHMA NOS W (AC) EXAC
C1176342|T047||SNOMEDCT_US|ASTHMA, UNSPECIFIED TYPE, WITH (ACUTE) EXACERBATION
