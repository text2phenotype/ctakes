// CUI|TUI|CODE|VOCAB|TXT|PREF TEXT
C000001|T109|1|DICT1|Drug|Drug annotation from dict 1
C000003|T109|3|DICT1|Proc|Procedure as a Drug from dict 1