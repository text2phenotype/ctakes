// CUI|TUI|CODE|VOCAB|TXT|PREF TEXT
C000001|T109|1|CUSTOM|aspirin|aspirin
C000002|T019|2|CUSTOM|oppenheims disease|Oppenheim's Disease
C000003|T033|3|CUSTOM|anisocorias|Anisocoria
C000004|T060|4|CUSTOM|aortography|Aortography
C000005|T021|5|CUSTOM|total body|Entire body as a whole
C000006|T034|6|CUSTOM|hemoglobin|Hemoglobin
C000007|T058|7|CUSTOM|ambulatory care|Ambulatory Care