C0085178|T037|283596007|SNOMEDCT_US|NEEDLESTICK INJURIES|NEEDLE STICK INJURY (DISORDER)
C0582072|T037|304235000|SNOMEDCT_US|SHARPS INJURIES|SHARPS INJURY (DISORDER)
C0561474|T037|283604006|SNOMEDCT_US|NEEDLE STICK INJURY OF NOSE|NEEDLE STICK INJURY OF NOSE (DISORDER)
C0561474|T037|283604006|SNOMEDCT_US|NEEDLE STICK INJURY OF NOSE |NEEDLE STICK INJURY OF NOSE (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|INJURIES, NEEDLE-STICK|NEEDLE STICK INJURY (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|INJURY, NEEDLE-STICK|NEEDLE STICK INJURY (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|INJURY, NEEDLESTICK|NEEDLE STICK INJURY (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|NEEDLE STICK INJURIES|NEEDLE STICK INJURY (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|NEEDLE STICKS|NEEDLE STICK INJURY (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|NEEDLE-STICK|NEEDLE STICK INJURY (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|NEEDLE-STICK INJURY|NEEDLE STICK INJURY (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|NEEDLESTICK|NEEDLE STICK INJURY (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|NEEDLESTICK INJURIES|NEEDLE STICK INJURY (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|NEEDLESTICK INJURY|NEEDLE STICK INJURY (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|NEEDLESTICK INJ|NEEDLE STICK INJURY (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|INJ NEEDLESTICK|NEEDLE STICK INJURY (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|NEEDLESTICKS|NEEDLE STICK INJURY (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|NEEDLE-STICK INJURIES|NEEDLE STICK INJURY (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|NEEDLE-STICKS|NEEDLE STICK INJURY (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|INJURIES, NEEDLESTICK|NEEDLE STICK INJURY (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|NEEDLESTICK INJURIES [DISEASE/FINDING]|NEEDLE STICK INJURY (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|INJURY;NEEDLE STICK|NEEDLE STICK INJURY (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|NEEDLE STICK|NEEDLE STICK INJURY (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|NEEDLE PRICK INJURY|NEEDLE STICK INJURY (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|NEEDLE STICK INJURY|NEEDLE STICK INJURY (DISORDER)
C0085178|T037|283596007|SNOMEDCT_US|NEEDLE STICK INJURY |NEEDLE STICK INJURY (DISORDER)
C2116782|T037||SNOMEDCT_US|PUNCTURE BY NEEDLE
C2116782|T037||SNOMEDCT_US|PUNCTURE BY NEEDLE (PHYSICAL FINDING)
C0582071|T037|304234001|SNOMEDCT_US|NEEDLE STICK INJURY WITH CONTAMINATED NEEDLE|NEEDLE STICK INJURY WITH CONTAMINATED NEEDLE (DISORDER)
C0582071|T037|304234001|SNOMEDCT_US|NEEDLE STICK INJURY WITH DIRTY NEEDLE|NEEDLE STICK INJURY WITH CONTAMINATED NEEDLE (DISORDER)
C0582071|T037|304234001|SNOMEDCT_US|NEEDLE STICK INJURY WITH CONTAMINATED NEEDLE |NEEDLE STICK INJURY WITH CONTAMINATED NEEDLE (DISORDER)
C0561467|T037|283597003|SNOMEDCT_US|NEEDLE STICK INJURY OF HEAD AND NECK|NEEDLE STICK INJURY OF HEAD AND NECK (DISORDER)
C0561467|T037|283597003|SNOMEDCT_US|NEEDLE STICK INJURY OF HEAD AND NECK |NEEDLE STICK INJURY OF HEAD AND NECK (DISORDER)
C0561500|T037|283630005|SNOMEDCT_US|NEEDLE STICK INJURY OF LOWER LIMB|NEEDLE STICK INJURY OF LOWER LIMB (DISORDER)
C0561500|T037|283630005|SNOMEDCT_US|NEEDLE STICK INJURY OF LOWER LIMB |NEEDLE STICK INJURY OF LOWER LIMB (DISORDER)
C0561479|T037|283609001|SNOMEDCT_US|NEEDLE STICK INJURY OF UPPER LIMB|NEEDLE STICK INJURY OF UPPER LIMB (DISORDER)
C0561479|T037|283609001|SNOMEDCT_US|NEEDLE STICK INJURY OF UPPER LIMB |NEEDLE STICK INJURY OF UPPER LIMB (DISORDER)
C0561491|T037|283621002|SNOMEDCT_US|NEEDLE STICK INJURY OF TRUNK|NEEDLE STICK INJURY OF TRUNK (DISORDER)
C0561491|T037|283621002|SNOMEDCT_US|NEEDLE STICK INJURY OF TRUNK |NEEDLE STICK INJURY OF TRUNK (DISORDER)
C0582072|T037|304235000|SNOMEDCT_US|SHARPS INJURY|SHARPS INJURY (DISORDER)
C0582072|T037|304235000|SNOMEDCT_US|SHARPS INJURY |SHARPS INJURY (DISORDER)
C0582072|T037|304235000|SNOMEDCT_US|INJURIES, SHARPS|SHARPS INJURY (DISORDER)
C0582072|T037|304235000|SNOMEDCT_US|INJURY, SHARPS|SHARPS INJURY (DISORDER)
C0582072|T037|304235000|SNOMEDCT_US|SHARPS INJURIES|SHARPS INJURY (DISORDER)
