C2062763|T053||SNOMEDCT_US|BENZODIAZEPINE ABUSE
C0418282|T053|242832005|SNOMEDCT_US|INTENTIONAL BENZODIAZEPINE OVERDOSE|INTENTIONAL BENZODIAZEPINE OVERDOSE (DISORDER)
C0747951|T053||SNOMEDCT_US|PRESCRIPTION DRUG ABUSE BENZODIAZEPINE
C0747952|T053||SNOMEDCT_US|PRESCRIPTION DRUG ABUSE BENZODIAZEPINE DEPENDENCE
C0747953|T053||SNOMEDCT_US|PRESCRIPTION DRUG ABUSE BENZODIAZEPINE POTENTIAL
C0747954|T053||SNOMEDCT_US|PRESCRIPTION DRUG ABUSE BENZODIAZEPINE REMISSION
C0747955|T053||SNOMEDCT_US|PRESCRIPTION DRUG ABUSE BENZODIAZEPINE WITHDRAWAL
C2104566|T053||SNOMEDCT_US|CONTINUOUS BENZODIAZEPINE ABUSE 
C2104566|T053||SNOMEDCT_US|CONTINUOUS BENZODIAZEPINE ABUSE
C2104567|T053||SNOMEDCT_US|EPISODIC BENZODIAZEPINE ABUSE 
C2104567|T053||SNOMEDCT_US|EPISODIC BENZODIAZEPINE ABUSE
C2104568|T053||SNOMEDCT_US|BENZODIAZEPINE ABUSE IN REMISSION 
C2104568|T053||SNOMEDCT_US|BENZODIAZEPINE ABUSE IN REMISSION
C0572936|T053|296056007|SNOMEDCT_US|INTENTIONAL FLUNITRAZEPAM OVERDOSE|INTENTIONAL FLUNITRAZEPAM OVERDOSE (DISORDER)
C0572936|T053|296056007|SNOMEDCT_US|INTENTIONAL FLUNITRAZEPAM OVERDOSE |INTENTIONAL FLUNITRAZEPAM OVERDOSE (DISORDER)
C0572989|T053|296112009|SNOMEDCT_US|INTENTIONAL PRAZEPAM OVERDOSE|INTENTIONAL PRAZEPAM OVERDOSE (DISORDER)
C0572989|T053|296112009|SNOMEDCT_US|INTENTIONAL PRAZEPAM OVERDOSE |INTENTIONAL PRAZEPAM OVERDOSE (DISORDER)
C0572977|T053|296100005|SNOMEDCT_US|INTENTIONAL KETAZOLAM OVERDOSE|INTENTIONAL KETAZOLAM OVERDOSE (DISORDER)
C0572977|T053|296100005|SNOMEDCT_US|INTENTIONAL KETAZOLAM OVERDOSE |INTENTIONAL KETAZOLAM OVERDOSE (DISORDER)
C0572950|T053|296072004|SNOMEDCT_US|INTENTIONAL NITRAZEPAM OVERDOSE|INTENTIONAL NITRAZEPAM OVERDOSE (DISORDER)
C0572950|T053|296072004|SNOMEDCT_US|INTENTIONAL NITRAZEPAM OVERDOSE |INTENTIONAL NITRAZEPAM OVERDOSE (DISORDER)
C0572969|T053|296092006|SNOMEDCT_US|INTENTIONAL CLOBAZAM OVERDOSE|INTENTIONAL CLOBAZAM OVERDOSE (DISORDER)
C0572969|T053|296092006|SNOMEDCT_US|INTENTIONAL CLOBAZAM OVERDOSE |INTENTIONAL CLOBAZAM OVERDOSE (DISORDER)
C0572962|T053|296085001|SNOMEDCT_US|INTENTIONAL BROMAZEPAM OVERDOSE|INTENTIONAL BROMAZEPAM OVERDOSE (DISORDER)
C0572962|T053|296085001|SNOMEDCT_US|INTENTIONAL BROMAZEPAM OVERDOSE |INTENTIONAL BROMAZEPAM OVERDOSE (DISORDER)
C0572939|T053|296060005|SNOMEDCT_US|INTENTIONAL FLURAZEPAM OVERDOSE|INTENTIONAL FLURAZEPAM OVERDOSE (DISORDER)
C0572939|T053|296060005|SNOMEDCT_US|INTENTIONAL FLURAZEPAM OVERDOSE |INTENTIONAL FLURAZEPAM OVERDOSE (DISORDER)
C0572947|T053|296068003|SNOMEDCT_US|INTENTIONAL LORMETAZEPAM OVERDOSE|INTENTIONAL LORMETAZEPAM OVERDOSE (DISORDER)
C0572947|T053|296068003|SNOMEDCT_US|INTENTIONAL LORMETAZEPAM OVERDOSE |INTENTIONAL LORMETAZEPAM OVERDOSE (DISORDER)
C0572943|T053|296064001|SNOMEDCT_US|INTENTIONAL LOPRAZOLAM OVERDOSE|INTENTIONAL LOPRAZOLAM OVERDOSE (DISORDER)
C0572943|T053|296064001|SNOMEDCT_US|INTENTIONAL LOPRAZOLAM OVERDOSE |INTENTIONAL LOPRAZOLAM OVERDOSE (DISORDER)
C0572981|T053|296104001|SNOMEDCT_US|INTENTIONAL MEDAZEPAM OVERDOSE|INTENTIONAL MEDAZEPAM OVERDOSE (DISORDER)
C0572981|T053|296104001|SNOMEDCT_US|INTENTIONAL MEDAZEPAM OVERDOSE |INTENTIONAL MEDAZEPAM OVERDOSE (DISORDER)
C0418284|T053|242834006|SNOMEDCT_US|INTENTIONAL CHLORDIAZEPOXIDE OVERDOSE |INTENTIONAL CHLORDIAZEPOXIDE OVERDOSE (DISORDER)
C0418284|T053|242834006|SNOMEDCT_US|DELIBERATE OVERDOSE OF CHLORDIAZEPOXIDE|INTENTIONAL CHLORDIAZEPOXIDE OVERDOSE (DISORDER)
C0418284|T053|242834006|SNOMEDCT_US|INTENTIONAL CHLORDIAZEPOXIDE OVERDOSE|INTENTIONAL CHLORDIAZEPOXIDE OVERDOSE (DISORDER)
C0418284|T053|242834006|SNOMEDCT_US|DELIBERATE OVERDOSE OF CHLORDIAZEPOXIDE |INTENTIONAL CHLORDIAZEPOXIDE OVERDOSE (DISORDER)
C0572993|T053|296116007|SNOMEDCT_US|INTENTIONAL MIDAZOLAM OVERDOSE|INTENTIONAL MIDAZOLAM OVERDOSE (DISORDER)
C0572993|T053|296116007|SNOMEDCT_US|INTENTIONAL MIDAZOLAM OVERDOSE |INTENTIONAL MIDAZOLAM OVERDOSE (DISORDER)
C0418283|T053|242833000|SNOMEDCT_US|SELF-INFLICTED OVERDOSE OF DIAZEPAM|INTENTIONAL DIAZEPAM OVERDOSE (DISORDER)
C0418283|T053|242833000|SNOMEDCT_US|SELF-INFLICTED OVERDOSE OF DIAZEPAM |INTENTIONAL DIAZEPAM OVERDOSE (DISORDER)
C0418283|T053|242833000|SNOMEDCT_US|TOXICITY FROM DIAZEPAM DUE TO A SELF-INFLICTED OVERDOSE|INTENTIONAL DIAZEPAM OVERDOSE (DISORDER)
C0418283|T053|242833000|SNOMEDCT_US|INTENTIONAL DIAZEPAM OVERDOSE|INTENTIONAL DIAZEPAM OVERDOSE (DISORDER)
C0418283|T053|242833000|SNOMEDCT_US|DELIBERATE OVERDOSE OF DIAZEPAM |INTENTIONAL DIAZEPAM OVERDOSE (DISORDER)
C0418283|T053|242833000|SNOMEDCT_US|DELIBERATE OVERDOSE OF DIAZEPAM|INTENTIONAL DIAZEPAM OVERDOSE (DISORDER)
C0418283|T053|242833000|SNOMEDCT_US|INTENTIONAL DIAZEPAM OVERDOSE |INTENTIONAL DIAZEPAM OVERDOSE (DISORDER)
C0418285|T053|242835007|SNOMEDCT_US|DELIBERATE OVERDOSE OF TEMAZEPAM |INTENTIONAL TEMAZEPAM OVERDOSE (DISORDER)
C0418285|T053|242835007|SNOMEDCT_US|INTENTIONAL TEMAZEPAM OVERDOSE |INTENTIONAL TEMAZEPAM OVERDOSE (DISORDER)
C0418285|T053|242835007|SNOMEDCT_US|INTENTIONAL TEMAZEPAM OVERDOSE|INTENTIONAL TEMAZEPAM OVERDOSE (DISORDER)
C0418285|T053|242835007|SNOMEDCT_US|DELIBERATE OVERDOSE OF TEMAZEPAM|INTENTIONAL TEMAZEPAM OVERDOSE (DISORDER)
C0572954|T053|296076001|SNOMEDCT_US|INTENTIONAL TRIAZOLAM OVERDOSE|INTENTIONAL TRIAZOLAM OVERDOSE (DISORDER)
C0572954|T053|296076001|SNOMEDCT_US|INTENTIONAL TRIAZOLAM OVERDOSE |INTENTIONAL TRIAZOLAM OVERDOSE (DISORDER)
C0572958|T053|296081005|SNOMEDCT_US|INTENTIONAL ALPRAZOLAM OVERDOSE|INTENTIONAL ALPRAZOLAM OVERDOSE (DISORDER)
C0572958|T053|296081005|SNOMEDCT_US|INTENTIONAL ALPRAZOLAM OVERDOSE |INTENTIONAL ALPRAZOLAM OVERDOSE (DISORDER)
C0572973|T053|296096009|SNOMEDCT_US|INTENTIONAL POTASSIUM CLORAZEPATE OVERDOSE|INTENTIONAL DIPOTASSIUM CLORAZEPATE OVERDOSE
C0572973|T053|296096009|SNOMEDCT_US|INTENTIONAL POTASSIUM CLORAZEPATE OVERDOSE |INTENTIONAL DIPOTASSIUM CLORAZEPATE OVERDOSE
C0572973|T053|296096009|SNOMEDCT_US|INTENTIONAL DIPOTASSIUM CLORAZEPATE OVERDOSE|INTENTIONAL DIPOTASSIUM CLORAZEPATE OVERDOSE
C0572985|T053|296108003|SNOMEDCT_US|INTENTIONAL OXAZEPAM OVERDOSE|INTENTIONAL OXAZEPAM OVERDOSE (DISORDER)
C0572985|T053|296108003|SNOMEDCT_US|INTENTIONAL OXAZEPAM OVERDOSE |INTENTIONAL OXAZEPAM OVERDOSE (DISORDER)
C0573000|T053|296123008|SNOMEDCT_US|INTENTIONAL LORAZEPAM OVERDOSE|INTENTIONAL LORAZEPAM OVERDOSE (DISORDER)
C0573000|T053|296123008|SNOMEDCT_US|INTENTIONAL LORAZEPAM OVERDOSE |INTENTIONAL LORAZEPAM OVERDOSE (DISORDER)
C0572892|T053|296012007|SNOMEDCT_US|INTENTIONAL CLONAZEPAM OVERDOSE|INTENTIONAL CLONAZEPAM OVERDOSE (DISORDER)
C0572892|T053|296012007|SNOMEDCT_US|INTENTIONAL CLONAZEPAM OVERDOSE |INTENTIONAL CLONAZEPAM OVERDOSE (DISORDER)
