C0005437|T034|LP15448-1|LNC|BILIRUBIN|BILIRUBIN
C0201913|T034||LNC|BILIRUBIN, TOTAL MEASUREMENT
C0863174|T034||LNC|BLOOD BILIRUBIN MEASUREMENT
C0005437|T034|LP15448-1|LNC|BILIRUBIN, TOTAL|BILIRUBIN
C0005437|T034|LP15448-1|LNC|BILIRUBIN|BILIRUBIN
C0005437|T034|LP15448-1|LNC|BILIRUBIN [CHEMICAL/INGREDIENT]|BILIRUBIN
C0005437|T034|LP15448-1|LNC|CONJUGATED AND UNCONJUGATED BILIRUBIN|BILIRUBIN
C0005437|T034|LP15448-1|LNC|BILIRUBIN |BILIRUBIN
C0005437|T034|LP15448-1|LNC|BILIRUBIN, NOS|BILIRUBIN
C0005437|T034|LP15448-1|LNC|TOTAL BILIRUBIN|BILIRUBIN
C2924724|T034|LP100772-5|LNC|BILIRUBIN &#X7C; BLOOD ARTERIAL|BILIRUBIN &#X7C; BLOOD ARTERIAL
C1982578|T034|LP43561-7|LNC|BILIRUBIN &#X7C; BLD-SER-PLAS|BILIRUBIN &#X7C; BLD-SER-PLAS
C2924726|T034|LP100773-3|LNC|BILIRUBIN &#X7C; BLOOD VENOUS|BILIRUBIN &#X7C; BLOOD VENOUS
C2356967|T034|LP69695-2|LNC|BILIRUBIN.GLUCURONIDATED+BILIRUBIN.NON-GLUCURONIDATED &#X7C; BLD-SER-PLAS|BILIRUBIN.GLUCURONIDATED+BILIRUBIN.NON-GLUCURONIDATED &#X7C; BLD-SER-PLAS
C1291178|T034||LNC|BILIRUBIN COMPOUND 
C1291178|T034||LNC|BILIRUBIN COMPOUND
C1278039|T034||LNC|SERUM TOTAL BILIRUBIN
C1278039|T034||LNC|SERUM TOTAL BILIRUBIN MEASUREMENT
C1278039|T034||LNC|TOTAL SERUM BILIRUBIN LEVEL
C1278039|T034||LNC|SERUM TOTAL BILIRUBIN MEASUREMENT 
C1278039|T034||LNC|SERUM TOTAL BILIRUBIN LEVEL
C1278039|T034||LNC|SERUM TOTAL BILIRUBIN LEVEL 
C1278039|T034||LNC|SERUM BILIRUBIN TOTAL
C1278039|T034||LNC|SERUM TOTAL BILIRUBIN MEASUREMENT 
C0201913|T034||LNC|BILIRUBIN; TOTAL
C0201913|T034||LNC|TOTAL BILIRUBIN MEASUREMENT
C0201913|T034||LNC|BILIRUBIN TOTAL
C0201913|T034||LNC|MEASUREMENT OF TOTAL BILIRUBIN
C0201913|T034||LNC|TOTAL BILIRUBIN
C0201913|T034||LNC|TOTAL BILIRUBIN (& LEVEL) 
C0201913|T034||LNC|BILIRUBIN, TOTAL MEASUREMENT
C0201913|T034||LNC|BILIRUBIN, TOTAL MEASUREMENT 
C0201913|T034||LNC|TOTAL BILIRUBIN (& LEVEL)
C0201913|T034||LNC|BILIRUBIN
C0201913|T034||LNC|BILI
C0201913|T034||LNC|TOTAL BILIRUBIN LEVEL
C0201913|T034||LNC|BILIRUBIN, TOTAL MEASUREMENT  [AMBIGUOUS]
C0373554|T034||LNC|BILIRUBIN; FECES, QUALITATIVE
C0373554|T034||LNC|BILIRUBIN FECES QUALITATIVE
C0373554|T034||LNC|FECAL BILIRUBIN TEST
C0697273|T034||LNC|BILIRUBIN; DIRECT
C0697273|T034||LNC|BILIRUBIN CONJUGATED
C0697273|T034||LNC|BILIRUBIN DIRECT
C0697273|T034||LNC|CONJUGATED BILIRUBIN TEST
C1278036|T034||LNC|PLASMA TOTAL BILIRUBIN LEVEL 
C1278036|T034||LNC|PLASMA TOTAL BILIRUBIN LEVEL
C1278036|T034||LNC|PLASMA BILIRUBIN TOTAL
C1278036|T034||LNC|PLASMA TOTAL BILIRUBIN TEST
C1278036|T034||LNC|PLASMA TOTAL BILIRUBIN MEASUREMENT 
C1278036|T034||LNC|PLASMA TOTAL BILIRUBIN MEASUREMENT
C0428441|T034||LNC|BILIRUBIN
C0428441|T034||LNC|SERUM BILIRUBIN MEASUREMENT 
C0428441|T034||LNC|SERUM BILIRUBIN (& LEVEL) 
C0428441|T034||LNC|BILIRUBIN - SERUM
C0428441|T034||LNC|SERUM BILIRUBIN NOS 
C0428441|T034||LNC|SERUM BILIRUBIN NOS
C0428441|T034||LNC|SERUM BILIRUBIN LEVEL
C0428441|T034||LNC|SERUM BILIRUBIN (& LEVEL)
C0428441|T034||LNC|SERUM BILIRUBIN
C0428441|T034||LNC|SB - SERUM BILIRUBIN
C0428441|T034||LNC|SERUM BILIRUBIN MEASUREMENT 
C0428441|T034||LNC|SERUM BILIRUBIN MEASUREMENT
C0863174|T034||LNC|BLOOD BILIRUBIN
C0863174|T034||LNC|BLOOD BILIRUBIN MEASUREMENT
C0863174|T034||LNC|BILIRUBIN
C0863174|T034||LNC|T. BILI
C0863174|T034||LNC|T BILI
