// CUI|TUI|TTY|CODE|SAB|STR|PREF
C0004096|T047|BN|195979001|SNOMEDCT_US|ASTHMA|ASTHMA UNSPECIFIED (DISORDER)