C3160090|T121||RXNORM|HCV NS3/4A PROTEASE INHIBITORS [MOA]
C1738934|T121|1102129|RXNORM|BOCEPREVIR|BOCEPREVIR
C1876229|T121|1102261|RXNORM|TELAPREVIR|TELAPREVIR
C2605855|T121|1482790|RXNORM|SIMEPREVIR|SIMEPREVIR
C3154649|T121|1102132|RXNORM|BOCEPREVIR 200 MG ORAL CAPSULE|BOCEPREVIR 200 MG ORAL CAPSULE
C3154711|T121|1102280|RXNORM|TELAPREVIR 375 MG ORAL TABLET|TELAPREVIR 375 MG ORAL TABLET
C0697341|T121|856450|RXNORM|INDERAL 10 MG ORAL TABLET|INDERAL 10 MG ORAL TABLET
C0591636|T121|151890|RXNORM|INDERAL|INDERAL
C3226084|T121|1172017|RXNORM|INDERAL PILL|INDERAL PILL
C3226083|T121|1172016|RXNORM|INDERAL ORAL PRODUCT|INDERAL ORAL PRODUCT
C2710361|T121|856461|RXNORM|PROPRANOLOL HYDROCHLORIDE 120 MG [INDERAL]|PROPRANOLOL HYDROCHLORIDE 120 MG [INDERAL]
C2710374|T121|856482|RXNORM|PROPRANOLOL HYDROCHLORIDE 160 MG [INDERAL]|PROPRANOLOL HYDROCHLORIDE 160 MG [INDERAL]
C2710406|T121|856536|RXNORM|PROPRANOLOL HYDROCHLORIDE 60 MG [INDERAL]|PROPRANOLOL HYDROCHLORIDE 60 MG [INDERAL]
C2710422|T121|856570|RXNORM|PROPRANOLOL HYDROCHLORIDE 80 MG [INDERAL]|PROPRANOLOL HYDROCHLORIDE 80 MG [INDERAL]
C1577533|T121|491323|RXNORM|PROPRANOLOL EXTENDED RELEASE ORAL CAPSULE [INDERAL]|PROPRANOLOL EXTENDED RELEASE ORAL CAPSULE [INDERAL]
C0697868|T121|856483|RXNORM|24 HR PROPRANOLOL HYDROCHLORIDE 160 MG EXTENDED RELEASE ORAL CAPSULE [INDERAL]|24 HR INDERAL LA 160 MG EXTENDED RELEASE ORAL CAPSULE
C0697871|T121|856571|RXNORM|24 HR PROPRANOLOL HYDROCHLORIDE 80 MG EXTENDED RELEASE ORAL CAPSULE [INDERAL]|INDERAL XL 80 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C0709220|T121|856537|RXNORM|24 HR PROPRANOLOL HYDROCHLORIDE 60 MG EXTENDED RELEASE ORAL CAPSULE [INDERAL]|INDERAL LA 60 MG 24HR EXTENDED RELEASE ORAL CAPSULE
C0709222|T121|856462|RXNORM|24 HR PROPRANOLOL HYDROCHLORIDE 120 MG EXTENDED RELEASE ORAL CAPSULE [INDERAL]|INDERAL XL 120 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C0022957|T121|6218|RXNORM|LACTULOSE|LACTULOSE
C0994966|T121|756967|RXNORM|LACTULOSE ORAL SOLUTION [ENULOSE]|LACTULOSE ORAL SOLUTION [ENULOSE]
C1134051|T121|336731|RXNORM|LACTULOSE 667 MG/ML|LACTULOSE 667 MG/ML
C1178770|T121|360554|RXNORM|LACTULOSE 670 MG/ML|LACTULOSE 670 MG/ML
C1252332|T121|378092|RXNORM|LACTULOSE ORAL SOLUTION|LACTULOSE ORAL SOLUTION
C1589308|T121|544451|RXNORM|LACTULOSE ORAL SOLUTION [CONSTULOSE]|LACTULOSE ORAL SOLUTION [CONSTULOSE]
C1589310|T121|544454|RXNORM|LACTULOSE ORAL SOLUTION [GENERLAC]|LACTULOSE ORAL SOLUTION [GENERLAC]
C3216530|T121|1162200|RXNORM|LACTULOSE ORAL LIQUID PRODUCT|LACTULOSE ORAL LIQUID PRODUCT
C3216531|T121|1162201|RXNORM|LACTULOSE ORAL PRODUCT|LACTULOSE ORAL PRODUCT
C4306942|T121|1868578|RXNORM|LACTULOSE 10000 MG [KRISTALOSE]|LACTULOSE 10000 MG [KRISTALOSE]
C4306943|T121|1868572|RXNORM|LACTULOSE 20000 MG [KRISTALOSE]|LACTULOSE 20000 MG [KRISTALOSE]
C4307200|T121|1868576|RXNORM|LACTULOSE 10000 MG|LACTULOSE 10000 MG
C4307201|T121|1868568|RXNORM|LACTULOSE 20000 MG|LACTULOSE 20000 MG
C4307247|T121|1868570|RXNORM|LACTULOSE POWDER FOR ORAL SOLUTION|LACTULOSE POWDER FOR ORAL SOLUTION
C4307286|T121|1868569|RXNORM|LACTULOSE ORAL POWDER PRODUCT|LACTULOSE ORAL POWDER PRODUCT
C1589307|T121|544450|RXNORM|LACTULOSE 667 MG/ML [CONSTULOSE]|LACTULOSE 667 MG/ML [CONSTULOSE]
C1589309|T121|544453|RXNORM|LACTULOSE 667 MG/ML [GENERLAC]|LACTULOSE 667 MG/ML [GENERLAC]
C1600254|T121|567837|RXNORM|LACTULOSE 667 MG/ML [ENULOSE]|LACTULOSE 667 MG/ML [ENULOSE]
C4307030|T121|1868573|RXNORM|LACTULOSE POWDER FOR ORAL SOLUTION [KRISTALOSE]|LACTULOSE POWDER FOR ORAL SOLUTION [KRISTALOSE]
C0353982|T121|104148|RXNORM|LACTULOSE 670 MG/ML ORAL SOLUTION|LACTULOSE 3.35 GM PER 5 ML ORAL SOLUTION
C0708296|T121|755470|RXNORM|LACTULOSE 667 MG/ML ORAL SOLUTION [ENULOSE]|ENULOSE 10 GM PER 15 ML SYRUP
C0978083|T121|1251190|RXNORM|LACTULOSE 10000 MG POWDER FOR ORAL SOLUTION|LACTULOSE 10 GM GRANULES FOR ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 667 MG/ML ORAL SOLUTION|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1586235|T121|544452|RXNORM|LACTULOSE 667 MG/ML ORAL SOLUTION [CONSTULOSE]|CONSTULOSE 10 GM PER 15 ML SYRUP
C1586236|T121|544455|RXNORM|LACTULOSE 667 MG/ML ORAL SOLUTION [GENERLAC]|GENERLAC 667 MG/ML ORAL SOLUTION
C1613498|T121|1251196|RXNORM|LACTULOSE 20000 MG POWDER FOR ORAL SOLUTION [KRISTALOSE]|KRISTALOSE 20 GM POWDER FOR ORAL SOLUTION
C1620382|T121|1251192|RXNORM|LACTULOSE 10000 MG POWDER FOR ORAL SOLUTION [KRISTALOSE]|KRISTALOSE 10000 MG POWDER FOR ORAL SOLUTION
C1737835|T121|1251194|RXNORM|LACTULOSE 20000 MG POWDER FOR ORAL SOLUTION|LACTULOSE 20 GM GRANULES FOR ORAL SOLUTION
C0043031|T121|11289|RXNORM|WARFARIN|WARFARIN
C3154650|T121|1102133|RXNORM|VICTRELIS|VICTRELIS
C3154650|T121|1102133|RXNORM|VICRTELIS|VICTRELIS
C1738934|T121|1102129|RXNORM|N-(3-AMINO-1-(CYCLOBUTYLMETHYL)-2,3-DIOXOPROPYL)-3-(2-((((1,1-DIMETHYLETHYL)AMINO)CARBONYL)AMINO)-3,3-DIMETHYL-1-OXOBUTYL)-6,6-DIMETHYL-3-AZABICYCLO(3.1.0)HEXAN-2-CARBOXAMIDE|BOCEPREVIR
C1738934|T121|1102129|RXNORM|BOCEPREVIR|BOCEPREVIR
C1738934|T121|1102129|RXNORM|ANTIVIRALS BOCEPREVIR|BOCEPREVIR
C1738934|T121|1102129|RXNORM|ANTIVIRALS BOCEPREVIR |BOCEPREVIR
C1738934|T121|1102129|RXNORM|BOCEPREVIR |BOCEPREVIR
C1738934|T121|1102129|RXNORM|BOCEPREVIR |BOCEPREVIR
C1738934|T121|1102129|RXNORM|3-AZABICYCLO(3.1.0)HEXANE-2-CARBOXAMIDE, N-(3-AMINO-1-(CYCLOBUTYLMETHYL)-2,3-DIOXOPROPYL)-3-((2S)-2-((((1,1- DIMETHYLETHYL)AMINO)CARBONYL)AMINO)-3,3-DIMETHYL-1-OXOBUTYL)-6,6- DIMETHYL-, (1R,2S,5S)-|BOCEPREVIR
C3154649|T121|1102132|RXNORM|BOCEPREVIR CAP 200 MG|BOCEPREVIR 200 MG ORAL CAPSULE
C3154649|T121|1102132|RXNORM|BOCEPREVIR 200MG CAP|BOCEPREVIR 200 MG ORAL CAPSULE
C3154649|T121|1102132|RXNORM|BOCEPREVIR 200 MG ORAL CAPSULE|BOCEPREVIR 200 MG ORAL CAPSULE
C3154649|T121|1102132|RXNORM|BOCEPREVIR 200MG CAP [VA PRODUCT]|BOCEPREVIR 200 MG ORAL CAPSULE
C3154649|T121|1102132|RXNORM|BOCEPREVIR 200MG ORAL CAPSULE|BOCEPREVIR 200 MG ORAL CAPSULE
C3154649|T121|1102132|RXNORM|BOCEPREVIR 200MG CAPSULE |BOCEPREVIR 200 MG ORAL CAPSULE
C3154649|T121|1102132|RXNORM|BOCEPREVIR 200MG CAPSULE|BOCEPREVIR 200 MG ORAL CAPSULE
C1741239|T121||RXNORM|SCH-503034
C1741239|T121||RXNORM|SCH 503034
C1741239|T121||RXNORM|SCH503034
C3896865|T121||RXNORM|EBP 520
C3154701|T121|1102265|RXNORM|INCIVEK|INCIVEK
C1876229|T121|1102261|RXNORM|TELAPREVIR|TELAPREVIR
C1876229|T121|1102261|RXNORM|ANTIVIRAL TELAPREVIR|TELAPREVIR
C1876229|T121|1102261|RXNORM|ANTIVIRAL TELAPREVIR |TELAPREVIR
C1876229|T121|1102261|RXNORM|TELAPREVIR |TELAPREVIR
C1876229|T121|1102261|RXNORM|TELAPREVIR |TELAPREVIR
C3281323|T121||RXNORM|VRT-111950
C3281324|T121||RXNORM|MP-424
C3281325|T121||RXNORM|LY-570310
C1956374|T121||RXNORM|VX-950
C1956374|T121||RXNORM|VX 950
C1956374|T121||RXNORM|VX950 CPD
C3154711|T121|1102280|RXNORM|TELAPREVIR 375 MG ORAL TABLET|TELAPREVIR 375 MG ORAL TABLET
C3154711|T121|1102280|RXNORM|TELAPREVIR TAB 375 MG|TELAPREVIR 375 MG ORAL TABLET
C3154711|T121|1102280|RXNORM|TELAPREVIR 375MG TAB|TELAPREVIR 375 MG ORAL TABLET
C3154711|T121|1102280|RXNORM|TELAPREVIR 375MG TAB,28 [VA PRODUCT]|TELAPREVIR 375 MG ORAL TABLET
C3154711|T121|1102280|RXNORM|TELAPREVIR 375MG TAB,28|TELAPREVIR 375 MG ORAL TABLET
C3154711|T121|1102280|RXNORM|TELAPREVIR 375MG TAB [VA PRODUCT]|TELAPREVIR 375 MG ORAL TABLET
C3154711|T121|1102280|RXNORM|TELAPREVIR 375MG ORAL TABLET|TELAPREVIR 375 MG ORAL TABLET
C3154711|T121|1102280|RXNORM|TELAPREVIR 375MG TAB,UD|TELAPREVIR 375 MG ORAL TABLET
C3154711|T121|1102280|RXNORM|TELAPREVIR 375MG UD TAB|TELAPREVIR 375 MG ORAL TABLET
C3154711|T121|1102280|RXNORM|TELAPREVIR 375MG TAB,UD [VA PRODUCT]|TELAPREVIR 375 MG ORAL TABLET
C3154711|T121|1102280|RXNORM|TELAPREVIR 375MG TABLET|TELAPREVIR 375 MG ORAL TABLET
C3154711|T121|1102280|RXNORM|TELAPREVIR 375MG TABLET |TELAPREVIR 375 MG ORAL TABLET
C2605856|T121||RXNORM|435350, TMC
C2605856|T121||RXNORM|TMC435350
C2605856|T121||RXNORM|TMC-435350
C2605856|T121||RXNORM|TMC 435350
C2745868|T121||RXNORM|435, TMC
C2745868|T121||RXNORM|TMC435
C2745868|T121||RXNORM|TMC-435
C2745868|T121||RXNORM|TMC 435
C3696409|T121|1482802|RXNORM|OLYSIO|OLYSIO
C2605855|T121|1482790|RXNORM|SIMEPREVIR|SIMEPREVIR
C2605855|T121|1482790|RXNORM|SIMEPREVIR |SIMEPREVIR
C2605855|T121|1482790|RXNORM|ANTIVIRAL SIMEPREVIR|SIMEPREVIR
C2605855|T121|1482790|RXNORM|SIMEPREVIR |SIMEPREVIR
C2605855|T121|1482790|RXNORM|N-(17-(2-(4-ISOPROPYLTHIAZOLE-2-YL)-7-METHOXY-8-METHYLQUINOLIN-4-YLOXY)-13-METHYL-2,14-DIOXO-3,13-DIAZATRICYCLO(13.3.0.04,6)OCTADEC-7-ENE-4-CARBONYL)(CYCLOPROPYL)SULFONAMIDE|SIMEPREVIR
C2605855|T121|1482790|RXNORM|SIMEPREVIR [CHEMICAL/INGREDIENT]|SIMEPREVIR
C2605855|T121|1482790|RXNORM|SIMEPREVIR |SIMEPREVIR
C3696072|T121|1484518|RXNORM|SIMEPREVIR SODIUM|SIMEPREVIR SODIUM
C3696072|T121|1484518|RXNORM|SIMEPREVIR (AS SODIUM)|SIMEPREVIR SODIUM
C3696748|T121|1482798|RXNORM|SIMEPREVIR ORAL PRODUCT|SIMEPREVIR ORAL PRODUCT
C3696748|T121|1482798|RXNORM|ORAL FORM SIMEPREVIR |SIMEPREVIR ORAL PRODUCT
C3696748|T121|1482798|RXNORM|ORAL FORM SIMEPREVIR|SIMEPREVIR ORAL PRODUCT
C4075528|T121||RXNORM|SIMEPREVIR + SOFOSBUVIR 
C4075528|T121||RXNORM|SIMEPREVIR + SOFOSBUVIR
C3154653|T121|1102136|RXNORM|BOCEPREVIR 200 MG ORAL CAPSULE [VICTRELIS]|VICTRELIS 200 MG ORAL CAPSULE
C3154653|T121|1102136|RXNORM|VICTRELIS 200 MG ORAL CAPSULE|VICTRELIS 200 MG ORAL CAPSULE
C3154653|T121|1102136|RXNORM|VICTRELIS 200MG CAPSULE|VICTRELIS 200 MG ORAL CAPSULE
C3154653|T121|1102136|RXNORM|VICTRELIS, 200 MG ORAL CAPSULE|VICTRELIS 200 MG ORAL CAPSULE
C3154713|T121|1102282|RXNORM|TELAPREVIR 375 MG ORAL TABLET [INCIVEK]|INCIVEK 375 MG ORAL TABLET
C3154713|T121|1102282|RXNORM|INCIVEK 375 MG ORAL TABLET|INCIVEK 375 MG ORAL TABLET
C3154713|T121|1102282|RXNORM|INCIVEK 375MG TABLET|INCIVEK 375 MG ORAL TABLET
C3154713|T121|1102282|RXNORM|INCIVEK, 375 MG ORAL TABLET|INCIVEK 375 MG ORAL TABLET
C3154713|T121|1102282|RXNORM|INCIVEK 375 MG ORAL TABLET, TWICE DAILY|INCIVEK 375 MG ORAL TABLET
C0697341|T121|856450|RXNORM|INDERAL 10MG TABLET|INDERAL 10 MG ORAL TABLET
C0697341|T121|856450|RXNORM|INDERAL, 10 MG ORAL TABLET|INDERAL 10 MG ORAL TABLET
C0697341|T121|856450|RXNORM|INDERAL 10 MG ORAL TABLET|INDERAL 10 MG ORAL TABLET
C0697341|T121|856450|RXNORM|PROPRANOLOL HYDROCHLORIDE 10 MG ORAL TABLET [INDERAL]|INDERAL 10 MG ORAL TABLET
C0282321|T121|82084|RXNORM|HYDROCHLORIDE, PROPRANOLOL|PROPRANOLOL HYDROCHLORIDE
C0282321|T121|82084|RXNORM|PROPRANOLOL HYDROCHLORIDE|PROPRANOLOL HYDROCHLORIDE
C0282321|T121|82084|RXNORM|2-PROPANOL-1-[(1-METHYLETHYL)AMINO]-3-(1-NAPHTHALENYLOXY) HYDROCHLORIDE|PROPRANOLOL HYDROCHLORIDE
C0282321|T121|82084|RXNORM|PROPRANOLOL HYDROCHLORIDE PRODUCT|PROPRANOLOL HYDROCHLORIDE
C0282321|T121|82084|RXNORM|PROPRANOLOL HYDROCHLORIDE |PROPRANOLOL HYDROCHLORIDE
C0282321|T121|82084|RXNORM|PROPRANOLOL HYDROCHLORIDE [CHEMICAL/INGREDIENT]|PROPRANOLOL HYDROCHLORIDE
C0282321|T121|82084|RXNORM|PROPRANOLOL HYDROCHLORIDE [2]|PROPRANOLOL HYDROCHLORIDE
C0282321|T121|82084|RXNORM|PROPRANOLOL HYDROCHLORIDE [2] |PROPRANOLOL HYDROCHLORIDE
C0282321|T121|82084|RXNORM|PROPRANOLOL HYDROCHLORIDE |PROPRANOLOL HYDROCHLORIDE
C0282321|T121|82084|RXNORM|PROPRANOLOL HYDROCHLORIDE |PROPRANOLOL HYDROCHLORIDE
C0282321|T121|82084|RXNORM|PROPRANOLOL HYDROCHLORIDE [2] |PROPRANOLOL HYDROCHLORIDE
C0282321|T121|82084|RXNORM|PROPRANOLOL HYDROCHLORIDE PRODUCT |PROPRANOLOL HYDROCHLORIDE
C0282321|T121|82084|RXNORM|PROPRANOLOL HYDROCHLORIDE PRODUCT |PROPRANOLOL HYDROCHLORIDE
C0591636|T121|151890|RXNORM|INDERAL|INDERAL
C0697332|T121|200836|RXNORM|INDERAL 160 MG ORAL TABLET|INDERAL 160 MG ORAL TABLET
C0697332|T121|200836|RXNORM|PROPRANOLOL HYDROCHLORIDE 160 MG ORAL TABLET [INDERAL]|INDERAL 160 MG ORAL TABLET
C1271144|T121|387876|RXNORM|INDERAL 80 MG ORAL CAPSULE|INDERAL 80 MG ORAL CAPSULE
C1271144|T121|387876|RXNORM|PROPRANOLOL HYDROCHLORIDE 80 MG ORAL CAPSULE [INDERAL]|INDERAL 80 MG ORAL CAPSULE
C1271144|T121|387876|RXNORM|INDERAL 80MG CAPSULE|INDERAL 80 MG ORAL CAPSULE
C1271144|T121|387876|RXNORM|INDERAL 80MG CAPSULE |INDERAL 80 MG ORAL CAPSULE
C0709222|T121|856462|RXNORM|PROPRANOLOL HYDROCHLORIDE 120 MILLIGRAM IN 1 CAPSULE ORAL CAPSULE, EXTENDED RELEASE [INDERAL LA]|INDERAL XL 120 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C0709222|T121|856462|RXNORM|INDERAL LA 120MG EXTENDED-RELEASE CAPSULE|INDERAL XL 120 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C0709222|T121|856462|RXNORM|INDERAL LA, 120 MG ORAL CAPSULE, EXTENDED RELEASE|INDERAL XL 120 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C0709222|T121|856462|RXNORM|PROPRANOLOL HYDROCHLORIDE 120 MG ORAL CAPSULE, EXTENDED RELEASE [INDERAL LA]|INDERAL XL 120 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C0709222|T121|856462|RXNORM|PROPRANOLOL HYDROCHLORIDE 120 MG ORAL CAPSULE, EXTENDED RELEASE [INDERAL XL]|INDERAL XL 120 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C0709222|T121|856462|RXNORM|INDERAL XL, 120 MG ORAL CAPSULE, EXTENDED RELEASE|INDERAL XL 120 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C0709222|T121|856462|RXNORM|INDERAL XL 120MG EXTENDED-RELEASE CAPSULE|INDERAL XL 120 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C0709222|T121|856462|RXNORM|24 HR PROPRANOLOL HYDROCHLORIDE 120 MG EXTENDED RELEASE ORAL CAPSULE [INDERAL]|INDERAL XL 120 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C0709222|T121|856462|RXNORM|INDERAL LA 120 MG 24HR EXTENDED RELEASE ORAL CAPSULE|INDERAL XL 120 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C0709222|T121|856462|RXNORM|INDERAL XL 120 MG 24 HR EXTENDED RELEASE ORAL CAPSULE|INDERAL XL 120 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C2710362|T121|856464|RXNORM|INDERAL 120 MG EXTENDED RELEASE ORAL CAPSULE|INDERAL 120 MG EXTENDED RELEASE ORAL CAPSULE
C2710362|T121|856464|RXNORM|PROPRANOLOL HYDROCHLORIDE 120 MG EXTENDED RELEASE ORAL CAPSULE [INDERAL]|INDERAL 120 MG EXTENDED RELEASE ORAL CAPSULE
C0697868|T121|856483|RXNORM|PROPRANOLOL HYDROCHLORIDE 160 MILLIGRAM IN 1 CAPSULE ORAL CAPSULE, EXTENDED RELEASE [INDERAL LA]|24 HR INDERAL LA 160 MG EXTENDED RELEASE ORAL CAPSULE
C0697868|T121|856483|RXNORM|INDERAL LA 160MG EXTENDED-RELEASE CAPSULE|24 HR INDERAL LA 160 MG EXTENDED RELEASE ORAL CAPSULE
C0697868|T121|856483|RXNORM|INDERAL LA, 160 MG ORAL CAPSULE, EXTENDED RELEASE|24 HR INDERAL LA 160 MG EXTENDED RELEASE ORAL CAPSULE
C0697868|T121|856483|RXNORM|PROPRANOLOL HYDROCHLORIDE 160 MG ORAL CAPSULE, EXTENDED RELEASE [INDERAL LA]|24 HR INDERAL LA 160 MG EXTENDED RELEASE ORAL CAPSULE
C0697868|T121|856483|RXNORM|INDERAL LA 160 MG 24 HR EXTENDED RELEASE ORAL CAPSULE|24 HR INDERAL LA 160 MG EXTENDED RELEASE ORAL CAPSULE
C0697868|T121|856483|RXNORM|INDERAL LA 160 MG 24HR EXTENDED RELEASE ORAL CAPSULE|24 HR INDERAL LA 160 MG EXTENDED RELEASE ORAL CAPSULE
C0697868|T121|856483|RXNORM|24 HR INDERAL LA 160 MG EXTENDED RELEASE ORAL CAPSULE|24 HR INDERAL LA 160 MG EXTENDED RELEASE ORAL CAPSULE
C0697868|T121|856483|RXNORM|24 HR PROPRANOLOL HYDROCHLORIDE 160 MG EXTENDED RELEASE ORAL CAPSULE [INDERAL]|24 HR INDERAL LA 160 MG EXTENDED RELEASE ORAL CAPSULE
C2710375|T121|856485|RXNORM|PROPRANOLOL HYDROCHLORIDE 160 MG EXTENDED RELEASE ORAL CAPSULE [INDERAL]|INDERAL 160 MG EXTENDED RELEASE ORAL CAPSULE
C2710375|T121|856485|RXNORM|INDERAL 160 MG EXTENDED RELEASE ORAL CAPSULE|INDERAL 160 MG EXTENDED RELEASE ORAL CAPSULE
C0709233|T121|856508|RXNORM|INDERAL 20MG TABLET|INDERAL 20 MG ORAL TABLET
C0709233|T121|856508|RXNORM|INDERAL, 20 MG ORAL TABLET|INDERAL 20 MG ORAL TABLET
C0709233|T121|856508|RXNORM|PROPRANOLOL HYDROCHLORIDE 20 MG ORAL TABLET [INDERAL]|INDERAL 20 MG ORAL TABLET
C0709233|T121|856508|RXNORM|INDERAL 20 MG ORAL TABLET|INDERAL 20 MG ORAL TABLET
C0697330|T121|856521|RXNORM|INDERAL 40MG TABLET|INDERAL 40 MG ORAL TABLET
C0697330|T121|856521|RXNORM|INDERAL, 40 MG ORAL TABLET|INDERAL 40 MG ORAL TABLET
C0697330|T121|856521|RXNORM|PROPRANOLOL HYDROCHLORIDE 40 MG ORAL TABLET [INDERAL]|INDERAL 40 MG ORAL TABLET
C0697330|T121|856521|RXNORM|INDERAL 40 MG ORAL TABLET|INDERAL 40 MG ORAL TABLET
C0709220|T121|856537|RXNORM|PROPRANOLOL HYDROCHLORIDE 60 MILLIGRAM IN 1 CAPSULE ORAL CAPSULE, EXTENDED RELEASE [INDERAL LA]|INDERAL LA 60 MG 24HR EXTENDED RELEASE ORAL CAPSULE
C0709220|T121|856537|RXNORM|INDERAL LA 60MG EXTENDED-RELEASE CAPSULE|INDERAL LA 60 MG 24HR EXTENDED RELEASE ORAL CAPSULE
C0709220|T121|856537|RXNORM|INDERAL LA, 60 MG ORAL CAPSULE, EXTENDED RELEASE|INDERAL LA 60 MG 24HR EXTENDED RELEASE ORAL CAPSULE
C0709220|T121|856537|RXNORM|PROPRANOLOL HYDROCHLORIDE 60 MG ORAL CAPSULE, EXTENDED RELEASE [INDERAL LA]|INDERAL LA 60 MG 24HR EXTENDED RELEASE ORAL CAPSULE
C0709220|T121|856537|RXNORM|INDERAL LA 60 MG 24 HR EXTENDED RELEASE ORAL CAPSULE|INDERAL LA 60 MG 24HR EXTENDED RELEASE ORAL CAPSULE
C0709220|T121|856537|RXNORM|24 HR PROPRANOLOL HYDROCHLORIDE 60 MG EXTENDED RELEASE ORAL CAPSULE [INDERAL]|INDERAL LA 60 MG 24HR EXTENDED RELEASE ORAL CAPSULE
C0709220|T121|856537|RXNORM|24 HR INDERAL LA 60 MG EXTENDED RELEASE ORAL CAPSULE|INDERAL LA 60 MG 24HR EXTENDED RELEASE ORAL CAPSULE
C0709220|T121|856537|RXNORM|INDERAL LA 60 MG 24HR EXTENDED RELEASE ORAL CAPSULE|INDERAL LA 60 MG 24HR EXTENDED RELEASE ORAL CAPSULE
C2710407|T121|856539|RXNORM|INDERAL 60 MG EXTENDED RELEASE ORAL CAPSULE|INDERAL 60 MG EXTENDED RELEASE ORAL CAPSULE
C2710407|T121|856539|RXNORM|PROPRANOLOL HYDROCHLORIDE 60 MG EXTENDED RELEASE ORAL CAPSULE [INDERAL]|INDERAL 60 MG EXTENDED RELEASE ORAL CAPSULE
C0709234|T121|856557|RXNORM|INDERAL 60MG TABLET|INDERAL 60 MG ORAL TABLET
C0709234|T121|856557|RXNORM|INDERAL, 60 MG ORAL TABLET|INDERAL 60 MG ORAL TABLET
C0709234|T121|856557|RXNORM|INDERAL 60 MG ORAL TABLET|INDERAL 60 MG ORAL TABLET
C0709234|T121|856557|RXNORM|PROPRANOLOL HYDROCHLORIDE 60 MG ORAL TABLET [INDERAL]|INDERAL 60 MG ORAL TABLET
C0697871|T121|856571|RXNORM|PROPRANOLOL HYDROCHLORIDE 80 MILLIGRAM IN 1 CAPSULE ORAL CAPSULE, EXTENDED RELEASE [INDERAL LA]|INDERAL XL 80 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C0697871|T121|856571|RXNORM|INDERAL LA 80MG EXTENDED-RELEASE CAPSULE|INDERAL XL 80 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C0697871|T121|856571|RXNORM|INDERAL LA, 80 MG ORAL CAPSULE, EXTENDED RELEASE|INDERAL XL 80 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C0697871|T121|856571|RXNORM|PROPRANOLOL HYDROCHLORIDE 80 MG ORAL CAPSULE, EXTENDED RELEASE [INDERAL LA]|INDERAL XL 80 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C0697871|T121|856571|RXNORM|PROPRANOLOL HYDROCHLORIDE 80 MG ORAL CAPSULE, EXTENDED RELEASE [INDERAL XL]|INDERAL XL 80 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C0697871|T121|856571|RXNORM|INDERAL XL 80MG EXTENDED-RELEASE CAPSULE|INDERAL XL 80 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C0697871|T121|856571|RXNORM|INDERAL XL, 80 MG ORAL CAPSULE, EXTENDED RELEASE|INDERAL XL 80 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C0697871|T121|856571|RXNORM|24 HR PROPRANOLOL HYDROCHLORIDE 80 MG EXTENDED RELEASE ORAL CAPSULE [INDERAL]|INDERAL XL 80 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C0697871|T121|856571|RXNORM|INDERAL XL 80 MG 24 HR EXTENDED RELEASE ORAL CAPSULE|INDERAL XL 80 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C0697871|T121|856571|RXNORM|INDERAL LA 80 MG 24HR EXTENDED RELEASE ORAL CAPSULE|INDERAL XL 80 MG 24 HR EXTENDED RELEASE ORAL CAPSULE
C2710423|T121|856573|RXNORM|INDERAL 80 MG EXTENDED RELEASE ORAL CAPSULE|INDERAL 80 MG EXTENDED RELEASE ORAL CAPSULE
C2710423|T121|856573|RXNORM|PROPRANOLOL HYDROCHLORIDE 80 MG EXTENDED RELEASE ORAL CAPSULE [INDERAL]|INDERAL 80 MG EXTENDED RELEASE ORAL CAPSULE
C0697347|T121|856579|RXNORM|INDERAL 80MG TABLET|INDERAL 80 MG ORAL TABLET
C0697347|T121|856579|RXNORM|INDERAL, 80 MG ORAL TABLET|INDERAL 80 MG ORAL TABLET
C0697347|T121|856579|RXNORM|PROPRANOLOL HYDROCHLORIDE 80 MG ORAL TABLET [INDERAL]|INDERAL 80 MG ORAL TABLET
C0697347|T121|856579|RXNORM|INDERAL 80 MG ORAL TABLET|INDERAL 80 MG ORAL TABLET
C1306227|T121|393312|RXNORM|PROPRANOLOL ORAL CAPSULE [INDERAL]|PROPRANOLOL ORAL CAPSULE [INDERAL]
C1577533|T121|491323|RXNORM|PROPRANOLOL EXTENDED RELEASE ORAL CAPSULE [INDERAL]|PROPRANOLOL EXTENDED RELEASE ORAL CAPSULE [INDERAL]
C0306453|T121|92960|RXNORM|PROPRANOLOL ORAL TABLET [INDERAL]|PROPRANOLOL ORAL TABLET [INDERAL]
C0059478|T121||RXNORM|EPSILON-N-1-(1-DEOXYLACTULOSYL)LYSINE
C0701236|T121||RXNORM|NORMASE
C0701237|T121||RXNORM|AMIVALEX
C0719221|T121|215949|RXNORM|CEPHULAC|CEPHULAC
C0719324|T121|216045|RXNORM|CHOLAC|CHOLAC
C0719340|T121|216060|RXNORM|CHRONULAC|CHRONULAC
C0719488|T121|216200|RXNORM|CONSTILAC|CONSTILAC
C0719489|T121|216201|RXNORM|CONSTULOSE|CONSTULOSE
C0720231|T121|216928|RXNORM|ENULOSE|ENULOSE
C0720316|T121|217008|RXNORM|EVALOSE|EVALOSE
C0720632|T121|217314|RXNORM|GENERLAC|GENERLAC
C0720849|T121|217522|RXNORM|HEPTALAC|HEPTALAC
C0721265|T121|217928|RXNORM|KRISTALOSE|KRISTALOSE
C0116371|T121||RXNORM|EPSILON-(DEOXYLACTULOSE)LYSINE
C0125215|T121||RXNORM|LACTOSE-LYSINE
C0125227|T121||RXNORM|LACTULOSE-LYSINE
C0284752|T121||RXNORM|LACTULOSELYSINE
C0022957|T121|6218|RXNORM|LACTULOSE|LACTULOSE
C0022957|T121|6218|RXNORM|D-FRUCTOSE, 4-O-BETA-D-GALACTOPYRANOSYL-|LACTULOSE
C0022957|T121|6218|RXNORM|LACTULOSE |LACTULOSE
C0022957|T121|6218|RXNORM|LAXATIVES LACTULOSE|LACTULOSE
C0022957|T121|6218|RXNORM|4-O-BETA-D-GALACTOPYRANOSYL-D-FRUCTOFURANOSE|LACTULOSE
C0022957|T121|6218|RXNORM|LACTULOSE [CHEMICAL/INGREDIENT]|LACTULOSE
C0022957|T121|6218|RXNORM|LACTULOSE PRODUCT|LACTULOSE
C0022957|T121|6218|RXNORM|LACTULOSE |LACTULOSE
C0022957|T121|6218|RXNORM|LACTULOSE |LACTULOSE
C1737835|T121|1251194|RXNORM|LACTULOSE 20G POWDER FOR ORAL SOL/PWD [CONSTIPATION]|LACTULOSE 20 GM GRANULES FOR ORAL SOLUTION
C1737835|T121|1251194|RXNORM|LACTULOSE 20GM/PKT PWDR|LACTULOSE 20 GM GRANULES FOR ORAL SOLUTION
C1737835|T121|1251194|RXNORM|LACTULOSE ORAL CRYSTAL PACKET 20 GM|LACTULOSE 20 GM GRANULES FOR ORAL SOLUTION
C1737835|T121|1251194|RXNORM|LACTULOSE 20GM/PKT PWDR [VA PRODUCT]|LACTULOSE 20 GM GRANULES FOR ORAL SOLUTION
C1737835|T121|1251194|RXNORM|LACTULOSE 167 MG/ML ORAL SOLUTION|LACTULOSE 20 GM GRANULES FOR ORAL SOLUTION
C1737835|T121|1251194|RXNORM|LACTULOSE 20 GM PER 4 OZ. POWDER FOR ORAL SOLUTION|LACTULOSE 20 GM GRANULES FOR ORAL SOLUTION
C1737835|T121|1251194|RXNORM|LACTULOSE 20 G ORAL POWDER FOR RECONSTITUTION|LACTULOSE 20 GM GRANULES FOR ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 667 MG/ML ORAL SOLUTION|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE (ENCEPHALOPATHY) SOLUTION 10 GM/15ML|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE SOLUTION 10 GM/15ML|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10G/15ML ORAL SOLUTION [ENCEPHALOPATHY]|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10G/15ML ORAL SOLUTION [CONSTIPATION]|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10GM/15ML SYRUP|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10 GM/15 ML SOLUTION|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10 G IN 15 ML ORAL SOLUTION|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10 GM PER 15 ML ORAL SOLUTION|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10 G IN 15 ML ORAL SOLUTION [LACTULOSE]|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10GM/15ML SYRUP [VA PRODUCT]|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 20 G IN 30 ML ORAL SOLUTION|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10 G IN 15 ML RECTAL SOLUTION|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE, 10 G/15 ML ORAL AND RECTAL LIQUID|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10 G/15 ML ORAL AND RECTAL LIQUID|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10GM/15ML ORAL SOLN|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10GM/15ML SOLN,ORAL|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10GM/15ML SOLN,ORAL [VA PRODUCT]|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10G/15 ML SOLUTION |LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10G/15 ML SOLUTION|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|ACILAC 10G/15ML SOLUTION|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10G/15ML SOLUTION |LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10G/15ML SOLUTION|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10G/15ML SYRUP |LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10G/15ML SYRUP|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10 GM/15 ML ORAL SOLUTION|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10 GM/15 ML ORAL SYRUP|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE, 10 G/15 ML ORAL SYRUP|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C1298316|T121|391937|RXNORM|LACTULOSE 10 G/15 ML ORAL SYRUP|LACTULOSE 20 GM PER 30 ML ORAL SOLUTION
C3216531|T121|1162201|RXNORM|LACTULOSE ORAL PRODUCT|LACTULOSE ORAL PRODUCT
C3216531|T121|1162201|RXNORM|ORAL FORM LACTULOSE |LACTULOSE ORAL PRODUCT
C3216531|T121|1162201|RXNORM|ORAL FORM LACTULOSE|LACTULOSE ORAL PRODUCT
C0353982|T121|104148|RXNORM|LACTULOSE 670 MG/ML ORAL SOLUTION|LACTULOSE 3.35 GM PER 5 ML ORAL SOLUTION
C0353982|T121|104148|RXNORM|LACTULOSE 3.35 GM PER 5 ML ORAL SOLUTION|LACTULOSE 3.35 GM PER 5 ML ORAL SOLUTION
C0353982|T121|104148|RXNORM|LACTULOSE 3.35G/5ML ORAL SOLUTION|LACTULOSE 3.35 GM PER 5 ML ORAL SOLUTION
C0353982|T121|104148|RXNORM|LACTULOSE 3.35G/5ML ORAL SOLUTION |LACTULOSE 3.35 GM PER 5 ML ORAL SOLUTION
C0353982|T121|104148|RXNORM|LACTULOSE 3.35G/5ML ORAL SOLUTION |LACTULOSE 3.35 GM PER 5 ML ORAL SOLUTION
C0591418|T121|151674|RXNORM|DUPHALAC|DUPHALAC
C1589304|T121|544446|RXNORM|CATULAC|CATULAC
C1589311|T121|544456|RXNORM|RO-LACTULOSE|RO-LACTULOSE
C0605673|T121||RXNORM|CHOLAN-24-OIC ACID, 3,7,12-TRIOXO-, (5BETA)-, MIXT. WITH (3(S)-ENDO)-8-(2-(1,1'-BIPHENYL)-4-YL-2-OXOETHYL)-3-(3-HYDROXY-1-OXO-2-PHENYLPROPOXY)-8-METHYL-8-AZONIABICYCLO(3.2.1)OCTANE BROMIDE, 4-O-BETA-D-GALACTOPYRANOSYL-D-FRUCTOSE AND PANCREATIN
C0605673|T121||RXNORM|FZ 560
C0605673|T121||RXNORM|FZ-560
C0708296|T121|755470|RXNORM|LACTULOSE 10 GRAM IN 15 MILLILITER ORAL LIQUID [ENULOSE]|ENULOSE 10 GM PER 15 ML SYRUP
C0708296|T121|755470|RXNORM|LACTULOSE 10 GRAM IN 15 MILLILITER RECTAL LIQUID [ENULOSE]|ENULOSE 10 GM PER 15 ML SYRUP
C0708296|T121|755470|RXNORM|LACTULOSE 667 MG/ML ORAL SOLUTION [ENULOSE]|ENULOSE 10 GM PER 15 ML SYRUP
C0708296|T121|755470|RXNORM|ENULOSE 667 MG/ML ORAL SOLUTION|ENULOSE 10 GM PER 15 ML SYRUP
C0708296|T121|755470|RXNORM|ENULOSE 10 GM PER 15 ML SYRUP|ENULOSE 10 GM PER 15 ML SYRUP
C0708296|T121|755470|RXNORM|LACTULOSE 10 GM/15 ML ORAL SOLUTION [ENULOSE]|ENULOSE 10 GM PER 15 ML SYRUP
C0708296|T121|755470|RXNORM|LACTULOSE 10 GM/15 ML ORAL SYRUP [ENULOSE]|ENULOSE 10 GM PER 15 ML SYRUP
C0708296|T121|755470|RXNORM|LACTULOSE 10 G IN 15 ML RECTAL SOLUTION [ENULOSE]|ENULOSE 10 GM PER 15 ML SYRUP
C0708296|T121|755470|RXNORM|LACTULOSE 10 G IN 15 ML ORAL SOLUTION [ENULOSE]|ENULOSE 10 GM PER 15 ML SYRUP
C0708296|T121|755470|RXNORM|ENULOSE, 10 G/15 ML ORAL AND RECTAL LIQUID|ENULOSE 10 GM PER 15 ML SYRUP
C0708296|T121|755470|RXNORM|ENULOSE 10G/15ML SOLUTION|ENULOSE 10 GM PER 15 ML SYRUP
C0994966|T121|756967|RXNORM|LACTULOSE ORAL SOLUTION [ENULOSE]|LACTULOSE ORAL SOLUTION [ENULOSE]
C0994966|T121|756967|RXNORM|LACTULOSE 10GM/15ML SYRUP|LACTULOSE ORAL SOLUTION [ENULOSE]
C0994966|T121|756967|RXNORM|ENULOSE SYRUP|LACTULOSE ORAL SOLUTION [ENULOSE]
C0994966|T121|756967|RXNORM|ENULOSE SYRUP [VA PRODUCT]|LACTULOSE ORAL SOLUTION [ENULOSE]
C1589305|T121|544447|RXNORM|LACTULOSE 667 MG/ML [CATULAC]|LACTULOSE 667 MG/ML [CATULAC]
C1589307|T121|544450|RXNORM|LACTULOSE 667 MG/ML [CONSTULOSE]|LACTULOSE 667 MG/ML [CONSTULOSE]
C1589309|T121|544453|RXNORM|LACTULOSE 667 MG/ML [GENERLAC]|LACTULOSE 667 MG/ML [GENERLAC]
C1589312|T121|544457|RXNORM|LACTULOSE 667 MG/ML [RO-LACTULOSE]|LACTULOSE 667 MG/ML [RO-LACTULOSE]
C1600249|T121|567832|RXNORM|LACTULOSE 667 MG/ML [CEPHULAC]|LACTULOSE 667 MG/ML [CEPHULAC]
C1600250|T121|567833|RXNORM|LACTULOSE 667 MG/ML [CHOLAC]|LACTULOSE 667 MG/ML [CHOLAC]
C1600251|T121|567834|RXNORM|LACTULOSE 667 MG/ML [CHRONULAC]|LACTULOSE 667 MG/ML [CHRONULAC]
C1600252|T121|567835|RXNORM|LACTULOSE 667 MG/ML [CONSTILAC]|LACTULOSE 667 MG/ML [CONSTILAC]
C1600253|T121|567836|RXNORM|LACTULOSE 667 MG/ML [DUPHALAC]|LACTULOSE 667 MG/ML [DUPHALAC]
C1600254|T121|567837|RXNORM|LACTULOSE 667 MG/ML [ENULOSE]|LACTULOSE 667 MG/ML [ENULOSE]
C1600255|T121|567838|RXNORM|LACTULOSE 667 MG/ML [EVALOSE]|LACTULOSE 667 MG/ML [EVALOSE]
C1600256|T121|567839|RXNORM|LACTULOSE 667 MG/ML [HEPTALAC]|LACTULOSE 667 MG/ML [HEPTALAC]
C0978083|T121|1251190|RXNORM|LACTULOSE 10G POWDER FOR ORAL SOL/PWD [CONSTIPATION]|LACTULOSE 10 GM GRANULES FOR ORAL SOLUTION
C0978083|T121|1251190|RXNORM|LACTULOSE 10GM/PKT PWDR|LACTULOSE 10 GM GRANULES FOR ORAL SOLUTION
C0978083|T121|1251190|RXNORM|LACTULOSE ORAL CRYSTAL PACKET 10 GM|LACTULOSE 10 GM GRANULES FOR ORAL SOLUTION
C0978083|T121|1251190|RXNORM|LACTULOSE 10GM/PKT PWDR [VA PRODUCT]|LACTULOSE 10 GM GRANULES FOR ORAL SOLUTION
C0978083|T121|1251190|RXNORM|LACTULOSE 10 GM PER 4 OZ. POWDER FOR ORAL SOLUTION|LACTULOSE 10 GM GRANULES FOR ORAL SOLUTION
C0978083|T121|1251190|RXNORM|LACTULOSE 83.3 MG/ML ORAL SOLUTION|LACTULOSE 10 GM GRANULES FOR ORAL SOLUTION
C0978083|T121|1251190|RXNORM|LACTULOSE 10 G ORAL POWDER FOR RECONSTITUTION|LACTULOSE 10 GM GRANULES FOR ORAL SOLUTION
C1352027|T121|422759|RXNORM|LACTULOSE 660 MG/ML ORAL SOLUTION|LACTULOSE 660 MG/ML ORAL SOLUTION
C1238377|T121||RXNORM|LACTULOSE ORAL SOLUTION [KRISTALOSE]
C1589308|T121|544451|RXNORM|LACTULOSE ORAL SOLUTION [CONSTULOSE]|LACTULOSE ORAL SOLUTION [CONSTULOSE]
C1589310|T121|544454|RXNORM|LACTULOSE ORAL SOLUTION [GENERLAC]|LACTULOSE ORAL SOLUTION [GENERLAC]
C1589313|T121|544458|RXNORM|LACTULOSE ORAL SOLUTION [RO-LACTULOSE]|LACTULOSE ORAL SOLUTION [RO-LACTULOSE]
C1355127|T121|756118|RXNORM|LACTULOSE 606 MG/ML ORAL SOLUTION|LACTULOSE 606 MG/ML ORAL SOLUTION
C1355126|T121|756119|RXNORM|LACTULOSE 650 MG/ML ORAL SOLUTION|LACTULOSE 650 MG/ML ORAL SOLUTION
C1355125|T121|756120|RXNORM|LACTULOSE 666 MG/ML ORAL SOLUTION|LACTULOSE 666 MG/ML ORAL SOLUTION
C1589306|T121|756961|RXNORM|LACTULOSE ORAL SOLUTION [CATULAC]|LACTULOSE ORAL SOLUTION [CATULAC]
C2240661|T121|756962|RXNORM|LACTULOSE ORAL SOLUTION [CEPHULAC]|LACTULOSE ORAL SOLUTION [CEPHULAC]
C1239130|T121|756963|RXNORM|LACTULOSE ORAL SOLUTION [CHOLAC]|LACTULOSE ORAL SOLUTION [CHOLAC]
C2240662|T121|756964|RXNORM|LACTULOSE ORAL SOLUTION [CHRONULAC]|LACTULOSE ORAL SOLUTION [CHRONULAC]
C1239069|T121|756965|RXNORM|LACTULOSE ORAL SOLUTION [CONSTILAC]|LACTULOSE ORAL SOLUTION [CONSTILAC]
C2240663|T121|756966|RXNORM|LACTULOSE ORAL SOLUTION [DUPHALAC]|LACTULOSE ORAL SOLUTION [DUPHALAC]
C1239128|T121|756968|RXNORM|LACTULOSE ORAL SOLUTION [EVALOSE]|LACTULOSE ORAL SOLUTION [EVALOSE]
C1239126|T121|756969|RXNORM|LACTULOSE ORAL SOLUTION [HEPTALAC]|LACTULOSE ORAL SOLUTION [HEPTALAC]
C1586235|T121|544452|RXNORM|LACTULOSE 667 MG/ML ORAL SOLUTION [CONSTULOSE]|CONSTULOSE 10 GM PER 15 ML SYRUP
C1586235|T121|544452|RXNORM|CONSTULOSE 667 MG/ML ORAL SOLUTION|CONSTULOSE 10 GM PER 15 ML SYRUP
C1586235|T121|544452|RXNORM|CONSTULOSE 10 GM PER 15 ML SYRUP|CONSTULOSE 10 GM PER 15 ML SYRUP
C1586235|T121|544452|RXNORM|LACTULOSE 10 GM/15 ML ORAL SOLUTION [CONSTULOSE]|CONSTULOSE 10 GM PER 15 ML SYRUP
C1586235|T121|544452|RXNORM|LACTULOSE 10 GM/15 ML ORAL SYRUP [CONSTULOSE]|CONSTULOSE 10 GM PER 15 ML SYRUP
C1586235|T121|544452|RXNORM|LACTULOSE 10 G IN 15 ML ORAL SOLUTION [CONSTULOSE]|CONSTULOSE 10 GM PER 15 ML SYRUP
C1586235|T121|544452|RXNORM|CONSTULOSE 10G/15ML SOLUTION|CONSTULOSE 10 GM PER 15 ML SYRUP
C1586235|T121|544452|RXNORM|CONSTULOSE, 10 G/15 ML ORAL SYRUP|CONSTULOSE 10 GM PER 15 ML SYRUP
C1586236|T121|544455|RXNORM|GENERLAC 667 MG/ML ORAL SOLUTION|GENERLAC 667 MG/ML ORAL SOLUTION
C1586236|T121|544455|RXNORM|LACTULOSE 667 MG/ML ORAL SOLUTION [GENERLAC]|GENERLAC 667 MG/ML ORAL SOLUTION
C1586236|T121|544455|RXNORM|LACTULOSE 10 GM/15 ML ORAL SOLUTION [GENERLAC]|GENERLAC 667 MG/ML ORAL SOLUTION
C1586236|T121|544455|RXNORM|LACTULOSE 10 G IN 15 ML ORAL SOLUTION [GENERLAC]|GENERLAC 667 MG/ML ORAL SOLUTION
C1586236|T121|544455|RXNORM|GENERLAC 10 GM PER 15 ML ORAL SOLUTION|GENERLAC 667 MG/ML ORAL SOLUTION
C1586236|T121|544455|RXNORM|GENERLAC, 10 G/15 ML ORAL AND RECTAL LIQUID|GENERLAC 667 MG/ML ORAL SOLUTION
C1586236|T121|544455|RXNORM|GENERLAC 10G/15ML SOLUTION|GENERLAC 667 MG/ML ORAL SOLUTION
C3221021|T121|1166820|RXNORM|CEPHULAC ORAL LIQUID PRODUCT|CEPHULAC ORAL LIQUID PRODUCT
C3221216|T121|1167018|RXNORM|DUPHALAC ORAL LIQUID PRODUCT|DUPHALAC ORAL LIQUID PRODUCT
C3221248|T121|1167052|RXNORM|ENULOSE ORAL LIQUID PRODUCT|ENULOSE ORAL LIQUID PRODUCT
C3222920|T121|1168756|RXNORM|CONSTILAC ORAL LIQUID PRODUCT|CONSTILAC ORAL LIQUID PRODUCT
C3222922|T121|1168758|RXNORM|CONSTULOSE ORAL LIQUID PRODUCT|CONSTULOSE ORAL LIQUID PRODUCT
C3223259|T121|1169108|RXNORM|HEPTALAC ORAL LIQUID PRODUCT|HEPTALAC ORAL LIQUID PRODUCT
C3223942|T121|1169806|RXNORM|GENERLAC ORAL LIQUID PRODUCT|GENERLAC ORAL LIQUID PRODUCT
C3224342|T121|1170217|RXNORM|CHOLAC ORAL LIQUID PRODUCT|CHOLAC ORAL LIQUID PRODUCT
C3224366|T121|1170241|RXNORM|CHRONULAC ORAL LIQUID PRODUCT|CHRONULAC ORAL LIQUID PRODUCT
C3225241|T121|1171159|RXNORM|EVALOSE ORAL LIQUID PRODUCT|EVALOSE ORAL LIQUID PRODUCT
C3228268|T121||RXNORM|KRISTALOSE ORAL LIQUID PRODUCT
C3230348|T121|1176396|RXNORM|CATULAC ORAL LIQUID PRODUCT|CATULAC ORAL LIQUID PRODUCT
C3231581|T121|1177664|RXNORM|RO-LACTULOSE ORAL LIQUID PRODUCT|RO-LACTULOSE ORAL LIQUID PRODUCT
C1252332|T121|378092|RXNORM|LACTULOSE ORAL SOLUTION|LACTULOSE ORAL SOLUTION
C0787976|T121|247050|RXNORM|LACTULOSE 0.4 MG/MG ORAL GEL|LACTULOSE 0.4 MG/MG ORAL GEL
C1359419|T121|430151|RXNORM|LACTULOSE 2500 MG ORAL TABLET|LACTULOSE 2500 MG ORAL TABLET
C1363276|T121|434006|RXNORM|LACTULOSE 2865 MG CHEWABLE TABLET|LACTULOSE 2865 MG CHEWABLE TABLET
C3221022|T121|1166821|RXNORM|CEPHULAC ORAL PRODUCT|CEPHULAC ORAL PRODUCT
C3221217|T121|1167019|RXNORM|DUPHALAC ORAL PRODUCT|DUPHALAC ORAL PRODUCT
C3221249|T121|1167053|RXNORM|ENULOSE ORAL PRODUCT|ENULOSE ORAL PRODUCT
C3222921|T121|1168757|RXNORM|CONSTILAC ORAL PRODUCT|CONSTILAC ORAL PRODUCT
C3222923|T121|1168759|RXNORM|CONSTULOSE ORAL PRODUCT|CONSTULOSE ORAL PRODUCT
C3223260|T121|1169109|RXNORM|HEPTALAC ORAL PRODUCT|HEPTALAC ORAL PRODUCT
C3223943|T121|1169807|RXNORM|GENERLAC ORAL PRODUCT|GENERLAC ORAL PRODUCT
C3224343|T121|1170218|RXNORM|CHOLAC ORAL PRODUCT|CHOLAC ORAL PRODUCT
C3224367|T121|1170242|RXNORM|CHRONULAC ORAL PRODUCT|CHRONULAC ORAL PRODUCT
C3225242|T121|1171160|RXNORM|EVALOSE ORAL PRODUCT|EVALOSE ORAL PRODUCT
C3228269|T121|1174250|RXNORM|KRISTALOSE ORAL PRODUCT|KRISTALOSE ORAL PRODUCT
C3230349|T121|1176397|RXNORM|CATULAC ORAL PRODUCT|CATULAC ORAL PRODUCT
C3231582|T121|1177665|RXNORM|RO-LACTULOSE ORAL PRODUCT|RO-LACTULOSE ORAL PRODUCT
C1252272|T121|378034|RXNORM|LACTULOSE ORAL GEL|LACTULOSE ORAL GEL
C1370590|T121|440553|RXNORM|LACTULOSE ORAL TABLET|LACTULOSE ORAL TABLET
C1370592|T121|440555|RXNORM|LACTULOSE CHEWABLE TABLET|LACTULOSE CHEWABLE TABLET
C1620382|T121|1251192|RXNORM|LACTULOSE 10 GM/PACKET ORAL POWDER FOR SUSPENSION [KRISTALOSE]|KRISTALOSE 10000 MG POWDER FOR ORAL SOLUTION
C1620382|T121|1251192|RXNORM|KRISTALOSE 83.3 MG/ML ORAL SOLUTION|KRISTALOSE 10000 MG POWDER FOR ORAL SOLUTION
C1620382|T121|1251192|RXNORM|KRISTALOSE 10 GM PER 4 OZ. POWDER FOR ORAL SOLUTION|KRISTALOSE 10000 MG POWDER FOR ORAL SOLUTION
C1620382|T121|1251192|RXNORM|LACTULOSE 83.3 MG/ML ORAL SOLUTION [KRISTALOSE]|KRISTALOSE 10000 MG POWDER FOR ORAL SOLUTION
C1620382|T121|1251192|RXNORM|LACTULOSE 10 G IN 10 G ORAL POWDER, FOR SOLUTION [KRISTALOSE]|KRISTALOSE 10000 MG POWDER FOR ORAL SOLUTION
C1620382|T121|1251192|RXNORM|KRISTALOSE 10G POWDER FOR SOLUTION|KRISTALOSE 10000 MG POWDER FOR ORAL SOLUTION
C1620382|T121|1251192|RXNORM|KRISTALOSE, 10 G ORAL POWDER FOR RECONSTITUTION|KRISTALOSE 10000 MG POWDER FOR ORAL SOLUTION
C0708295|T121|755469|RXNORM|LACTULOSE 667 MG/ML ORAL SOLUTION [DUPHALAC]|DUPHALAC 10 GM PER 15 ML SYRUP
C0708295|T121|755469|RXNORM|DUPHALAC 667 MG/ML ORAL SOLUTION|DUPHALAC 10 GM PER 15 ML SYRUP
C0708295|T121|755469|RXNORM|DUPHALAC 10 GM PER 15 ML SYRUP|DUPHALAC 10 GM PER 15 ML SYRUP
C0708295|T121|755469|RXNORM|LACTULOSE 10 GM/15 ML ORAL SYRUP [DUPHALAC]|DUPHALAC 10 GM PER 15 ML SYRUP
C0708295|T121|755469|RXNORM|DUPHALAC, 10 G/15 ML ORAL SYRUP|DUPHALAC 10 GM PER 15 ML SYRUP
C1695496|T121|544459|RXNORM|LACTULOSE 667 MG/ML ORAL SOLUTION [RO-LACTULOSE]|RO-LACTULOSE 667 MG/ML ORAL SOLUTION
C1695496|T121|544459|RXNORM|RO-LACTULOSE 667 MG/ML ORAL SOLUTION|RO-LACTULOSE 667 MG/ML ORAL SOLUTION
C1586234|T121|755464|RXNORM|LACTULOSE 667 MG/ML ORAL SOLUTION [CATULAC]|CATULAC 667 MG/ML ORAL SOLUTION
C1586234|T121|755464|RXNORM|CATULAC 667 MG/ML ORAL SOLUTION|CATULAC 667 MG/ML ORAL SOLUTION
C0708290|T121|755465|RXNORM|CEPHULAC 10G/15ML SOLUTION|CEPHULAC 10 GM PER 15 ML SYRUP
C0708290|T121|755465|RXNORM|CEPHULAC 667 MG/ML ORAL SOLUTION|CEPHULAC 10 GM PER 15 ML SYRUP
C0708290|T121|755465|RXNORM|LACTULOSE 667 MG/ML ORAL SOLUTION [CEPHULAC]|CEPHULAC 10 GM PER 15 ML SYRUP
C0708290|T121|755465|RXNORM|CEPHULAC 10 GM PER 15 ML SYRUP|CEPHULAC 10 GM PER 15 ML SYRUP
C0708290|T121|755465|RXNORM|LACTULOSE 10 GM/15 ML ORAL SYRUP [CEPHULAC]|CEPHULAC 10 GM PER 15 ML SYRUP
C0708290|T121|755465|RXNORM|CEPHULAC, 10 G/15 ML ORAL SYRUP|CEPHULAC 10 GM PER 15 ML SYRUP
C0708291|T121|755466|RXNORM|CHOLAC 667 MG/ML ORAL SOLUTION|CHOLAC 10 GM PER 15 ML SYRUP
C0708291|T121|755466|RXNORM|LACTULOSE 667 MG/ML ORAL SOLUTION [CHOLAC]|CHOLAC 10 GM PER 15 ML SYRUP
C0708291|T121|755466|RXNORM|CHOLAC 10 GM PER 15 ML SYRUP|CHOLAC 10 GM PER 15 ML SYRUP
C0708291|T121|755466|RXNORM|LACTULOSE 10 GM/15 ML ORAL SYRUP [CHOLAC]|CHOLAC 10 GM PER 15 ML SYRUP
C0708291|T121|755466|RXNORM|CHOLAC 10G/15ML SOLUTION|CHOLAC 10 GM PER 15 ML SYRUP
C0708291|T121|755466|RXNORM|CHOLAC, 10 G/15 ML ORAL SYRUP|CHOLAC 10 GM PER 15 ML SYRUP
C0708292|T121|755467|RXNORM|CHRONULAC 10G/15ML SOLUTION|CHRONULAC 10 GM PER 15 ML SYRUP
C0708292|T121|755467|RXNORM|LACTULOSE 667 MG/ML ORAL SOLUTION [CHRONULAC]|CHRONULAC 10 GM PER 15 ML SYRUP
C0708292|T121|755467|RXNORM|CHRONULAC 667 MG/ML ORAL SOLUTION|CHRONULAC 10 GM PER 15 ML SYRUP
C0708292|T121|755467|RXNORM|CHRONULAC 10 GM PER 15 ML SYRUP|CHRONULAC 10 GM PER 15 ML SYRUP
C0708292|T121|755467|RXNORM|LACTULOSE 10 GM/15 ML ORAL SYRUP [CHRONULAC]|CHRONULAC 10 GM PER 15 ML SYRUP
C0708292|T121|755467|RXNORM|CHRONULAC, 10 G/15 ML ORAL SYRUP|CHRONULAC 10 GM PER 15 ML SYRUP
C0708293|T121|755468|RXNORM|LACTULOSE 667 MG/ML ORAL SOLUTION [CONSTILAC]|CONSTILAC 10 GM PER 15 ML SYRUP
C0708293|T121|755468|RXNORM|CONSTILAC 667 MG/ML ORAL SOLUTION|CONSTILAC 10 GM PER 15 ML SYRUP
C0708293|T121|755468|RXNORM|CONSTILAC 10 GM PER 15 ML SYRUP|CONSTILAC 10 GM PER 15 ML SYRUP
C0708293|T121|755468|RXNORM|LACTULOSE 10 GM/15 ML ORAL SYRUP [CONSTILAC]|CONSTILAC 10 GM PER 15 ML SYRUP
C0708293|T121|755468|RXNORM|CONSTILAC 10G/15ML SOLUTION|CONSTILAC 10 GM PER 15 ML SYRUP
C0708293|T121|755468|RXNORM|CONSTILAC, 10 G/15 ML ORAL SYRUP|CONSTILAC 10 GM PER 15 ML SYRUP
C0708297|T121|755471|RXNORM|EVALOSE 667 MG/ML ORAL SOLUTION|EVALOSE 10 GM PER 15 ML SYRUP
C0708297|T121|755471|RXNORM|LACTULOSE 667 MG/ML ORAL SOLUTION [EVALOSE]|EVALOSE 10 GM PER 15 ML SYRUP
C0708297|T121|755471|RXNORM|EVALOSE 10 GM PER 15 ML SYRUP|EVALOSE 10 GM PER 15 ML SYRUP
C0708297|T121|755471|RXNORM|LACTULOSE 10 GM/15 ML ORAL SYRUP [EVALOSE]|EVALOSE 10 GM PER 15 ML SYRUP
C0708297|T121|755471|RXNORM|EVALOSE, 10 G/15 ML ORAL SYRUP|EVALOSE 10 GM PER 15 ML SYRUP
C0708299|T121|755472|RXNORM|LACTULOSE 667 MG/ML ORAL SOLUTION [HEPTALAC]|HEPTALAC 667 MG/ML ORAL SOLUTION
C0708299|T121|755472|RXNORM|HEPTALAC 667 MG/ML ORAL SOLUTION|HEPTALAC 667 MG/ML ORAL SOLUTION
C0708299|T121|755472|RXNORM|LACTULOSE 10 GM/15 ML ORAL SOLUTION [HEPTALAC]|HEPTALAC 667 MG/ML ORAL SOLUTION
C0708299|T121|755472|RXNORM|LACTULOSE 10 GM/15 ML ORAL SYRUP [HEPTALAC]|HEPTALAC 667 MG/ML ORAL SOLUTION
C0708299|T121|755472|RXNORM|HEPTALAC, 10 G/15 ML ORAL SYRUP|HEPTALAC 667 MG/ML ORAL SOLUTION
C1613498|T121|1251196|RXNORM|LACTULOSE 20 GM/PACKET ORAL POWDER FOR SUSPENSION [KRISTALOSE]|KRISTALOSE 20 GM POWDER FOR ORAL SOLUTION
C1613498|T121|1251196|RXNORM|LACTULOSE 167 MG/ML ORAL SOLUTION [KRISTALOSE]|KRISTALOSE 20 GM POWDER FOR ORAL SOLUTION
C1613498|T121|1251196|RXNORM|KRISTALOSE 20 GM PER 4 OZ. POWDER FOR ORAL SOLUTION|KRISTALOSE 20 GM POWDER FOR ORAL SOLUTION
C1613498|T121|1251196|RXNORM|KRISTALOSE 167 MG/ML ORAL SOLUTION|KRISTALOSE 20 GM POWDER FOR ORAL SOLUTION
C1613498|T121|1251196|RXNORM|LACTULOSE 20 G IN 20 G ORAL POWDER, FOR SOLUTION [KRISTALOSE]|KRISTALOSE 20 GM POWDER FOR ORAL SOLUTION
C1613498|T121|1251196|RXNORM|KRISTALOSE 20G POWDER FOR SOLUTION|KRISTALOSE 20 GM POWDER FOR ORAL SOLUTION
C1613498|T121|1251196|RXNORM|KRISTALOSE, 20 G ORAL POWDER FOR RECONSTITUTION|KRISTALOSE 20 GM POWDER FOR ORAL SOLUTION
C0981135|T121|855288|RXNORM|WARFARIN SODIUM 1MG ORAL TABLET|WARFARIN SODIUM 1 MG ORAL TABLET
C0981135|T121|855288|RXNORM|WARFARIN SODIUM, 1 MG ORAL TABLET|WARFARIN SODIUM 1 MG ORAL TABLET
C0981135|T121|855288|RXNORM|WARFARIN 1 MG ORAL TABLET|WARFARIN SODIUM 1 MG ORAL TABLET
C0981135|T121|855288|RXNORM|WARFARIN (COUMADIN) NA 1MG TAB UD|WARFARIN SODIUM 1 MG ORAL TABLET
C0981135|T121|855288|RXNORM|WARFARIN (COUMADIN) NA 1MG TAB|WARFARIN SODIUM 1 MG ORAL TABLET
C0981135|T121|855288|RXNORM|WARFARIN SODIUM TAB 1 MG|WARFARIN SODIUM 1 MG ORAL TABLET
C0981135|T121|855288|RXNORM|WARFARIN SODIUM 1 MG ORAL TABLET|WARFARIN SODIUM 1 MG ORAL TABLET
C0981135|T121|855288|RXNORM|WARFARIN NA (GOLDEN STATE) 1MG TAB|WARFARIN SODIUM 1 MG ORAL TABLET
C0981135|T121|855288|RXNORM|WARFARIN NA 1MG TAB|WARFARIN SODIUM 1 MG ORAL TABLET
C0981135|T121|855288|RXNORM|WARFARIN NA (GOLDEN STATE) 1MG TAB [VA PRODUCT]|WARFARIN SODIUM 1 MG ORAL TABLET
C0981135|T121|855288|RXNORM|WARFARIN NA 1MG TAB,UD|WARFARIN SODIUM 1 MG ORAL TABLET
C0981135|T121|855288|RXNORM|WARFARIN NA 1MG TAB,UD [VA PRODUCT]|WARFARIN SODIUM 1 MG ORAL TABLET
C0981135|T121|855288|RXNORM|WARFARIN NA 1MG TAB [VA PRODUCT]|WARFARIN SODIUM 1 MG ORAL TABLET
C0981135|T121|855288|RXNORM|WARFARIN SODIUM 1 MG ORAL TABLET [WARFARIN SODIUM]|WARFARIN SODIUM 1 MG ORAL TABLET
C0981135|T121|855288|RXNORM|WARFARIN NA (EXELAN) 1MG TAB|WARFARIN SODIUM 1 MG ORAL TABLET
C0981135|T121|855288|RXNORM|WARFARIN NA (EXELAN) 1MG TAB [VA PRODUCT]|WARFARIN SODIUM 1 MG ORAL TABLET
C0981135|T121|855288|RXNORM|WARFARIN SODIUM 1MG TABLET|WARFARIN SODIUM 1 MG ORAL TABLET
C0981135|T121|855288|RXNORM|WARFARIN SODIUM 1MG TABLET |WARFARIN SODIUM 1 MG ORAL TABLET
C0981135|T121|855288|RXNORM|WARFARIN SODIUM 1MG TABLET |WARFARIN SODIUM 1 MG ORAL TABLET
C0690746|T121|855324|RXNORM|WARFARIN SODIUM 4MG ORAL TABLET|WARFARIN SODIUM 4 MG ORAL TABLET
C0690746|T121|855324|RXNORM|WARFARIN NA 4MG TAB,UD|WARFARIN SODIUM 4 MG ORAL TABLET
C0690746|T121|855324|RXNORM|WARFARIN SODIUM, 4 MG ORAL TABLET|WARFARIN SODIUM 4 MG ORAL TABLET
C0690746|T121|855324|RXNORM|WARFARIN 4 MG ORAL TABLET|WARFARIN SODIUM 4 MG ORAL TABLET
C0690746|T121|855324|RXNORM|WARFARIN (COUMADIN) NA 4MG TAB UD|WARFARIN SODIUM 4 MG ORAL TABLET
C0690746|T121|855324|RXNORM|WARFARIN (COUMADIN) NA 4MG TAB|WARFARIN SODIUM 4 MG ORAL TABLET
C0690746|T121|855324|RXNORM|WARFARIN SODIUM TAB 4 MG|WARFARIN SODIUM 4 MG ORAL TABLET
C0690746|T121|855324|RXNORM|WARFARIN SODIUM 4 MG ORAL TABLET|WARFARIN SODIUM 4 MG ORAL TABLET
C0690746|T121|855324|RXNORM|WARFARIN NA (GOLDEN STATE) 4MG TAB|WARFARIN SODIUM 4 MG ORAL TABLET
C0690746|T121|855324|RXNORM|WARFARIN NA 4MG TAB [VA PRODUCT]|WARFARIN SODIUM 4 MG ORAL TABLET
C0690746|T121|855324|RXNORM|WARFARIN NA (GOLDEN STATE) 4MG TAB [VA PRODUCT]|WARFARIN SODIUM 4 MG ORAL TABLET
C0690746|T121|855324|RXNORM|WARFARIN NA 4MG TAB|WARFARIN SODIUM 4 MG ORAL TABLET
C0690746|T121|855324|RXNORM|WARFARIN NA 4MG TAB,UD [VA PRODUCT]|WARFARIN SODIUM 4 MG ORAL TABLET
C0690746|T121|855324|RXNORM|WARFARIN SODIUM 4 MG ORAL TABLET [WARFARIN SODIUM]|WARFARIN SODIUM 4 MG ORAL TABLET
C0690746|T121|855324|RXNORM|WARFARIN NA (EXELAN) 4MG TAB|WARFARIN SODIUM 4 MG ORAL TABLET
C0690746|T121|855324|RXNORM|WARFARIN NA (EXELAN) 4MG TAB [VA PRODUCT]|WARFARIN SODIUM 4 MG ORAL TABLET
C0690746|T121|855324|RXNORM|WARFARIN SODIUM 4MG TABLET |WARFARIN SODIUM 4 MG ORAL TABLET
C0690746|T121|855324|RXNORM|WARFARIN SODIUM 4MG TABLET|WARFARIN SODIUM 4 MG ORAL TABLET
C0981139|T121|855308|RXNORM|WARFARIN 2MG/ML POWDER FOR INJECTION SOLUTION |WARFARIN SODIUM 2 MG/ML INJECTABLE SOLUTION
C0981139|T121|855308|RXNORM|WARFARIN 2MG/ML POWDER FOR INJECTION SOLUTION|WARFARIN SODIUM 2 MG/ML INJECTABLE SOLUTION
C0981139|T121|855308|RXNORM|WARFARIN 5 MG INTRAVENOUS POWDER FOR INJECTION|WARFARIN SODIUM 2 MG/ML INJECTABLE SOLUTION
C0981139|T121|855308|RXNORM|WARFARIN SODIUM 5MG/VIL INJ|WARFARIN SODIUM 2 MG/ML INJECTABLE SOLUTION
C0981139|T121|855308|RXNORM|WARFARIN SODIUM FOR INJ 5 MG|WARFARIN SODIUM 2 MG/ML INJECTABLE SOLUTION
C0981139|T121|855308|RXNORM|WARFARIN SODIUM 2 MG/ML INJECTABLE SOLUTION|WARFARIN SODIUM 2 MG/ML INJECTABLE SOLUTION
C0981139|T121|855308|RXNORM|WARFARIN NA 5MG/VIL INJ|WARFARIN SODIUM 2 MG/ML INJECTABLE SOLUTION
C0981139|T121|855308|RXNORM|WARFARIN NA 5MG/VIL INJ [VA PRODUCT]|WARFARIN SODIUM 2 MG/ML INJECTABLE SOLUTION
C0981139|T121|855308|RXNORM|WARFARIN 5MG LYOPHILISATE FOR SOLUTION FOR INJECTION|WARFARIN SODIUM 2 MG/ML INJECTABLE SOLUTION
C0981139|T121|855308|RXNORM|WARFARIN SODIUM 5 MG INTRAVENOUS POWDER FOR SOLUTION|WARFARIN SODIUM 2 MG/ML INJECTABLE SOLUTION
C0981141|T121|855344|RXNORM|WARFARIN SODIUM 7.5MG ORAL TABLET|WARFARIN SODIUM 7.5 MG ORAL TABLET
C0981141|T121|855344|RXNORM|WARFARIN SODIUM, 7.5 MG ORAL TABLET|WARFARIN SODIUM 7.5 MG ORAL TABLET
C0981141|T121|855344|RXNORM|WARFARIN 7.5 MG ORAL TABLET|WARFARIN SODIUM 7.5 MG ORAL TABLET
C0981141|T121|855344|RXNORM|WARFARIN (COUMADIN) NA 7.5MG TAB|WARFARIN SODIUM 7.5 MG ORAL TABLET
C0981141|T121|855344|RXNORM|WARFARIN (COUMADIN) NA 7.5MG TAB UD|WARFARIN SODIUM 7.5 MG ORAL TABLET
C0981141|T121|855344|RXNORM|WARFARIN SODIUM TAB 7.5 MG|WARFARIN SODIUM 7.5 MG ORAL TABLET
C0981141|T121|855344|RXNORM|WARFARIN SODIUM 7.5 MG ORAL TABLET|WARFARIN SODIUM 7.5 MG ORAL TABLET
C0981141|T121|855344|RXNORM|WARFARIN NA (GOLDEN STATE) 7.5MG TAB|WARFARIN SODIUM 7.5 MG ORAL TABLET
C0981141|T121|855344|RXNORM|WARFARIN NA 7.5MG TAB,UD [VA PRODUCT]|WARFARIN SODIUM 7.5 MG ORAL TABLET
C0981141|T121|855344|RXNORM|WARFARIN SODIUM 7.5 MG ORAL TABLET [WARFARIN SODIUM]|WARFARIN SODIUM 7.5 MG ORAL TABLET
C0981141|T121|855344|RXNORM|WARFARIN NA (GOLDEN STATE) 7.5MG TAB [VA PRODUCT]|WARFARIN SODIUM 7.5 MG ORAL TABLET
C0981141|T121|855344|RXNORM|WARFARIN NA 7.5MG TAB,UD|WARFARIN SODIUM 7.5 MG ORAL TABLET
C0981141|T121|855344|RXNORM|WARFARIN NA 7.5MG TAB [VA PRODUCT]|WARFARIN SODIUM 7.5 MG ORAL TABLET
C0981141|T121|855344|RXNORM|WARFARIN NA 7.5MG TAB|WARFARIN SODIUM 7.5 MG ORAL TABLET
C0981141|T121|855344|RXNORM|WARFARIN NA (EXELAN) 7.5MG TAB|WARFARIN SODIUM 7.5 MG ORAL TABLET
C0981141|T121|855344|RXNORM|WARFARIN NA (EXELAN) 7.5MG TAB [VA PRODUCT]|WARFARIN SODIUM 7.5 MG ORAL TABLET
C0981141|T121|855344|RXNORM|WARFARIN SODIUM 7.5MG TABLET |WARFARIN SODIUM 7.5 MG ORAL TABLET
C0981141|T121|855344|RXNORM|WARFARIN SODIUM 7.5MG TABLET|WARFARIN SODIUM 7.5 MG ORAL TABLET
C0981794|T121|855318|RXNORM|WARFARIN SODIUM 3MG ORAL TABLET|WARFARIN SODIUM 3 MG ORAL TABLET
C0981794|T121|855318|RXNORM|WARFARIN SODIUM, 3 MG ORAL TABLET|WARFARIN SODIUM 3 MG ORAL TABLET
C0981794|T121|855318|RXNORM|WARFARIN 3 MG ORAL TABLET|WARFARIN SODIUM 3 MG ORAL TABLET
C0981794|T121|855318|RXNORM|WARFARIN (COUMADIN) NA 3MG TAB|WARFARIN SODIUM 3 MG ORAL TABLET
C0981794|T121|855318|RXNORM|WARFARIN (COUMADIN) NA 3MG TAB UD|WARFARIN SODIUM 3 MG ORAL TABLET
C0981794|T121|855318|RXNORM|WARFARIN SODIUM TAB 3 MG|WARFARIN SODIUM 3 MG ORAL TABLET
C0981794|T121|855318|RXNORM|WARFARIN SODIUM 3 MG ORAL TABLET|WARFARIN SODIUM 3 MG ORAL TABLET
C0981794|T121|855318|RXNORM|WARFARIN NA (GOLDEN STATE) 3MG TAB|WARFARIN SODIUM 3 MG ORAL TABLET
C0981794|T121|855318|RXNORM|WARFARIN NA (GOLDEN STATE) 3MG TAB [VA PRODUCT]|WARFARIN SODIUM 3 MG ORAL TABLET
C0981794|T121|855318|RXNORM|WARFARIN NA 3MG TAB [VA PRODUCT]|WARFARIN SODIUM 3 MG ORAL TABLET
C0981794|T121|855318|RXNORM|WARFARIN NA 3MG TAB,UD|WARFARIN SODIUM 3 MG ORAL TABLET
C0981794|T121|855318|RXNORM|WARFARIN SODIUM 3 MG ORAL TABLET [WARFARIN SODIUM]|WARFARIN SODIUM 3 MG ORAL TABLET
C0981794|T121|855318|RXNORM|WARFARIN NA 3MG TAB|WARFARIN SODIUM 3 MG ORAL TABLET
C0981794|T121|855318|RXNORM|WARFARIN NA 3MG TAB,UD [VA PRODUCT]|WARFARIN SODIUM 3 MG ORAL TABLET
C0981794|T121|855318|RXNORM|WARFARIN NA (EXELAN) 3MG TAB|WARFARIN SODIUM 3 MG ORAL TABLET
C0981794|T121|855318|RXNORM|WARFARIN NA (EXELAN) 3MG TAB [VA PRODUCT]|WARFARIN SODIUM 3 MG ORAL TABLET
C0981794|T121|855318|RXNORM|WARFARIN SODIUM 3MG TABLET|WARFARIN SODIUM 3 MG ORAL TABLET
C0981794|T121|855318|RXNORM|WARFARIN SODIUM 3MG TABLET |WARFARIN SODIUM 3 MG ORAL TABLET
C0981794|T121|855318|RXNORM|WARFARIN SODIUM 3MG TABLET |WARFARIN SODIUM 3 MG ORAL TABLET
C0981140|T121|855338|RXNORM|WARFARIN SODIUM 6MG ORAL TABLET|WARFARIN SODIUM 6 MG ORAL TABLET
C0981140|T121|855338|RXNORM|WARFARIN SODIUM, 6 MG ORAL TABLET|WARFARIN SODIUM 6 MG ORAL TABLET
C0981140|T121|855338|RXNORM|WARFARIN 6 MG ORAL TABLET|WARFARIN SODIUM 6 MG ORAL TABLET
C0981140|T121|855338|RXNORM|WARFARIN (COUMADIN) NA 6MG TAB|WARFARIN SODIUM 6 MG ORAL TABLET
C0981140|T121|855338|RXNORM|WARFARIN (COUMADIN) NA 6MG TAB UD|WARFARIN SODIUM 6 MG ORAL TABLET
C0981140|T121|855338|RXNORM|WARFARIN SODIUM TAB 6 MG|WARFARIN SODIUM 6 MG ORAL TABLET
C0981140|T121|855338|RXNORM|WARFARIN SODIUM 6 MG ORAL TABLET|WARFARIN SODIUM 6 MG ORAL TABLET
C0981140|T121|855338|RXNORM|WARFARIN NA (GOLDEN STATE) 6MG TAB|WARFARIN SODIUM 6 MG ORAL TABLET
C0981140|T121|855338|RXNORM|WARFARIN NA (GOLDEN STATE) 6MG TAB [VA PRODUCT]|WARFARIN SODIUM 6 MG ORAL TABLET
C0981140|T121|855338|RXNORM|WARFARIN NA 6MG TAB|WARFARIN SODIUM 6 MG ORAL TABLET
C0981140|T121|855338|RXNORM|WARFARIN NA 6MG TAB,UD [VA PRODUCT]|WARFARIN SODIUM 6 MG ORAL TABLET
C0981140|T121|855338|RXNORM|WARFARIN NA 6MG TAB [VA PRODUCT]|WARFARIN SODIUM 6 MG ORAL TABLET
C0981140|T121|855338|RXNORM|WARFARIN NA 6MG TAB,UD|WARFARIN SODIUM 6 MG ORAL TABLET
C0981140|T121|855338|RXNORM|WARFARIN SODIUM 6 MG ORAL TABLET [WARFARIN SODIUM]|WARFARIN SODIUM 6 MG ORAL TABLET
C0981140|T121|855338|RXNORM|WARFARIN NA (EXELAN) 6MG TAB|WARFARIN SODIUM 6 MG ORAL TABLET
C0981140|T121|855338|RXNORM|WARFARIN NA (EXELAN) 6MG TAB [VA PRODUCT]|WARFARIN SODIUM 6 MG ORAL TABLET
C0981140|T121|855338|RXNORM|WARFARIN SODIUM 6MG TABLET |WARFARIN SODIUM 6 MG ORAL TABLET
C0981140|T121|855338|RXNORM|WARFARIN SODIUM 6MG TABLET|WARFARIN SODIUM 6 MG ORAL TABLET
C0981793|T121|855332|RXNORM|WARFARIN SODIUM 5MG ORAL TABLET|WARFARIN SODIUM 5 MG ORAL TABLET
C0981793|T121|855332|RXNORM|WARFARIN SODIUM, 5 MG ORAL TABLET|WARFARIN SODIUM 5 MG ORAL TABLET
C0981793|T121|855332|RXNORM|WARFARIN 5 MG ORAL TABLET|WARFARIN SODIUM 5 MG ORAL TABLET
C0981793|T121|855332|RXNORM|WARFARIN (COUMADIN) NA 5MG TAB UD|WARFARIN SODIUM 5 MG ORAL TABLET
C0981793|T121|855332|RXNORM|WARFARIN (COUMADIN) NA 5MG TAB|WARFARIN SODIUM 5 MG ORAL TABLET
C0981793|T121|855332|RXNORM|WARFARIN SODIUM TAB 5 MG|WARFARIN SODIUM 5 MG ORAL TABLET
C0981793|T121|855332|RXNORM|WARFARIN SODIUM 5 MG ORAL TABLET|WARFARIN SODIUM 5 MG ORAL TABLET
C0981793|T121|855332|RXNORM|WARFARIN NA (GOLDEN STATE) 5MG TAB|WARFARIN SODIUM 5 MG ORAL TABLET
C0981793|T121|855332|RXNORM|WARFARIN NA 5MG TAB,UD|WARFARIN SODIUM 5 MG ORAL TABLET
C0981793|T121|855332|RXNORM|WARFARIN NA 5MG TAB,UD [VA PRODUCT]|WARFARIN SODIUM 5 MG ORAL TABLET
C0981793|T121|855332|RXNORM|WARFARIN SODIUM 5 MG ORAL TABLET [WARFARIN SODIUM]|WARFARIN SODIUM 5 MG ORAL TABLET
C0981793|T121|855332|RXNORM|WARFARIN NA 5MG TAB|WARFARIN SODIUM 5 MG ORAL TABLET
C0981793|T121|855332|RXNORM|WARFARIN NA (GOLDEN STATE) 5MG TAB [VA PRODUCT]|WARFARIN SODIUM 5 MG ORAL TABLET
C0981793|T121|855332|RXNORM|WARFARIN NA 5MG TAB [VA PRODUCT]|WARFARIN SODIUM 5 MG ORAL TABLET
C0981793|T121|855332|RXNORM|WARFARIN NA (EXELAN) 5MG TAB|WARFARIN SODIUM 5 MG ORAL TABLET
C0981793|T121|855332|RXNORM|WARFARIN NA (EXELAN) 5MG TAB [VA PRODUCT]|WARFARIN SODIUM 5 MG ORAL TABLET
C0981793|T121|855332|RXNORM|WARFARIN SODIUM 5MG TABLET|WARFARIN SODIUM 5 MG ORAL TABLET
C0981793|T121|855332|RXNORM|WARFARIN SODIUM 5MG TABLET |WARFARIN SODIUM 5 MG ORAL TABLET
C0981793|T121|855332|RXNORM|WARFARIN SODIUM 5MG TABLET |WARFARIN SODIUM 5 MG ORAL TABLET
C0917972|T121||RXNORM|ATHROMBIN-K
C0981136|T121|855312|RXNORM|WARFARIN SODIUM 2.5MG ORAL TABLET|WARFARIN SODIUM 2.5 MG ORAL TABLET
C0981136|T121|855312|RXNORM|WARFARIN SODIUM, 2.5 MG ORAL TABLET|WARFARIN SODIUM 2.5 MG ORAL TABLET
C0981136|T121|855312|RXNORM|WARFARIN 2.5 MG ORAL TABLET|WARFARIN SODIUM 2.5 MG ORAL TABLET
C0981136|T121|855312|RXNORM|WARFARIN (COUMADIN) NA 2.5MG TAB|WARFARIN SODIUM 2.5 MG ORAL TABLET
C0981136|T121|855312|RXNORM|WARFARIN (COUMADIN) NA 2.5MG TAB UD|WARFARIN SODIUM 2.5 MG ORAL TABLET
C0981136|T121|855312|RXNORM|WARFARIN SODIUM TAB 2.5 MG|WARFARIN SODIUM 2.5 MG ORAL TABLET
C0981136|T121|855312|RXNORM|WARFARIN SODIUM 2.5 MG ORAL TABLET|WARFARIN SODIUM 2.5 MG ORAL TABLET
C0981136|T121|855312|RXNORM|WARFARIN NA (GOLDEN STATE) 2.5MG TAB|WARFARIN SODIUM 2.5 MG ORAL TABLET
C0981136|T121|855312|RXNORM|WARFARIN NA 2.5MG TAB,UD|WARFARIN SODIUM 2.5 MG ORAL TABLET
C0981136|T121|855312|RXNORM|WARFARIN NA 2.5MG TAB,UD [VA PRODUCT]|WARFARIN SODIUM 2.5 MG ORAL TABLET
C0981136|T121|855312|RXNORM|WARFARIN SODIUM 2.5 MG ORAL TABLET [WARFARIN SODIUM]|WARFARIN SODIUM 2.5 MG ORAL TABLET
C0981136|T121|855312|RXNORM|WARFARIN NA (GOLDEN STATE) 2.5MG TAB [VA PRODUCT]|WARFARIN SODIUM 2.5 MG ORAL TABLET
C0981136|T121|855312|RXNORM|WARFARIN NA 2.5MG TAB [VA PRODUCT]|WARFARIN SODIUM 2.5 MG ORAL TABLET
C0981136|T121|855312|RXNORM|WARFARIN NA 2.5MG TAB|WARFARIN SODIUM 2.5 MG ORAL TABLET
C0981136|T121|855312|RXNORM|WARFARIN NA (EXELAN) 2.5MG TAB [VA PRODUCT]|WARFARIN SODIUM 2.5 MG ORAL TABLET
C0981136|T121|855312|RXNORM|WARFARIN NA (EXELAN) 2.5MG TAB|WARFARIN SODIUM 2.5 MG ORAL TABLET
C0981136|T121|855312|RXNORM|WARFARIN SODIUM 2.5MG TABLET |WARFARIN SODIUM 2.5 MG ORAL TABLET
C0981136|T121|855312|RXNORM|WARFARIN SODIUM 2.5MG TABLET|WARFARIN SODIUM 2.5 MG ORAL TABLET
C0043031|T121|11289|RXNORM|WARFARIN|WARFARIN
C0043031|T121|11289|RXNORM|2H-1-BENZOPYRAN-2-ONE, 4-HYDROXY-3-(3-OXO-1-PHENYLBUTYL)-|WARFARIN
C0043031|T121|11289|RXNORM|4-HYDROXY-3-(3-OXO-1-PHENYLBUTYL)-2H-1-BENZOPYRAN-2-ONE|WARFARIN
C0043031|T121|11289|RXNORM|3-(ALPHA-ACETONYLBENZYL)-4-HYDROXYCOUMARIN|WARFARIN
C0043031|T121|11289|RXNORM|3-ALPHA-PHENYL-BETA-ACETYLETHYL-4-HYDROXYCOUMARIN|WARFARIN
C0043031|T121|11289|RXNORM|1-(4'-HYDROXY-3'-COUMARINYL)-1-PHENYL-3-BUTANONE|WARFARIN
C0043031|T121|11289|RXNORM|WARFARIN [CHEMICAL/INGREDIENT]|WARFARIN
C0043031|T121|11289|RXNORM|3-(.ALPHA.-ACETONYLBENZYL)-4-HYDROXYCOUMARIN|WARFARIN
C0043031|T121|11289|RXNORM|3-(.ALPHA.-PHENYL-.BETA.-ACETYLETHYL)-4-HYDROXYCOUMARIN|WARFARIN
C0043031|T121|11289|RXNORM|WARFARIN |WARFARIN
C0043031|T121|11289|RXNORM|ANTICOAGULANTS WARFARIN|WARFARIN
C0043031|T121|11289|RXNORM|WARFARIN |WARFARIN
C0043031|T121|11289|RXNORM|WARFARIN |WARFARIN
C0043031|T121|11289|RXNORM|WARF|WARFARIN
C0981134|T121|855296|RXNORM|WARFARIN SODIUM 10MG ORAL TABLET|WARFARIN SODIUM 10 MG ORAL TABLET
C0981134|T121|855296|RXNORM|WARFARIN SODIUM, 10 MG ORAL TABLET|WARFARIN SODIUM 10 MG ORAL TABLET
C0981134|T121|855296|RXNORM|WARFARIN 10 MG ORAL TABLET|WARFARIN SODIUM 10 MG ORAL TABLET
C0981134|T121|855296|RXNORM|WARFARIN (COUMADIN) NA 10MG TAB|WARFARIN SODIUM 10 MG ORAL TABLET
C0981134|T121|855296|RXNORM|WARFARIN (COUMADIN) NA 10MG TAB UD|WARFARIN SODIUM 10 MG ORAL TABLET
C0981134|T121|855296|RXNORM|WARFARIN SODIUM TAB 10 MG|WARFARIN SODIUM 10 MG ORAL TABLET
C0981134|T121|855296|RXNORM|WARFARIN SODIUM 10 MG ORAL TABLET|WARFARIN SODIUM 10 MG ORAL TABLET
C0981134|T121|855296|RXNORM|WARFARIN NA (GOLDEN STATE) 10MG TAB|WARFARIN SODIUM 10 MG ORAL TABLET
C0981134|T121|855296|RXNORM|WARFARIN NA 10MG TAB,UD|WARFARIN SODIUM 10 MG ORAL TABLET
C0981134|T121|855296|RXNORM|WARFARIN NA 10MG TAB|WARFARIN SODIUM 10 MG ORAL TABLET
C0981134|T121|855296|RXNORM|WARFARIN NA 10MG TAB,UD [VA PRODUCT]|WARFARIN SODIUM 10 MG ORAL TABLET
C0981134|T121|855296|RXNORM|WARFARIN SODIUM 10 MG ORAL TABLET [WARFARIN SODIUM]|WARFARIN SODIUM 10 MG ORAL TABLET
C0981134|T121|855296|RXNORM|WARFARIN NA 10MG TAB [VA PRODUCT]|WARFARIN SODIUM 10 MG ORAL TABLET
C0981134|T121|855296|RXNORM|WARFARIN NA (GOLDEN STATE) 10MG TAB [VA PRODUCT]|WARFARIN SODIUM 10 MG ORAL TABLET
C0981134|T121|855296|RXNORM|WARFARIN SODIUM 10 MG ORAL TABLET [PANWARFIN]|WARFARIN SODIUM 10 MG ORAL TABLET
C0981134|T121|855296|RXNORM|WARFARIN NA (EXELAN) 10MG TAB|WARFARIN SODIUM 10 MG ORAL TABLET
C0981134|T121|855296|RXNORM|WARFARIN NA (EXELAN) 10MG TAB [VA PRODUCT]|WARFARIN SODIUM 10 MG ORAL TABLET
C0981134|T121|855296|RXNORM|WARFARIN SODIUM 10MG TABLET |WARFARIN SODIUM 10 MG ORAL TABLET
C0981134|T121|855296|RXNORM|WARFARIN SODIUM 10MG TABLET|WARFARIN SODIUM 10 MG ORAL TABLET
C1584930|T121|855302|RXNORM|WARFARIN SODIUM 2MG ORAL TABLET|WARFARIN SODIUM 2 MG ORAL TABLET
C1584930|T121|855302|RXNORM|WARFARIN SODIUM, 2 MG ORAL TABLET|WARFARIN SODIUM 2 MG ORAL TABLET
C1584930|T121|855302|RXNORM|WARFARIN 2 MG ORAL TABLET|WARFARIN SODIUM 2 MG ORAL TABLET
C1584930|T121|855302|RXNORM|WARFARIN (COUMADIN) NA 2MG TAB|WARFARIN SODIUM 2 MG ORAL TABLET
C1584930|T121|855302|RXNORM|WARFARIN (COUMADIN) NA 2MG TAB UD|WARFARIN SODIUM 2 MG ORAL TABLET
C1584930|T121|855302|RXNORM|WARFARIN SODIUM TAB 2 MG|WARFARIN SODIUM 2 MG ORAL TABLET
C1584930|T121|855302|RXNORM|WARFARIN SODIUM 2 MG ORAL TABLET|WARFARIN SODIUM 2 MG ORAL TABLET
C1584930|T121|855302|RXNORM|WARFARIN NA (GOLDEN STATE) 2MG TAB|WARFARIN SODIUM 2 MG ORAL TABLET
C1584930|T121|855302|RXNORM|WARFARIN NA 2MG TAB [VA PRODUCT]|WARFARIN SODIUM 2 MG ORAL TABLET
C1584930|T121|855302|RXNORM|WARFARIN NA 2MG TAB|WARFARIN SODIUM 2 MG ORAL TABLET
C1584930|T121|855302|RXNORM|WARFARIN SODIUM 2 MG ORAL TABLET [WARFARIN SODIUM]|WARFARIN SODIUM 2 MG ORAL TABLET
C1584930|T121|855302|RXNORM|WARFARIN NA 2MG TAB,UD|WARFARIN SODIUM 2 MG ORAL TABLET
C1584930|T121|855302|RXNORM|WARFARIN NA (GOLDEN STATE) 2MG TAB [VA PRODUCT]|WARFARIN SODIUM 2 MG ORAL TABLET
C1584930|T121|855302|RXNORM|WARFARIN NA 2MG TAB,UD [VA PRODUCT]|WARFARIN SODIUM 2 MG ORAL TABLET
C1584930|T121|855302|RXNORM|WARFARIN NA (EXELAN) 2MG TAB|WARFARIN SODIUM 2 MG ORAL TABLET
C1584930|T121|855302|RXNORM|WARFARIN NA (EXELAN) 2MG TAB [VA PRODUCT]|WARFARIN SODIUM 2 MG ORAL TABLET
C1584930|T121|855302|RXNORM|WARFARIN SODIUM 2MG TABLET |WARFARIN SODIUM 2 MG ORAL TABLET
C1584930|T121|855302|RXNORM|WARFARIN SODIUM 2MG TABLET|WARFARIN SODIUM 2 MG ORAL TABLET
C1584930|T121|855302|RXNORM|WARFAREN SODIUM 2MG TABLET USP|WARFARIN SODIUM 2 MG ORAL TABLET
C0376218|T121|114194|RXNORM|SODIUM, WARFARIN|WARFARIN SODIUM
C0376218|T121|114194|RXNORM|WARFARIN SODIUM|WARFARIN SODIUM
C0376218|T121|114194|RXNORM|WARFARIN SODIUM |WARFARIN SODIUM
C0376218|T121|114194|RXNORM|WARFARIN SODIUM [CHEMICAL/INGREDIENT]|WARFARIN SODIUM
C0376218|T121|114194|RXNORM|WARFARIN SODIUM |WARFARIN SODIUM
C0376218|T121|114194|RXNORM|PROTHROMADIN|WARFARIN SODIUM
C0376218|T121|114194|RXNORM|SODIUM WARFARIN|WARFARIN SODIUM
C0376218|T121|114194|RXNORM|TINTORANE|WARFARIN SODIUM
C1572765|T121||RXNORM|WARFARIN SODIUM ISOPROPANOL COMPLEX
C1601608|T121|540210|RXNORM|WARFIN|WARFIN
C0163698|T121||RXNORM|2H-1-BENZOPYRAN-2-ONE, 3-(1-(4-AZIDOPHENYL)-3-OXOBUTYL)-4-HYDROXY-
C0163698|T121||RXNORM|AZIDOWARFARIN
C0298589|T121||RXNORM|WARFARIN HEXADECYL ETHER
C0265374|T121||RXNORM|DYSMORPHISM DUE TO WARFARIN
C0265374|T121||RXNORM|FOETAL WARFARIN SYNDROME
C0265374|T121||RXNORM|CONGENITAL WARFARIN SYNDROME
C0265374|T121||RXNORM|WARFARIN SYNDROME
C0265374|T121||RXNORM|FETAL ANTICOAGULANT SYNDROME
C0265374|T121||RXNORM|COUMARIN SYNDROME
C0265374|T121||RXNORM|WARFARIN EMBRYOPATHY
C0265374|T121||RXNORM|DISALA SYNDROME
C0265374|T121||RXNORM|FETAL WARFARIN SYNDROME
C0265374|T121||RXNORM|FETAL WARFARIN SYNDROME 
C0265374|T121||RXNORM|FETAL COUMADIN SYNDROME
C0265374|T121||RXNORM|DYSMORPHISM; WARFARIN
C0265374|T121||RXNORM|WARFARIN; DYSMORPHISM
C0282378|T121|82118|RXNORM|POTASSIUM, WARFARIN|WARFARIN POTASSIUM
C0282378|T121|82118|RXNORM|WARFARIN POTASSIUM|WARFARIN POTASSIUM
C0282378|T121|82118|RXNORM|WARFARIN POTASSIUM (DISCONTINUED) |WARFARIN POTASSIUM
C0282378|T121|82118|RXNORM|WARFARIN POTASSIUM (DISCONTINUED)|WARFARIN POTASSIUM
C0282378|T121|82118|RXNORM|POTASSIUM WARFARIN|WARFARIN POTASSIUM
C0282378|T121|82118|RXNORM|POTASSIUM WARFARIN |WARFARIN POTASSIUM
C0588999|T121||RXNORM|WARFARIN - RODENTICIDE
C0588999|T121||RXNORM|WARFARIN - RODENTICIDE 
C1975542|T121||RXNORM|WARFARIN &#X7C; URINE
C2966895|T121||RXNORM|WARFARIN &#X7C; XXX
C0366686|T121||RXNORM|WARFARIN:MASS:PT:DOSE:QN
C0366686|T121||RXNORM|WARFARIN [MASS] OF DOSE
C0366686|T121||RXNORM|WARFARIN DOSE
C0366686|T121||RXNORM|WARFARIN:MASS:POINT IN TIME:DOSE MED OR SUBSTANCE:QUANTITATIVE
C1975540|T121||RXNORM|WARFARIN &#X7C; BLD-SER-PLAS
C1975541|T121||RXNORM|WARFARIN &#X7C; GASTRIC FLUID
C0647187|T121||RXNORM|3'-HYDROXYWARFARIN
C0648649|T121||RXNORM|N-ACETYL-GAMMA-GLUTAMYL-4'-AMINOWARFARIN
C0648649|T121||RXNORM|AGAW
C0049626|T121||RXNORM|4,6-DIHYDROXY-3-(3-OXO-1-PHENYLBUTYL)-2H-1- BENZOPYRAN-2-ONE
C0049626|T121||RXNORM|6-HYDROXYWARFARIN
C0639160|T121||RXNORM|6-METHYL-6,12-METHANO-6H,12H,13H-BENZOPYRAN(4,3-D)BENZODIOXOCIN-13-ONE
C0639160|T121||RXNORM|MMBBD
C0207897|T121||RXNORM|4'-AMINOWARFARIN
C0207897|T121||RXNORM|3-(1-(4-AMINOPHENYL)-3-OXOBUTYL)-4-HYDROXY-2H-1-BENZOPYRAN-2-ONE
C0529816|T121||RXNORM|8-HYDROXYWARFARIN
C0637401|T121||RXNORM|4-HYDROXY-3-(1-(4-HYDROXYPHENYL)-3-OXOBUTYL)-2H-1-BENZOPYRAN-2-ONE
C0637401|T121||RXNORM|4'-HYDROXYWARFARIN
C2363289|T121||RXNORM|COUMAFURYL
C2363289|T121||RXNORM|COUMAFURYL 
C2363289|T121||RXNORM|COUMAFURYL 
C0627500|T121||RXNORM|MS-WARFARIN
C0627500|T121||RXNORM|METHYLSULFINYLWARFARIN
C0642757|T121||RXNORM|4-HYDROXY-3-(2-HYDROXY-3-OXO-1-PHENYLBUTYL)-2H-1-BENZOPYRAN-2-ONE
C0642757|T121||RXNORM|10-HYDROXYWARFARIN
C0255975|T121||RXNORM|7-HYDROXYWARFARIN
C0255975|T121||RXNORM|2H-1-BENZOPYRAN-2-ONE, 4,7-DIHYDROXY-3-(3-OXO-1-PHENYLBUTYL)-
C1276897|T121|855350|RXNORM|WARFARIN SODIUM 0.5 MG ORAL TABLET|WARFARIN SODIUM 0.5 MG ORAL TABLET
C1276897|T121|855350|RXNORM|WARFARIN SODIUM 0.5MG TABLET |WARFARIN SODIUM 0.5 MG ORAL TABLET
C1276897|T121|855350|RXNORM|WARFARIN SODIUM 0.5MG TABLET|WARFARIN SODIUM 0.5 MG ORAL TABLET
C1276897|T121|855350|RXNORM|WARFARIN SODIUM 0.5MG TABLET |WARFARIN SODIUM 0.5 MG ORAL TABLET
C1527323|T121||RXNORM|RODEX
C1527323|T121||RXNORM|RODEX BRAND OF WARFARIN
C1520121|T121||RXNORM|CO-RAX
C1520122|T121||RXNORM|COMPOUND 42
C1520123|T121||RXNORM|WARF COMPOUND 42
C0699129|T121|202421|RXNORM|COUMADIN|COUMADIN
C0699129|T121|202421|RXNORM|MAREVAN|COUMADIN
C0699129|T121|202421|RXNORM|BRISTOL-MYERS SQUIBB BRAND OF WARFARIN SODIUM|COUMADIN
C0699129|T121|202421|RXNORM|GOLDSHIELD BRAND OF WARFARIN SODIUM|COUMADIN
C0699129|T121|202421|RXNORM|BOOTS BRAND OF WARFARIN SODIUM|COUMADIN
C1564392|T121||RXNORM|GENPHARM BRAND OF WARFARIN SODIUM
C1564392|T121||RXNORM|GEN-WARFARIN
C1564393|T121||RXNORM|ALDO BRAND OF WARFARIN SODIUM
C1564393|T121||RXNORM|ALDOCUMAR
C1564394|T121||RXNORM|COUMADINE
C1564394|T121||RXNORM|BAILLY BRAND OF WARFARIN SODIUM
C1564395|T121||RXNORM|APO-WARFARIN
C1564395|T121||RXNORM|APOTEX BRAND OF WARFARIN SODIUM
C1564396|T121||RXNORM|ESTEDI BRAND OF WARFARIN SODIUM
C1564396|T121||RXNORM|TEDICUMAR
C1564397|T121||RXNORM|WARFANT
C1564397|T121||RXNORM|ANTIGEN BRAND OF WARFARIN SODIUM
C1330361|T121|405155|RXNORM|JANTOVEN|JANTOVEN
C1601605|T121|540205|RXNORM|NARFARIN|NARFARIN
C1601620|T121|540226|RXNORM|MARFARIN|MARFARIN
C0605881|T121||RXNORM|ACTOSIN P
C0605881|T121||RXNORM|PINDONE, WARFARIN DRUG COMBINATION
C0605881|T121||RXNORM|PINDONE - WARFARIN
C0699130|T121||RXNORM|PANWARFIN
C1996947|T121||RXNORM|PARENTERAL FORM WARFARIN
C1996947|T121||RXNORM|PARENTERAL FORM WARFARIN 
C1998178|T121||RXNORM|ORAL FORM WARFARIN
C1998178|T121||RXNORM|ORAL FORM WARFARIN 
