C0010294|T034|LP14355-9|LNC|CREATININE|CREATININE
C0201975|T034||LNC|CREATININE
C1561535|T034||LNC|CREATININE
C0201975|T034||LNC|CREATININE MEASUREMENT
C0239150|T034||LNC|INTERPERTATION
C0428279|T034||LNC|FINDING OF CREATININE LEVEL
C0428279|T034||LNC|CREATININE LEVEL
C0428279|T034||LNC|CREATININE LEVEL IN BLOOD
C0555149|T034||LNC|CREATININE IN SAMPLE 
C0742904|T034||LNC|CREATININE RISING
C0201975|T034||LNC|CREATININE MEASUREMENT
C0201976|T034||LNC|CREATININE MEASUREMENT, SERUM 
C0236408|T034||LNC|CHEM-7 CREATININE MEASUREMENT
C0010294|T034|LP14355-9|LNC|CREATININE|CREATININE
C0010294|T034|LP14355-9|LNC|CREATININE [CHEMICAL/INGREDIENT]|CREATININE
C0010294|T034|LP14355-9|LNC|CREATININE |CREATININE
C0201976|T034||LNC|SERUM CREATININE
C0201976|T034||LNC|SERUM CREATININE MEASUREMENT
C0201976|T034||LNC|CREATININE MEASUREMENT, SERUM 
C0201976|T034||LNC|SERUM CREATININE LEVEL
C0201976|T034||LNC|SERUM CREATININE MEASUREMENT 
C0201976|T034||LNC|CREATININE.SERUM
C0201976|T034||LNC|SERUM CREATININE (& LEVEL) 
C0201976|T034||LNC|CREATININE - SERUM
C0201976|T034||LNC|SERUM CREATININE NOS 
C0201976|T034||LNC|SERUM CREATININE NOS
C0201976|T034||LNC|SERUM CREATININE (& LEVEL)
C0201976|T034||LNC|SERUM CREATININE TEST
C0201976|T034||LNC|CREATININE MEASUREMENT, SERUM
C1318439|T034||LNC|CREATININE LEVEL
C0201975|T034||LNC|CREATININE MEASUREMENT
C0201975|T034||LNC|CREATININE; BLOOD
C0201975|T034||LNC|BLOOD CREATININE
C0201975|T034||LNC|CREATININE
C0201975|T034||LNC|TEST;CREATININE
C0201975|T034||LNC|CREATININE BLOOD
C0201975|T034||LNC|BLOOD CREATININE LEVEL
C0201975|T034||LNC|MEASUREMENT OF CREATININE
C0201975|T034||LNC|CR
C0201975|T034||LNC|LAB-BASED CHEM MEASUREMENTS CREATININE
C0201975|T034||LNC|MEASUREMENT OF CREATININE 
C0201975|T034||LNC|CREAT
C0201975|T034||LNC|BLOOD CREATININE LEVEL 
C0201975|T034||LNC|CREATININE MEASUREMENT 
C0201975|T034||LNC|CREATININE MEASUREMENT, NOS
C0201975|T034||LNC|ASSAY OF CREATININE
C0201975|T034||LNC|CREATININE TEST
C2981751|T034||LNC|SERUM CREATININE ASSAY
C1278055|T034||LNC|PLASMA CREATININE MEASUREMENT
C1278055|T034||LNC|PLASMA CREATININE LEVEL
C1278055|T034||LNC|PLASMA CREATININE LEVEL 
C1278055|T034||LNC|PLASMA CREATININE
C1278055|T034||LNC|PLASMA CREATININE MEASUREMENT 
C1278055|T034||LNC|PLASMA CREATININE MEASUREMENT 
C3694999|T034||LNC|CREATININE CONCENTRATION (SERUM OR PLASMA)
C3694999|T034||LNC|SERUM OR PLASMA CREATININE CONCENTRATION 
C3694999|T034||LNC|SERUM OR PLASMA CREATININE CONCENTRATION
C3694393|T034||LNC|LAB-BASED CHEM MEASUREMENTS CREATININE CLEARANCE - GLOMERULAR FILTRATION 
C3694393|T034||LNC|LAB-BASED CHEM MEASUREMENTS CREATININE CLEARANCE - GLOMERULAR FILTRATION
C0428279|T034||LNC|FINDING OF CREATININE LEVEL
C0428279|T034||LNC|LAB-BASED CHEM MEASUREMENTS CREATININE LEVEL FINDING
C0428279|T034||LNC|CREATININE LEVEL FINDING 
C0428279|T034||LNC|CREATININE LEVEL FINDING
C0428279|T034||LNC|CREATININE LEVEL
C0428279|T034||LNC|CREATININE LEVEL - FINDING
C0428279|T034||LNC|FINDING OF CREATININE LEVEL 
C1278053|T034||LNC|UNCOMMON CORRECTION, BUT I SUPPOSE YOU CAN KEEP IT
C1278053|T034||LNC|CORRECTED PLASMA CREATININE LEVEL 
C1278053|T034||LNC|CORRECTED PLASMA CREATININE MEASUREMENT 
C1278053|T034||LNC|CORRECTED PLASMA CREATININE MEASUREMENT
C0852810|T034||LNC|CREATININE BLOOD DECREASED
C0239150|T034||LNC|CREATININE LOW
C0239150|T034||LNC|CREATININE DECREASED
C0555149|T034||LNC|CREATININE IN SAMPLE 
C0555149|T034||LNC|CREATININE IN SAMPLE
C0600061|T034||LNC|SERUM CREATININE
C0600061|T034||LNC|SERUM CREATININE LEVEL
C0600061|T034||LNC|FINDING OF SERUM CREATININE LEVEL
C0600061|T034||LNC|SERUM CREATININE LEVEL FINDING
C0600061|T034||LNC|SERUM CREATININE LEVEL FINDING 
C0600061|T034||LNC|FINDING OF SERUM CREATININE LEVEL 
C0600061|T034||LNC|SERUM CREATININE LEVEL - FINDING
C2114518|T034||LNC|PREVIOUSLY (LESS THAN 3 MONTHS) NORMAL CREATININE NOW RISING DAILY
C2114518|T034||LNC|PREVIOUSLY (LESS THAN 3 MONTHS) NORMAL CREATININE NOW RISING DAILY 
C2114518|T034||LNC|PREVIOUSLY (< 3 MONTHS) NORMAL CREATININE NOW RISING DAILY
C2114518|T034||LNC|PREVIOUSLY (< 3MO.) NORMAL CREATININE NOW RISING DAILY
C2114518|T034||LNC|A PREVIOUSLY (< 3MO.) NORMAL CREATININE IS NOW RISING DAILY
C1278054|T034||LNC|CORRECTED SERUM CREATININE LEVEL 
C1278054|T034||LNC|CORRECTED SERUM CREATININE LEVEL
C1278054|T034||LNC|CORRECTED SERUM CREATININE MEASUREMENT 
C1278054|T034||LNC|CORRECTED SERUM CREATININE MEASUREMENT
