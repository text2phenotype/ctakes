C0003962|T047|158530005|SNOMEDCT_US|ASCITES|[D]ASCITES (SITUATION)
C0741240|T047||SNOMEDCT_US|ASCITES FLUID INFECTION
C0741242|T047||SNOMEDCT_US|ASCITES NEW ONSET
C0741245|T047||SNOMEDCT_US|ASCITES UNKNOWN ORIGIN
C0003964|T047|409615008|SNOMEDCT_US|PERITONEAL FLUID |ASCITIC FLUID (SUBSTANCE)
C0401037|T047|236004002|SNOMEDCT_US|HEPATIC ASCITES|HEPATIC ASCITES (DISORDER)
C0003962|T047|158530005|SNOMEDCT_US|ASCITES|[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|[D]ASCITES (CONTEXT-DEPENDENT CATEGORY)|[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|[D]ASCITES NOS (CONTEXT-DEPENDENT CATEGORY)|[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|ABDOMINAL DROPSY|[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|HYDROPS ABDOMINIS|[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|PERITONEAL DROPSY|[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|PERITONEAL EXUDATE|[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|HYDROPERITONIA|[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|ABDOMINAL ASCITES|[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|ASCITES (PHYSICAL FINDING)|[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|ASCITES |[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|ABDOMEN ASCITES|[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|ASCITES WAS DISCOVERED|[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|ASCITES NOS|[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|ASCITES [DISEASE/FINDING]|[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|[D]ASCITES |[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|[D]ASCITES NOS |[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|ASCITES |[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|[D]ASCITES NOS|[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|[D]ASCITES|[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|HYDROPERITONEUM|[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|INCREASING ABDOMINAL DISTENTION OR ASCITES|[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|ABDOMINIS; HYDROPS|[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|HYDROPS; ABDOMINIS|[D]ASCITES (SITUATION)
C0003962|T047|158530005|SNOMEDCT_US|ASCITES, NOS|[D]ASCITES (SITUATION)
C2227708|T047||SNOMEDCT_US|ABDOMINAL X-RAY, AP VIEW: ASCITES 
C2227708|T047||SNOMEDCT_US|ABDOMINAL X-RAY, AP VIEW: ASCITES
C1955521|T047||SNOMEDCT_US|OTHER ASCITES
C1955521|T047||SNOMEDCT_US|ASCITES NEC
C2142846|T047||SNOMEDCT_US|PSEUDOCHYLOUS ASCITES
C2142846|T047||SNOMEDCT_US|PSEUDOCHYLOUS ASCITES 
C0426682|T047|27144005|SNOMEDCT_US|ASCITES FLUID WAVE|FLUID THRILL IN ABDOMEN (FINDING)
C0426682|T047|27144005|SNOMEDCT_US|ABDOMINAL FLUID WAVE (PHYSICAL FINDING)|FLUID THRILL IN ABDOMEN (FINDING)
C0426682|T047|27144005|SNOMEDCT_US|FINDING OF FLUID THRILL OF ABDOMEN |FLUID THRILL IN ABDOMEN (FINDING)
C0426682|T047|27144005|SNOMEDCT_US|FINDING OF FLUID THRILL OF ABDOMEN|FLUID THRILL IN ABDOMEN (FINDING)
C0426682|T047|27144005|SNOMEDCT_US|OBSERVATION OF FLUID THRILL OF ABDOMEN|FLUID THRILL IN ABDOMEN (FINDING)
C0426682|T047|27144005|SNOMEDCT_US|FLUID THRILL IN ABDOMEN |FLUID THRILL IN ABDOMEN (FINDING)
C0277979|T047|53073005|SNOMEDCT_US|SHIFTING ABDOMINAL DULLNESS FINDING|SHIFTING DULLNESS (FINDING)
C0277979|T047|53073005|SNOMEDCT_US|ASCITES SHIFTING DULLNESS|SHIFTING DULLNESS (FINDING)
C0277979|T047|53073005|SNOMEDCT_US|ABDOMINAL SHIFTING DULLNESS|SHIFTING DULLNESS (FINDING)
C0277979|T047|53073005|SNOMEDCT_US|SHIFTING DULLNESS OF ABDOMEN|SHIFTING DULLNESS (FINDING)
C0277979|T047|53073005|SNOMEDCT_US|ABDOMINAL SHIFTING DULLNESS (PHYSICAL FINDING)|SHIFTING DULLNESS (FINDING)
C0277979|T047|53073005|SNOMEDCT_US|ASCITES WITH SHIFTING DULLNESS WAS DISCOVERED|SHIFTING DULLNESS (FINDING)
C0277979|T047|53073005|SNOMEDCT_US|SHIFTING DULLNESS |SHIFTING DULLNESS (FINDING)
C0277979|T047|53073005|SNOMEDCT_US|SHIFTING DULLNESS|SHIFTING DULLNESS (FINDING)
C0277979|T047|53073005|SNOMEDCT_US|SHIFTING ABDOMINAL DULLNESS|SHIFTING DULLNESS (FINDING)
C0277979|T047|53073005|SNOMEDCT_US|SHIFTING ABDOMINAL DULLNESS (OBSERVABLE ENTITY)|SHIFTING DULLNESS (FINDING)
C0277979|T047|53073005|SNOMEDCT_US|SHIFTING ABDOMINAL DULLNESS FINDING |SHIFTING DULLNESS (FINDING)
C0426679|T047|249557007|SNOMEDCT_US|ABDOMINAL PUDDLE SIGN|PUDDLE SIGN (FINDING)
C0426679|T047|249557007|SNOMEDCT_US|ABDOMINAL PUDDLE SIGN (PHYSICAL FINDING)|PUDDLE SIGN (FINDING)
C0426679|T047|249557007|SNOMEDCT_US|ASCITES PUDDLE SIGN|PUDDLE SIGN (FINDING)
C0426679|T047|249557007|SNOMEDCT_US|PUDDLE SIGN|PUDDLE SIGN (FINDING)
C0426679|T047|249557007|SNOMEDCT_US|PUDDLE SIGN |PUDDLE SIGN (FINDING)
C2022430|T047||SNOMEDCT_US|ECHOCARDIOGRAPHY: ASCITES 
C2022430|T047||SNOMEDCT_US|ECHOCARDIOGRAPHY: ASCITES
C2321829|T047||SNOMEDCT_US|SAMPLE TEMPLATE ASCITES 
C2321829|T047||SNOMEDCT_US|SAMPLE TEMPLATE ASCITES
C3532188|T047|470758004|SNOMEDCT_US|REFRACTORY ASCITES|REFRACTORY ASCITES (DISORDER)
C3532188|T047|470758004|SNOMEDCT_US|REFRACTORY ASCITES |REFRACTORY ASCITES (DISORDER)
C0585187|T047|307311001|SNOMEDCT_US|INFECTED ASCITES|INFECTED ASCITES (DISORDER)
C0585187|T047|307311001|SNOMEDCT_US|INFECTED ASCITES |INFECTED ASCITES (DISORDER)
C0267773|T047|18037001|SNOMEDCT_US|BILIARY ASCITES|BILE ASCITES (DISORDER)
C0267773|T047|18037001|SNOMEDCT_US|BILE ASCITES|BILE ASCITES (DISORDER)
C0267773|T047|18037001|SNOMEDCT_US|BILE ASCITES |BILE ASCITES (DISORDER)
C0031144|T047|78609007|SNOMEDCT_US|CHRONIC PERITONEAL EFFUSION |CHRONIC PERITONEAL EFFUSION
C0031144|T047|78609007|SNOMEDCT_US|CHRONIC PERITONEAL EFFUSION|CHRONIC PERITONEAL EFFUSION
C0031144|T047|78609007|SNOMEDCT_US|CHRONIC PERITONEAL EFFUSION |CHRONIC PERITONEAL EFFUSION
C0031144|T047|78609007|SNOMEDCT_US|PERITONEAL EFFUSION|CHRONIC PERITONEAL EFFUSION
C0031144|T047|78609007|SNOMEDCT_US|PERITONEAL EFFUSION (CHRONIC)|CHRONIC PERITONEAL EFFUSION
C0008732|T047|52985009|SNOMEDCT_US|CHYLOUS ASCITES|CHYLOUS ASCITES (DISORDER)
C0008732|T047|52985009|SNOMEDCT_US|ASCITES, CHYLOUS|CHYLOUS ASCITES (DISORDER)
C0008732|T047|52985009|SNOMEDCT_US|CHYLOPERITONEUM|CHYLOUS ASCITES (DISORDER)
C0008732|T047|52985009|SNOMEDCT_US|CHYLOUS ASCITES |CHYLOUS ASCITES (DISORDER)
C0008732|T047|52985009|SNOMEDCT_US|CHYLOUS ASCITES [DISEASE/FINDING]|CHYLOUS ASCITES (DISORDER)
C0008732|T047|52985009|SNOMEDCT_US|ASCITES CHYLOUS|CHYLOUS ASCITES (DISORDER)
C0008732|T047|52985009|SNOMEDCT_US|CHYLOUS ASCITES |CHYLOUS ASCITES (DISORDER)
C0008732|T047|52985009|SNOMEDCT_US|ASCITES; CHYLOUS|CHYLOUS ASCITES (DISORDER)
C0008732|T047|52985009|SNOMEDCT_US|CHYLOUS; ASCITES|CHYLOUS ASCITES (DISORDER)
C0401038|T047|236006000|SNOMEDCT_US|HYPOALBUMINAEMIC ASCITES|METABOLIC ASCITES (DISORDER)
C0401038|T047|236006000|SNOMEDCT_US|HYPOALBUMINEMIC ASCITES|METABOLIC ASCITES (DISORDER)
C0401037|T047|236004002|SNOMEDCT_US|HEPATIC ASCITES|HEPATIC ASCITES (DISORDER)
C0401037|T047|236004002|SNOMEDCT_US|HEPATIC ASCITES |HEPATIC ASCITES (DISORDER)
C3670559|T047||SNOMEDCT_US|FIBRINOUS PERITONEAL EFFUSION
C3670559|T047||SNOMEDCT_US|FIBRINOUS ASCITES
C3670559|T047||SNOMEDCT_US|FIBRINOUS ASCITES 
C3670560|T047||SNOMEDCT_US|MODIFIED TRANSUDATIVE PERITONEAL EFFUSION
C3670560|T047||SNOMEDCT_US|MODIFIED TRANSUDATIVE ASCITES 
C3670560|T047||SNOMEDCT_US|MODIFIED TRANSUDATIVE ASCITES
C3670560|T047||SNOMEDCT_US|MODIFIED TRANSUDATE ASCITES
C0519092|T047||SNOMEDCT_US|TRANSUDATE ASCITES
C0519092|T047||SNOMEDCT_US|TRANSUDATIVE PERITONEAL EFFUSION
C0519092|T047||SNOMEDCT_US|TRANSUDATIVE ASCITES 
C0519092|T047||SNOMEDCT_US|TRANSUDATIVE ASCITES
C4038874|T047|1082601000119104|SNOMEDCT_US|ASCITES DUE TO ALCOHOLIC CIRRHOSIS |ASCITES DUE TO ALCOHOLIC CIRRHOSIS (DISORDER)
C4038874|T047|1082601000119104|SNOMEDCT_US|ASCITES DUE TO ALCOHOLIC CIRRHOSIS|ASCITES DUE TO ALCOHOLIC CIRRHOSIS (DISORDER)
C4038944|T047|1082611000119101|SNOMEDCT_US|ASCITES DUE TO ALCOHOLIC HEPATITIS|ASCITES DUE TO ALCOHOLIC HEPATITIS (DISORDER)
C4038944|T047|1082611000119101|SNOMEDCT_US|ASCITES DUE TO ALCOHOLIC HEPATITIS |ASCITES DUE TO ALCOHOLIC HEPATITIS (DISORDER)
C3665480|T047|207253004|SNOMEDCT_US|[D]FLUID IN PERITONEAL CAVITY (CONTEXT-DEPENDENT CATEGORY)|[D]FLUID IN PERITONEAL CAVITY (SITUATION)
C3665480|T047|207253004|SNOMEDCT_US|FLUID IN PERITONEAL CAVITY|[D]FLUID IN PERITONEAL CAVITY (SITUATION)
C3665480|T047|207253004|SNOMEDCT_US|[D]FLUID IN PERITONEAL CAVITY |[D]FLUID IN PERITONEAL CAVITY (SITUATION)
C3665480|T047|207253004|SNOMEDCT_US|[D]FLUID IN PERITONEAL CAVITY|[D]FLUID IN PERITONEAL CAVITY (SITUATION)
C3665480|T047|207253004|SNOMEDCT_US|FLUID IN PERITONEAL CAVITY |[D]FLUID IN PERITONEAL CAVITY (SITUATION)
C1385680|T047||SNOMEDCT_US|EFFUSION; ABDOMEN
C1385680|T047||SNOMEDCT_US|ABDOMEN; EFFUSION
C1390873|T047||SNOMEDCT_US|ABDOMEN; UPSET, FLUID
C1390873|T047||SNOMEDCT_US|UPSET; ABDOMEN, FLUID
C1390876|T047||SNOMEDCT_US|DISTENSION; ABDOMEN, FLUID
C1390876|T047||SNOMEDCT_US|ABDOMEN; DISTENSION, FLUID
C1390885|T047||SNOMEDCT_US|EFFUSION; PERITONEAL CAVITY
C1390885|T047||SNOMEDCT_US|PERITONEAL CAVITY; EFFUSION
C0003964|T047|409615008|SNOMEDCT_US|ASCITIC FLUID|ASCITIC FLUID (SUBSTANCE)
C0003964|T047|409615008|SNOMEDCT_US|ASCITIC FLUIDS|ASCITIC FLUID (SUBSTANCE)
C0003964|T047|409615008|SNOMEDCT_US|EFFUSION, PERITONEAL|ASCITIC FLUID (SUBSTANCE)
C0003964|T047|409615008|SNOMEDCT_US|EFFUSIONS, PERITONEAL|ASCITIC FLUID (SUBSTANCE)
C0003964|T047|409615008|SNOMEDCT_US|FLUID, ASCITIC|ASCITIC FLUID (SUBSTANCE)
C0003964|T047|409615008|SNOMEDCT_US|FLUID, PERITONEAL|ASCITIC FLUID (SUBSTANCE)
C0003964|T047|409615008|SNOMEDCT_US|FLUIDS, ASCITIC|ASCITIC FLUID (SUBSTANCE)
C0003964|T047|409615008|SNOMEDCT_US|FLUIDS, PERITONEAL|ASCITIC FLUID (SUBSTANCE)
C0003964|T047|409615008|SNOMEDCT_US|PERITONEAL EFFUSIONS|ASCITIC FLUID (SUBSTANCE)
C0003964|T047|409615008|SNOMEDCT_US|PERITONEAL FLUIDS|ASCITIC FLUID (SUBSTANCE)
C0003964|T047|409615008|SNOMEDCT_US|PERITONEAL FLUID|ASCITIC FLUID (SUBSTANCE)
C0003964|T047|409615008|SNOMEDCT_US|PERITONEAL FLUID |ASCITIC FLUID (SUBSTANCE)
C0003964|T047|409615008|SNOMEDCT_US|PERITONEAL FLUID |ASCITIC FLUID (SUBSTANCE)
C0003964|T047|409615008|SNOMEDCT_US|PERITONEAL EFFUSION|ASCITIC FLUID (SUBSTANCE)
C0003964|T047|409615008|SNOMEDCT_US|FLUID, ASCITES|ASCITIC FLUID (SUBSTANCE)
C0003964|T047|409615008|SNOMEDCT_US|EFFUSION; PERITONEAL|ASCITIC FLUID (SUBSTANCE)
C0003964|T047|409615008|SNOMEDCT_US|PERITONEAL; EFFUSION|ASCITIC FLUID (SUBSTANCE)
C0003964|T047|409615008|SNOMEDCT_US|ASCITIC FLUID |ASCITIC FLUID (SUBSTANCE)
C0437001|T047|140519000|SNOMEDCT_US|ON EXAMINATION - ASCITES|O/E - ASCITES (FINDING)
C0437001|T047|140519000|SNOMEDCT_US|O/E - ASCITES|O/E - ASCITES (FINDING)
C0437001|T047|140519000|SNOMEDCT_US|O/E - ASCITES NOS |O/E - ASCITES (FINDING)
C0437001|T047|140519000|SNOMEDCT_US|ON EXAMINATION - ASCITES NOS|O/E - ASCITES (FINDING)
C0437001|T047|140519000|SNOMEDCT_US|O/E - ASCITES NOS|O/E - ASCITES (FINDING)
C0437001|T047|140519000|SNOMEDCT_US|ON EXAMINATION - ASCITES NOS |O/E - ASCITES (FINDING)
C0437001|T047|140519000|SNOMEDCT_US|O/E - ASCITES |O/E - ASCITES (FINDING)
C0437001|T047|140519000|SNOMEDCT_US|ON EXAMINATION - ASCITES (CONTEXT-DEPENDENT CATEGORY)|O/E - ASCITES (FINDING)
C0437001|T047|140519000|SNOMEDCT_US|ON EXAMINATION - ASCITES NOS (CONTEXT-DEPENDENT CATEGORY)|O/E - ASCITES (FINDING)
C0437001|T047|140519000|SNOMEDCT_US|ON EXAMINATION - ASCITES |O/E - ASCITES (FINDING)
C4038684|T047|1092801000119102|SNOMEDCT_US|HEPATIC ASCITES CO-OCCURRENT WITH CHRONIC ACTIVE HEPATITIS DUE TO TOXIC LIVER DISEASE|HEPATIC ASCITES CO-OCCURRENT WITH CHRONIC ACTIVE HEPATITIS DUE TO TOXIC LIVER DISEASE (DISORDER)
C4038684|T047|1092801000119102|SNOMEDCT_US|HEPATIC ASCITES CO-OCCURRENT WITH CHRONIC ACTIVE HEPATITIS DUE TO TOXIC LIVER DISEASE |HEPATIC ASCITES CO-OCCURRENT WITH CHRONIC ACTIVE HEPATITIS DUE TO TOXIC LIVER DISEASE (DISORDER)
C4040413|T047|1085021000119106|SNOMEDCT_US|HEPATIC ASCITES DUE TO CHRONIC ALCOHOLIC HEPATITIS |HEPATIC ASCITES DUE TO CHRONIC ALCOHOLIC HEPATITIS (DISORDER)
C4040413|T047|1085021000119106|SNOMEDCT_US|HEPATIC ASCITES DUE TO CHRONIC ALCOHOLIC HEPATITIS|HEPATIC ASCITES DUE TO CHRONIC ALCOHOLIC HEPATITIS (DISORDER)
