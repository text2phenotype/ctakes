C2239176|T191|187769009|SNOMEDCT_US|LIVER CARCINOMA|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|LIVER CELL CARCINOMA|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|CARCINOMA, HEPATOCELLULAR|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|CARCINOMAS, HEPATOCELLULAR|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|HEPATOCELLULAR CARCINOMAS|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|HEPATOMA|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|HEPATOMAS|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|HEPATOCELLULAR CARCINOMA|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|CARCINOMA OF LIVER |PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|HEPATOCELLULAR CARCINOMA OF LIVER |PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|HEPATOCELLULAR CARCINOMA OF LIVER|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|LIVER NEOPLASM MALIGNANT CARCINOMA|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|CARCINOMA OF LIVER|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|LIVER CARCINOMA|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|LIVER CELL CANCER (HEPATOCELLULAR CARCINOMA)|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|CARCINOMA, HEPATOCELLULAR [DISEASE/FINDING]|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|CANCERS, ADULT LIVER|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|ADULT LIVER CANCER|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|CANCER, ADULT LIVER|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|ADULT LIVER CANCERS|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|LIVER CANCERS, ADULT|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|LIVER CANCER, ADULT|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|LIVER CELL CARCINOMA, ADULT|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|LIVER CELL CARCINOMAS|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|CELL CARCINOMA, LIVER|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|CELL CARCINOMAS, LIVER|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|CARCINOMA, LIVER CELL|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|CARCINOMAS, LIVER CELL|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|HEPATIC CELL CARCINOMA|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|PRIMARY CARCINOMA OF LIVER|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|LIVER NEOPLASM MALIGNANT CARCINOMA PRIMARY|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|PRIMARY CARCINOMA OF LIVER |PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|HCC|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|CARCINOMA, HEPATOCELLULAR, MALIGNANT|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|[M]HEPATOCELLULAR CARCINOMA NOS|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|CARCINOMA OF THE LIVER CELLS|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|PRIMARY CARCINOMA OF THE LIVER CELLS|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|CARCINOMA OF LIVER CELLS|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|PRIMARY CARCINOMA OF LIVER CELLS|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|LIVER CELL CARCINOMA (CLINICAL)|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|HEPATOCELLULAR CARCINOMA (CLINICAL)|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|CARCINOMA LIVER|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|CARCINOMA HEPATOCELLULAR|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|HEPATOCARCINOMA|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|HEPATOMA, MALIGNANT|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|MALIGNANT HEPATOMA|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|LCC - LIVER CELL CARCINOMA|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|HCC - HEPATOCELLULAR CARCINOMA|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|HEPATOCELLULAR CARCINOMA (MORPHOLOGIC ABNORMALITY)|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|LIVER CELL CARCINOMA |PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|PRIMARY CARCINOMA OF LIVER |PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|CARCINOMA; HEPATIC CELL|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|CARCINOMA; HEPATOCELLULAR|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|HEPATIC CELL; CARCINOMA|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|HEPATOCELLULAR; CARCINOMA|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|HEPATOCELLULAR CARCINOMA, NOS|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|HEPATOMA, NOS|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|CARCINOMA OF LIVER, SPECIFIED AS PRIMARY|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2239176|T191|187769009|SNOMEDCT_US|CARCINOMA OF LIVER CELL|PRIMARY CARCINOMA OF LIVER (DISORDER)
C2205336|T191||SNOMEDCT_US|MALIGNANT EPITHELIOMA OF LIVER
C2205336|T191||SNOMEDCT_US|LIVER NEOPLASM MALIGNANT CARCINOMA EPITHELIOMA
C2205336|T191||SNOMEDCT_US|MALIGNANT EPITHELIOMA OF LIVER 
C2111635|T191||SNOMEDCT_US|LARGE CELL CARCINOMA OF LIVER
C2111635|T191||SNOMEDCT_US|LARGE CELL CARCINOMA OF LIVER 
C2012092|T191||SNOMEDCT_US|GLASSY CELL CARCINOMA OF LIVER 
C2012092|T191||SNOMEDCT_US|GLASSY CELL CARCINOMA OF LIVER
C2205337|T191||SNOMEDCT_US|ANAPLASTIC CARCINOMA OF LIVER 
C2205337|T191||SNOMEDCT_US|ANAPLASTIC CARCINOMA OF LIVER
C2205337|T191||SNOMEDCT_US|LIVER NEOPLASM MALIGNANT CARCINOMA ANAPLASTIC
C2082443|T191||SNOMEDCT_US|PLEOMORPHIC CARCINOMA OF LIVER
C2082443|T191||SNOMEDCT_US|PLEOMORPHIC CARCINOMA OF LIVER 
C2011254|T191||SNOMEDCT_US|GIANT CELL CARCINOMA OF LIVER 
C2011254|T191||SNOMEDCT_US|GIANT CELL CARCINOMA OF LIVER
C2018394|T191||SNOMEDCT_US|SPINDLE CELL CARCINOMA OF LIVER
C2018394|T191||SNOMEDCT_US|SPINDLE CELL CARCINOMA OF LIVER 
C2011218|T191||SNOMEDCT_US|GIANT CELL AND SPINDLE CELL CARCINOMA OF LIVER 
C2011218|T191||SNOMEDCT_US|LIVER NEOPLASM MALIGNANT CARCINOMA GIANT CELL & SPINDLE CELL
C2011218|T191||SNOMEDCT_US|GIANT CELL AND SPINDLE CELL CARCINOMA OF LIVER
C2142923|T191||SNOMEDCT_US|PSEUDOSARCOMATOUS CARCINOMA OF LIVER 
C2142923|T191||SNOMEDCT_US|PSEUDOSARCOMATOUS CARCINOMA OF LIVER
C2111805|T191||SNOMEDCT_US|POLYGONAL CELL CARCINOMA OF LIVER 
C2111805|T191||SNOMEDCT_US|POLYGONAL CELL CARCINOMA OF LIVER
C2076526|T191||SNOMEDCT_US|MORE LIKELY CHOLANGIOCARCINOMA, BUT MIGHT BE HCC
C2076526|T191||SNOMEDCT_US|INFILTRATING DUCTAL CARCINOMA OF LIVER
C2106546|T191||SNOMEDCT_US|COMEDOCARCINOMA OF LIVER
C2106546|T191||SNOMEDCT_US|LIVER NEOPLASM MALIGNANT CARCINOMA COMEDOCARCINOMA
C2106546|T191||SNOMEDCT_US|COMEDOCARCINOMA OF LIVER 
C2078053|T191||SNOMEDCT_US|I'M NOT SURE IF THIS IS A TYPE OF HCC
C2078053|T191||SNOMEDCT_US|INTRACYSTIC CARCINOMA OF LIVER
C2047535|T191||SNOMEDCT_US|HYPERSECRETORY CYSTIC CARCINOMA OF LIVER 
C2047535|T191||SNOMEDCT_US|LIVER NEOPLASM MALIGNANT CARCINOMA CYSTIC HYPERSECRETORY
C2047535|T191||SNOMEDCT_US|HYPERSECRETORY CYSTIC CARCINOMA OF LIVER
C2064401|T191||SNOMEDCT_US|UNDIFFERENTIATED CARCINOMA OF LIVER 
C2064401|T191||SNOMEDCT_US|UNDIFFERENTIATED CARCINOMA OF LIVER
C2064401|T191||SNOMEDCT_US|UNDIFFERENTIATED LIVER CARCINOMA
C2064401|T191||SNOMEDCT_US|UNDIFFERENTIATED PRIMARY LIVER CARCINOMA
C0334287|T191|253018005|SNOMEDCT_US|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA OF LIVER |FIBROLAMELLAR HEPATOCELLULAR CARCINOMA (DISORDER)
C0334287|T191|253018005|SNOMEDCT_US|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA OF LIVER|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA (DISORDER)
C0334287|T191|253018005|SNOMEDCT_US|FIBROLAMELLAR VARIANT OF HEPATOCELLULAR CARCINOMA|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA (DISORDER)
C0334287|T191|253018005|SNOMEDCT_US|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA (DISORDER)
C0334287|T191|253018005|SNOMEDCT_US|HEPATOCELLULAR CARCINOMA (FIBROLAMELLAR VARIANT)|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA (DISORDER)
C0334287|T191|253018005|SNOMEDCT_US|FLC|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA (DISORDER)
C0334287|T191|253018005|SNOMEDCT_US|FIBROLAMELLAR CARCINOMA|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA (DISORDER)
C0334287|T191|253018005|SNOMEDCT_US|[M]HEPATOCELLULAR CARCINOMA, FIBROLAMELLAR|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA (DISORDER)
C0334287|T191|253018005|SNOMEDCT_US|[M] HEPATOCELLULAR CARCINOMA, FIBROLAMELLAR|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA (DISORDER)
C0334287|T191|253018005|SNOMEDCT_US|HEPATOCELLULAR CARCINOMA, FIBROLAMELLAR|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA (DISORDER)
C0334287|T191|253018005|SNOMEDCT_US|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA |FIBROLAMELLAR HEPATOCELLULAR CARCINOMA (DISORDER)
C0334287|T191|253018005|SNOMEDCT_US|HEPATOCELLULAR CARCINOMA, FIBROLAMELLAR (MORPHOLOGIC ABNORMALITY)|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA (DISORDER)
C0334287|T191|253018005|SNOMEDCT_US|CARCINOMA; HEPATOCELLULAR, FIBROLAMELLAR|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA (DISORDER)
C0334287|T191|253018005|SNOMEDCT_US|FIBROLAMELLAR; HEPATOCELLULAR CARCINOMA|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA (DISORDER)
C0334287|T191|253018005|SNOMEDCT_US|HEPATOCELLULAR; CARCINOMA, FIBROLAMELLAR|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA (DISORDER)
C0334287|T191|253018005|SNOMEDCT_US|FIBROLAMELLAR CARCINOMA OF LIVER CELLS|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA (DISORDER)
C0334287|T191|253018005|SNOMEDCT_US|FIBROLAMELLAR CARCINOMA OF THE LIVER CELLS|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA (DISORDER)
C0334287|T191|253018005|SNOMEDCT_US|HEPATOCELLULAR FIBROLAMELLAR CARCINOMA|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA (DISORDER)
C0334287|T191|253018005|SNOMEDCT_US|LIVER CELL FIBROLAMELLAR CARCINOMA|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA (DISORDER)
C0334287|T191|253018005|SNOMEDCT_US|ONCOCYTIC HEPATOCELLULAR TUMOR|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA (DISORDER)
C0334287|T191|253018005|SNOMEDCT_US|POLYGONAL CELL TYPE HEPATOCELLULAR CARCINOMA WITH FIBROUS STROMA|FIBROLAMELLAR HEPATOCELLULAR CARCINOMA (DISORDER)
C2205338|T191||SNOMEDCT_US|SCIRRHOUS HEPATOCELLULAR CARCINOMA OF LIVER 
C2205338|T191||SNOMEDCT_US|SCIRRHOUS HEPATOCELLULAR CARCINOMA OF LIVER
C1266019|T191|128648009|SNOMEDCT_US|SPINDLE CELL HEPATOCELLULAR CARCINOMA OF LIVER|HEPATOCELLULAR CARCINOMA, SARCOMATOID
C1266019|T191|128648009|SNOMEDCT_US|SPINDLE CELL HEPATOCELLULAR CARCINOMA OF LIVER |HEPATOCELLULAR CARCINOMA, SARCOMATOID
C1266019|T191|128648009|SNOMEDCT_US|HEPATOCELLULAR CARCINOMA, SARCOMATOID|HEPATOCELLULAR CARCINOMA, SARCOMATOID
C1266019|T191|128648009|SNOMEDCT_US|HEPATOCELLULAR CARCINOMA, SPINDLE CELL VARIANT (MORPHOLOGIC ABNORMALITY)|HEPATOCELLULAR CARCINOMA, SARCOMATOID
C1266019|T191|128648009|SNOMEDCT_US|HEPATOCELLULAR CARCINOMA, SPINDLE CELL VARIANT|HEPATOCELLULAR CARCINOMA, SARCOMATOID
C1266020|T191|128649001|SNOMEDCT_US|CLEAR CELL HEPATOCELLULAR CARCINOMA OF LIVER |HEPATOCELLULAR CARCINOMA, CLEAR CELL TYPE (MORPHOLOGIC ABNORMALITY)
C1266020|T191|128649001|SNOMEDCT_US|CLEAR CELL HEPATOCELLULAR CARCINOMA OF LIVER|HEPATOCELLULAR CARCINOMA, CLEAR CELL TYPE (MORPHOLOGIC ABNORMALITY)
C1266020|T191|128649001|SNOMEDCT_US|HEPATOCELLULAR CARCINOMA, CLEAR CELL TYPE (MORPHOLOGIC ABNORMALITY)|HEPATOCELLULAR CARCINOMA, CLEAR CELL TYPE (MORPHOLOGIC ABNORMALITY)
C1266020|T191|128649001|SNOMEDCT_US|HEPATOCELLULAR CARCINOMA, CLEAR CELL TYPE|HEPATOCELLULAR CARCINOMA, CLEAR CELL TYPE (MORPHOLOGIC ABNORMALITY)
C2082477|T191||SNOMEDCT_US|PLEOMORPHIC HEPATOCELLULAR CARCINOMA OF LIVER
C2082477|T191||SNOMEDCT_US|PLEOMORPHIC HEPATOCELLULAR CARCINOMA OF LIVER 
C0221287|T191|274902006|SNOMEDCT_US|HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA|COMBINED HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA (DISORDER)
C0221287|T191|274902006|SNOMEDCT_US|LIVER NEOPLASM HEPATOCELLULAR CARCINOMA & CHOLANGIOCARCINOMA|COMBINED HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA (DISORDER)
C0221287|T191|274902006|SNOMEDCT_US|HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA |COMBINED HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA (DISORDER)
C0221287|T191|274902006|SNOMEDCT_US|MIXED HEPATOCELLULAR CHOLANGIOCARCINOMA|COMBINED HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA (DISORDER)
C0221287|T191|274902006|SNOMEDCT_US|[M]COMBINED HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA|COMBINED HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA (DISORDER)
C0221287|T191|274902006|SNOMEDCT_US|COMBINED HEPATOCELLULAR AND CHOLANGIOCARCINOMA|COMBINED HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA (DISORDER)
C0221287|T191|274902006|SNOMEDCT_US|HEPATOCHOLANGIOCARCINOMA|COMBINED HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA (DISORDER)
C0221287|T191|274902006|SNOMEDCT_US|MIXED HEPATOCELLULAR AND BILE DUCT CARCINOMA|COMBINED HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA (DISORDER)
C0221287|T191|274902006|SNOMEDCT_US|COMBINED HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA|COMBINED HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA (DISORDER)
C0221287|T191|274902006|SNOMEDCT_US|COMBINED HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA |COMBINED HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA (DISORDER)
C0221287|T191|274902006|SNOMEDCT_US|COMBINED HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA (MORPHOLOGIC ABNORMALITY)|COMBINED HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA (DISORDER)
C0221287|T191|274902006|SNOMEDCT_US|CHOLANGIOCARCINOMA; WITH HEPATOCELLULAR CARCINOMA|COMBINED HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA (DISORDER)
C0221287|T191|274902006|SNOMEDCT_US|CHOLANGIOHEPATOMA|COMBINED HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA (DISORDER)
C0221287|T191|274902006|SNOMEDCT_US|HEPATOCELLULAR CARCINOMA; CHOLANGIOCARCINOMA|COMBINED HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA (DISORDER)
C0221287|T191|274902006|SNOMEDCT_US|LIVER AND INTRAHEPATIC BILIARY TRACT CARCINOMA|COMBINED HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA (DISORDER)
C0221287|T191|274902006|SNOMEDCT_US|CARCINOMA OF LIVER AND INTRAHEPATIC BILIARY TRACT|COMBINED HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA (DISORDER)
C0221287|T191|274902006|SNOMEDCT_US|CARCINOMA OF THE LIVER AND INTRAHEPATIC BILIARY TRACT|COMBINED HEPATOCELLULAR CARCINOMA AND CHOLANGIOCARCINOMA (DISORDER)
C0279607|T191||SNOMEDCT_US|HEPATOMA, ADULT PRIMARY
C0279607|T191||SNOMEDCT_US|ADULT PRIMARY HEPATOCELLULAR CARCINOMA
C0279607|T191||SNOMEDCT_US|HEPATOCELLULAR CARCINOMA, ADULT PRIMARY
C0279607|T191||SNOMEDCT_US|ADULT HEPATOCELLULAR CARCINOMA
C0279607|T191||SNOMEDCT_US|ADULT HEPATOMA
C0279607|T191||SNOMEDCT_US|ADULT LIVER CARCINOMA
C0279607|T191||SNOMEDCT_US|ADULT PRIMARY CARCINOMA OF LIVER CELL
C0279607|T191||SNOMEDCT_US|ADULT PRIMARY CARCINOMA OF THE LIVER CELL
C0279607|T191||SNOMEDCT_US|ADULT PRIMARY HEPATOMA
C0279607|T191||SNOMEDCT_US|ADULT PRIMARY LIVER CARCINOMA
C0279607|T191||SNOMEDCT_US|ADULT PRIMARY LIVER CELL CARCINOMA
C2983709|T191||SNOMEDCT_US|HEPATOCELLULAR CARCINOMA BY AJCC V6 STAGE
C2984092|T191||SNOMEDCT_US|HEPATOCELLULAR CARCINOMA BY AJCC V7 STAGE
C3273019|T191||SNOMEDCT_US|EARLY HEPATOCELLULAR CARCINOMA
C3273032|T191||SNOMEDCT_US|LYMPHOEPITHELIOMA-LIKE HEPATOCELLULAR CARCINOMA
C3273033|T191||SNOMEDCT_US|WELL DIFFERENTIATED HEPATOCELLULAR CARCINOMA
C3273034|T191||SNOMEDCT_US|MODERATELY DIFFERENTIATED HEPATOCELLULAR CARCINOMA
C3273035|T191||SNOMEDCT_US|POORLY DIFFERENTIATED HEPATOCELLULAR CARCINOMA
C0345904|T191|363361004|SNOMEDCT_US|MALIGNANT NEOPLASM OF LIVER, UNSPECIFIED|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|MALIGNANT NEOPLASM OF LIVER|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|LIVER CANCER|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|LIVER CANCER |MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|LIVER NEOPLASM MALIGNANT|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|MALIGNANT NEOPLASM OF LIVER |MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|HEPATIC NEOPLASMS MALIGNANT|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|CANCER, HEPATIC|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|CANCERS, HEPATIC|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|HEPATIC CANCERS|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|CANCERS, LIVER|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|LIVER CANCERS|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|MALIGNANT TUMOR OF LIVER|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|MALIGNANT NEO LIVER NOS|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|MALIGNANT NEOPLASM OF LIVER, NOT SPECIFIED AS PRIMARY OR SECONDARY|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|HEPATIC CANCER|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|CANCER, LIVER|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|MALIG NEOPLASM OF LIVER, NOT SPECIFIED AS PRIMARY OR SEC|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|CANCERS, HEPATOCELLULAR|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|HEPATOCELLULAR CANCERS|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|MALIGNANT NEOPLASM OF LIVER UNSPECIFIED |MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|MALIGNANT TUMOR OF LIVER |MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|MALIGNANT NEOPLASM OF LIVER UNSPECIFIED|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|MALIGNANT TUMOUR OF LIVER|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|LIVER--CANCER|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|CANCER, HEPATOCELLULAR|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|HEPATIC NEOPLASM MALIGNANT NOS|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|MALIGNANT HEPATIC NEOPLASM|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|MALIGNANT LIVER TUMOR|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|HEPATIC TUMOUR MALIGNANT|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|LIVER, CANCER OF|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|MALIGNANT LIVER TUMOUR|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|HEPATIC NEOPLASM MALIGNANT|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|HEPATIC TUMOR MALIGNANT|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|HEPATOCELLULAR CANCER|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|CANCER OF THE LIVER|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|CA - LIVER CANCER|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|MALIGNANT NEOPLASM OF LIVER |MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|MALIGNANT NEOPLASM OF LIVER, NOS|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|CANCER OF LIVER|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|NEOPLASM MALIG;LIVER|MALIGNANT TUMOR OF LIVER (DISORDER)
C0345904|T191|363361004|SNOMEDCT_US|MALIGNANT NEOSPLASM OF THE LIVER|MALIGNANT TUMOR OF LIVER (DISORDER)
C0564703|T191|286888000|SNOMEDCT_US|CA LIVER/BILIARY SYSTEM NOS |CARCINOMA LIVER/BILIARY SYSTEM NOS (DISORDER)
C0564703|T191|286888000|SNOMEDCT_US|CARCINOMA LIVER/BILIARY SYSTEM NOS|CARCINOMA LIVER/BILIARY SYSTEM NOS (DISORDER)
C0564703|T191|286888000|SNOMEDCT_US|CA LIVER/BILIARY SYSTEM|CARCINOMA LIVER/BILIARY SYSTEM NOS (DISORDER)
C0564703|T191|286888000|SNOMEDCT_US|CARCINOMA LIVER/BILIARY SYSTEM NOS |CARCINOMA LIVER/BILIARY SYSTEM NOS (DISORDER)
C0564703|T191|286888000|SNOMEDCT_US|CA LIVER/BILIARY SYSTEM NOS|CARCINOMA LIVER/BILIARY SYSTEM NOS (DISORDER)
C0564703|T191|286888000|SNOMEDCT_US|CARCINOMA OF LIVER AND BILIARY SYSTEM |CARCINOMA LIVER/BILIARY SYSTEM NOS (DISORDER)
C0564703|T191|286888000|SNOMEDCT_US|NEOPLASM MALIGNANT CARCINOMA OF LIVER AND BILIARY SYSTEM|CARCINOMA LIVER/BILIARY SYSTEM NOS (DISORDER)
C0564703|T191|286888000|SNOMEDCT_US|CARCINOMA OF LIVER AND BILIARY SYSTEM|CARCINOMA LIVER/BILIARY SYSTEM NOS (DISORDER)
C0564703|T191|286888000|SNOMEDCT_US|CARCINOMA LIVER/BILIARY SYSTEM|CARCINOMA LIVER/BILIARY SYSTEM NOS (DISORDER)
C0564703|T191|286888000|SNOMEDCT_US|CARCINOMA LIVER AND/OR BILIARY SYSTEM |CARCINOMA LIVER/BILIARY SYSTEM NOS (DISORDER)
C0564703|T191|286888000|SNOMEDCT_US|CARCINOMA LIVER AND/OR BILIARY SYSTEM|CARCINOMA LIVER/BILIARY SYSTEM NOS (DISORDER)
C0564703|T191|286888000|SNOMEDCT_US|CARCINOMA LIVER/BILIARY SYSTEM |CARCINOMA LIVER/BILIARY SYSTEM NOS (DISORDER)
C2676033|T191||SNOMEDCT_US|HEPATOBLASTOMA CAUSED BY SOMATIC MUTATION
C1969388|T191||SNOMEDCT_US|HEPATOCELLULAR CARCINOMA, SOMATIC 
C1969388|T191||SNOMEDCT_US|HEPATOCELLULAR CARCINOMA, SOMATIC
C3898888|T191||SNOMEDCT_US|HEPATOCELLULAR CARCINOMA BARCELONA CLINIC LIVER CANCER STAGING
C3898888|T191||SNOMEDCT_US|HEPATOCELLULAR CARCINOMA BY BCLC STAGE
C3898888|T191||SNOMEDCT_US|BCLC STAGING FOR HEPATOCELLULAR CARCINOMA
C3898888|T191||SNOMEDCT_US|HEPATOCELLULAR CARCINOMA BY BARCELONA CLINIC LIVER CANCER STAGE
C3898888|T191||SNOMEDCT_US|HEPATOCELLULAR CARCINOMA BCLC STAGING
C3898888|T191||SNOMEDCT_US|BARCELONA CLINIC LIVER CANCER STAGING FOR HEPATOCELLULAR CARCINOMA
C4030880|T191||SNOMEDCT_US|BIOPSY OF LIVER SHOWED CARCINOMA
C4030880|T191||SNOMEDCT_US|BIOPSY OF LIVER SHOWED CARCINOMA 
C4030854|T191||SNOMEDCT_US|BIOPSY OF LIVER SHOWED CARCINOMA PRIMARY
C4030854|T191||SNOMEDCT_US|BIOPSY OF LIVER SHOWED CARCINOMA PRIMARY 
C0744869|T191|708973006|SNOMEDCT_US|METASTATIC HEPATOCELLULAR CARCINOMA (MORPHOLOGIC ABNORMALITY)|METASTATIC HEPATOCELLULAR CARCINOMA (MORPHOLOGIC ABNORMALITY)
C0744869|T191|708973006|SNOMEDCT_US|METASTATIC HEPATOCELLULAR CARCINOMA|METASTATIC HEPATOCELLULAR CARCINOMA (MORPHOLOGIC ABNORMALITY)
C0348340|T191|190088005|SNOMEDCT_US|OTHER SPECIFIED CARCINOMAS OF LIVER|[X]OTHER SPECIFIED CARCINOMAS OF LIVER (DISORDER)
C0348340|T191|190088005|SNOMEDCT_US|[X]OTHER SPECIFIED CARCINOMAS OF LIVER|[X]OTHER SPECIFIED CARCINOMAS OF LIVER (DISORDER)
C0348340|T191|190088005|SNOMEDCT_US|OTHER SPECIFIED CARCINOMA OF LIVER|[X]OTHER SPECIFIED CARCINOMAS OF LIVER (DISORDER)
C0348340|T191|190088005|SNOMEDCT_US|OTHER SPECIFIED CARCINOMA OF LIVER |[X]OTHER SPECIFIED CARCINOMAS OF LIVER (DISORDER)
C0348340|T191|190088005|SNOMEDCT_US|[X]OTHER SPECIFIED CARCINOMAS OF LIVER |[X]OTHER SPECIFIED CARCINOMAS OF LIVER (DISORDER)
C1391911|T191||SNOMEDCT_US|BILE DUCT; CARCINOMA, WITH HEPATOCELLULAR CARCINOMA
C1391911|T191||SNOMEDCT_US|CARCINOMA; BILE DUCT, WITH HEPATOCELLULAR CARCINOMA
C1391911|T191||SNOMEDCT_US|CARCINOMA; HEPATOCELLULAR, WITH BILE DUCT CARCINOMA
C1391911|T191||SNOMEDCT_US|HEPATOCELLULAR; CARCINOMA, WITH BILE DUCT CARCINOMA
C1391914|T191||SNOMEDCT_US|CARCINOMA; HEPATOCHOLANGIOLITIC
C1391914|T191||SNOMEDCT_US|HEPATOCHOLANGIOLITIC; CARCINOMA
C1336811|T191||SNOMEDCT_US|TRANSPLANT-RELATED HEPATOCELLULAR CARCINOMA
C1333067|T191||SNOMEDCT_US|CLEAR CELL CARCINOMA OF LIVER CELLS
C1333067|T191||SNOMEDCT_US|CLEAR CELL CARCINOMA OF THE LIVER CELLS
C1333067|T191||SNOMEDCT_US|CLEAR CELL HEPATOCELLULAR CARCINOMA
C1333067|T191||SNOMEDCT_US|HEPATOCELLULAR CLEAR CELL CARCINOMA
C1333067|T191||SNOMEDCT_US|LIVER CELL CLEAR CELL CARCINOMA
C0279606|T191||SNOMEDCT_US|CHILDHOOD HEPATOCELLULAR CARCINOMA
C0279606|T191||SNOMEDCT_US|CARCINOMA, HEPATOCELLULAR, CHILDHOOD
C0279606|T191||SNOMEDCT_US|HEPATOCELLULAR CARCINOMA, CHILDHOOD
C0279606|T191||SNOMEDCT_US|PEDIATRIC HEPATOCELLULAR CARCINOMA
C0279606|T191||SNOMEDCT_US|CHILDHOOD HEPATOMA
C0279606|T191||SNOMEDCT_US|CHILDHOOD LIVER CELL CARCINOMA
C0279606|T191||SNOMEDCT_US|PEDIATRIC CARCINOMA OF LIVER CELL
C0279606|T191||SNOMEDCT_US|PEDIATRIC CARCINOMA OF THE LIVER CELL
C0279606|T191||SNOMEDCT_US|PEDIATRIC HEPATOMA
C0279606|T191||SNOMEDCT_US|PEDIATRIC LIVER CELL CARCINOMA
C0279606|T191||SNOMEDCT_US|CHILDHOOD CARCINOMA OF LIVER CELL
C0279606|T191||SNOMEDCT_US|CHILDHOOD CARCINOMA OF THE LIVER CELL
C1112459|T191||SNOMEDCT_US|LIVER CELL CARCINOMA NON-RESECTABLE
C1112459|T191||SNOMEDCT_US|HEPATOCELLULAR CARCINOMA NON-RESECTABLE
C1112459|T191||SNOMEDCT_US|NON-RESECTABLE HEPATOCELLULAR CARCINOMA
C0861876|T191||SNOMEDCT_US|LIVER CARCINOMA RECURRENT
C0861876|T191||SNOMEDCT_US|CARCINOMA LIVER RECURRENT
C0861876|T191||SNOMEDCT_US|HEPATOMA RECURRENT
C0861876|T191||SNOMEDCT_US|HEPATOCELLULAR CARCINOMA RECURRENT
C0861876|T191||SNOMEDCT_US|LIVER CELL CARCINOMA RECURRENT
C0861876|T191||SNOMEDCT_US|MALIGNANT HEPATOMA RECURRENT
C0861876|T191||SNOMEDCT_US|HEPATOCELLULAR CARCINOMA, RECURRENT
C0861876|T191||SNOMEDCT_US|RECURRENT CARCINOMA OF LIVER CELL
C0861876|T191||SNOMEDCT_US|RECURRENT CARCINOMA OF THE LIVER CELL
C0861876|T191||SNOMEDCT_US|RECURRENT HEPATOCELLULAR CARCINOMA
C0861876|T191||SNOMEDCT_US|RECURRENT HEPATOMA
C0861876|T191||SNOMEDCT_US|RECURRENT LIVER CELL CARCINOMA
C0861876|T191||SNOMEDCT_US|RELAPSED CARCINOMA OF LIVER CELL
C0861876|T191||SNOMEDCT_US|RELAPSED CARCINOMA OF THE LIVER CELL
C0861876|T191||SNOMEDCT_US|RELAPSED HEPATOCELLULAR CARCINOMA
C0861876|T191||SNOMEDCT_US|RELAPSED HEPATOMA
C0861876|T191||SNOMEDCT_US|RELAPSED LIVER CELL CARCINOMA
C1332222|T191||SNOMEDCT_US|AFLATOXINS-RELATED HEPATOCELLULAR CARCINOMA
C1710014|T191||SNOMEDCT_US|SARCOMATOID HEPATOCELLULAR CARCINOMA
C1710014|T191||SNOMEDCT_US|SARCOMATOUS HEPATOCELLULAR CARCINOMA
C1709568|T191||SNOMEDCT_US|PLEOMORPHIC HEPATOCELLULAR CARCINOMA
C1266018|T191|128646008|SNOMEDCT_US|SCLEROSING HEPATOCELLULAR CARCINOMA|SCLEROSING HEPATIC CARCINOMA
C1266018|T191|128646008|SNOMEDCT_US|SCIRRHOUS HEPATOCELLULAR CARCINOMA|SCLEROSING HEPATIC CARCINOMA
C1266018|T191|128646008|SNOMEDCT_US|HEPATOCELLULAR CARCINOMA, SCIRRHOUS (MORPHOLOGIC ABNORMALITY)|SCLEROSING HEPATIC CARCINOMA
C1266018|T191|128646008|SNOMEDCT_US|HEPATOCELLULAR CARCINOMA, SCIRRHOUS|SCLEROSING HEPATIC CARCINOMA
C1266018|T191|128646008|SNOMEDCT_US|SCLEROSING HEPATIC CARCINOMA|SCLEROSING HEPATIC CARCINOMA
C1332228|T191||SNOMEDCT_US|ALCOHOL-RELATED HEPATOCELLULAR CARCINOMA
C1333979|T191||SNOMEDCT_US|HEPATITIS VIRUS RELATED HEPATOCELLULAR CARCINOMA
C1333979|T191||SNOMEDCT_US|HEPATITIS VIRUS-RELATED HEPATOCELLULAR CARCINOMA
C0863194|T191||SNOMEDCT_US|CARCINOMA LIVER RESECTABLE
C0863194|T191||SNOMEDCT_US|LIVER CELL CARCINOMA RESECTABLE
C0863194|T191||SNOMEDCT_US|MALIGNANT HEPATOMA RESECTABLE
C0863194|T191||SNOMEDCT_US|HEPATOMA RESECTABLE
C0863194|T191||SNOMEDCT_US|LIVER CARCINOMA RESECTABLE
C0863194|T191||SNOMEDCT_US|HEPATOCELLULAR CARCINOMA RESECTABLE
C0863194|T191||SNOMEDCT_US|HEPATOCELLULAR CARCINOMA, RESECTABLE
C0863194|T191||SNOMEDCT_US|RESECTABLE CARCINOMA OF LIVER CELL
C0863194|T191||SNOMEDCT_US|RESECTABLE CARCINOMA OF THE LIVER CELL
C0863194|T191||SNOMEDCT_US|RESECTABLE HEPATOCELLULAR CARCINOMA
C0863194|T191||SNOMEDCT_US|RESECTABLE HEPATOMA
C0863194|T191||SNOMEDCT_US|RESECTABLE LIVER CELL CARCINOMA
C2111636|T191||SNOMEDCT_US|LARGE CELL CARCINOMA OF LIVER WITH RHABDOID PHENOTYPE
C2111636|T191||SNOMEDCT_US|LARGE CELL CARCINOMA OF LIVER WITH RHABDOID PHENOTYPE 
C2075624|T191||SNOMEDCT_US|LIVER NEOPLASM MALIGNANT CLEAR CELL TYPE
C2075624|T191||SNOMEDCT_US|CLEAR CELL TYPE NEOPLASM OF LIVER 
C2075624|T191||SNOMEDCT_US|CLEAR CELL TYPE NEOPLASM OF LIVER
C2111730|T191||SNOMEDCT_US|THIS MORE LIKELY REFERS TO A DIFFERENT TYPE OF CANCER, BUT THERE ARE CASE REPORTS OF HCC STAINING NEUROENDOCRINE-LIKE, SO WILL LEAVE IT ON
C2111730|T191||SNOMEDCT_US|LARGE CELL NEUROENDOCRINE CARCINOMA OF LIVER 
