C1990758|T034|LP54274-3|LNC|INR PLATELET POOR PLASMA|INR &#X7C; PLATELET POOR PLASMA
C0005790|T034|LP7788-5|LNC| THIS WOULD BE A FULL PANEL (PT/PTT/INR)|COAG
C0525032|T034|LP20762-8|LNC|INTERNATIONAL NORMALIZED RATIO|INR
C0525032|T034|LP20762-8|LNC|INR|INR
C0525032|T034|LP20762-8|LNC|LOINC LP20762-8|INR
C0525032|T034|LP20762-8|LNC|LOINC 20762-8|INR
C2360882|T034|52129-4|LNC|COAGULATION TISSUE FACTOR INDUCED.INR^POST HEPARIN ADSORPTION:RELTIME:PT:PPP:QN:COAG|INR IN PLATELET POOR PLASMA BY COAGULATION ASSAY --POST HEPARIN ADSORPTION
C2360882|T034|52129-4|LNC|THIS IS STANDARD PROTOOL|INR IN PLATELET POOR PLASMA BY COAGULATION ASSAY --POST HEPARIN ADSORPTION
C2360882|T034|52129-4|LNC|INR P HEPARIN ADSORPTION PPP|INR IN PLATELET POOR PLASMA BY COAGULATION ASSAY --POST HEPARIN ADSORPTION
C2360882|T034|52129-4|LNC|COAGULATION TISSUE FACTOR INDUCED.INR^POST HEPARIN ADSORPTION:RELATIVE TIME:POINT IN TIME:PLATELET POOR PLASMA:QUANTITATIVE:COAGULATION ASSAY|INR IN PLATELET POOR PLASMA BY COAGULATION ASSAY --POST HEPARIN ADSORPTION
C0482691|T034|6301-6|LNC|INR IN PLATELET POOR PLASMA BY COAGULATION ASSAY|INR PPP
C0482691|T034|6301-6|LNC|INR PPP|INR PPP
C0482691|T034|6301-6|LNC|COAGULATION TISSUE FACTOR INDUCED.INR:RELTIME:PT:PPP:QN:COAG|INR PPP
C0482691|T034|6301-6|LNC|COAGULATION TISSUE FACTOR INDUCED.INR:RELATIVE TIME:POINT IN TIME:PLATELET POOR PLASMA:QUANTITATIVE:COAGULATION ASSAY|INR PPP
C0525032|T034|LP20762-8|LNC|INTERNATIONAL NORMALIZED RATIO|INR
C0525032|T034|LP20762-8|LNC|INTERNATIONAL NORMALIZED RATIOS|INR
C0525032|T034|LP20762-8|LNC|NORMALIZED RATIO, INTERNATIONAL|INR
C0525032|T034|LP20762-8|LNC|NORMALIZED RATIOS, INTERNATIONAL|INR
C0525032|T034|LP20762-8|LNC|RATIO, INTERNATIONAL NORMALIZED|INR
C0525032|T034|LP20762-8|LNC|RATIOS, INTERNATIONAL NORMALIZED|INR
C0525032|T034|LP20762-8|LNC|INR|INR
C0525032|T034|LP20762-8|LNC|INTERNATIONAL NORMALIZED RATIO (INR)|INR
C0525032|T034|LP20762-8|LNC|INTERNATIONAL NORMALIZED RATIO (INR) |INR
C0525032|T034|LP20762-8|LNC|INTERNATIONAL NORMALISED RATIO|INR
C0525032|T034|LP20762-8|LNC|COAGULATION STUDIES: INR|INR
C0525032|T034|LP20762-8|LNC|INTERNATIONAL NORMALISED RATIO |INR
C0525032|T034|LP20762-8|LNC|PROTHROMBIN INTL. NORMALIZED RATIO|INR
C0525032|T034|LP20762-8|LNC|INR (INTERNATIONAL NORMALISED RATIO)|INR
C0525032|T034|LP20762-8|LNC|INR (INTERNATIONAL NORMALIZED RATIO)|INR
C0525032|T034|LP20762-8|LNC|INTERNATIONAL NORMALIZED RATIO (QUALIFIER VALUE)|INR
C0525032|T034|LP20762-8|LNC|INR - INTERNATIONALISED RATIO|INR
C0525032|T034|LP20762-8|LNC|INTERNATIONALISED RATIO|INR
C0525032|T034|LP20762-8|LNC|INTERNATIONAL NORMALIZED RATIO (OBSERVABLE ENTITY)|INR
C0525032|T034|LP20762-8|LNC|INR - INTERNATIONALIZED RATIO|INR
C0525032|T034|LP20762-8|LNC|INTERNATIONALIZED RATIO|INR
C0486259|T034|5895-7|LNC|COAGULATION TISSUE FACTOR INDUCED.INR:TRTO:PT:PLAS:QN:COAG|DEPRECATED INR PLAS
C0486259|T034|5895-7|LNC|DEPRECATED INR PLAS|DEPRECATED INR PLAS
C0486259|T034|5895-7|LNC|COAGULATION TISSUE FACTOR INDUCED.INR:TIME RATIO:POINT IN TIME:PLASMA:QUANTITATIVE:COAGULATION ASSAY|DEPRECATED INR PLAS
C0482772|T034|3289-6|LNC|PROTHROMBIN.ACTIVITY ACTUAL/NORMAL:RELTIME:PT:PPP:QN:COAG|PROTHROM ACT/NOR PPP
C0482772|T034|3289-6|LNC|PROTHROM ACT/NOR PPP|PROTHROM ACT/NOR PPP
C0482772|T034|3289-6|LNC|PROTHROMBIN ACTIVITY ACTUAL/NORMAL IN PLATELET POOR PLASMA BY COAGULATION ASSAY|PROTHROM ACT/NOR PPP
C0482772|T034|3289-6|LNC|PROTHROMBIN.ACTIVITY ACTUAL/NORMAL:RELATIVE TIME:POINT IN TIME:PLATELET POOR PLASMA:QUANTITATIVE:COAGULATION ASSAY|PROTHROM ACT/NOR PPP
C0943508|T034|27813-5|LNC|PROTHROMBIN AG ACTUAL/NORMAL IN PLATELET POOR PLASMA BY IMMUNOLOGIC METHOD|PROTHROMBIN AG ACTUAL/NORMAL IN PLATELET POOR PLASMA BY IMMUNOASSAY
C0943508|T034|27813-5|LNC|PROTHROM AG ACT/NOR PPP IMM|PROTHROMBIN AG ACTUAL/NORMAL IN PLATELET POOR PLASMA BY IMMUNOASSAY
C0943508|T034|27813-5|LNC|PROTHROMBIN AG ACTUAL/NORMAL:RELMCNC:PT:PPP:QN:IMM|PROTHROMBIN AG ACTUAL/NORMAL IN PLATELET POOR PLASMA BY IMMUNOASSAY
C0943508|T034|27813-5|LNC|PROTHROMBIN ANTIGEN ACTUAL/NORMAL:RELATIVE MASS CONCENTRATION:POINT IN TIME:PLATELET POOR PLASMA:QUANTITATIVE:IMM|PROTHROMBIN AG ACTUAL/NORMAL IN PLATELET POOR PLASMA BY IMMUNOASSAY
C1543007|T034|38875-1|LNC|INR IN PLATELET POOR PLASMA OR BLOOD BY COAGULATION ASSAY|INR PPP/BLD
C1543007|T034|38875-1|LNC|COAGULATION TISSUE FACTOR INDUCED.INR:RELTIME:PT:PPP/BLD:QN:COAG|INR PPP/BLD
C1543007|T034|38875-1|LNC|COAGULATION TISSUE FACTOR INDUCED.INR:RELATIVE TIME:POINT IN TIME:PLATELET POOR PLASMA/WHOLE BLOOD:QUANTITATIVE:COAGULATION ASSAY|INR PPP/BLD
C1543007|T034|38875-1|LNC|INR PPP/BLD|INR PPP/BLD
C1369580|T034|34714-6|LNC|INR BLD|INR BLD
C1369580|T034|34714-6|LNC|INR IN BLOOD BY COAGULATION ASSAY|INR BLD
C1369580|T034|34714-6|LNC|COAGULATION TISSUE FACTOR INDUCED.INR:RELTIME:PT:BLD:QN:COAG|INR BLD
C1369580|T034|34714-6|LNC|COAGULATION TISSUE FACTOR INDUCED.INR:RELATIVE TIME:POINT IN TIME:WHOLE BLOOD:QUANTITATIVE:COAGULATION ASSAY|INR BLD
C2584422|T034||LNC|INTERNATIONAL NORMALIZED RATIO RESULT OBTAINED USING PORTABLE INTERNATIONAL NORMALIZED RATIO MONITORING DEVICE (OBSERVABLE ENTITY)
C2584422|T034||LNC|INTERNATIONAL NORMALIZED RATIO RESULT OBTAINED USING PORTABLE INTERNATIONAL NORMALIZED RATIO MONITORING DEVICE
C2584422|T034||LNC|INTERNATIONAL NORMALISED RATIO RESULT OBTAINED USING PORTABLE INTERNATIONAL NORMALISED RATIO MONITORING DEVICE
C1254541|T034||LNC|CALCULATION OF INTERNATIONAL NORMALISED RATIO (INR)
C1254541|T034||LNC|CALCULATION OF INTERNATIONAL NORMALIZED RATIO (INR)
C1254541|T034||LNC|CALCULATION OF INTERNATIONAL NORMALISED RATIO
C1254541|T034||LNC|CALCULATION OF INTERNATIONAL NORMALIZED RATIO
C1254541|T034||LNC|CALCULATION OF INTERNATIONAL NORMALIZED RATIO 
C1254541|T034||LNC|INTERNATIONAL NORMALIZED RATIO (INR) CALCULATIONS
C3838119|T034||LNC|COAGULATION STUDIES: INR IN BLOOD OR PLATELET-POOR PLASMA 
C3838119|T034||LNC|COAGULATION STUDIES: INR IN BLOOD OR PLATELET-POOR PLASMA
