C0017725|T034|LP32534-7|LNC|GLUCOSE|GLUCOSE
C0364479|T034|2339-0|LNC|GLUCOSE|GLUCOSE [MASS/VOLUME] IN BLOOD
C0364479|T034|2339-0|LNC|GLUCOSE:MCNC:PT:BLD:QN|GLUCOSE [MASS/VOLUME] IN BLOOD
C0337438|T034||LNC|GLUCOSE
C0337438|T034||LNC|GLUCOSE MEASUREMENT
C0337438|T034||LNC|TEST;GLUCOSE
C0337438|T034||LNC|MEASUREMENT OF GLUCOSE
C0337438|T034||LNC|GLUCOSE MEASUREMENT 
C0337438|T034||LNC|GLUCOSE MEASUREMENT, NOS
C0337438|T034||LNC|GLUCOSE TEST
C0523658|T034||LNC|ASSAY GLUCOSE BLOOD QUANT
C0523658|T034||LNC|GLUCOSE; QUANTITATIVE, BLOOD (EXCEPT REAGENT STRIP)
C0523658|T034||LNC|GLUCOSE QUANTITATIVE BLOOD XCPT REAGENT STRIP
C0523658|T034||LNC|GLUCOSE MEASUREMENT, QUANTITATIVE
C0523658|T034||LNC|GLUCOSE MEASUREMENT, QUANTITATIVE 
C0202045|T034||LNC|GLUCOSE MEASUREMENT, FASTING
C0428568|T034||LNC|FASTING BLOOD GLUCOSE MEASUREMENT
C0005802|T034||LNC|BLOOD GLUCOSE
C0005802|T034||LNC|SUGAR, BLOOD
C0005802|T034||LNC|BLOOD SUGAR
C0005802|T034||LNC|BLOOD GLUCOSE [CHEMICAL/INGREDIENT]
C0005802|T034||LNC|GLUCOSE, BLOOD
C0017725|T034|LP32534-7|LNC|GLUCOSE|GLUCOSE
C0017725|T034|LP32534-7|LNC|GLUCOSE [CHEMICAL/INGREDIENT]|GLUCOSE
C0017725|T034|LP32534-7|LNC|GLUCOSE [ENDOCRINE]|GLUCOSE
C0017725|T034|LP32534-7|LNC|GLUCOSE [ENDOCRINE] |GLUCOSE
C0017725|T034|LP32534-7|LNC|GLUCOSE |GLUCOSE
C0017725|T034|LP32534-7|LNC|GLUCOSE PREPARATION |GLUCOSE
C0017725|T034|LP32534-7|LNC|GLUCOSE, NOS|GLUCOSE
C0017725|T034|LP32534-7|LNC|GLUCOSE [ENDOCRINE] |GLUCOSE
C1644627|T034|41604-0|LNC|GLUCOSE P FAST BLDC GLUCOMTR-MCNC|FASTING GLUCOSE [MASS/VOLUME] IN CAPILLARY BLOOD BY GLUCOMETER
C1644627|T034|41604-0|LNC|GLUCOSE^POST CFST:MCNC:PT:BLDC:QN:GLUCOMETER|FASTING GLUCOSE [MASS/VOLUME] IN CAPILLARY BLOOD BY GLUCOMETER
C1644627|T034|41604-0|LNC|FASTING GLUCOSE [MASS/VOLUME] IN CAPILLARY BLOOD BY GLUCOMETER|FASTING GLUCOSE [MASS/VOLUME] IN CAPILLARY BLOOD BY GLUCOMETER
C1644627|T034|41604-0|LNC|GLUCOSE^POST CALORIE FAST:MASS CONCENTRATION:POINT IN TIME:BLOOD CAPILLARY:QUANTITATIVE:GLUCOMETER|FASTING GLUCOSE [MASS/VOLUME] IN CAPILLARY BLOOD BY GLUCOMETER
C0363687|T034|1556-0|LNC|GLUCOSE^POST CFST:MCNC:PT:BLDC:QN|FASTING GLUCOSE [MASS/VOLUME] IN CAPILLARY BLOOD
C0363687|T034|1556-0|LNC|FASTING GLUCOSE [MASS/VOLUME] IN CAPILLARY BLOOD|FASTING GLUCOSE [MASS/VOLUME] IN CAPILLARY BLOOD
C0363687|T034|1556-0|LNC|GLUCOSE P FAST BLDC-MCNC|FASTING GLUCOSE [MASS/VOLUME] IN CAPILLARY BLOOD
C0363687|T034|1556-0|LNC|GLUCOSE^POST CALORIE FAST:MASS CONCENTRATION:POINT IN TIME:BLOOD CAPILLARY:QUANTITATIVE|FASTING GLUCOSE [MASS/VOLUME] IN CAPILLARY BLOOD
C2706820|T034|54257-1|LNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --PRE DOSE INSULIN IV|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --PRE DOSE INSULIN IV
C2706820|T034|54257-1|LNC|GLUCOSE PRE INS IV SERPL-SCNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --PRE DOSE INSULIN IV
C2706820|T034|54257-1|LNC|GLUCOSE^PRE DOSE INSULIN INTRAVENOUS:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --PRE DOSE INSULIN IV
C1988482|T034|LP51365-2|LNC|GLUCOSE &#X7C; BLOOD ARTERIAL|GLUCOSE &#X7C; BLOOD ARTERIAL
C2361582|T034|53094-9|LNC|GLUCOSE^POST MEAL:SCNC:PT:SER/PLAS:QN|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --POST MEAL
C2361582|T034|53094-9|LNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --POST MEAL|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --POST MEAL
C2361582|T034|53094-9|LNC|GLUCOSE^POST MEAL:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --POST MEAL
C0484599|T034|10450-5|LNC|GLUCOSE^POST 10H CFST:MCNC:PT:SER/PLAS:QN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --10 HOURS FASTING
C0484599|T034|10450-5|LNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --10 HOURS FASTING|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --10 HOURS FASTING
C0484599|T034|10450-5|LNC|GLUCOSE^POST 10H CALORIE FAST:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --10 HOURS FASTING
C0484599|T034|10450-5|LNC|GLUCOSE P 10H FAST SERPL-MCNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --10 HOURS FASTING
C0799333|T034|16168-7|LNC|GLUCOSE^3 PM SPECIMEN:MCNC:PT:SER/PLAS:QN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --3 PM SPECIMEN
C0799333|T034|16168-7|LNC|GLUCOSE 3 PM SERPL-MCNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --3 PM SPECIMEN
C0799333|T034|16168-7|LNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --3 PM SPECIMEN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --3 PM SPECIMEN
C0799333|T034|16168-7|LNC|GLUCOSE^3 PM SPECIMEN:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --3 PM SPECIMEN
C0799334|T034|16169-5|LNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --4 PM SPECIMEN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --4 PM SPECIMEN
C0799334|T034|16169-5|LNC|GLUCOSE^4 PM SPECIMEN:MCNC:PT:SER/PLAS:QN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --4 PM SPECIMEN
C0799334|T034|16169-5|LNC|GLUCOSE 4 PM SERPL-MCNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --4 PM SPECIMEN
C0799334|T034|16169-5|LNC|GLUCOSE^4 PM SPECIMEN:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --4 PM SPECIMEN
C0797943|T034|14769-4|LNC|GLUCOSE^PRE 12H CFST:SCNC:PT:SER/PLAS:QN|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --PRE 12 HOUR FAST
C0797943|T034|14769-4|LNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --PRE 12 HOUR FAST|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --PRE 12 HOUR FAST
C0797943|T034|14769-4|LNC|GLUCOSE^PRE 12 HOURS CALORIE FAST:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --PRE 12 HOUR FAST
C0797943|T034|14769-4|LNC|GLUCOSE PRE 12H FAST SERPL-SCNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --PRE 12 HOUR FAST
C2923563|T034|59814-4|LNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --7 AM SPECIMEN|GLUCOSE^7 AM SPECIMEN:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE
C2923563|T034|59814-4|LNC|GLUCOSE^7 AM SPECIMEN:SCNC:PT:SER/PLAS:QN|GLUCOSE^7 AM SPECIMEN:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE
C2923563|T034|59814-4|LNC|GLUCOSE 7 AM SERPL-SCNC|GLUCOSE^7 AM SPECIMEN:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE
C2923563|T034|59814-4|LNC|GLUCOSE^7 AM SPECIMEN:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE^7 AM SPECIMEN:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE
C1716223|T034|45056-9|LNC|GLUCOSE^8 PM SPECIMEN:SCNC:PT:SER/PLAS:QN|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --8 PM SPECIMEN
C1716223|T034|45056-9|LNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --8 PM SPECIMEN|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --8 PM SPECIMEN
C1716223|T034|45056-9|LNC|GLUCOSE 8 PM SERPL-SCNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --8 PM SPECIMEN
C1716223|T034|45056-9|LNC|GLUCOSE^8 PM SPECIMEN:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --8 PM SPECIMEN
C1988485|T034|LP51830-5|LNC|GLUCOSE &#X7C; BLOOD VENOUS|GLUCOSE &#X7C; BLOOD VENOUS
C2706825|T034|54262-1|LNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --3 HOURS PRE DOSE INSULIN IV|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --3 HOURS PRE DOSE INSULIN IV
C2706825|T034|54262-1|LNC|GLUCOSE^3H PRE DOSE INSULIN IV:SCNC:PT:SER/PLAS:QN|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --3 HOURS PRE DOSE INSULIN IV
C2706825|T034|54262-1|LNC|GLUCOSE^3 HOURS PRE DOSE INSULIN INTRAVENOUS:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --3 HOURS PRE DOSE INSULIN IV
C2706825|T034|54262-1|LNC|GLUCOSE 3H PRE INS IV SERPL-SCNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --3 HOURS PRE DOSE INSULIN IV
C1988483|T034|LP43629-2|LNC|GLUCOSE &#X7C; BLOOD CAPILLARY|GLUCOSE &#X7C; BLOOD CAPILLARY
C1716203|T034|45052-8|LNC|GLUCOSE 12 AM SERPL-SCNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --12 AM SPECIMEN
C1716203|T034|45052-8|LNC|GLUCOSE^12 AM SPECIMEN:SCNC:PT:SER/PLAS:QN|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --12 AM SPECIMEN
C1716203|T034|45052-8|LNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --12 AM SPECIMEN|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --12 AM SPECIMEN
C1716203|T034|45052-8|LNC|GLUCOSE^12 AM SPECIMEN:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --12 AM SPECIMEN
C1716205|T034|45054-4|LNC|GLUCOSE^12 PM SPECIMEN:SCNC:PT:SER/PLAS:QN|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --12 PM SPECIMEN
C1716205|T034|45054-4|LNC|GLUCOSE 12 PM SERPL-SCNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --12 PM SPECIMEN
C1716205|T034|45054-4|LNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --12 PM SPECIMEN|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --12 PM SPECIMEN
C1716205|T034|45054-4|LNC|GLUCOSE^12 PM SPECIMEN:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --12 PM SPECIMEN
C1952717|T034|48986-4|LNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --8 AM SPECIMEN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --8 AM SPECIMEN
C1952717|T034|48986-4|LNC|GLUCOSE^8 AM SPECIMEN:MCNC:PT:SER/PLAS:QN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --8 AM SPECIMEN
C1952717|T034|48986-4|LNC|GLUCOSE 8 AM SERPL-MCNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --8 AM SPECIMEN
C1952717|T034|48986-4|LNC|GLUCOSE^8 AM SPECIMEN:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --8 AM SPECIMEN
C0482544|T034|1558-6|LNC|FASTING GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA|FASTING GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA
C0482544|T034|1558-6|LNC|GLUCOSE P FAST SERPL-MCNC|FASTING GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA
C0482544|T034|1558-6|LNC|GLUCOSE^POST CALORIE FAST:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|FASTING GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA
C2607838|T034|35184-1|LNC|GLUCOSE [MASS OR MOLECULES/VOLUME] IN SERUM OR PLASMA --POST CFST|FASTING GLUCOSE [MASS OR MOLES/VOLUME] IN SERUM OR PLASMA
C2607838|T034|35184-1|LNC|GLUCOSE P FAST SERPL-MSCNC|FASTING GLUCOSE [MASS OR MOLES/VOLUME] IN SERUM OR PLASMA
C2607838|T034|35184-1|LNC|GLUCOSE^POST CFST:MSCNC:PT:SER/PLAS:QN|FASTING GLUCOSE [MASS OR MOLES/VOLUME] IN SERUM OR PLASMA
C2607838|T034|35184-1|LNC|FASTING GLUCOSE [MASS OR MOLES/VOLUME] IN SERUM OR PLASMA|FASTING GLUCOSE [MASS OR MOLES/VOLUME] IN SERUM OR PLASMA
C2607838|T034|35184-1|LNC|GLUCOSE^POST CALORIE FAST:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|FASTING GLUCOSE [MASS OR MOLES/VOLUME] IN SERUM OR PLASMA
C1952721|T034|48989-8|LNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --6 PM SPECIMEN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --6 PM SPECIMEN
C1952721|T034|48989-8|LNC|GLUCOSE^6 PM SPECIMEN:MCNC:PT:SER/PLAS:QN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --6 PM SPECIMEN
C1952721|T034|48989-8|LNC|GLUCOSE 6 PM SERPL-MCNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --6 PM SPECIMEN
C1952721|T034|48989-8|LNC|GLUCOSE^6 PM SPECIMEN:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --6 PM SPECIMEN
C1954699|T034|48992-2|LNC|GLUCOSE^12 AM SPECIMEN:MCNC:PT:SER/PLAS:QN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --12 AM SPECIMEN
C1954699|T034|48992-2|LNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --12 AM SPECIMEN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --12 AM SPECIMEN
C1954699|T034|48992-2|LNC|GLUCOSE 12 AM SERPL-MCNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --12 AM SPECIMEN
C1954699|T034|48992-2|LNC|GLUCOSE^12 AM SPECIMEN:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --12 AM SPECIMEN
C2706819|T034|54256-3|LNC|GLUCOSE 8M P GC SERPL-SCNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --8 MINUTES POST DOSE GLUCAGON
C2706819|T034|54256-3|LNC|GLUCOSE^8M POST DOSE GLUCAGON:SCNC:PT:SER/PLAS:QN|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --8 MINUTES POST DOSE GLUCAGON
C2706819|T034|54256-3|LNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --8 MINUTES POST DOSE GLUCAGON|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --8 MINUTES POST DOSE GLUCAGON
C2706819|T034|54256-3|LNC|GLUCOSE^8 MINUTES POST DOSE GLUCAGON:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --8 MINUTES POST DOSE GLUCAGON
C2706827|T034|54264-7|LNC|GLUCOSE^45M POST DOSE INSULIN INTRAVENOUS:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --45 MINUTES POST DOSE INSULIN IV
C2706827|T034|54264-7|LNC|GLUCOSE^45M POST DOSE INSULIN IV:SCNC:PT:SER/PLAS:QN|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --45 MINUTES POST DOSE INSULIN IV
C2706827|T034|54264-7|LNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --45 MINUTES POST DOSE INSULIN IV|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --45 MINUTES POST DOSE INSULIN IV
C2706827|T034|54264-7|LNC|GLUCOSE 45M P INS IV SERPL-SCNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --45 MINUTES POST DOSE INSULIN IV
C2598578|T034|53474-3|LNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --4 AM SPECIMEN|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --4 AM SPECIMEN
C2598578|T034|53474-3|LNC|GLUCOSE^4 AM SPECIMEN:SCNC:PT:SER/PLAS:QN|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --4 AM SPECIMEN
C2598578|T034|53474-3|LNC|GLUCOSE 4 AM SPECIMEN SERPL-SCNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --4 AM SPECIMEN
C2598578|T034|53474-3|LNC|GLUCOSE^4 AM SPECIMEN:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --4 AM SPECIMEN
C0799332|T034|16167-9|LNC|GLUCOSE 2 PM SERPL-MCNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --2 PM SPECIMEN
C0799332|T034|16167-9|LNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --2 PM SPECIMEN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --2 PM SPECIMEN
C0799332|T034|16167-9|LNC|GLUCOSE^2 PM SPECIMEN:MCNC:PT:SER/PLAS:QN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --2 PM SPECIMEN
C0799332|T034|16167-9|LNC|GLUCOSE^2 PM SPECIMEN:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --2 PM SPECIMEN
C0363685|T034|1554-5|LNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --12 HOURS FASTING|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --12 HOURS FASTING
C0363685|T034|1554-5|LNC|GLUCOSE^POST 12H CFST:MCNC:PT:SER/PLAS:QN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --12 HOURS FASTING
C0363685|T034|1554-5|LNC|GLUCOSE^POST 12 HOURS CALORIE FAST:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --12 HOURS FASTING
C0363685|T034|1554-5|LNC|GLUCOSE P 12H FAST SERPL-MCNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --12 HOURS FASTING
C0797934|T034|14760-3|LNC|GLUCOSE^2H POST MEAL:SCNC:PT:BLDC:QN|GLUCOSE [MOLES/VOLUME] IN CAPILLARY BLOOD --2 HOURS POST MEAL
C0797934|T034|14760-3|LNC|GLUCOSE [MOLES/VOLUME] IN CAPILLARY BLOOD --2 HOURS POST MEAL|GLUCOSE [MOLES/VOLUME] IN CAPILLARY BLOOD --2 HOURS POST MEAL
C0797934|T034|14760-3|LNC|GLUCOSE^2 HOURS POST MEAL:SUBSTANCE CONCENTRATION:POINT IN TIME:BLOOD CAPILLARY:QUANTITATIVE|GLUCOSE [MOLES/VOLUME] IN CAPILLARY BLOOD --2 HOURS POST MEAL
C0797934|T034|14760-3|LNC|GLUCOSE 2H P MEAL BLDC-SCNC|GLUCOSE [MOLES/VOLUME] IN CAPILLARY BLOOD --2 HOURS POST MEAL
C0797945|T034|14771-0|LNC|FASTING GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA|FASTING GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA
C0797945|T034|14771-0|LNC|GLUCOSE^POST CFST:SCNC:PT:SER/PLAS:QN|FASTING GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA
C0797945|T034|14771-0|LNC|GLUCOSE P FAST SERPL-SCNC|FASTING GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA
C0797945|T034|14771-0|LNC|GLUCOSE^POST CALORIE FAST:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|FASTING GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA
C2923561|T034|59812-8|LNC|GLUCOSE^11 AM SPECIMEN:SCNC:PT:SER/PLAS:QN|GLUCOSE^11 AM SPECIMEN:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE
C2923561|T034|59812-8|LNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --11 AM SPECIMEN|GLUCOSE^11 AM SPECIMEN:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE
C2923561|T034|59812-8|LNC|GLUCOSE 11 AM SERPL-SCNC|GLUCOSE^11 AM SPECIMEN:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE
C2923561|T034|59812-8|LNC|GLUCOSE^11 AM SPECIMEN:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE^11 AM SPECIMEN:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE
C1988481|T034|LP42107-0|LNC|GLUCOSE &#X7C; BLD-SER-PLAS|GLUCOSE &#X7C; BLD-SER-PLAS
C1952722|T034|48990-6|LNC|GLUCOSE 8 PM SERPL-MCNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --8 PM SPECIMEN
C1952722|T034|48990-6|LNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --8 PM SPECIMEN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --8 PM SPECIMEN
C1952722|T034|48990-6|LNC|GLUCOSE^8 PM SPECIMEN:MCNC:PT:SER/PLAS:QN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --8 PM SPECIMEN
C1952722|T034|48990-6|LNC|GLUCOSE^8 PM SPECIMEN:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --8 PM SPECIMEN
C1954698|T034|48991-4|LNC|GLUCOSE 10 PM SERPL-MCNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --10 PM SPECIMEN
C1954698|T034|48991-4|LNC|GLUCOSE^10 PM SPECIMEN:MCNC:PT:SER/PLAS:QN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --10 PM SPECIMEN
C1954698|T034|48991-4|LNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --10 PM SPECIMEN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --10 PM SPECIMEN
C1954698|T034|48991-4|LNC|GLUCOSE^10 PM SPECIMEN:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --10 PM SPECIMEN
C1716206|T034|45055-1|LNC|GLUCOSE^4 PM SPECIMEN:SCNC:PT:SER/PLAS:QN|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --4 PM SPECIMEN
C1716206|T034|45055-1|LNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --4 PM SPECIMEN|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --4 PM SPECIMEN
C1716206|T034|45055-1|LNC|GLUCOSE 4 PM SERPL-SCNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --4 PM SPECIMEN
C1716206|T034|45055-1|LNC|GLUCOSE^4 PM SPECIMEN:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --4 PM SPECIMEN
C2361537|T034|53049-3|LNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --PRE-MEAL|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --PRE-MEAL
C2361537|T034|53049-3|LNC|GLUCOSE^PRE-MEAL:MCNC:PT:SER/PLAS:QN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --PRE-MEAL
C2361537|T034|53049-3|LNC|GLUCOSE PRE-MEAL SERPL-MCNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --PRE-MEAL
C2361537|T034|53049-3|LNC|GLUCOSE^PRE-MEAL:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --PRE-MEAL
C2923562|T034|59813-6|LNC|GLUCOSE^7 AM SPECIMEN:SCNC:PT:BLDC:QN:GLUCOMETER|GLUCOSE^7 AM SPECIMEN:SUBSTANCE CONCENTRATION:POINT IN TIME:BLOOD CAPILLARY:QUANTITATIVE:GLUCOMETER
C2923562|T034|59813-6|LNC|GLUCOSE [MOLES/VOLUME] IN CAPILLARY BLOOD BY GLUCOMETER --7 AM SPECIMEN|GLUCOSE^7 AM SPECIMEN:SUBSTANCE CONCENTRATION:POINT IN TIME:BLOOD CAPILLARY:QUANTITATIVE:GLUCOMETER
C2923562|T034|59813-6|LNC|GLUCOSE 7 AM BLDC GLUCOMTR-SCNC|GLUCOSE^7 AM SPECIMEN:SUBSTANCE CONCENTRATION:POINT IN TIME:BLOOD CAPILLARY:QUANTITATIVE:GLUCOMETER
C2923562|T034|59813-6|LNC|GLUCOSE^7 AM SPECIMEN:SUBSTANCE CONCENTRATION:POINT IN TIME:BLOOD CAPILLARY:QUANTITATIVE:GLUCOMETER|GLUCOSE^7 AM SPECIMEN:SUBSTANCE CONCENTRATION:POINT IN TIME:BLOOD CAPILLARY:QUANTITATIVE:GLUCOMETER
C0484581|T034|10449-7|LNC|GLUCOSE^1H POST MEAL:MCNC:PT:SER/PLAS:QN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --1 HOUR POST MEAL
C0484581|T034|10449-7|LNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --1 HOUR POST MEAL|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --1 HOUR POST MEAL
C0484581|T034|10449-7|LNC|GLUCOSE^1 HOUR POST MEAL:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --1 HOUR POST MEAL
C0484581|T034|10449-7|LNC|GLUCOSE 1H P MEAL SERPL-MCNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --1 HOUR POST MEAL
C0799330|T034|16165-3|LNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --10 AM SPECIMEN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --10 AM SPECIMEN
C0799330|T034|16165-3|LNC|GLUCOSE 10 AM SERPL-MCNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --10 AM SPECIMEN
C0799330|T034|16165-3|LNC|GLUCOSE^10 AM SPECIMEN:MCNC:PT:SER/PLAS:QN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --10 AM SPECIMEN
C0799330|T034|16165-3|LNC|GLUCOSE^10 AM SPECIMEN:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --10 AM SPECIMEN
C0797935|T034|14761-1|LNC|GLUCOSE^2H POST MEAL:SCNC:PT:SER/PLAS:QN|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --2 HOURS POST MEAL
C0797935|T034|14761-1|LNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --2 HOURS POST MEAL|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --2 HOURS POST MEAL
C0797935|T034|14761-1|LNC|GLUCOSE^2 HOURS POST MEAL:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --2 HOURS POST MEAL
C0797935|T034|14761-1|LNC|GLUCOSE 2H P MEAL SERPL-SCNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --2 HOURS POST MEAL
C0797942|T034|14768-6|LNC|GLUCOSE BS SERPL-SCNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --BASELINE
C0797942|T034|14768-6|LNC|GLUCOSE^BASELINE:SCNC:PT:SER/PLAS:QN|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --BASELINE
C0797942|T034|14768-6|LNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --BASELINE|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --BASELINE
C0797942|T034|14768-6|LNC|GLUCOSE^BASELINE:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --BASELINE
C1544263|T034|40287-5|LNC|GLUCOSE^1H POST MEAL:SCNC:PT:SER/PLAS:QN|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --1 HOUR POST MEAL
C1544263|T034|40287-5|LNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --1 HOUR POST MEAL|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --1 HOUR POST MEAL
C1544263|T034|40287-5|LNC|GLUCOSE^1 HOUR POST MEAL:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --1 HOUR POST MEAL
C1544263|T034|40287-5|LNC|GLUCOSE 1H P MEAL SERPL-SCNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --1 HOUR POST MEAL
C0800049|T034|16915-1|LNC|GLUCOSE^POST MEAL:MCNC:PT:SER/PLAS:QN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --POST MEAL
C0800049|T034|16915-1|LNC|GLUCOSE P MEAL SERPL-MCNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --POST MEAL
C0800049|T034|16915-1|LNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --POST MEAL|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --POST MEAL
C0800049|T034|16915-1|LNC|GLUCOSE^POST MEAL:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --POST MEAL
C0363688|T034|1557-8|LNC|GLUCOSE^POST CFST:MCNC:PT:BLDV:QN|FASTING GLUCOSE [MASS/VOLUME] IN VENOUS BLOOD
C0363688|T034|1557-8|LNC|GLUCOSE P FAST BLDV-MCNC|FASTING GLUCOSE [MASS/VOLUME] IN VENOUS BLOOD
C0363688|T034|1557-8|LNC|FASTING GLUCOSE [MASS/VOLUME] IN VENOUS BLOOD|FASTING GLUCOSE [MASS/VOLUME] IN VENOUS BLOOD
C0363688|T034|1557-8|LNC|GLUCOSE^POST CALORIE FAST:MASS CONCENTRATION:POINT IN TIME:BLOOD VENOUS:QUANTITATIVE|FASTING GLUCOSE [MASS/VOLUME] IN VENOUS BLOOD
C1544179|T034|40193-5|LNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --PRE-MEAL|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --PRE-MEAL
C1544179|T034|40193-5|LNC|GLUCOSE PRE-MEAL SERPL-SCNC|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --PRE-MEAL
C1544179|T034|40193-5|LNC|GLUCOSE^PRE-MEAL:SCNC:PT:SER/PLAS:QN|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --PRE-MEAL
C1544179|T034|40193-5|LNC|GLUCOSE^PRE-MEAL:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MOLES/VOLUME] IN SERUM OR PLASMA --PRE-MEAL
C1954701|T034|48994-8|LNC|GLUCOSE 6 AM SERPL-MCNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --6 AM SPECIMEN
C1954701|T034|48994-8|LNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --6 AM SPECIMEN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --6 AM SPECIMEN
C1954701|T034|48994-8|LNC|GLUCOSE^6 AM SPECIMEN:MCNC:PT:SER/PLAS:QN|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --6 AM SPECIMEN
C1954701|T034|48994-8|LNC|GLUCOSE^6 AM SPECIMEN:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA --6 AM SPECIMEN
C2602566|T034|LP71758-4|LNC|ESTIMATED AVERAGE GLUCOSE &#X7C; BLD-SER-PLAS|ESTIMATED AVERAGE GLUCOSE &#X7C; BLD-SER-PLAS
C4036718|T034|77677-3|LNC|GLUCOSE^2H POST MEAL:SCNC:PT:SER/PLAS/BLD:QN|GLUCOSE [MOLES/VOLUME] IN SERUM, PLASMA OR BLOOD --2 HOURS POST MEAL
C4036718|T034|77677-3|LNC|GLUCOSE^2 HOURS POST MEAL:SUBSTANCE CONCENTRATION:POINT IN TIME:SERUM/PLASMA/WHOLE BLOOD:QUANTITATIVE|GLUCOSE [MOLES/VOLUME] IN SERUM, PLASMA OR BLOOD --2 HOURS POST MEAL
C4036718|T034|77677-3|LNC|GLUCOSE [MOLES/VOLUME] IN SERUM, PLASMA OR BLOOD --2 HOURS POST MEAL|GLUCOSE [MOLES/VOLUME] IN SERUM, PLASMA OR BLOOD --2 HOURS POST MEAL
C4036718|T034|77677-3|LNC|GLUCOSE 2H P MEAL SERPLBLD-SCNC|GLUCOSE [MOLES/VOLUME] IN SERUM, PLASMA OR BLOOD --2 HOURS POST MEAL
C0364479|T034|2339-0|LNC|GLUCOSE:MCNC:PT:BLD:QN|GLUCOSE [MASS/VOLUME] IN BLOOD
C0364479|T034|2339-0|LNC|GLUCOSE [MASS/VOLUME] IN BLOOD|GLUCOSE [MASS/VOLUME] IN BLOOD
C0364479|T034|2339-0|LNC|GLUCOSE BLD-MCNC|GLUCOSE [MASS/VOLUME] IN BLOOD
C0364479|T034|2339-0|LNC|GLUCOSE:MASS CONCENTRATION:POINT IN TIME:WHOLE BLOOD:QUANTITATIVE|GLUCOSE [MASS/VOLUME] IN BLOOD
C0523660|T034||LNC|GLUCOSE MEASUREMENT, POST GLUCOSE DOSE
C0523660|T034||LNC|GLUCOSE MEASUREMENT, POST GLUCOSE DOSE 
C0337438|T034||LNC|GLUCOSE
C0337438|T034||LNC|GLUCOSE MEASUREMENT
C0337438|T034||LNC|TEST;GLUCOSE
C0337438|T034||LNC|MEASUREMENT OF GLUCOSE
C0337438|T034||LNC|GLUC
C0337438|T034||LNC|GLUCOSE MEASUREMENT 
C0337438|T034||LNC|GLUCOSE MEASUREMENT, NOS
C0337438|T034||LNC|GLUCOSE TEST
C0392201|T034||LNC|BLOOD GLUCOSE
C0392201|T034||LNC|BLOOD GLUCOSE TESTS 
C0392201|T034||LNC|BLOOD GLUCOSE TESTS
C0392201|T034||LNC|BLOOD GLUCOSE MEASUREMENT
C0392201|T034||LNC|BLOOD GLUCOSE LEVEL
C0392201|T034||LNC|BLOOD GLUCOSE MEASUREMENT 
C0392201|T034||LNC|BLOOD GLUCOSE (SUGAR) LEVEL
C0392201|T034||LNC|MEASUREMENT OF GLUCOSE IN BLOOD
C0392201|T034||LNC|BLOOD SUGAR
C0392201|T034||LNC|GLUCOSE MEASUREMENT, BLOOD
C0392201|T034||LNC|BLOOD SUGAR LEVEL
C0392201|T034||LNC|BS - BLOOD GLUCOSE LEVEL
C0392201|T034||LNC|GLUCOSE MEASUREMENT, BLOOD 
C0202048|T034||LNC|GLUCOSE MEASUREMENT BY MONITORING DEVICE
C0202048|T034||LNC|GLUCOSE MEASUREMENT BY MONITORING DEVICE 
C0202048|T034||LNC|GLUCOSE MEASUREMENT BY MONITORING DEVICE  [AMBIGUOUS]
C0204885|T034||LNC|WARD GLUCOMETER TEST
C0204885|T034||LNC|WARD GLUCOMETER TEST 
C0202041|T034||LNC|SERUM GLUCOSE
C0202041|T034||LNC|SERUM GLUCOSE MEASUREMENT
C0202041|T034||LNC|SERUM GLUCOSE TEST
C0202041|T034||LNC|GLUCOSE MEASUREMENT, SERUM
C0202041|T034||LNC|GLUCOSE MEASUREMENT, SERUM 
C0202042|T034||LNC|PLASMA GLUCOSE MEASUREMENT
C0202042|T034||LNC|PLASMA GLUCOSE MEASUREMENT 
C0202042|T034||LNC|PLASMA GLUCOSE
C0202042|T034||LNC|PLASMA GLUCOSE LEVEL
C0202042|T034||LNC|PLASMA GLUCOSE LEVEL 
C0202042|T034||LNC|GLUCOSE MEASUREMENT, PLASMA
C0202042|T034||LNC|GLUCOSE MEASUREMENT, PLASMA 
C0373621|T034||LNC|GLUCOSE TEST
C0523658|T034||LNC|ASSAY GLUCOSE BLOOD QUANT
C0523658|T034||LNC|GLUCOSE; QUANTITATIVE, BLOOD (EXCEPT REAGENT STRIP)
C0523658|T034||LNC|GLUCOSE QUANTITATIVE BLOOD XCPT REAGENT STRIP
C0523658|T034||LNC|GLUCOSE MEASUREMENT, QUANTITATIVE
C0523658|T034||LNC|GLUCOSE MEASUREMENT, QUANTITATIVE 
C0373620|T034||LNC|GLUCOSE; BLOOD, REAGENT STRIP
C0373620|T034||LNC|BLOOD GLUCOSE DETERMINATION BY REAGENT STRIP 
C0373620|T034||LNC|BLOOD GLUCOSE DETERMINATION BY REAGENT STRIP
C0373620|T034||LNC|BLOOD GLUCOSE LEVEL BY REAGENT STRIP
C0373620|T034||LNC|GLUCOSE BLOOD REAGENT STRIP
C0373620|T034||LNC|BLOOD GLUCOSE (SUGAR) MEASUREMENT USING REAGENT STRIP
C0373620|T034||LNC|MEASUREMENT OF GLUCOSE IN BLOOD USING REAGENT STRIP
C0373620|T034||LNC|REAGENT STRIP/BLOOD GLUCOSE
C4064987|T034||LNC|GLUCOSE IN SERUM OR PLASMA 
C4064987|T034||LNC|GLUCOSE IN SERUM OR PLASMA
C0202045|T034||LNC|GLUCOSE MEASUREMENT, FASTING
C0202045|T034||LNC|GLUCOSE MEASUREMENT, FASTING 
C0202045|T034||LNC|FASTING GLUCOSE TEST
C0202045|T034||LNC|TEST;GLUCOSE;FASTING
C0202046|T034||LNC|GLUCOSE MEASUREMENT, RANDOM
C0202046|T034||LNC|GLUCOSE MEASUREMENT, RANDOM 
C0202046|T034||LNC|RANDOM GLUCOSE TEST
C0202046|T034||LNC|TEST;GLUCOSE;RANDOM
C0427743|T034||LNC|GLUCOSE CONCENTRATION
C0427743|T034||LNC|GLUCOSE CONCENTRATION, TEST STRIP MEASUREMENT 
C0427743|T034||LNC|GLUCOSE CONCENTRATION, TEST STRIP MEASUREMENT
C1295145|T034||LNC|GLUCOSE MEASUREMENT ESTIMATED FROM GLYCATED HAEMOGLOBIN
C1295145|T034||LNC|GLUCOSE MEASUREMENT ESTIMATED FROM GLYCATED HEMOGLOBIN 
C1295145|T034||LNC|GLUCOSE MEASUREMENT ESTIMATED FROM GLYCATED HEMOGLOBIN
C2732716|T034||LNC|QUANTITATIVE MEASUREMENT OF MASS CONCENTRATION OF GLUCOSE IN POSTCALORIE FASTING SERUM OR PLASMA SPECIMEN
C2732716|T034||LNC|QUANTITATIVE MEASUREMENT OF MASS CONCENTRATION OF GLUCOSE IN POSTCALORIE FASTING SERUM OR PLASMA
C2732716|T034||LNC|QUANTITATIVE MEASUREMENT OF MASS CONCENTRATION OF GLUCOSE IN POSTCALORIE FASTING SERUM OR PLASMA SPECIMEN 
C0428568|T034||LNC|FASTING BLOOD GLUCOSE MEASUREMENT 
C0428568|T034||LNC|FASTING BLOOD GLUCOSE MEASUREMENT
C0428568|T034||LNC|BLOOD GLUCOSE FASTING
C0428568|T034||LNC|FASTING BLOOD GLUCOSE
C0428568|T034||LNC|FASTING BLOOD GLUCOSE (& LEVEL)
C0428568|T034||LNC|FASTING BLOOD GLUCOSE (& LEVEL) 
C0428568|T034||LNC|FASTING BLOOD GLUCOSE LEVEL
C0428568|T034||LNC|FASTING BLOOD GLUCOSE LEVEL 
C0428568|T034||LNC|FBS - FASTING BLOOD SUGAR
C0428568|T034||LNC|FBG - FASTING BLOOD GLUCOSE
C0428568|T034||LNC|FASTING BLOOD GLUCOSE MEASUREMENT 
C2238123|T034||LNC|FASTING WHOLE BLOOD GLUCOSE MEASUREMENT
C2238123|T034||LNC|FASTING WHOLE BLOOD GLUCOSE MEASUREMENT 
C2238123|T034||LNC|GLUCOSE, FASTING, WHOLE BLOOD
C2238123|T034||LNC|FASTING WHOLE BLOOD GLUCOSE
C2238123|T034||LNC|WHOLE BLOOD FASTING GLUCOSE
C2317664|T034||LNC|FASTING FINGERSTICK BLOOD GLUCOSE
C2317664|T034||LNC|FASTING FINGERSTICK BLOOD GLUCOSE MEASUREMENT
C2317664|T034||LNC|FINGERSTICK BLOOD GLUCOSE FASTING
C2317664|T034||LNC|FASTING FINGERSTICK BLOOD GLUCOSE MEASUREMENT 
C4028983|T034||LNC|FOOTSTICK BLOOD GLUCOSE FASTING 
C4028983|T034||LNC|FOOTSTICK BLOOD GLUCOSE FASTING
