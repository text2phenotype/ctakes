C0524662|T053|191818005|SNOMEDCT_US|OPIATE ADDICTION|UNSPECIFIED OPIOID DEPENDENCE (DISORDER)
C0494376|T053|268686000|SNOMEDCT_US|MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF OPIOIDS, DEPENDENCE SYNDROME|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF OPIOIDS: DEPENDENCE SYNDROME (DISORDER)
C0261864|T053||SNOMEDCT_US|OPIATE ANTAGONISTS CAUSING ADVERSE EFFECTS IN THERAPEUTIC USE
C0261817|T053||SNOMEDCT_US|OTHER OPIATES AND RELATED NARCOTICS CAUSING ADVERSE EFFECTS IN THERAPEUTIC USE
C0747024|T053||SNOMEDCT_US|OPIATE ABUSE OPIUM
C0025605|T053|387286002|SNOMEDCT_US|METHADONE|METHADONE (SUBSTANCE)
C2874436|T053||SNOMEDCT_US|OPIOID DEPENDENCE, UNCOMPLICATED
C2874436|T053||SNOMEDCT_US|OPIOID DEPENDENCE UNCOMPLICATED
C2874436|T053||SNOMEDCT_US|OPIOID DEPENDENCE UNCOMPLICATED 
C0338781|T053|191821007|SNOMEDCT_US|OPIOID DEPENDENCE IN REMISSION |OPIOID DEPENDENCE IN REMISSION (DISORDER)
C0338781|T053|191821007|SNOMEDCT_US|OPIOID DEPENDENCE IN REMISSION|OPIOID DEPENDENCE IN REMISSION (DISORDER)
C0338781|T053|191821007|SNOMEDCT_US|OPIOID DEPENDENCE, IN REMISSION|OPIOID DEPENDENCE IN REMISSION (DISORDER)
C0338781|T053|191821007|SNOMEDCT_US|OPIOID DEPENDENCE IN REMISSION |OPIOID DEPENDENCE IN REMISSION (DISORDER)
C2874441|T053||SNOMEDCT_US|OPIOID DEPENDENCE WITH INTOXICATION
C2874441|T053||SNOMEDCT_US|OPIOID DEPENDENCE WITH INTOXICATION, UNSPECIFIED
C2874441|T053||SNOMEDCT_US|OPIOID DEPENDENCE WITH INTOXICATION 
C2874442|T053||SNOMEDCT_US|OPIOID DEPENDENCE WITH WITHDRAWAL
C2874442|T053||SNOMEDCT_US|OPIOID DEPENDENCE WITH WITHDRAWAL 
C2874443|T053||SNOMEDCT_US|OPIOID DEPENDENCE WITH OPIOID-INDUCED MOOD DISORDER
C2874443|T053||SNOMEDCT_US|OPIOID DEPENDENCE WITH OPIOID-INDUCED MOOD DISORDER 
C2874447|T053||SNOMEDCT_US|OPIOID DEPENDENCE WITH OPIOID-INDUCED PSYCHOTIC DISORDER
C2874447|T053||SNOMEDCT_US|OPIOID DEPENDENCE WITH OPIOID-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED
C2874447|T053||SNOMEDCT_US|OPIOID DEPENDENCE W OPIOID-INDUCED PSYCHOTIC DISORDER, UNSP
C2874447|T053||SNOMEDCT_US|OPIOID DEPENDENCE WITH OPIOID-INDUCED PSYCHOTIC DISORDER 
C2874448|T053||SNOMEDCT_US|OPIOID DEPENDENCE WITH OTHER OPIOID-INDUCED DISORDER
C2874451|T053||SNOMEDCT_US|OPIOID DEPENDENCE WITH UNSPECIFIED OPIOID-INDUCED DISORDER
C0338779|T053|191819002|SNOMEDCT_US|OPIOID DEPENDENCE WITH CONTINUOUS USE |CONTINUOUS OPIOID DEPENDENCE (DISORDER)
C0338779|T053|191819002|SNOMEDCT_US|OPIOID DEPENDENCE WITH CONTINUOUS USE|CONTINUOUS OPIOID DEPENDENCE (DISORDER)
C0338779|T053|191819002|SNOMEDCT_US|CONTINUOUS OPIOID DEPENDENCE|CONTINUOUS OPIOID DEPENDENCE (DISORDER)
C0338779|T053|191819002|SNOMEDCT_US|CONTINUOUS OPIOID DEPENDENCE |CONTINUOUS OPIOID DEPENDENCE (DISORDER)
C0338780|T053|191820008|SNOMEDCT_US|OPIOID DEPENDENCE WITH EPISODIC USE|EPISODIC OPIOID DEPENDENCE (DISORDER)
C0338780|T053|191820008|SNOMEDCT_US|OPIOID DEPENDENCE WITH EPISODIC USE |EPISODIC OPIOID DEPENDENCE (DISORDER)
C0338780|T053|191820008|SNOMEDCT_US|EPISODIC OPIOID DEPENDENCE|EPISODIC OPIOID DEPENDENCE (DISORDER)
C0338780|T053|191820008|SNOMEDCT_US|EPISODIC OPIOID DEPENDENCE |EPISODIC OPIOID DEPENDENCE (DISORDER)
C0338734|T053|191865004|SNOMEDCT_US|OPIOID DEPENDENCE IN COMBINATION WITH ANOTHER DRUG |COMBINED OPIOID WITH NON-OPIOID DRUG DEPENDENCE
C0338734|T053|191865004|SNOMEDCT_US|OPIOID DEPENDENCE IN COMBINATION WITH ANOTHER DRUG|COMBINED OPIOID WITH NON-OPIOID DRUG DEPENDENCE
C0338734|T053|191865004|SNOMEDCT_US|COMBINED OPIOID WITH NON-OPIOID DRUG DEPENDENCE |COMBINED OPIOID WITH NON-OPIOID DRUG DEPENDENCE
C0338734|T053|191865004|SNOMEDCT_US|COMBINED OPIOID WITH OTHER DRUG DEPENDENCE |COMBINED OPIOID WITH NON-OPIOID DRUG DEPENDENCE
C0338734|T053|191865004|SNOMEDCT_US|COMBINED OPIOID WITH NON-OPIOID DRUG DEPENDENCE|COMBINED OPIOID WITH NON-OPIOID DRUG DEPENDENCE
C0338734|T053|191865004|SNOMEDCT_US|COMBINED OPIOID WITH OTHER DRUG DEPENDENCE, UNSPECIFIED|COMBINED OPIOID WITH NON-OPIOID DRUG DEPENDENCE
C0338734|T053|191865004|SNOMEDCT_US|COMBINED OPIOID WITH OTHER DRUG DEPENDENCE, UNSPECIFIED |COMBINED OPIOID WITH NON-OPIOID DRUG DEPENDENCE
C0338734|T053|191865004|SNOMEDCT_US|COMBINED OPIOID WITH OTHER DRUG DEPENDENCE NOS|COMBINED OPIOID WITH NON-OPIOID DRUG DEPENDENCE
C0338734|T053|191865004|SNOMEDCT_US|COMBINED OPIOID WITH OTHER DRUG DEPENDENCE NOS |COMBINED OPIOID WITH NON-OPIOID DRUG DEPENDENCE
C0338734|T053|191865004|SNOMEDCT_US|COMBINED OPIOID WITH OTHER DRUG DEPENDENCE|COMBINED OPIOID WITH NON-OPIOID DRUG DEPENDENCE
C3472691|T053|1081000119105|SNOMEDCT_US|OPIOID DEPENDENCE, ON AGONIST THERAPY |OPIOID DEPENDENCE, ON AGONIST THERAPY (DISORDER)
C3472691|T053|1081000119105|SNOMEDCT_US|OPIOID DEPENDENCE, ON AGONIST THERAPY|OPIOID DEPENDENCE, ON AGONIST THERAPY (DISORDER)
C3472691|T053|1081000119105|SNOMEDCT_US|OPIOID DEPENDENCE, ON AGONIST THERAPY |OPIOID DEPENDENCE, ON AGONIST THERAPY (DISORDER)
C0524662|T053|191818005|SNOMEDCT_US|OPIOID DEPENDENCE|UNSPECIFIED OPIOID DEPENDENCE (DISORDER)
C0524662|T053|191818005|SNOMEDCT_US|DEPENDENCE, OPIATE|UNSPECIFIED OPIOID DEPENDENCE (DISORDER)
C0524662|T053|191818005|SNOMEDCT_US|OPIATE ADDICTION|UNSPECIFIED OPIOID DEPENDENCE (DISORDER)
C0524662|T053|191818005|SNOMEDCT_US|OPIOID DEPENDENCE |UNSPECIFIED OPIOID DEPENDENCE (DISORDER)
C0524662|T053|191818005|SNOMEDCT_US|ADDICTION, OPIATE|UNSPECIFIED OPIOID DEPENDENCE (DISORDER)
C0524662|T053|191818005|SNOMEDCT_US|OPIOID DEPENDENCE-UNSPEC|UNSPECIFIED OPIOID DEPENDENCE (DISORDER)
C0524662|T053|191818005|SNOMEDCT_US|OPIOID TYPE DEPENDENCE, UNSPECIFIED USE|UNSPECIFIED OPIOID DEPENDENCE (DISORDER)
C0524662|T053|191818005|SNOMEDCT_US|OPIOID TYPE DEPENDENCE, UNSPECIFIED|UNSPECIFIED OPIOID DEPENDENCE (DISORDER)
C0524662|T053|191818005|SNOMEDCT_US|[X]DRUG ADDICTION - OPIOIDS|UNSPECIFIED OPIOID DEPENDENCE (DISORDER)
C0524662|T053|191818005|SNOMEDCT_US|UNSPECIFIED OPIOID DEPENDENCE|UNSPECIFIED OPIOID DEPENDENCE (DISORDER)
C0524662|T053|191818005|SNOMEDCT_US|UNSPECIFIED OPIOID DEPENDENCE |UNSPECIFIED OPIOID DEPENDENCE (DISORDER)
C0524662|T053|191818005|SNOMEDCT_US|OPIOID TYPE DRUG DEPENDENCE|UNSPECIFIED OPIOID DEPENDENCE (DISORDER)
C0524662|T053|191818005|SNOMEDCT_US|DEPENDENCE ON OPIATES|UNSPECIFIED OPIOID DEPENDENCE (DISORDER)
C0524662|T053|191818005|SNOMEDCT_US|OPIOID TYPE DEPENDENCE|UNSPECIFIED OPIOID DEPENDENCE (DISORDER)
C0524662|T053|191818005|SNOMEDCT_US|NARCOTISM|UNSPECIFIED OPIOID DEPENDENCE (DISORDER)
C0524662|T053|191818005|SNOMEDCT_US|OPIOID DEPENDENCE |UNSPECIFIED OPIOID DEPENDENCE (DISORDER)
C0524662|T053|191818005|SNOMEDCT_US|DEPENDENCE; OPIATE|UNSPECIFIED OPIOID DEPENDENCE (DISORDER)
C0524662|T053|191818005|SNOMEDCT_US|DEPENDENCE; OPIOIDS|UNSPECIFIED OPIOID DEPENDENCE (DISORDER)
C0524662|T053|191818005|SNOMEDCT_US|OPIOIDS; DEPENDENCE|UNSPECIFIED OPIOID DEPENDENCE (DISORDER)
C0524662|T053|191818005|SNOMEDCT_US|OPIATE DEPENDENCE|UNSPECIFIED OPIOID DEPENDENCE (DISORDER)
C3509112|T053||SNOMEDCT_US|OPIOID DEPENDENCE WITH OPIOID-INDUCED DISORDER
C3509112|T053||SNOMEDCT_US|OPIOID DEPENDENCE WITH OPIOID-INDUCED DISORDER 
C0338782|T053|191822000|SNOMEDCT_US|OPIOID DRUG DEPENDENCE NOS |OPIOID DRUG DEPENDENCE NOS (DISORDER)
C0338782|T053|191822000|SNOMEDCT_US|OPIOID DRUG DEPENDENCE NOS|OPIOID DRUG DEPENDENCE NOS (DISORDER)
C0019337|T053|231477003|SNOMEDCT_US|HEROIN DEPENDENCE|HEROIN DEPENDENCE (DISORDER)
C0019337|T053|231477003|SNOMEDCT_US|ADDICTION, HEROIN|HEROIN DEPENDENCE (DISORDER)
C0019337|T053|231477003|SNOMEDCT_US|DEPENDENCE, HEROIN|HEROIN DEPENDENCE (DISORDER)
C0019337|T053|231477003|SNOMEDCT_US|HEROIN ADDICTION|HEROIN DEPENDENCE (DISORDER)
C0019337|T053|231477003|SNOMEDCT_US|HEROIN DEPENDENCE [DISEASE/FINDING]|HEROIN DEPENDENCE (DISORDER)
C0019337|T053|231477003|SNOMEDCT_US|ADDICTION;DRUG(S);HEROIN|HEROIN DEPENDENCE (DISORDER)
C0019337|T053|231477003|SNOMEDCT_US|[X]HEROIN ADDICTION|HEROIN DEPENDENCE (DISORDER)
C0019337|T053|231477003|SNOMEDCT_US|HEROIN DEPENDENCE |HEROIN DEPENDENCE (DISORDER)
C0019337|T053|231477003|SNOMEDCT_US|OPIOID DEPENDENCE HEROIN|HEROIN DEPENDENCE (DISORDER)
C0019337|T053|231477003|SNOMEDCT_US|HEROIN DEPENDENCE |HEROIN DEPENDENCE (DISORDER)
C0019337|T053|231477003|SNOMEDCT_US|DEPENDENCE; HEROIN|HEROIN DEPENDENCE (DISORDER)
C0019337|T053|231477003|SNOMEDCT_US|HEROIN; DEPENDENCE|HEROIN DEPENDENCE (DISORDER)
C1960518|T053|426001001|SNOMEDCT_US|FENTANYL DEPENDENCE |FENTANYL DEPENDENCE (DISORDER)
C1960518|T053|426001001|SNOMEDCT_US|FENTANYL DEPENDENCE|FENTANYL DEPENDENCE (DISORDER)
C1960518|T053|426001001|SNOMEDCT_US|FENTANYL DEPENDENCE |FENTANYL DEPENDENCE (DISORDER)
C1960518|T053|426001001|SNOMEDCT_US|OPIOID DEPENDENCE FENTANYL|FENTANYL DEPENDENCE (DISORDER)
C0026552|T053|231479000|SNOMEDCT_US|MORPHINE DEPENDENCE|MORPHINE DEPENDENCE (DISORDER)
C0026552|T053|231479000|SNOMEDCT_US|ADDICTION, MORPHINE|MORPHINE DEPENDENCE (DISORDER)
C0026552|T053|231479000|SNOMEDCT_US|DEPENDENCE, MORPHINE|MORPHINE DEPENDENCE (DISORDER)
C0026552|T053|231479000|SNOMEDCT_US|MORPHINE ADDICTION|MORPHINE DEPENDENCE (DISORDER)
C0026552|T053|231479000|SNOMEDCT_US|MORPHINE DEPENDENCE [DISEASE/FINDING]|MORPHINE DEPENDENCE (DISORDER)
C0026552|T053|231479000|SNOMEDCT_US|OPIOID DEPENDENCE MORPHINE|MORPHINE DEPENDENCE (DISORDER)
C0026552|T053|231479000|SNOMEDCT_US|MORPHINE DEPENDENCE |MORPHINE DEPENDENCE (DISORDER)
C0026552|T053|231479000|SNOMEDCT_US|MORPHINE DEPENDENCE |MORPHINE DEPENDENCE (DISORDER)
C0026552|T053|231479000|SNOMEDCT_US|DEPENDENCE; MORPHINE|MORPHINE DEPENDENCE (DISORDER)
C0026552|T053|231479000|SNOMEDCT_US|MORPHINE; DEPENDENCE|MORPHINE DEPENDENCE (DISORDER)
C0026552|T053|231479000|SNOMEDCT_US|MORPHINISM|MORPHINE DEPENDENCE (DISORDER)
C0338776|T053|231478008|SNOMEDCT_US|METHADONE DEPENDENCE|METHADONE DEPENDENCE (DISORDER)
C0338776|T053|231478008|SNOMEDCT_US|OPIOID DEPENDENCE METHADONE|METHADONE DEPENDENCE (DISORDER)
C0338776|T053|231478008|SNOMEDCT_US|METHADONE DEPENDENCE |METHADONE DEPENDENCE (DISORDER)
C0338776|T053|231478008|SNOMEDCT_US|METHADONE DEPENDENCE |METHADONE DEPENDENCE (DISORDER)
C0338776|T053|231478008|SNOMEDCT_US|DEPENDENCE; METHADONE|METHADONE DEPENDENCE (DISORDER)
C0338776|T053|231478008|SNOMEDCT_US|METHADONE; DEPENDENCE|METHADONE DEPENDENCE (DISORDER)
C0338777|T053|231480002|SNOMEDCT_US|OPIUM DEPENDENCE|OPIUM DEPENDENCE (DISORDER)
C0338777|T053|231480002|SNOMEDCT_US|OPIUM DEPENDENCE |OPIUM DEPENDENCE (DISORDER)
C0338777|T053|231480002|SNOMEDCT_US|OPIOID DEPENDENCE OPIUM|OPIUM DEPENDENCE (DISORDER)
C0338777|T053|231480002|SNOMEDCT_US|OPIUM DEPENDENCE |OPIUM DEPENDENCE (DISORDER)
C0338777|T053|231480002|SNOMEDCT_US|DEPENDENCE; OPIUM|OPIUM DEPENDENCE (DISORDER)
C3840144|T053|703845008|SNOMEDCT_US|BUPRENORPHINE DEPENDENCE |BUPRENORPHINE DEPENDENCE (DISORDER)
C3840144|T053|703845008|SNOMEDCT_US|BUPRENORPHINE DEPENDENCE|BUPRENORPHINE DEPENDENCE (DISORDER)
C0154478|T053||SNOMEDCT_US|OPIOID DEPENDENCE-CONTIN
C0154478|T053||SNOMEDCT_US|OPIOID TYPE DEPENDENCE, CONTINUOUS
C0154478|T053||SNOMEDCT_US|OPIOID TYPE DEPENDENCE, CONTINUOUS USE
C0154479|T053||SNOMEDCT_US|OPIOID DEPENDENCE-EPISOD
C0154479|T053||SNOMEDCT_US|OPIOID TYPE DEPENDENCE, EPISODIC
C0154479|T053||SNOMEDCT_US|OPIOID TYPE DEPENDENCE, EPISODIC USE
C0154480|T053||SNOMEDCT_US|OPIOID DEPENDENCE-REMISS
C0154480|T053||SNOMEDCT_US|OPIOID TYPE DEPENDENCE, IN REMISSION
C0494376|T053|268686000|SNOMEDCT_US|MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF OPIOIDS, DEPENDENCE SYNDROME|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF OPIOIDS: DEPENDENCE SYNDROME (DISORDER)
C0494376|T053|268686000|SNOMEDCT_US|MENTAL AND BEHAVIOURAL DISORDERS DUE TO USE OF OPIOIDS, DEPENDENCE SYNDROME|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF OPIOIDS: DEPENDENCE SYNDROME (DISORDER)
C0494376|T053|268686000|SNOMEDCT_US|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF OPIOIDS: DEPENDENCE SYNDROME|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF OPIOIDS: DEPENDENCE SYNDROME (DISORDER)
C0494376|T053|268686000|SNOMEDCT_US|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF OPIOIDS: DEPENDENCE SYNDROME |[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF OPIOIDS: DEPENDENCE SYNDROME (DISORDER)
C0494376|T053|268686000|SNOMEDCT_US|[X]MENTAL AND BEHAVIOURAL DISORDERS DUE TO USE OF OPIOIDS: DEPENDENCE SYNDROME|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF OPIOIDS: DEPENDENCE SYNDROME (DISORDER)
C0494376|T053|268686000|SNOMEDCT_US|OPIUMISM|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF OPIOIDS: DEPENDENCE SYNDROME (DISORDER)
C0865342|T053||SNOMEDCT_US|OPIUM ALKALOIDS AND THEIR DERIVATIVES DEPENDENCE
C1386557|T053||SNOMEDCT_US|CODEINE; DEPENDENCE
C1386557|T053||SNOMEDCT_US|DEPENDENCE; CODEINE
C1386560|T053||SNOMEDCT_US|DEPENDENCE; DEXTROMETHORPHAN
C1386560|T053||SNOMEDCT_US|DEXTROMETHORPHAN; DEPENDENCE
C1386561|T053||SNOMEDCT_US|DEPENDENCE; DEXTROMORAMIDE
C1386561|T053||SNOMEDCT_US|DEXTROMORAMIDE; DEPENDENCE
C1386562|T053||SNOMEDCT_US|DEPENDENCE; DEXTRORPHAN
C1386562|T053||SNOMEDCT_US|DEXTRORPHAN; DEPENDENCE
C1386566|T053||SNOMEDCT_US|DEPENDENCE; ETHYLMORPHINE
C1386566|T053||SNOMEDCT_US|ETHYLMORPHINE; DEPENDENCE
C1386570|T053||SNOMEDCT_US|DEPENDENCE; DRUG, SYNTHETIC, WITH MORPHINE-LIKE EFFECT
C1386577|T053||SNOMEDCT_US|DEPENDENCE; LAUDANUM
C1386577|T053||SNOMEDCT_US|LAUDANUM; DEPENDENCE
C1386588|T053||SNOMEDCT_US|DEPENDENCE; METHYL MORPHINE
C1386588|T053||SNOMEDCT_US|METHYL MORPHINE; DEPENDENCE
C1386594|T053||SNOMEDCT_US|DEPENDENCE; PAREGORIC
C1386594|T053||SNOMEDCT_US|PAREGORIC; DEPENDENCE
C1404354|T053||SNOMEDCT_US|MORPHINOMANIA
C0025607|T053||SNOMEDCT_US|METHADYL ACETATE
C0025607|T053||SNOMEDCT_US|METHADYLACETATE
C0025607|T053||SNOMEDCT_US|ACETYLMETHADOL
C0699057|T053||SNOMEDCT_US|BRAND OF METHADONE
C0699057|T053||SNOMEDCT_US|ROXANE BRAND OF METHADONE HYDROCHLORIDE
C0699061|T053||SNOMEDCT_US|AMIDONE
C0699061|T053||SNOMEDCT_US|AMIDINE
C0699061|T053||SNOMEDCT_US|AMIDONE BRAND OF METHADONE
C0730805|T053||SNOMEDCT_US|PINADONE
C0730805|T053||SNOMEDCT_US|PINEWOOD BRAND OF METHADONE HYDROCHLORIDE
C0788510|T053||SNOMEDCT_US|NORMETHADONE 10 MG/ML / OXILOFRINE 20 MG/ML ORAL SOLUTION
C0116497|T053||SNOMEDCT_US|ERYTHRO-5-METHYLMETHADONE
C0145747|T053||SNOMEDCT_US|THREO-5-METHYLMETHADONE
C0592779|T053||SNOMEDCT_US|METHADOSE
C0592779|T053||SNOMEDCT_US|MALLINCKRODT BRAND OF METHADONE HYDROCHLORIDE
C0592779|T053||SNOMEDCT_US|ROSEMONT BRAND OF METHADONE HYDROCHLORIDE
C0594373|T053||SNOMEDCT_US|METHEX
C0594373|T053||SNOMEDCT_US|GENERICS BRAND OF METHADONE HYDROCHLORIDE
C0025605|T053|387286002|SNOMEDCT_US|METHADONE|METHADONE (SUBSTANCE)
C0025605|T053|387286002|SNOMEDCT_US|3-HEPTANONE, 6-(DIMETHYLAMINO)-4,4-DIPHENYL-|METHADONE (SUBSTANCE)
C0025605|T053|387286002|SNOMEDCT_US|METHADONE [CHEMICAL/INGREDIENT]|METHADONE (SUBSTANCE)
C0025605|T053|387286002|SNOMEDCT_US|METHADONE |METHADONE (SUBSTANCE)
C0025605|T053|387286002|SNOMEDCT_US|METHADONE |METHADONE (SUBSTANCE)
C0981584|T053|322591003|SNOMEDCT_US|METHADONE HYDROCHLORIDE 5MG ORAL TABLET|METHADONE HYDROCHLORIDE 5MG TABLET (SUBSTANCE)
C0981584|T053|322591003|SNOMEDCT_US|METHADONE HYDROCHLORIDE, 5 MG ORAL TABLET|METHADONE HYDROCHLORIDE 5MG TABLET (SUBSTANCE)
C0981584|T053|322591003|SNOMEDCT_US|METHADONE 5 MG ORAL TABLET|METHADONE HYDROCHLORIDE 5MG TABLET (SUBSTANCE)
C0981584|T053|322591003|SNOMEDCT_US|METHADONE HCL 5MG EFFERVSC TAB|METHADONE HYDROCHLORIDE 5MG TABLET (SUBSTANCE)
C0981584|T053|322591003|SNOMEDCT_US|METHADONE HCL 5MG TAB|METHADONE HYDROCHLORIDE 5MG TABLET (SUBSTANCE)
C0981584|T053|322591003|SNOMEDCT_US|METHADONE HCL TAB 5 MG|METHADONE HYDROCHLORIDE 5MG TABLET (SUBSTANCE)
C0981584|T053|322591003|SNOMEDCT_US|METHADONE HYDROCHLORIDE 5 MG ORAL TABLET|METHADONE HYDROCHLORIDE 5MG TABLET (SUBSTANCE)
C0981584|T053|322591003|SNOMEDCT_US|METHADONE HCL 5MG TAB [VA PRODUCT]|METHADONE HYDROCHLORIDE 5MG TABLET (SUBSTANCE)
C0981584|T053|322591003|SNOMEDCT_US|METHADONE HCL 5MG TAB,EFFERVSC|METHADONE HYDROCHLORIDE 5MG TABLET (SUBSTANCE)
C0981584|T053|322591003|SNOMEDCT_US|METHADONE HCL 5MG TAB,EFFERVSC [VA PRODUCT]|METHADONE HYDROCHLORIDE 5MG TABLET (SUBSTANCE)
C0981584|T053|322591003|SNOMEDCT_US|METHADONE HCL 5 MG ORAL TABLET|METHADONE HYDROCHLORIDE 5MG TABLET (SUBSTANCE)
C0981584|T053|322591003|SNOMEDCT_US|METHADONE HYDROCHLORIDE 5MG TABLET|METHADONE HYDROCHLORIDE 5MG TABLET (SUBSTANCE)
C0981584|T053|322591003|SNOMEDCT_US|METHADONE HYDROCHLORIDE 5MG TABLET |METHADONE HYDROCHLORIDE 5MG TABLET (SUBSTANCE)
C0981584|T053|322591003|SNOMEDCT_US|METHADONE HYDROCHLORIDE 5MG TABLET |METHADONE HYDROCHLORIDE 5MG TABLET (SUBSTANCE)
C0721688|T053|23883005|SNOMEDCT_US|METHADONE HYDROCHLORIDE|METHADONE HYDROCHLORIDE (SUBSTANCE)
C0721688|T053|23883005|SNOMEDCT_US|METHADONE HYDROCHLORIDE |METHADONE HYDROCHLORIDE (SUBSTANCE)
C0721688|T053|23883005|SNOMEDCT_US|HYDROCHLORIDE, METHADONE|METHADONE HYDROCHLORIDE (SUBSTANCE)
C0721688|T053|23883005|SNOMEDCT_US|METHADONE HYDROCHLORIDE [CHEMICAL/INGREDIENT]|METHADONE HYDROCHLORIDE (SUBSTANCE)
C0721688|T053|23883005|SNOMEDCT_US|METHADONE HCL [ANALGESIC]|METHADONE HYDROCHLORIDE (SUBSTANCE)
C0721688|T053|23883005|SNOMEDCT_US|METHADONE HCL [COUGH] |METHADONE HYDROCHLORIDE (SUBSTANCE)
C0721688|T053|23883005|SNOMEDCT_US|METHADONE HCL [ANALGESIC] |METHADONE HYDROCHLORIDE (SUBSTANCE)
C0721688|T053|23883005|SNOMEDCT_US|METHADONE HCL [COUGH]|METHADONE HYDROCHLORIDE (SUBSTANCE)
C0721688|T053|23883005|SNOMEDCT_US|METHADONE HYDROCHLORIDE |METHADONE HYDROCHLORIDE (SUBSTANCE)
C0721688|T053|23883005|SNOMEDCT_US|METHADONE HCL [ANALGESIC] |METHADONE HYDROCHLORIDE (SUBSTANCE)
C0721688|T053|23883005|SNOMEDCT_US|METHADONE HCL [COUGH] |METHADONE HYDROCHLORIDE (SUBSTANCE)
C2093101|T053||SNOMEDCT_US|METHADONE HYDROCHLORIDE (DOLOPHINE) INJECTION
C2093101|T053||SNOMEDCT_US|METHADONE HYDROCHLORIDE INJECTION
C2093101|T053||SNOMEDCT_US|METHADONE HYDROCHLORIDE INJECTION 
C1992369|T053||SNOMEDCT_US|METHADONE &#X7C; BLD-SER-PLAS
C1992375|T053||SNOMEDCT_US|METHADONE &#X7C; STOOL
C1992378|T053||SNOMEDCT_US|METHADONE &#X7C; XXX
C1992373|T053||SNOMEDCT_US|METHADONE &#X7C; MECONIUM
C1626306|T053||SNOMEDCT_US|METHADONE+METABOLITE
C1992383|T053||SNOMEDCT_US|METHADONE.R &#X7C; BLD-SER-PLAS
C1992377|T053||SNOMEDCT_US|METHADONE &#X7C; VITREOUS FLUID
C1992374|T053||SNOMEDCT_US|METHADONE &#X7C; MILK
C1992368|T053||SNOMEDCT_US|METHADONE &#124; BILE FLUID
C1992368|T053||SNOMEDCT_US|METHADONE &#X7C; BILE FLUID
C3534187|T053||SNOMEDCT_US|METHADONE &#X7C; SALIVA
C0366544|T053||SNOMEDCT_US|METHADONE DOSE
C0366544|T053||SNOMEDCT_US|METHADONE:MASS:PT:DOSE:QN
C0366544|T053||SNOMEDCT_US|METHADONE [MASS] OF DOSE
C0366544|T053||SNOMEDCT_US|METHADONE:MASS:POINT IN TIME:DOSE MED OR SUBSTANCE:QUANTITATIVE
C1992376|T053||SNOMEDCT_US|METHADONE &#X7C; URINE
C0046103|T053|725546006|SNOMEDCT_US|1,5-DIMETHYL-3,3-DIPHENYL-2-ETHYLIDENEPYRROLIDINE|2-ETHYLIDENE-1,5-DIMETHYL-3,3-DIPHENYLPYRROLIDINE (SUBSTANCE)
C0046103|T053|725546006|SNOMEDCT_US|2-ETHYLIDENE-1,5-DIMETHYL-3,3-DIPHENYLPYRROLIDINE|2-ETHYLIDENE-1,5-DIMETHYL-3,3-DIPHENYLPYRROLIDINE (SUBSTANCE)
C0046103|T053|725546006|SNOMEDCT_US|EDPP|2-ETHYLIDENE-1,5-DIMETHYL-3,3-DIPHENYLPYRROLIDINE (SUBSTANCE)
C0046103|T053|725546006|SNOMEDCT_US|2-ET-1,5-DIME-3,3-DPP|2-ETHYLIDENE-1,5-DIMETHYL-3,3-DIPHENYLPYRROLIDINE (SUBSTANCE)
C0046103|T053|725546006|SNOMEDCT_US|EDDP-3,3|2-ETHYLIDENE-1,5-DIMETHYL-3,3-DIPHENYLPYRROLIDINE (SUBSTANCE)
C1992371|T053||SNOMEDCT_US|METHADONE &#X7C; GASTRIC FLUID
C1992372|T053||SNOMEDCT_US|METHADONE &#X7C; HAIR
C0628179|T053||SNOMEDCT_US|6-DIMETHYLAMINO-4-(4-HYDROXYPHENYL)-4-PHENYLHEPTAN-3-ONE
C0628179|T053||SNOMEDCT_US|PARA-HYDROXYMETHADONE
C0624343|T053||SNOMEDCT_US|2-FORMAMIDO-4,4-DIPHENYL-5-HEPTANONE
C0069008|T053||SNOMEDCT_US|6-DIMETHYLAMINO-4,4-DIPHENYLHEXAN-3-ONE
C0069008|T053||SNOMEDCT_US|NOR-METHADONE
C0069008|T053||SNOMEDCT_US|NORMETHADONE
C0360477|T053|350295000|SNOMEDCT_US|ORAL METHADONE|ORAL FORM METHADONE (PRODUCT)
C0360477|T053|350295000|SNOMEDCT_US|METHADONE ORAL PRODUCT|ORAL FORM METHADONE (PRODUCT)
C0360477|T053|350295000|SNOMEDCT_US|ORAL FORM METHADONE |ORAL FORM METHADONE (PRODUCT)
C0360477|T053|350295000|SNOMEDCT_US|ORAL FORM METHADONE|ORAL FORM METHADONE (PRODUCT)
C0360477|T053|350295000|SNOMEDCT_US|ORAL METHADONE |ORAL FORM METHADONE (PRODUCT)
C0360477|T053|350295000|SNOMEDCT_US|ORAL METHADONE |ORAL FORM METHADONE (PRODUCT)
C0360478|T053|350296004|SNOMEDCT_US|PARENTERAL METHADONE|PARENTERAL FORM METHADONE (PRODUCT)
C0360478|T053|350296004|SNOMEDCT_US|PARENTERAL FORM METHADONE |PARENTERAL FORM METHADONE (PRODUCT)
C0360478|T053|350296004|SNOMEDCT_US|PARENTERAL FORM METHADONE|PARENTERAL FORM METHADONE (PRODUCT)
C0360478|T053|350296004|SNOMEDCT_US|PARENTERAL METHADONE |PARENTERAL FORM METHADONE (PRODUCT)
C0360478|T053|350296004|SNOMEDCT_US|PARENTERAL METHADONE |PARENTERAL FORM METHADONE (PRODUCT)
C0684217|T053||SNOMEDCT_US|PHYSEPTONE
C0684217|T053||SNOMEDCT_US|MARTINDALE BRAND OF METHADONE HYDROCHLORIDE
C0684217|T053||SNOMEDCT_US|PHYMET
C0684217|T053||SNOMEDCT_US|GLAXOSMITHKLINE BRAND OF METHADONE HYDROCHLORIDE
C1563840|T053||SNOMEDCT_US|BIOMET BRAND OF METHADONE HYDROCHLORIDE
C1563840|T053||SNOMEDCT_US|BIODONE
C1563841|T053||SNOMEDCT_US|PHARMASCIENCE BRAND OF METHADONE HYDROCHLORIDE
C1563841|T053||SNOMEDCT_US|METADOL
C1563842|T053||SNOMEDCT_US|ESTEVE BRAND OF METHADONE HYDROCHLORIDE
C1563842|T053||SNOMEDCT_US|METASEDIN
C1563843|T053||SNOMEDCT_US|ADDICARE BRAND OF METHADONE HYDROCHLORIDE
C1563843|T053||SNOMEDCT_US|METHADDICT
C1563844|T053||SNOMEDCT_US|YAMANOUCHI BRAND OF METHADONE HYDROCHLORIDE
C1563844|T053||SNOMEDCT_US|SYMORON
C0731186|T053||SNOMEDCT_US|MARTINDALE METHADONE DTF
